magic
tech sky130A
magscale 1 2
timestamp 1733616469
<< viali >>
rect 3341 43401 3375 43435
rect 3985 43401 4019 43435
rect 4445 43401 4479 43435
rect 5181 43401 5215 43435
rect 5917 43401 5951 43435
rect 6653 43401 6687 43435
rect 7389 43401 7423 43435
rect 8125 43401 8159 43435
rect 9137 43401 9171 43435
rect 9597 43401 9631 43435
rect 10333 43401 10367 43435
rect 11069 43401 11103 43435
rect 11805 43401 11839 43435
rect 12541 43401 12575 43435
rect 13277 43401 13311 43435
rect 13829 43401 13863 43435
rect 1501 43265 1535 43299
rect 2053 43265 2087 43299
rect 2697 43265 2731 43299
rect 3157 43265 3191 43299
rect 3801 43265 3835 43299
rect 4353 43265 4387 43299
rect 4997 43265 5031 43299
rect 5733 43265 5767 43299
rect 6469 43265 6503 43299
rect 7205 43265 7239 43299
rect 7941 43265 7975 43299
rect 8953 43265 8987 43299
rect 9413 43265 9447 43299
rect 10149 43265 10183 43299
rect 10977 43265 11011 43299
rect 11621 43265 11655 43299
rect 12449 43265 12483 43299
rect 13093 43265 13127 43299
rect 13553 43265 13587 43299
rect 2237 43129 2271 43163
rect 1593 43061 1627 43095
rect 2789 43061 2823 43095
rect 2881 42857 2915 42891
rect 3249 42857 3283 42891
rect 4077 42857 4111 42891
rect 4813 42857 4847 42891
rect 6285 42857 6319 42891
rect 7021 42857 7055 42891
rect 7757 42857 7791 42891
rect 8493 42857 8527 42891
rect 9229 42857 9263 42891
rect 9873 42857 9907 42891
rect 10701 42857 10735 42891
rect 11437 42857 11471 42891
rect 12173 42857 12207 42891
rect 13645 42857 13679 42891
rect 13461 42721 13495 42755
rect 3433 42653 3467 42687
rect 4261 42653 4295 42687
rect 4997 42653 5031 42687
rect 6469 42653 6503 42687
rect 7205 42653 7239 42687
rect 7941 42653 7975 42687
rect 8677 42653 8711 42687
rect 9413 42653 9447 42687
rect 10057 42653 10091 42687
rect 10885 42653 10919 42687
rect 11621 42653 11655 42687
rect 12357 42653 12391 42687
rect 13829 42653 13863 42687
rect 1409 42585 1443 42619
rect 9689 42585 9723 42619
rect 13185 42585 13219 42619
rect 10333 42517 10367 42551
rect 1961 42313 1995 42347
rect 4077 42313 4111 42347
rect 4721 42313 4755 42347
rect 13369 42313 13403 42347
rect 13829 42313 13863 42347
rect 2145 42177 2179 42211
rect 4261 42177 4295 42211
rect 4905 42177 4939 42211
rect 13553 42177 13587 42211
rect 13737 42177 13771 42211
rect 13093 42109 13127 42143
rect 13093 41769 13127 41803
rect 13645 41769 13679 41803
rect 13277 41565 13311 41599
rect 13829 41565 13863 41599
rect 1409 41089 1443 41123
rect 1593 40885 1627 40919
rect 1501 40069 1535 40103
rect 13461 40001 13495 40035
rect 13829 40001 13863 40035
rect 1685 39865 1719 39899
rect 13277 39797 13311 39831
rect 14105 39797 14139 39831
rect 9505 39593 9539 39627
rect 7757 39525 7791 39559
rect 8953 39525 8987 39559
rect 7941 39389 7975 39423
rect 8585 39389 8619 39423
rect 9137 39389 9171 39423
rect 9689 39389 9723 39423
rect 12909 39389 12943 39423
rect 1501 39321 1535 39355
rect 1869 39321 1903 39355
rect 13369 39321 13403 39355
rect 13737 39321 13771 39355
rect 8401 39253 8435 39287
rect 13093 39253 13127 39287
rect 12449 39049 12483 39083
rect 12633 38913 12667 38947
rect 12909 38913 12943 38947
rect 13093 38913 13127 38947
rect 13645 38913 13679 38947
rect 12725 38709 12759 38743
rect 13369 38709 13403 38743
rect 13921 38709 13955 38743
rect 12357 38505 12391 38539
rect 12081 38437 12115 38471
rect 1409 38301 1443 38335
rect 12265 38301 12299 38335
rect 12541 38301 12575 38335
rect 12817 38301 12851 38335
rect 12909 38301 12943 38335
rect 13369 38233 13403 38267
rect 13737 38233 13771 38267
rect 1593 38165 1627 38199
rect 12633 38165 12667 38199
rect 13093 38165 13127 38199
rect 11529 37961 11563 37995
rect 11897 37961 11931 37995
rect 12173 37961 12207 37995
rect 12449 37961 12483 37995
rect 13185 37893 13219 37927
rect 13737 37893 13771 37927
rect 1409 37825 1443 37859
rect 11161 37825 11195 37859
rect 11713 37825 11747 37859
rect 12081 37825 12115 37859
rect 12357 37825 12391 37859
rect 12633 37825 12667 37859
rect 12725 37825 12759 37859
rect 13553 37825 13587 37859
rect 1593 37621 1627 37655
rect 10977 37621 11011 37655
rect 12909 37621 12943 37655
rect 14013 37621 14047 37655
rect 10333 37417 10367 37451
rect 12265 37349 12299 37383
rect 10517 37213 10551 37247
rect 11897 37213 11931 37247
rect 12173 37213 12207 37247
rect 12449 37213 12483 37247
rect 12725 37213 12759 37247
rect 13001 37213 13035 37247
rect 13369 37145 13403 37179
rect 13553 37145 13587 37179
rect 11713 37077 11747 37111
rect 11989 37077 12023 37111
rect 12541 37077 12575 37111
rect 13645 37077 13679 37111
rect 1593 36873 1627 36907
rect 12265 36873 12299 36907
rect 13737 36805 13771 36839
rect 1409 36737 1443 36771
rect 1961 36737 1995 36771
rect 11897 36737 11931 36771
rect 12173 36737 12207 36771
rect 12449 36737 12483 36771
rect 12725 36737 12759 36771
rect 13185 36737 13219 36771
rect 13553 36737 13587 36771
rect 1777 36601 1811 36635
rect 11713 36601 11747 36635
rect 11989 36533 12023 36567
rect 12909 36533 12943 36567
rect 14013 36533 14047 36567
rect 1961 36329 1995 36363
rect 11897 36329 11931 36363
rect 11345 36261 11379 36295
rect 1777 36193 1811 36227
rect 2145 36125 2179 36159
rect 11529 36125 11563 36159
rect 11805 36125 11839 36159
rect 12081 36125 12115 36159
rect 12817 36125 12851 36159
rect 1501 36057 1535 36091
rect 12265 36057 12299 36091
rect 12633 36057 12667 36091
rect 13185 36057 13219 36091
rect 13369 36057 13403 36091
rect 13737 36057 13771 36091
rect 11621 35989 11655 36023
rect 10241 35785 10275 35819
rect 10609 35785 10643 35819
rect 10885 35785 10919 35819
rect 11161 35785 11195 35819
rect 13185 35717 13219 35751
rect 9505 35649 9539 35683
rect 10425 35649 10459 35683
rect 10793 35649 10827 35683
rect 11069 35649 11103 35683
rect 11345 35649 11379 35683
rect 11805 35649 11839 35683
rect 12081 35649 12115 35683
rect 12173 35649 12207 35683
rect 12633 35649 12667 35683
rect 13737 35649 13771 35683
rect 14105 35649 14139 35683
rect 9321 35513 9355 35547
rect 11621 35513 11655 35547
rect 12357 35513 12391 35547
rect 11897 35445 11931 35479
rect 12909 35445 12943 35479
rect 13461 35445 13495 35479
rect 5549 35241 5583 35275
rect 8953 35241 8987 35275
rect 9505 35241 9539 35275
rect 10793 35241 10827 35275
rect 11069 35241 11103 35275
rect 1409 35037 1443 35071
rect 5733 35037 5767 35071
rect 9137 35037 9171 35071
rect 9689 35037 9723 35071
rect 10977 35037 11011 35071
rect 11253 35037 11287 35071
rect 11529 35037 11563 35071
rect 11803 35027 11837 35061
rect 13093 35037 13127 35071
rect 13369 34969 13403 35003
rect 1593 34901 1627 34935
rect 12541 34901 12575 34935
rect 12909 34901 12943 34935
rect 13645 34901 13679 34935
rect 1593 34697 1627 34731
rect 5549 34697 5583 34731
rect 10609 34697 10643 34731
rect 12725 34697 12759 34731
rect 1409 34561 1443 34595
rect 5733 34561 5767 34595
rect 10793 34561 10827 34595
rect 10977 34561 11011 34595
rect 11345 34561 11379 34595
rect 11955 34561 11989 34595
rect 13277 34561 13311 34595
rect 13829 34561 13863 34595
rect 14197 34561 14231 34595
rect 11713 34493 11747 34527
rect 13369 34357 13403 34391
rect 10425 34153 10459 34187
rect 10977 34153 11011 34187
rect 11253 34153 11287 34187
rect 11529 34153 11563 34187
rect 10701 34085 10735 34119
rect 13277 34017 13311 34051
rect 10057 33949 10091 33983
rect 10333 33949 10367 33983
rect 10609 33949 10643 33983
rect 10885 33945 10919 33979
rect 11161 33949 11195 33983
rect 11437 33949 11471 33983
rect 11713 33949 11747 33983
rect 11897 33881 11931 33915
rect 12265 33881 12299 33915
rect 12449 33881 12483 33915
rect 13001 33881 13035 33915
rect 13553 33881 13587 33915
rect 9873 33813 9907 33847
rect 10149 33813 10183 33847
rect 12725 33813 12759 33847
rect 13829 33813 13863 33847
rect 10425 33609 10459 33643
rect 1409 33473 1443 33507
rect 10609 33473 10643 33507
rect 10885 33473 10919 33507
rect 11345 33473 11379 33507
rect 11803 33483 11837 33517
rect 13185 33473 13219 33507
rect 13737 33473 13771 33507
rect 11529 33405 11563 33439
rect 11161 33337 11195 33371
rect 1593 33269 1627 33303
rect 10701 33269 10735 33303
rect 12541 33269 12575 33303
rect 13461 33269 13495 33303
rect 14013 33269 14047 33303
rect 10425 33065 10459 33099
rect 11529 32929 11563 32963
rect 13277 32929 13311 32963
rect 1409 32861 1443 32895
rect 10333 32861 10367 32895
rect 10609 32861 10643 32895
rect 10885 32861 10919 32895
rect 11771 32861 11805 32895
rect 11069 32793 11103 32827
rect 13001 32793 13035 32827
rect 13553 32793 13587 32827
rect 13921 32793 13955 32827
rect 1593 32725 1627 32759
rect 10149 32725 10183 32759
rect 10701 32725 10735 32759
rect 11345 32725 11379 32759
rect 12541 32725 12575 32759
rect 10517 32521 10551 32555
rect 13461 32521 13495 32555
rect 13001 32453 13035 32487
rect 9379 32385 9413 32419
rect 10701 32385 10735 32419
rect 10977 32385 11011 32419
rect 11771 32385 11805 32419
rect 13645 32385 13679 32419
rect 13829 32385 13863 32419
rect 9137 32317 9171 32351
rect 11529 32317 11563 32351
rect 10149 32181 10183 32215
rect 11253 32181 11287 32215
rect 12541 32181 12575 32215
rect 13277 32181 13311 32215
rect 14105 32181 14139 32215
rect 9505 31977 9539 32011
rect 10793 31977 10827 32011
rect 11161 31977 11195 32011
rect 12633 31977 12667 32011
rect 9965 31909 9999 31943
rect 10241 31909 10275 31943
rect 7481 31841 7515 31875
rect 1409 31773 1443 31807
rect 7755 31773 7789 31807
rect 9689 31773 9723 31807
rect 10149 31773 10183 31807
rect 10425 31773 10459 31807
rect 10701 31773 10735 31807
rect 10977 31773 11011 31807
rect 11345 31773 11379 31807
rect 11713 31773 11747 31807
rect 13277 31773 13311 31807
rect 12081 31705 12115 31739
rect 12357 31705 12391 31739
rect 12909 31705 12943 31739
rect 13461 31705 13495 31739
rect 13829 31705 13863 31739
rect 1593 31637 1627 31671
rect 8493 31637 8527 31671
rect 10517 31637 10551 31671
rect 9873 31433 9907 31467
rect 9965 31433 9999 31467
rect 13553 31433 13587 31467
rect 10977 31365 11011 31399
rect 1409 31297 1443 31331
rect 8953 31297 8987 31331
rect 9229 31297 9263 31331
rect 10149 31297 10183 31331
rect 10701 31297 10735 31331
rect 12909 31297 12943 31331
rect 13737 31297 13771 31331
rect 8033 31229 8067 31263
rect 8217 31229 8251 31263
rect 9070 31229 9104 31263
rect 11713 31229 11747 31263
rect 11897 31229 11931 31263
rect 12357 31229 12391 31263
rect 12633 31229 12667 31263
rect 12750 31229 12784 31263
rect 8677 31161 8711 31195
rect 10517 31161 10551 31195
rect 1593 31093 1627 31127
rect 11253 31093 11287 31127
rect 14013 31093 14047 31127
rect 8309 30889 8343 30923
rect 12449 30821 12483 30855
rect 13645 30821 13679 30855
rect 7297 30753 7331 30787
rect 8953 30753 8987 30787
rect 10425 30753 10459 30787
rect 7539 30685 7573 30719
rect 9211 30685 9245 30719
rect 10699 30685 10733 30719
rect 11805 30685 11839 30719
rect 11989 30685 12023 30719
rect 12725 30685 12759 30719
rect 12842 30685 12876 30719
rect 13001 30685 13035 30719
rect 13921 30685 13955 30719
rect 9965 30549 9999 30583
rect 11437 30549 11471 30583
rect 13737 30549 13771 30583
rect 10885 30277 10919 30311
rect 13829 30277 13863 30311
rect 1409 30209 1443 30243
rect 10241 30209 10275 30243
rect 13185 30209 13219 30243
rect 14105 30209 14139 30243
rect 9045 30141 9079 30175
rect 9229 30141 9263 30175
rect 9689 30141 9723 30175
rect 9965 30141 9999 30175
rect 10082 30141 10116 30175
rect 11989 30141 12023 30175
rect 12173 30141 12207 30175
rect 12633 30141 12667 30175
rect 12909 30141 12943 30175
rect 13026 30141 13060 30175
rect 13921 30073 13955 30107
rect 1593 30005 1627 30039
rect 2145 29801 2179 29835
rect 6101 29665 6135 29699
rect 12633 29665 12667 29699
rect 1409 29597 1443 29631
rect 1961 29597 1995 29631
rect 6359 29567 6393 29601
rect 10333 29597 10367 29631
rect 10607 29597 10641 29631
rect 12875 29597 12909 29631
rect 9873 29529 9907 29563
rect 10241 29529 10275 29563
rect 12173 29529 12207 29563
rect 1593 29461 1627 29495
rect 7113 29461 7147 29495
rect 11345 29461 11379 29495
rect 12265 29461 12299 29495
rect 13645 29461 13679 29495
rect 7113 29121 7147 29155
rect 7387 29121 7421 29155
rect 8767 29121 8801 29155
rect 10147 29121 10181 29155
rect 12047 29121 12081 29155
rect 13553 29121 13587 29155
rect 8493 29053 8527 29087
rect 9873 29053 9907 29087
rect 11805 29053 11839 29087
rect 9505 28985 9539 29019
rect 13829 28985 13863 29019
rect 8125 28917 8159 28951
rect 10885 28917 10919 28951
rect 12817 28917 12851 28951
rect 1593 28713 1627 28747
rect 11529 28645 11563 28679
rect 12725 28645 12759 28679
rect 7113 28577 7147 28611
rect 11805 28577 11839 28611
rect 13185 28577 13219 28611
rect 1409 28509 1443 28543
rect 7355 28509 7389 28543
rect 10885 28509 10919 28543
rect 11069 28509 11103 28543
rect 11922 28509 11956 28543
rect 12081 28509 12115 28543
rect 12909 28441 12943 28475
rect 13461 28441 13495 28475
rect 8125 28373 8159 28407
rect 10517 28373 10551 28407
rect 13737 28373 13771 28407
rect 8861 28169 8895 28203
rect 14197 28169 14231 28203
rect 11621 28101 11655 28135
rect 1409 28033 1443 28067
rect 7021 28033 7055 28067
rect 8217 28033 8251 28067
rect 9137 28033 9171 28067
rect 9990 28033 10024 28067
rect 10149 28033 10183 28067
rect 10977 28033 11011 28067
rect 12541 28033 12575 28067
rect 13553 28033 13587 28067
rect 7205 27965 7239 27999
rect 7665 27965 7699 27999
rect 7941 27965 7975 27999
rect 8079 27965 8113 27999
rect 8953 27965 8987 27999
rect 9873 27965 9907 27999
rect 12357 27965 12391 27999
rect 13001 27965 13035 27999
rect 13277 27965 13311 27999
rect 13394 27965 13428 27999
rect 9597 27897 9631 27931
rect 1593 27829 1627 27863
rect 10793 27829 10827 27863
rect 11253 27829 11287 27863
rect 11897 27829 11931 27863
rect 2881 27557 2915 27591
rect 8493 27557 8527 27591
rect 11621 27489 11655 27523
rect 2697 27421 2731 27455
rect 7481 27421 7515 27455
rect 7723 27421 7757 27455
rect 10241 27421 10275 27455
rect 10499 27391 10533 27425
rect 11879 27391 11913 27425
rect 13093 27353 13127 27387
rect 13461 27353 13495 27387
rect 11253 27285 11287 27319
rect 12633 27285 12667 27319
rect 1593 27081 1627 27115
rect 2789 27081 2823 27115
rect 8217 27081 8251 27115
rect 14197 27081 14231 27115
rect 11621 27013 11655 27047
rect 1501 26945 1535 26979
rect 2973 26945 3007 26979
rect 4905 26945 4939 26979
rect 5179 26945 5213 26979
rect 6377 26945 6411 26979
rect 7573 26945 7607 26979
rect 10115 26955 10149 26989
rect 12357 26945 12391 26979
rect 6561 26877 6595 26911
rect 7297 26877 7331 26911
rect 7414 26877 7448 26911
rect 9873 26877 9907 26911
rect 12541 26877 12575 26911
rect 13001 26877 13035 26911
rect 13277 26877 13311 26911
rect 13394 26877 13428 26911
rect 13553 26877 13587 26911
rect 5917 26809 5951 26843
rect 7021 26809 7055 26843
rect 10885 26741 10919 26775
rect 11897 26741 11931 26775
rect 8217 26537 8251 26571
rect 12357 26537 12391 26571
rect 13645 26537 13679 26571
rect 6009 26469 6043 26503
rect 7021 26469 7055 26503
rect 11161 26469 11195 26503
rect 4997 26401 5031 26435
rect 7414 26401 7448 26435
rect 10701 26401 10735 26435
rect 11437 26401 11471 26435
rect 11575 26401 11609 26435
rect 5271 26333 5305 26367
rect 6377 26333 6411 26367
rect 6561 26333 6595 26367
rect 7297 26333 7331 26367
rect 7573 26333 7607 26367
rect 10517 26333 10551 26367
rect 11713 26333 11747 26367
rect 12633 26333 12667 26367
rect 12891 26303 12925 26337
rect 1501 26265 1535 26299
rect 1685 26265 1719 26299
rect 14197 25993 14231 26027
rect 7187 25887 7221 25921
rect 8567 25887 8601 25921
rect 9689 25857 9723 25891
rect 9963 25857 9997 25891
rect 11621 25857 11655 25891
rect 13277 25857 13311 25891
rect 6929 25789 6963 25823
rect 8309 25789 8343 25823
rect 12357 25789 12391 25823
rect 12541 25789 12575 25823
rect 13394 25789 13428 25823
rect 13553 25789 13587 25823
rect 12981 25721 13015 25755
rect 7941 25653 7975 25687
rect 9321 25653 9355 25687
rect 10701 25653 10735 25687
rect 11897 25653 11931 25687
rect 7481 25449 7515 25483
rect 10793 25449 10827 25483
rect 12357 25449 12391 25483
rect 9597 25381 9631 25415
rect 1685 25313 1719 25347
rect 6469 25313 6503 25347
rect 9137 25313 9171 25347
rect 9873 25313 9907 25347
rect 11345 25313 11379 25347
rect 13093 25313 13127 25347
rect 1409 25245 1443 25279
rect 6711 25245 6745 25279
rect 8953 25245 8987 25279
rect 9990 25245 10024 25279
rect 10149 25245 10183 25279
rect 11587 25245 11621 25279
rect 12817 25177 12851 25211
rect 13553 25177 13587 25211
rect 13829 25109 13863 25143
rect 13461 24905 13495 24939
rect 1501 24769 1535 24803
rect 6635 24799 6669 24833
rect 10425 24769 10459 24803
rect 10977 24769 11011 24803
rect 11345 24769 11379 24803
rect 11989 24769 12023 24803
rect 12723 24769 12757 24803
rect 6377 24701 6411 24735
rect 12452 24701 12486 24735
rect 1685 24633 1719 24667
rect 7389 24565 7423 24599
rect 10701 24565 10735 24599
rect 12265 24565 12299 24599
rect 7665 24361 7699 24395
rect 5457 24293 5491 24327
rect 6469 24293 6503 24327
rect 9965 24293 9999 24327
rect 4445 24225 4479 24259
rect 6009 24225 6043 24259
rect 6745 24225 6779 24259
rect 7021 24225 7055 24259
rect 8953 24225 8987 24259
rect 10517 24225 10551 24259
rect 11897 24225 11931 24259
rect 4719 24157 4753 24191
rect 5825 24157 5859 24191
rect 6862 24157 6896 24191
rect 9227 24157 9261 24191
rect 10775 24127 10809 24161
rect 12139 24157 12173 24191
rect 13369 24089 13403 24123
rect 13737 24089 13771 24123
rect 11529 24021 11563 24055
rect 12909 24021 12943 24055
rect 9229 23817 9263 23851
rect 12173 23817 12207 23851
rect 14197 23817 14231 23851
rect 11897 23749 11931 23783
rect 1501 23681 1535 23715
rect 7573 23681 7607 23715
rect 10115 23691 10149 23725
rect 12357 23681 12391 23715
rect 13415 23681 13449 23715
rect 7389 23613 7423 23647
rect 8309 23613 8343 23647
rect 8447 23613 8481 23647
rect 8585 23613 8619 23647
rect 9873 23613 9907 23647
rect 12541 23613 12575 23647
rect 13001 23613 13035 23647
rect 13277 23613 13311 23647
rect 13553 23613 13587 23647
rect 1685 23545 1719 23579
rect 8033 23545 8067 23579
rect 10885 23477 10919 23511
rect 12449 23273 12483 23307
rect 13645 23273 13679 23307
rect 8401 23205 8435 23239
rect 11253 23205 11287 23239
rect 7389 23137 7423 23171
rect 11529 23137 11563 23171
rect 11667 23137 11701 23171
rect 7663 23069 7697 23103
rect 10609 23069 10643 23103
rect 10793 23069 10827 23103
rect 11805 23069 11839 23103
rect 12621 23069 12655 23103
rect 12891 23039 12925 23073
rect 1501 23001 1535 23035
rect 1685 23001 1719 23035
rect 7849 22729 7883 22763
rect 14105 22729 14139 22763
rect 11989 22661 12023 22695
rect 6837 22593 6871 22627
rect 7111 22593 7145 22627
rect 9011 22593 9045 22627
rect 12691 22593 12725 22627
rect 13921 22593 13955 22627
rect 8769 22525 8803 22559
rect 12449 22525 12483 22559
rect 9781 22389 9815 22423
rect 12265 22389 12299 22423
rect 13461 22389 13495 22423
rect 10425 22117 10459 22151
rect 9965 22049 9999 22083
rect 10701 22049 10735 22083
rect 11621 22049 11655 22083
rect 13645 22049 13679 22083
rect 5549 21981 5583 22015
rect 5791 21981 5825 22015
rect 7481 21981 7515 22015
rect 7723 21981 7757 22015
rect 9781 21981 9815 22015
rect 10818 21981 10852 22015
rect 10977 21981 11011 22015
rect 11713 21981 11747 22015
rect 11987 21981 12021 22015
rect 1501 21913 1535 21947
rect 13369 21913 13403 21947
rect 1593 21845 1627 21879
rect 6561 21845 6595 21879
rect 8493 21845 8527 21879
rect 12725 21845 12759 21879
rect 9413 21641 9447 21675
rect 1685 21573 1719 21607
rect 11897 21573 11931 21607
rect 1501 21505 1535 21539
rect 4905 21505 4939 21539
rect 5163 21505 5197 21539
rect 7573 21505 7607 21539
rect 8493 21505 8527 21539
rect 8769 21505 8803 21539
rect 10701 21505 10735 21539
rect 11713 21505 11747 21539
rect 12357 21505 12391 21539
rect 13553 21505 13587 21539
rect 7757 21437 7791 21471
rect 8610 21437 8644 21471
rect 9505 21437 9539 21471
rect 9689 21437 9723 21471
rect 10149 21437 10183 21471
rect 10425 21437 10459 21471
rect 10563 21437 10597 21471
rect 12541 21437 12575 21471
rect 13001 21437 13035 21471
rect 13277 21437 13311 21471
rect 13394 21437 13428 21471
rect 8217 21369 8251 21403
rect 11529 21369 11563 21403
rect 5917 21301 5951 21335
rect 11345 21301 11379 21335
rect 12173 21301 12207 21335
rect 14197 21301 14231 21335
rect 3249 21097 3283 21131
rect 7297 21097 7331 21131
rect 10793 21097 10827 21131
rect 11621 21097 11655 21131
rect 12725 20961 12759 20995
rect 13277 20961 13311 20995
rect 3065 20893 3099 20927
rect 6377 20893 6411 20927
rect 9781 20893 9815 20927
rect 10023 20893 10057 20927
rect 11345 20893 11379 20927
rect 12449 20893 12483 20927
rect 13921 20893 13955 20927
rect 6285 20825 6319 20859
rect 6745 20825 6779 20859
rect 11897 20825 11931 20859
rect 12265 20825 12299 20859
rect 13001 20825 13035 20859
rect 13553 20825 13587 20859
rect 6009 20757 6043 20791
rect 7113 20757 7147 20791
rect 8033 20553 8067 20587
rect 11161 20553 11195 20587
rect 13645 20553 13679 20587
rect 7279 20447 7313 20481
rect 10039 20447 10073 20481
rect 11345 20417 11379 20451
rect 11529 20417 11563 20451
rect 11713 20417 11747 20451
rect 12155 20447 12189 20481
rect 13369 20417 13403 20451
rect 1409 20349 1443 20383
rect 1685 20349 1719 20383
rect 7021 20349 7055 20383
rect 9781 20349 9815 20383
rect 11897 20349 11931 20383
rect 10793 20281 10827 20315
rect 11621 20213 11655 20247
rect 12909 20213 12943 20247
rect 1593 20009 1627 20043
rect 13921 20009 13955 20043
rect 6377 19941 6411 19975
rect 8953 19873 8987 19907
rect 10793 19873 10827 19907
rect 11069 19873 11103 19907
rect 11253 19873 11287 19907
rect 12725 19873 12759 19907
rect 13118 19873 13152 19907
rect 4629 19805 4663 19839
rect 7021 19805 7055 19839
rect 7481 19805 7515 19839
rect 7755 19805 7789 19839
rect 9227 19805 9261 19839
rect 10701 19805 10735 19839
rect 10977 19805 11011 19839
rect 11805 19805 11839 19839
rect 12081 19805 12115 19839
rect 12265 19805 12299 19839
rect 13001 19805 13035 19839
rect 13277 19805 13311 19839
rect 1501 19737 1535 19771
rect 4896 19737 4930 19771
rect 6193 19737 6227 19771
rect 11253 19737 11287 19771
rect 11437 19737 11471 19771
rect 6009 19669 6043 19703
rect 6837 19669 6871 19703
rect 8493 19669 8527 19703
rect 9965 19669 9999 19703
rect 13553 19465 13587 19499
rect 14105 19465 14139 19499
rect 11805 19397 11839 19431
rect 6377 19329 6411 19363
rect 6651 19329 6685 19363
rect 7757 19329 7791 19363
rect 7941 19329 7975 19363
rect 8585 19329 8619 19363
rect 10977 19329 11011 19363
rect 12799 19359 12833 19393
rect 13921 19329 13955 19363
rect 8769 19261 8803 19295
rect 9229 19261 9263 19295
rect 9505 19261 9539 19295
rect 9622 19261 9656 19295
rect 9781 19261 9815 19295
rect 11253 19261 11287 19295
rect 12081 19261 12115 19295
rect 12541 19261 12575 19295
rect 7389 19193 7423 19227
rect 7849 19125 7883 19159
rect 10425 19125 10459 19159
rect 1593 18921 1627 18955
rect 9965 18921 9999 18955
rect 12173 18921 12207 18955
rect 7941 18853 7975 18887
rect 6745 18785 6779 18819
rect 7297 18785 7331 18819
rect 8953 18785 8987 18819
rect 10333 18785 10367 18819
rect 6377 18717 6411 18751
rect 6469 18717 6503 18751
rect 6561 18717 6595 18751
rect 7021 18717 7055 18751
rect 7113 18717 7147 18751
rect 7389 18717 7423 18751
rect 7849 18717 7883 18751
rect 8125 18717 8159 18751
rect 9195 18717 9229 18751
rect 10575 18717 10609 18751
rect 12449 18717 12483 18751
rect 12723 18717 12757 18751
rect 1501 18649 1535 18683
rect 5181 18649 5215 18683
rect 7481 18649 7515 18683
rect 11897 18649 11931 18683
rect 5273 18581 5307 18615
rect 6193 18581 6227 18615
rect 6745 18581 6779 18615
rect 7297 18581 7331 18615
rect 7665 18581 7699 18615
rect 11345 18581 11379 18615
rect 13461 18581 13495 18615
rect 5917 18377 5951 18411
rect 6653 18377 6687 18411
rect 6929 18377 6963 18411
rect 12081 18377 12115 18411
rect 1685 18309 1719 18343
rect 11805 18309 11839 18343
rect 1501 18241 1535 18275
rect 4793 18241 4827 18275
rect 6469 18241 6503 18275
rect 6653 18241 6687 18275
rect 6837 18241 6871 18275
rect 10055 18241 10089 18275
rect 11345 18241 11379 18275
rect 12357 18241 12391 18275
rect 13415 18241 13449 18275
rect 13553 18241 13587 18275
rect 4537 18173 4571 18207
rect 9781 18173 9815 18207
rect 12541 18173 12575 18207
rect 13001 18173 13035 18207
rect 13277 18173 13311 18207
rect 14197 18173 14231 18207
rect 10793 18037 10827 18071
rect 11161 18037 11195 18071
rect 6101 17833 6135 17867
rect 11529 17833 11563 17867
rect 12725 17833 12759 17867
rect 1409 17629 1443 17663
rect 1683 17629 1717 17663
rect 5089 17629 5123 17663
rect 5363 17629 5397 17663
rect 6469 17629 6503 17663
rect 6743 17629 6777 17663
rect 10517 17629 10551 17663
rect 10701 17629 10735 17663
rect 10793 17629 10827 17663
rect 11253 17629 11287 17663
rect 11713 17629 11747 17663
rect 11955 17629 11989 17663
rect 13093 17629 13127 17663
rect 13369 17629 13403 17663
rect 2421 17493 2455 17527
rect 7481 17493 7515 17527
rect 10609 17493 10643 17527
rect 10885 17493 10919 17527
rect 8677 17289 8711 17323
rect 14105 17289 14139 17323
rect 11805 17221 11839 17255
rect 12081 17221 12115 17255
rect 1501 17153 1535 17187
rect 1961 17153 1995 17187
rect 7874 17153 7908 17187
rect 9011 17153 9045 17187
rect 10517 17153 10551 17187
rect 10793 17153 10827 17187
rect 11253 17153 11287 17187
rect 11529 17153 11563 17187
rect 12783 17153 12817 17187
rect 14013 17153 14047 17187
rect 1685 17085 1719 17119
rect 6837 17085 6871 17119
rect 7021 17085 7055 17119
rect 7481 17085 7515 17119
rect 7757 17085 7791 17119
rect 8033 17085 8067 17119
rect 8769 17085 8803 17119
rect 11621 17085 11655 17119
rect 11805 17085 11839 17119
rect 12357 17085 12391 17119
rect 12541 17085 12575 17119
rect 1777 16949 1811 16983
rect 9781 16949 9815 16983
rect 10701 16949 10735 16983
rect 10977 16949 11011 16983
rect 11069 16949 11103 16983
rect 13553 16949 13587 16983
rect 1593 16745 1627 16779
rect 7757 16745 7791 16779
rect 11069 16745 11103 16779
rect 13921 16745 13955 16779
rect 9873 16677 9907 16711
rect 11345 16677 11379 16711
rect 6745 16609 6779 16643
rect 9229 16609 9263 16643
rect 9413 16609 9447 16643
rect 10287 16609 10321 16643
rect 12081 16609 12115 16643
rect 12725 16609 12759 16643
rect 13001 16609 13035 16643
rect 13277 16609 13311 16643
rect 7019 16541 7053 16575
rect 10149 16541 10183 16575
rect 10425 16541 10459 16575
rect 11161 16541 11195 16575
rect 11437 16541 11471 16575
rect 12265 16541 12299 16575
rect 13139 16541 13173 16575
rect 1501 16473 1535 16507
rect 11805 16473 11839 16507
rect 11621 16405 11655 16439
rect 11897 16405 11931 16439
rect 10057 16201 10091 16235
rect 12817 16201 12851 16235
rect 14105 16201 14139 16235
rect 13461 16133 13495 16167
rect 1409 16065 1443 16099
rect 1667 16095 1701 16129
rect 6837 16065 6871 16099
rect 7111 16065 7145 16099
rect 9287 16065 9321 16099
rect 12047 16065 12081 16099
rect 13829 16065 13863 16099
rect 9045 15997 9079 16031
rect 11805 15997 11839 16031
rect 2421 15861 2455 15895
rect 7849 15861 7883 15895
rect 13553 15861 13587 15895
rect 11989 15657 12023 15691
rect 1685 15589 1719 15623
rect 10793 15589 10827 15623
rect 7481 15521 7515 15555
rect 10333 15521 10367 15555
rect 11069 15521 11103 15555
rect 11345 15521 11379 15555
rect 12081 15521 12115 15555
rect 7723 15453 7757 15487
rect 10149 15453 10183 15487
rect 11186 15453 11220 15487
rect 12323 15453 12357 15487
rect 13737 15453 13771 15487
rect 1501 15385 1535 15419
rect 8493 15317 8527 15351
rect 13093 15317 13127 15351
rect 13829 15317 13863 15351
rect 9965 15113 9999 15147
rect 11897 15113 11931 15147
rect 14197 15113 14231 15147
rect 1501 15045 1535 15079
rect 2145 14977 2179 15011
rect 5147 14977 5181 15011
rect 6619 14977 6653 15011
rect 8125 14977 8159 15011
rect 9045 14977 9079 15011
rect 9321 14977 9355 15011
rect 10299 14977 10333 15011
rect 11713 14977 11747 15011
rect 12081 14977 12115 15011
rect 12265 14977 12299 15011
rect 12541 14977 12575 15011
rect 13277 14977 13311 15011
rect 4905 14909 4939 14943
rect 6377 14909 6411 14943
rect 8309 14909 8343 14943
rect 8769 14909 8803 14943
rect 9162 14909 9196 14943
rect 10057 14909 10091 14943
rect 12357 14909 12391 14943
rect 13001 14909 13035 14943
rect 13394 14909 13428 14943
rect 13553 14909 13587 14943
rect 1593 14773 1627 14807
rect 1961 14773 1995 14807
rect 5917 14773 5951 14807
rect 7389 14773 7423 14807
rect 11069 14773 11103 14807
rect 7665 14569 7699 14603
rect 13553 14569 13587 14603
rect 6469 14501 6503 14535
rect 11989 14501 12023 14535
rect 1409 14433 1443 14467
rect 5825 14433 5859 14467
rect 6862 14433 6896 14467
rect 7021 14433 7055 14467
rect 10333 14433 10367 14467
rect 10793 14433 10827 14467
rect 11087 14433 11121 14467
rect 12541 14433 12575 14467
rect 1651 14365 1685 14399
rect 6009 14365 6043 14399
rect 6745 14365 6779 14399
rect 10149 14365 10183 14399
rect 11207 14365 11241 14399
rect 11345 14365 11379 14399
rect 12291 14365 12325 14399
rect 12815 14365 12849 14399
rect 2421 14229 2455 14263
rect 12449 14229 12483 14263
rect 10517 14025 10551 14059
rect 1501 13957 1535 13991
rect 13921 13957 13955 13991
rect 7205 13889 7239 13923
rect 8125 13889 8159 13923
rect 8263 13889 8297 13923
rect 8401 13889 8435 13923
rect 9045 13889 9079 13923
rect 9779 13899 9813 13933
rect 11803 13889 11837 13923
rect 7389 13821 7423 13855
rect 7849 13821 7883 13855
rect 9505 13821 9539 13855
rect 11529 13821 11563 13855
rect 12909 13821 12943 13855
rect 13185 13821 13219 13855
rect 14105 13821 14139 13855
rect 1593 13685 1627 13719
rect 12541 13685 12575 13719
rect 7113 13481 7147 13515
rect 10793 13481 10827 13515
rect 13093 13481 13127 13515
rect 13829 13481 13863 13515
rect 8493 13413 8527 13447
rect 9597 13413 9631 13447
rect 13369 13413 13403 13447
rect 6101 13345 6135 13379
rect 8953 13345 8987 13379
rect 9990 13345 10024 13379
rect 11437 13345 11471 13379
rect 11897 13345 11931 13379
rect 12173 13345 12207 13379
rect 12311 13345 12345 13379
rect 12449 13345 12483 13379
rect 2145 13277 2179 13311
rect 6359 13247 6393 13281
rect 7481 13277 7515 13311
rect 7755 13277 7789 13311
rect 9137 13277 9171 13311
rect 9873 13277 9907 13311
rect 10149 13277 10183 13311
rect 11253 13277 11287 13311
rect 13185 13277 13219 13311
rect 1501 13209 1535 13243
rect 13737 13209 13771 13243
rect 1593 13141 1627 13175
rect 1961 13141 1995 13175
rect 8033 12937 8067 12971
rect 9873 12937 9907 12971
rect 14197 12937 14231 12971
rect 1409 12801 1443 12835
rect 1667 12831 1701 12865
rect 7021 12801 7055 12835
rect 7295 12801 7329 12835
rect 9103 12801 9137 12835
rect 10793 12801 10827 12835
rect 12081 12801 12115 12835
rect 12541 12801 12575 12835
rect 8861 12733 8895 12767
rect 10517 12733 10551 12767
rect 12357 12733 12391 12767
rect 13277 12733 13311 12767
rect 13415 12733 13449 12767
rect 13553 12733 13587 12767
rect 12265 12665 12299 12699
rect 13001 12665 13035 12699
rect 2421 12597 2455 12631
rect 11529 12393 11563 12427
rect 13185 12393 13219 12427
rect 4353 12257 4387 12291
rect 7113 12257 7147 12291
rect 10517 12257 10551 12291
rect 12173 12257 12207 12291
rect 2145 12189 2179 12223
rect 4627 12189 4661 12223
rect 5733 12189 5767 12223
rect 6007 12189 6041 12223
rect 7387 12189 7421 12223
rect 10759 12189 10793 12223
rect 11897 12189 11931 12223
rect 12415 12189 12449 12223
rect 13737 12189 13771 12223
rect 1501 12121 1535 12155
rect 1593 12053 1627 12087
rect 1961 12053 1995 12087
rect 5365 12053 5399 12087
rect 6745 12053 6779 12087
rect 8125 12053 8159 12087
rect 12081 12053 12115 12087
rect 13829 12053 13863 12087
rect 13645 11849 13679 11883
rect 1501 11713 1535 11747
rect 4905 11713 4939 11747
rect 5163 11743 5197 11777
rect 7923 11743 7957 11777
rect 10517 11713 10551 11747
rect 10793 11713 10827 11747
rect 11713 11713 11747 11747
rect 12891 11743 12925 11777
rect 14013 11713 14047 11747
rect 7665 11645 7699 11679
rect 11989 11645 12023 11679
rect 12633 11645 12667 11679
rect 1593 11509 1627 11543
rect 5917 11509 5951 11543
rect 8677 11509 8711 11543
rect 14197 11509 14231 11543
rect 7849 11305 7883 11339
rect 11161 11237 11195 11271
rect 6653 11169 6687 11203
rect 12357 11169 12391 11203
rect 12449 11169 12483 11203
rect 6009 11101 6043 11135
rect 6193 11101 6227 11135
rect 6929 11101 6963 11135
rect 7067 11101 7101 11135
rect 7205 11101 7239 11135
rect 10517 11101 10551 11135
rect 10701 11101 10735 11135
rect 11437 11101 11471 11135
rect 11575 11101 11609 11135
rect 11713 11101 11747 11135
rect 12707 11071 12741 11105
rect 13461 10965 13495 10999
rect 1961 10761 1995 10795
rect 7297 10761 7331 10795
rect 8125 10761 8159 10795
rect 11069 10761 11103 10795
rect 11713 10761 11747 10795
rect 11989 10761 12023 10795
rect 12265 10761 12299 10795
rect 14197 10761 14231 10795
rect 8401 10693 8435 10727
rect 8493 10693 8527 10727
rect 9229 10693 9263 10727
rect 1501 10625 1535 10659
rect 2145 10625 2179 10659
rect 6377 10625 6411 10659
rect 6653 10625 6687 10659
rect 6837 10625 6871 10659
rect 7205 10625 7239 10659
rect 8861 10625 8895 10659
rect 10315 10655 10349 10689
rect 11529 10625 11563 10659
rect 11805 10625 11839 10659
rect 12081 10625 12115 10659
rect 13277 10625 13311 10659
rect 13394 10625 13428 10659
rect 10057 10557 10091 10591
rect 12357 10557 12391 10591
rect 12541 10557 12575 10591
rect 13001 10557 13035 10591
rect 13553 10557 13587 10591
rect 1593 10421 1627 10455
rect 6469 10421 6503 10455
rect 6745 10421 6779 10455
rect 9413 10421 9447 10455
rect 2973 10217 3007 10251
rect 5733 10217 5767 10251
rect 10793 10217 10827 10251
rect 12725 10217 12759 10251
rect 6377 10149 6411 10183
rect 9597 10149 9631 10183
rect 5917 10081 5951 10115
rect 6837 10081 6871 10115
rect 7297 10081 7331 10115
rect 7849 10081 7883 10115
rect 9137 10081 9171 10115
rect 11529 10081 11563 10115
rect 12817 10081 12851 10115
rect 1409 10013 1443 10047
rect 1683 10013 1717 10047
rect 2789 10013 2823 10047
rect 5641 10013 5675 10047
rect 6285 10013 6319 10047
rect 6561 10013 6595 10047
rect 6653 10013 6687 10047
rect 7573 10013 7607 10047
rect 7690 10013 7724 10047
rect 8953 10013 8987 10047
rect 9873 10013 9907 10047
rect 10011 10013 10045 10047
rect 10149 10013 10183 10047
rect 10885 10013 10919 10047
rect 11069 10013 11103 10047
rect 11805 10013 11839 10047
rect 11922 10013 11956 10047
rect 12081 10013 12115 10047
rect 13093 10013 13127 10047
rect 2421 9877 2455 9911
rect 5917 9877 5951 9911
rect 6101 9877 6135 9911
rect 8493 9877 8527 9911
rect 14197 9605 14231 9639
rect 1667 9567 1701 9601
rect 9413 9537 9447 9571
rect 10149 9537 10183 9571
rect 10266 9537 10300 9571
rect 10425 9537 10459 9571
rect 12081 9537 12115 9571
rect 12357 9537 12391 9571
rect 13277 9537 13311 9571
rect 13415 9537 13449 9571
rect 1409 9469 1443 9503
rect 9229 9469 9263 9503
rect 12541 9469 12575 9503
rect 13553 9469 13587 9503
rect 9873 9401 9907 9435
rect 11069 9401 11103 9435
rect 13001 9401 13035 9435
rect 2421 9333 2455 9367
rect 12173 9333 12207 9367
rect 11345 9129 11379 9163
rect 12449 9129 12483 9163
rect 13921 9129 13955 9163
rect 8493 9061 8527 9095
rect 9689 8993 9723 9027
rect 10149 8993 10183 9027
rect 10701 8993 10735 9027
rect 11437 8993 11471 9027
rect 13093 8993 13127 9027
rect 2237 8925 2271 8959
rect 2513 8925 2547 8959
rect 2605 8925 2639 8959
rect 7481 8925 7515 8959
rect 7739 8925 7773 8959
rect 9505 8925 9539 8959
rect 10425 8925 10459 8959
rect 10542 8925 10576 8959
rect 11679 8925 11713 8959
rect 12817 8925 12851 8959
rect 13737 8925 13771 8959
rect 1501 8857 1535 8891
rect 2697 8857 2731 8891
rect 1593 8789 1627 8823
rect 2053 8789 2087 8823
rect 2329 8789 2363 8823
rect 6653 8585 6687 8619
rect 10747 8585 10781 8619
rect 13553 8585 13587 8619
rect 14105 8585 14139 8619
rect 1501 8517 1535 8551
rect 4905 8449 4939 8483
rect 5163 8479 5197 8513
rect 6377 8449 6411 8483
rect 6745 8449 6779 8483
rect 7021 8449 7055 8483
rect 7205 8449 7239 8483
rect 9873 8449 9907 8483
rect 10241 8449 10275 8483
rect 10517 8449 10551 8483
rect 11805 8449 11839 8483
rect 12541 8449 12575 8483
rect 12783 8449 12817 8483
rect 14013 8449 14047 8483
rect 6653 8381 6687 8415
rect 7113 8381 7147 8415
rect 8585 8381 8619 8415
rect 10425 8381 10459 8415
rect 11529 8381 11563 8415
rect 1685 8313 1719 8347
rect 5917 8313 5951 8347
rect 6469 8313 6503 8347
rect 6837 8313 6871 8347
rect 8493 8313 8527 8347
rect 9965 8245 9999 8279
rect 6377 8041 6411 8075
rect 13645 8041 13679 8075
rect 6653 7973 6687 8007
rect 6929 7905 6963 7939
rect 7573 7905 7607 7939
rect 7849 7905 7883 7939
rect 7987 7905 8021 7939
rect 8125 7905 8159 7939
rect 10241 7905 10275 7939
rect 10517 7905 10551 7939
rect 10634 7905 10668 7939
rect 11713 7905 11747 7939
rect 12633 7905 12667 7939
rect 1409 7837 1443 7871
rect 1683 7837 1717 7871
rect 6561 7837 6595 7871
rect 6837 7837 6871 7871
rect 7113 7837 7147 7871
rect 9597 7837 9631 7871
rect 9781 7837 9815 7871
rect 10793 7837 10827 7871
rect 11437 7837 11471 7871
rect 11989 7837 12023 7871
rect 12907 7837 12941 7871
rect 2421 7701 2455 7735
rect 8769 7701 8803 7735
rect 1961 7497 1995 7531
rect 9045 7497 9079 7531
rect 13001 7497 13035 7531
rect 1501 7429 1535 7463
rect 11713 7429 11747 7463
rect 2145 7361 2179 7395
rect 7205 7361 7239 7395
rect 7389 7361 7423 7395
rect 8263 7361 8297 7395
rect 9229 7361 9263 7395
rect 9505 7361 9539 7395
rect 10425 7361 10459 7395
rect 10542 7361 10576 7395
rect 12231 7361 12265 7395
rect 13645 7361 13679 7395
rect 7849 7293 7883 7327
rect 8125 7293 8159 7327
rect 8401 7293 8435 7327
rect 9689 7293 9723 7327
rect 10701 7293 10735 7327
rect 11989 7293 12023 7327
rect 13369 7293 13403 7327
rect 10149 7225 10183 7259
rect 1593 7157 1627 7191
rect 9413 7157 9447 7191
rect 11345 7157 11379 7191
rect 11805 7157 11839 7191
rect 7849 6953 7883 6987
rect 11989 6885 12023 6919
rect 8953 6817 8987 6851
rect 9597 6817 9631 6851
rect 9873 6817 9907 6851
rect 10159 6817 10193 6851
rect 6837 6749 6871 6783
rect 7111 6749 7145 6783
rect 9137 6749 9171 6783
rect 9990 6749 10024 6783
rect 10977 6749 11011 6783
rect 11251 6749 11285 6783
rect 13277 6749 13311 6783
rect 1501 6681 1535 6715
rect 12817 6681 12851 6715
rect 12909 6681 12943 6715
rect 13645 6681 13679 6715
rect 1593 6613 1627 6647
rect 10793 6613 10827 6647
rect 12541 6613 12575 6647
rect 13829 6613 13863 6647
rect 8953 6409 8987 6443
rect 14105 6409 14139 6443
rect 12817 6341 12851 6375
rect 13093 6341 13127 6375
rect 13553 6341 13587 6375
rect 13921 6341 13955 6375
rect 1667 6303 1701 6337
rect 7941 6273 7975 6307
rect 8183 6273 8217 6307
rect 9505 6273 9539 6307
rect 10358 6273 10392 6307
rect 10517 6273 10551 6307
rect 11713 6273 11747 6307
rect 13185 6273 13219 6307
rect 1409 6205 1443 6239
rect 9321 6205 9355 6239
rect 10241 6205 10275 6239
rect 11989 6205 12023 6239
rect 9965 6137 9999 6171
rect 2421 6069 2455 6103
rect 11161 6069 11195 6103
rect 2329 5865 2363 5899
rect 8309 5865 8343 5899
rect 7297 5729 7331 5763
rect 10609 5729 10643 5763
rect 10793 5729 10827 5763
rect 11253 5729 11287 5763
rect 11529 5729 11563 5763
rect 11646 5729 11680 5763
rect 12541 5729 12575 5763
rect 2237 5661 2271 5695
rect 2513 5661 2547 5695
rect 7571 5661 7605 5695
rect 11805 5661 11839 5695
rect 12783 5661 12817 5695
rect 1501 5593 1535 5627
rect 12449 5593 12483 5627
rect 1593 5525 1627 5559
rect 2053 5525 2087 5559
rect 13553 5525 13587 5559
rect 10333 5321 10367 5355
rect 12541 5321 12575 5355
rect 13921 5321 13955 5355
rect 1501 5253 1535 5287
rect 2053 5253 2087 5287
rect 1961 5185 1995 5219
rect 9579 5215 9613 5249
rect 11771 5195 11805 5229
rect 13151 5185 13185 5219
rect 9321 5117 9355 5151
rect 11529 5117 11563 5151
rect 12909 5117 12943 5151
rect 1593 4981 1627 5015
rect 9965 4777 9999 4811
rect 11345 4777 11379 4811
rect 12449 4777 12483 4811
rect 13645 4777 13679 4811
rect 8953 4641 8987 4675
rect 10333 4641 10367 4675
rect 12173 4641 12207 4675
rect 9227 4573 9261 4607
rect 10575 4573 10609 4607
rect 11989 4573 12023 4607
rect 12633 4573 12667 4607
rect 12891 4543 12925 4577
rect 12357 4505 12391 4539
rect 12357 4165 12391 4199
rect 13093 4165 13127 4199
rect 14013 4165 14047 4199
rect 1409 4097 1443 4131
rect 10517 4097 10551 4131
rect 13645 4097 13679 4131
rect 10793 4029 10827 4063
rect 12541 4029 12575 4063
rect 13829 4029 13863 4063
rect 1593 3893 1627 3927
rect 13185 3893 13219 3927
rect 14105 3893 14139 3927
rect 13829 3689 13863 3723
rect 13737 3485 13771 3519
rect 6561 2057 6595 2091
rect 7205 2057 7239 2091
rect 7941 2057 7975 2091
rect 8677 2057 8711 2091
rect 9413 2057 9447 2091
rect 10149 2057 10183 2091
rect 10885 2057 10919 2091
rect 13461 2057 13495 2091
rect 14013 2057 14047 2091
rect 2881 1989 2915 2023
rect 13369 1989 13403 2023
rect 2053 1921 2087 1955
rect 6469 1921 6503 1955
rect 7113 1921 7147 1955
rect 7849 1921 7883 1955
rect 8585 1921 8619 1955
rect 9321 1921 9355 1955
rect 10057 1921 10091 1955
rect 10793 1921 10827 1955
rect 11621 1921 11655 1955
rect 12265 1921 12299 1955
rect 12909 1921 12943 1955
rect 13737 1921 13771 1955
rect 14197 1921 14231 1955
rect 11805 1853 11839 1887
rect 13921 1853 13955 1887
rect 12357 1717 12391 1751
rect 13001 1717 13035 1751
rect 6009 1513 6043 1547
rect 7297 1513 7331 1547
rect 7941 1513 7975 1547
rect 8953 1513 8987 1547
rect 9413 1513 9447 1547
rect 10149 1513 10183 1547
rect 10885 1513 10919 1547
rect 11621 1513 11655 1547
rect 12357 1513 12391 1547
rect 13093 1513 13127 1547
rect 13369 1513 13403 1547
rect 3433 1377 3467 1411
rect 1409 1309 1443 1343
rect 2237 1309 2271 1343
rect 2697 1309 2731 1343
rect 3801 1309 3835 1343
rect 4629 1309 4663 1343
rect 5273 1309 5307 1343
rect 6193 1309 6227 1343
rect 6377 1309 6411 1343
rect 6653 1309 6687 1343
rect 7481 1309 7515 1343
rect 8125 1309 8159 1343
rect 9137 1309 9171 1343
rect 9597 1309 9631 1343
rect 10333 1309 10367 1343
rect 11069 1309 11103 1343
rect 11805 1309 11839 1343
rect 12541 1309 12575 1343
rect 13001 1309 13035 1343
rect 13277 1309 13311 1343
rect 13553 1309 13587 1343
rect 4077 1241 4111 1275
rect 4445 1241 4479 1275
rect 5089 1241 5123 1275
rect 13737 1241 13771 1275
rect 12817 1173 12851 1207
rect 13829 1173 13863 1207
<< metal1 >>
rect 1104 43546 14696 43568
rect 1104 43494 4308 43546
rect 4360 43494 4372 43546
rect 4424 43494 4436 43546
rect 4488 43494 4500 43546
rect 4552 43494 4564 43546
rect 4616 43494 7666 43546
rect 7718 43494 7730 43546
rect 7782 43494 7794 43546
rect 7846 43494 7858 43546
rect 7910 43494 7922 43546
rect 7974 43494 11024 43546
rect 11076 43494 11088 43546
rect 11140 43494 11152 43546
rect 11204 43494 11216 43546
rect 11268 43494 11280 43546
rect 11332 43494 14382 43546
rect 14434 43494 14446 43546
rect 14498 43494 14510 43546
rect 14562 43494 14574 43546
rect 14626 43494 14638 43546
rect 14690 43494 14696 43546
rect 1104 43472 14696 43494
rect 474 43392 480 43444
rect 532 43432 538 43444
rect 3329 43435 3387 43441
rect 3329 43432 3341 43435
rect 532 43404 3341 43432
rect 532 43392 538 43404
rect 3329 43401 3341 43404
rect 3375 43401 3387 43435
rect 3329 43395 3387 43401
rect 3418 43392 3424 43444
rect 3476 43432 3482 43444
rect 3973 43435 4031 43441
rect 3973 43432 3985 43435
rect 3476 43404 3985 43432
rect 3476 43392 3482 43404
rect 3973 43401 3985 43404
rect 4019 43401 4031 43435
rect 3973 43395 4031 43401
rect 4154 43392 4160 43444
rect 4212 43432 4218 43444
rect 4433 43435 4491 43441
rect 4433 43432 4445 43435
rect 4212 43404 4445 43432
rect 4212 43392 4218 43404
rect 4433 43401 4445 43404
rect 4479 43401 4491 43435
rect 4433 43395 4491 43401
rect 4890 43392 4896 43444
rect 4948 43432 4954 43444
rect 5169 43435 5227 43441
rect 5169 43432 5181 43435
rect 4948 43404 5181 43432
rect 4948 43392 4954 43404
rect 5169 43401 5181 43404
rect 5215 43401 5227 43435
rect 5169 43395 5227 43401
rect 5626 43392 5632 43444
rect 5684 43432 5690 43444
rect 5905 43435 5963 43441
rect 5905 43432 5917 43435
rect 5684 43404 5917 43432
rect 5684 43392 5690 43404
rect 5905 43401 5917 43404
rect 5951 43401 5963 43435
rect 5905 43395 5963 43401
rect 6362 43392 6368 43444
rect 6420 43432 6426 43444
rect 6641 43435 6699 43441
rect 6641 43432 6653 43435
rect 6420 43404 6653 43432
rect 6420 43392 6426 43404
rect 6641 43401 6653 43404
rect 6687 43401 6699 43435
rect 6641 43395 6699 43401
rect 7098 43392 7104 43444
rect 7156 43432 7162 43444
rect 7377 43435 7435 43441
rect 7377 43432 7389 43435
rect 7156 43404 7389 43432
rect 7156 43392 7162 43404
rect 7377 43401 7389 43404
rect 7423 43401 7435 43435
rect 7377 43395 7435 43401
rect 8018 43392 8024 43444
rect 8076 43432 8082 43444
rect 8113 43435 8171 43441
rect 8113 43432 8125 43435
rect 8076 43404 8125 43432
rect 8076 43392 8082 43404
rect 8113 43401 8125 43404
rect 8159 43401 8171 43435
rect 8113 43395 8171 43401
rect 8570 43392 8576 43444
rect 8628 43432 8634 43444
rect 9125 43435 9183 43441
rect 9125 43432 9137 43435
rect 8628 43404 9137 43432
rect 8628 43392 8634 43404
rect 9125 43401 9137 43404
rect 9171 43401 9183 43435
rect 9125 43395 9183 43401
rect 9306 43392 9312 43444
rect 9364 43432 9370 43444
rect 9585 43435 9643 43441
rect 9585 43432 9597 43435
rect 9364 43404 9597 43432
rect 9364 43392 9370 43404
rect 9585 43401 9597 43404
rect 9631 43401 9643 43435
rect 9585 43395 9643 43401
rect 10042 43392 10048 43444
rect 10100 43432 10106 43444
rect 10321 43435 10379 43441
rect 10321 43432 10333 43435
rect 10100 43404 10333 43432
rect 10100 43392 10106 43404
rect 10321 43401 10333 43404
rect 10367 43401 10379 43435
rect 10321 43395 10379 43401
rect 10778 43392 10784 43444
rect 10836 43432 10842 43444
rect 11057 43435 11115 43441
rect 11057 43432 11069 43435
rect 10836 43404 11069 43432
rect 10836 43392 10842 43404
rect 11057 43401 11069 43404
rect 11103 43401 11115 43435
rect 11057 43395 11115 43401
rect 11514 43392 11520 43444
rect 11572 43432 11578 43444
rect 11793 43435 11851 43441
rect 11793 43432 11805 43435
rect 11572 43404 11805 43432
rect 11572 43392 11578 43404
rect 11793 43401 11805 43404
rect 11839 43401 11851 43435
rect 11793 43395 11851 43401
rect 12250 43392 12256 43444
rect 12308 43432 12314 43444
rect 12529 43435 12587 43441
rect 12529 43432 12541 43435
rect 12308 43404 12541 43432
rect 12308 43392 12314 43404
rect 12529 43401 12541 43404
rect 12575 43401 12587 43435
rect 12529 43395 12587 43401
rect 12986 43392 12992 43444
rect 13044 43432 13050 43444
rect 13265 43435 13323 43441
rect 13265 43432 13277 43435
rect 13044 43404 13277 43432
rect 13044 43392 13050 43404
rect 13265 43401 13277 43404
rect 13311 43401 13323 43435
rect 13265 43395 13323 43401
rect 13817 43435 13875 43441
rect 13817 43401 13829 43435
rect 13863 43432 13875 43435
rect 15194 43432 15200 43444
rect 13863 43404 15200 43432
rect 13863 43401 13875 43404
rect 13817 43395 13875 43401
rect 15194 43392 15200 43404
rect 15252 43392 15258 43444
rect 1489 43299 1547 43305
rect 1489 43265 1501 43299
rect 1535 43296 1547 43299
rect 1762 43296 1768 43308
rect 1535 43268 1768 43296
rect 1535 43265 1547 43268
rect 1489 43259 1547 43265
rect 1762 43256 1768 43268
rect 1820 43256 1826 43308
rect 2038 43256 2044 43308
rect 2096 43256 2102 43308
rect 2685 43299 2743 43305
rect 2685 43265 2697 43299
rect 2731 43296 2743 43299
rect 3050 43296 3056 43308
rect 2731 43268 3056 43296
rect 2731 43265 2743 43268
rect 2685 43259 2743 43265
rect 3050 43256 3056 43268
rect 3108 43256 3114 43308
rect 3142 43256 3148 43308
rect 3200 43256 3206 43308
rect 3786 43256 3792 43308
rect 3844 43256 3850 43308
rect 4338 43256 4344 43308
rect 4396 43256 4402 43308
rect 4982 43256 4988 43308
rect 5040 43256 5046 43308
rect 5718 43256 5724 43308
rect 5776 43256 5782 43308
rect 6454 43256 6460 43308
rect 6512 43256 6518 43308
rect 7190 43256 7196 43308
rect 7248 43256 7254 43308
rect 7926 43256 7932 43308
rect 7984 43256 7990 43308
rect 8938 43256 8944 43308
rect 8996 43256 9002 43308
rect 9214 43256 9220 43308
rect 9272 43296 9278 43308
rect 9401 43299 9459 43305
rect 9401 43296 9413 43299
rect 9272 43268 9413 43296
rect 9272 43256 9278 43268
rect 9401 43265 9413 43268
rect 9447 43265 9459 43299
rect 9401 43259 9459 43265
rect 10134 43256 10140 43308
rect 10192 43256 10198 43308
rect 10962 43256 10968 43308
rect 11020 43256 11026 43308
rect 11606 43256 11612 43308
rect 11664 43256 11670 43308
rect 12434 43256 12440 43308
rect 12492 43256 12498 43308
rect 13078 43256 13084 43308
rect 13136 43256 13142 43308
rect 13538 43256 13544 43308
rect 13596 43256 13602 43308
rect 1946 43120 1952 43172
rect 2004 43160 2010 43172
rect 2225 43163 2283 43169
rect 2225 43160 2237 43163
rect 2004 43132 2237 43160
rect 2004 43120 2010 43132
rect 2225 43129 2237 43132
rect 2271 43129 2283 43163
rect 2225 43123 2283 43129
rect 1394 43052 1400 43104
rect 1452 43092 1458 43104
rect 1581 43095 1639 43101
rect 1581 43092 1593 43095
rect 1452 43064 1593 43092
rect 1452 43052 1458 43064
rect 1581 43061 1593 43064
rect 1627 43061 1639 43095
rect 1581 43055 1639 43061
rect 2774 43052 2780 43104
rect 2832 43052 2838 43104
rect 1104 43002 14536 43024
rect 1104 42950 2629 43002
rect 2681 42950 2693 43002
rect 2745 42950 2757 43002
rect 2809 42950 2821 43002
rect 2873 42950 2885 43002
rect 2937 42950 5987 43002
rect 6039 42950 6051 43002
rect 6103 42950 6115 43002
rect 6167 42950 6179 43002
rect 6231 42950 6243 43002
rect 6295 42950 9345 43002
rect 9397 42950 9409 43002
rect 9461 42950 9473 43002
rect 9525 42950 9537 43002
rect 9589 42950 9601 43002
rect 9653 42950 12703 43002
rect 12755 42950 12767 43002
rect 12819 42950 12831 43002
rect 12883 42950 12895 43002
rect 12947 42950 12959 43002
rect 13011 42950 14536 43002
rect 1104 42928 14536 42950
rect 2869 42891 2927 42897
rect 2869 42857 2881 42891
rect 2915 42888 2927 42891
rect 3142 42888 3148 42900
rect 2915 42860 3148 42888
rect 2915 42857 2927 42860
rect 2869 42851 2927 42857
rect 3142 42848 3148 42860
rect 3200 42848 3206 42900
rect 3237 42891 3295 42897
rect 3237 42857 3249 42891
rect 3283 42888 3295 42891
rect 3786 42888 3792 42900
rect 3283 42860 3792 42888
rect 3283 42857 3295 42860
rect 3237 42851 3295 42857
rect 3786 42848 3792 42860
rect 3844 42848 3850 42900
rect 4065 42891 4123 42897
rect 4065 42857 4077 42891
rect 4111 42888 4123 42891
rect 4338 42888 4344 42900
rect 4111 42860 4344 42888
rect 4111 42857 4123 42860
rect 4065 42851 4123 42857
rect 4338 42848 4344 42860
rect 4396 42848 4402 42900
rect 4801 42891 4859 42897
rect 4801 42857 4813 42891
rect 4847 42888 4859 42891
rect 4982 42888 4988 42900
rect 4847 42860 4988 42888
rect 4847 42857 4859 42860
rect 4801 42851 4859 42857
rect 4982 42848 4988 42860
rect 5040 42848 5046 42900
rect 6273 42891 6331 42897
rect 6273 42857 6285 42891
rect 6319 42888 6331 42891
rect 6454 42888 6460 42900
rect 6319 42860 6460 42888
rect 6319 42857 6331 42860
rect 6273 42851 6331 42857
rect 6454 42848 6460 42860
rect 6512 42848 6518 42900
rect 7009 42891 7067 42897
rect 7009 42857 7021 42891
rect 7055 42888 7067 42891
rect 7190 42888 7196 42900
rect 7055 42860 7196 42888
rect 7055 42857 7067 42860
rect 7009 42851 7067 42857
rect 7190 42848 7196 42860
rect 7248 42848 7254 42900
rect 7745 42891 7803 42897
rect 7745 42857 7757 42891
rect 7791 42888 7803 42891
rect 7926 42888 7932 42900
rect 7791 42860 7932 42888
rect 7791 42857 7803 42860
rect 7745 42851 7803 42857
rect 7926 42848 7932 42860
rect 7984 42848 7990 42900
rect 8481 42891 8539 42897
rect 8481 42857 8493 42891
rect 8527 42888 8539 42891
rect 8938 42888 8944 42900
rect 8527 42860 8944 42888
rect 8527 42857 8539 42860
rect 8481 42851 8539 42857
rect 8938 42848 8944 42860
rect 8996 42848 9002 42900
rect 9214 42848 9220 42900
rect 9272 42848 9278 42900
rect 9861 42891 9919 42897
rect 9861 42857 9873 42891
rect 9907 42888 9919 42891
rect 10134 42888 10140 42900
rect 9907 42860 10140 42888
rect 9907 42857 9919 42860
rect 9861 42851 9919 42857
rect 10134 42848 10140 42860
rect 10192 42848 10198 42900
rect 10689 42891 10747 42897
rect 10689 42857 10701 42891
rect 10735 42888 10747 42891
rect 10962 42888 10968 42900
rect 10735 42860 10968 42888
rect 10735 42857 10747 42860
rect 10689 42851 10747 42857
rect 10962 42848 10968 42860
rect 11020 42848 11026 42900
rect 11425 42891 11483 42897
rect 11425 42857 11437 42891
rect 11471 42888 11483 42891
rect 11606 42888 11612 42900
rect 11471 42860 11612 42888
rect 11471 42857 11483 42860
rect 11425 42851 11483 42857
rect 11606 42848 11612 42860
rect 11664 42848 11670 42900
rect 12161 42891 12219 42897
rect 12161 42857 12173 42891
rect 12207 42888 12219 42891
rect 12434 42888 12440 42900
rect 12207 42860 12440 42888
rect 12207 42857 12219 42860
rect 12161 42851 12219 42857
rect 12434 42848 12440 42860
rect 12492 42848 12498 42900
rect 13078 42848 13084 42900
rect 13136 42888 13142 42900
rect 13633 42891 13691 42897
rect 13633 42888 13645 42891
rect 13136 42860 13645 42888
rect 13136 42848 13142 42860
rect 13633 42857 13645 42860
rect 13679 42857 13691 42891
rect 13633 42851 13691 42857
rect 13449 42755 13507 42761
rect 13449 42721 13461 42755
rect 13495 42752 13507 42755
rect 14274 42752 14280 42764
rect 13495 42724 14280 42752
rect 13495 42721 13507 42724
rect 13449 42715 13507 42721
rect 14274 42712 14280 42724
rect 14332 42712 14338 42764
rect 3418 42644 3424 42696
rect 3476 42644 3482 42696
rect 4062 42644 4068 42696
rect 4120 42684 4126 42696
rect 4249 42687 4307 42693
rect 4249 42684 4261 42687
rect 4120 42656 4261 42684
rect 4120 42644 4126 42656
rect 4249 42653 4261 42656
rect 4295 42653 4307 42687
rect 4249 42647 4307 42653
rect 4982 42644 4988 42696
rect 5040 42644 5046 42696
rect 6454 42644 6460 42696
rect 6512 42644 6518 42696
rect 7190 42644 7196 42696
rect 7248 42644 7254 42696
rect 7926 42644 7932 42696
rect 7984 42644 7990 42696
rect 8662 42644 8668 42696
rect 8720 42644 8726 42696
rect 9401 42687 9459 42693
rect 9401 42653 9413 42687
rect 9447 42653 9459 42687
rect 9401 42647 9459 42653
rect 1394 42576 1400 42628
rect 1452 42576 1458 42628
rect 3602 42576 3608 42628
rect 3660 42616 3666 42628
rect 9416 42616 9444 42647
rect 10042 42644 10048 42696
rect 10100 42644 10106 42696
rect 10873 42687 10931 42693
rect 10873 42684 10885 42687
rect 10336 42656 10885 42684
rect 9677 42619 9735 42625
rect 9677 42616 9689 42619
rect 3660 42588 9689 42616
rect 3660 42576 3666 42588
rect 9677 42585 9689 42588
rect 9723 42585 9735 42619
rect 9677 42579 9735 42585
rect 10336 42560 10364 42656
rect 10873 42653 10885 42656
rect 10919 42653 10931 42687
rect 10873 42647 10931 42653
rect 11609 42687 11667 42693
rect 11609 42653 11621 42687
rect 11655 42653 11667 42687
rect 11609 42647 11667 42653
rect 10318 42508 10324 42560
rect 10376 42508 10382 42560
rect 11624 42548 11652 42647
rect 12342 42644 12348 42696
rect 12400 42644 12406 42696
rect 13814 42644 13820 42696
rect 13872 42644 13878 42696
rect 13170 42576 13176 42628
rect 13228 42576 13234 42628
rect 15562 42548 15568 42560
rect 11624 42520 15568 42548
rect 15562 42508 15568 42520
rect 15620 42508 15626 42560
rect 1104 42458 14696 42480
rect 1104 42406 4308 42458
rect 4360 42406 4372 42458
rect 4424 42406 4436 42458
rect 4488 42406 4500 42458
rect 4552 42406 4564 42458
rect 4616 42406 7666 42458
rect 7718 42406 7730 42458
rect 7782 42406 7794 42458
rect 7846 42406 7858 42458
rect 7910 42406 7922 42458
rect 7974 42406 11024 42458
rect 11076 42406 11088 42458
rect 11140 42406 11152 42458
rect 11204 42406 11216 42458
rect 11268 42406 11280 42458
rect 11332 42406 14382 42458
rect 14434 42406 14446 42458
rect 14498 42406 14510 42458
rect 14562 42406 14574 42458
rect 14626 42406 14638 42458
rect 14690 42406 14696 42458
rect 1104 42384 14696 42406
rect 1949 42347 2007 42353
rect 1949 42313 1961 42347
rect 1995 42344 2007 42347
rect 2038 42344 2044 42356
rect 1995 42316 2044 42344
rect 1995 42313 2007 42316
rect 1949 42307 2007 42313
rect 2038 42304 2044 42316
rect 2096 42304 2102 42356
rect 4062 42304 4068 42356
rect 4120 42304 4126 42356
rect 4709 42347 4767 42353
rect 4709 42313 4721 42347
rect 4755 42344 4767 42347
rect 4982 42344 4988 42356
rect 4755 42316 4988 42344
rect 4755 42313 4767 42316
rect 4709 42307 4767 42313
rect 4982 42304 4988 42316
rect 5040 42304 5046 42356
rect 5626 42304 5632 42356
rect 5684 42344 5690 42356
rect 12342 42344 12348 42356
rect 5684 42316 12348 42344
rect 5684 42304 5690 42316
rect 12342 42304 12348 42316
rect 12400 42304 12406 42356
rect 13357 42347 13415 42353
rect 13357 42313 13369 42347
rect 13403 42344 13415 42347
rect 13538 42344 13544 42356
rect 13403 42316 13544 42344
rect 13403 42313 13415 42316
rect 13357 42307 13415 42313
rect 13538 42304 13544 42316
rect 13596 42304 13602 42356
rect 13722 42304 13728 42356
rect 13780 42344 13786 42356
rect 13817 42347 13875 42353
rect 13817 42344 13829 42347
rect 13780 42316 13829 42344
rect 13780 42304 13786 42316
rect 13817 42313 13829 42316
rect 13863 42313 13875 42347
rect 13817 42307 13875 42313
rect 3970 42236 3976 42288
rect 4028 42276 4034 42288
rect 10318 42276 10324 42288
rect 4028 42248 10324 42276
rect 4028 42236 4034 42248
rect 10318 42236 10324 42248
rect 10376 42236 10382 42288
rect 2130 42168 2136 42220
rect 2188 42168 2194 42220
rect 4246 42168 4252 42220
rect 4304 42168 4310 42220
rect 4890 42168 4896 42220
rect 4948 42168 4954 42220
rect 13541 42211 13599 42217
rect 13541 42177 13553 42211
rect 13587 42177 13599 42211
rect 13541 42171 13599 42177
rect 13081 42143 13139 42149
rect 13081 42109 13093 42143
rect 13127 42140 13139 42143
rect 13556 42140 13584 42171
rect 13722 42168 13728 42220
rect 13780 42168 13786 42220
rect 13127 42112 15516 42140
rect 13127 42109 13139 42112
rect 13081 42103 13139 42109
rect 15488 42084 15516 42112
rect 15470 42032 15476 42084
rect 15528 42032 15534 42084
rect 1104 41914 14536 41936
rect 1104 41862 2629 41914
rect 2681 41862 2693 41914
rect 2745 41862 2757 41914
rect 2809 41862 2821 41914
rect 2873 41862 2885 41914
rect 2937 41862 5987 41914
rect 6039 41862 6051 41914
rect 6103 41862 6115 41914
rect 6167 41862 6179 41914
rect 6231 41862 6243 41914
rect 6295 41862 9345 41914
rect 9397 41862 9409 41914
rect 9461 41862 9473 41914
rect 9525 41862 9537 41914
rect 9589 41862 9601 41914
rect 9653 41862 12703 41914
rect 12755 41862 12767 41914
rect 12819 41862 12831 41914
rect 12883 41862 12895 41914
rect 12947 41862 12959 41914
rect 13011 41862 14536 41914
rect 1104 41840 14536 41862
rect 13081 41803 13139 41809
rect 13081 41769 13093 41803
rect 13127 41800 13139 41803
rect 13170 41800 13176 41812
rect 13127 41772 13176 41800
rect 13127 41769 13139 41772
rect 13081 41763 13139 41769
rect 13170 41760 13176 41772
rect 13228 41760 13234 41812
rect 13633 41803 13691 41809
rect 13633 41769 13645 41803
rect 13679 41800 13691 41803
rect 13722 41800 13728 41812
rect 13679 41772 13728 41800
rect 13679 41769 13691 41772
rect 13633 41763 13691 41769
rect 13722 41760 13728 41772
rect 13780 41760 13786 41812
rect 13265 41599 13323 41605
rect 13265 41565 13277 41599
rect 13311 41565 13323 41599
rect 13265 41559 13323 41565
rect 13817 41599 13875 41605
rect 13817 41565 13829 41599
rect 13863 41596 13875 41599
rect 14734 41596 14740 41608
rect 13863 41568 14740 41596
rect 13863 41565 13875 41568
rect 13817 41559 13875 41565
rect 13280 41528 13308 41559
rect 14734 41556 14740 41568
rect 14792 41556 14798 41608
rect 13998 41528 14004 41540
rect 13280 41500 14004 41528
rect 13998 41488 14004 41500
rect 14056 41488 14062 41540
rect 1104 41370 14696 41392
rect 1104 41318 4308 41370
rect 4360 41318 4372 41370
rect 4424 41318 4436 41370
rect 4488 41318 4500 41370
rect 4552 41318 4564 41370
rect 4616 41318 7666 41370
rect 7718 41318 7730 41370
rect 7782 41318 7794 41370
rect 7846 41318 7858 41370
rect 7910 41318 7922 41370
rect 7974 41318 11024 41370
rect 11076 41318 11088 41370
rect 11140 41318 11152 41370
rect 11204 41318 11216 41370
rect 11268 41318 11280 41370
rect 11332 41318 14382 41370
rect 14434 41318 14446 41370
rect 14498 41318 14510 41370
rect 14562 41318 14574 41370
rect 14626 41318 14638 41370
rect 14690 41318 14696 41370
rect 1104 41296 14696 41318
rect 750 41080 756 41132
rect 808 41120 814 41132
rect 1397 41123 1455 41129
rect 1397 41120 1409 41123
rect 808 41092 1409 41120
rect 808 41080 814 41092
rect 1397 41089 1409 41092
rect 1443 41089 1455 41123
rect 1397 41083 1455 41089
rect 1581 40919 1639 40925
rect 1581 40885 1593 40919
rect 1627 40916 1639 40919
rect 6362 40916 6368 40928
rect 1627 40888 6368 40916
rect 1627 40885 1639 40888
rect 1581 40879 1639 40885
rect 6362 40876 6368 40888
rect 6420 40876 6426 40928
rect 1104 40826 14536 40848
rect 1104 40774 2629 40826
rect 2681 40774 2693 40826
rect 2745 40774 2757 40826
rect 2809 40774 2821 40826
rect 2873 40774 2885 40826
rect 2937 40774 5987 40826
rect 6039 40774 6051 40826
rect 6103 40774 6115 40826
rect 6167 40774 6179 40826
rect 6231 40774 6243 40826
rect 6295 40774 9345 40826
rect 9397 40774 9409 40826
rect 9461 40774 9473 40826
rect 9525 40774 9537 40826
rect 9589 40774 9601 40826
rect 9653 40774 12703 40826
rect 12755 40774 12767 40826
rect 12819 40774 12831 40826
rect 12883 40774 12895 40826
rect 12947 40774 12959 40826
rect 13011 40774 14536 40826
rect 1104 40752 14536 40774
rect 1104 40282 14696 40304
rect 1104 40230 4308 40282
rect 4360 40230 4372 40282
rect 4424 40230 4436 40282
rect 4488 40230 4500 40282
rect 4552 40230 4564 40282
rect 4616 40230 7666 40282
rect 7718 40230 7730 40282
rect 7782 40230 7794 40282
rect 7846 40230 7858 40282
rect 7910 40230 7922 40282
rect 7974 40230 11024 40282
rect 11076 40230 11088 40282
rect 11140 40230 11152 40282
rect 11204 40230 11216 40282
rect 11268 40230 11280 40282
rect 11332 40230 14382 40282
rect 14434 40230 14446 40282
rect 14498 40230 14510 40282
rect 14562 40230 14574 40282
rect 14626 40230 14638 40282
rect 14690 40230 14696 40282
rect 1104 40208 14696 40230
rect 1486 40060 1492 40112
rect 1544 40060 1550 40112
rect 7466 39992 7472 40044
rect 7524 40032 7530 40044
rect 13449 40035 13507 40041
rect 13449 40032 13461 40035
rect 7524 40004 13461 40032
rect 7524 39992 7530 40004
rect 13449 40001 13461 40004
rect 13495 40001 13507 40035
rect 13449 39995 13507 40001
rect 13814 39992 13820 40044
rect 13872 39992 13878 40044
rect 1673 39899 1731 39905
rect 1673 39865 1685 39899
rect 1719 39896 1731 39899
rect 4706 39896 4712 39908
rect 1719 39868 4712 39896
rect 1719 39865 1731 39868
rect 1673 39859 1731 39865
rect 4706 39856 4712 39868
rect 4764 39856 4770 39908
rect 13262 39788 13268 39840
rect 13320 39788 13326 39840
rect 14090 39788 14096 39840
rect 14148 39788 14154 39840
rect 1104 39738 14536 39760
rect 1104 39686 2629 39738
rect 2681 39686 2693 39738
rect 2745 39686 2757 39738
rect 2809 39686 2821 39738
rect 2873 39686 2885 39738
rect 2937 39686 5987 39738
rect 6039 39686 6051 39738
rect 6103 39686 6115 39738
rect 6167 39686 6179 39738
rect 6231 39686 6243 39738
rect 6295 39686 9345 39738
rect 9397 39686 9409 39738
rect 9461 39686 9473 39738
rect 9525 39686 9537 39738
rect 9589 39686 9601 39738
rect 9653 39686 12703 39738
rect 12755 39686 12767 39738
rect 12819 39686 12831 39738
rect 12883 39686 12895 39738
rect 12947 39686 12959 39738
rect 13011 39686 14536 39738
rect 1104 39664 14536 39686
rect 6362 39584 6368 39636
rect 6420 39624 6426 39636
rect 6730 39624 6736 39636
rect 6420 39596 6736 39624
rect 6420 39584 6426 39596
rect 6730 39584 6736 39596
rect 6788 39624 6794 39636
rect 9493 39627 9551 39633
rect 6788 39596 8708 39624
rect 6788 39584 6794 39596
rect 7745 39559 7803 39565
rect 7745 39525 7757 39559
rect 7791 39525 7803 39559
rect 7745 39519 7803 39525
rect 7760 39488 7788 39519
rect 7760 39460 8616 39488
rect 4706 39380 4712 39432
rect 4764 39420 4770 39432
rect 8588 39429 8616 39460
rect 7929 39423 7987 39429
rect 7929 39420 7941 39423
rect 4764 39392 7941 39420
rect 4764 39380 4770 39392
rect 7929 39389 7941 39392
rect 7975 39389 7987 39423
rect 7929 39383 7987 39389
rect 8573 39423 8631 39429
rect 8573 39389 8585 39423
rect 8619 39389 8631 39423
rect 8680 39420 8708 39596
rect 9493 39593 9505 39627
rect 9539 39624 9551 39627
rect 13814 39624 13820 39636
rect 9539 39596 13820 39624
rect 9539 39593 9551 39596
rect 9493 39587 9551 39593
rect 13814 39584 13820 39596
rect 13872 39584 13878 39636
rect 8941 39559 8999 39565
rect 8941 39525 8953 39559
rect 8987 39525 8999 39559
rect 8941 39519 8999 39525
rect 8956 39488 8984 39519
rect 8956 39460 9720 39488
rect 9692 39429 9720 39460
rect 9125 39423 9183 39429
rect 9125 39420 9137 39423
rect 8680 39392 9137 39420
rect 8573 39383 8631 39389
rect 9125 39389 9137 39392
rect 9171 39389 9183 39423
rect 9125 39383 9183 39389
rect 9677 39423 9735 39429
rect 9677 39389 9689 39423
rect 9723 39389 9735 39423
rect 9677 39383 9735 39389
rect 12894 39380 12900 39432
rect 12952 39380 12958 39432
rect 750 39312 756 39364
rect 808 39352 814 39364
rect 1489 39355 1547 39361
rect 1489 39352 1501 39355
rect 808 39324 1501 39352
rect 808 39312 814 39324
rect 1489 39321 1501 39324
rect 1535 39321 1547 39355
rect 1489 39315 1547 39321
rect 1857 39355 1915 39361
rect 1857 39321 1869 39355
rect 1903 39352 1915 39355
rect 7466 39352 7472 39364
rect 1903 39324 7472 39352
rect 1903 39321 1915 39324
rect 1857 39315 1915 39321
rect 7466 39312 7472 39324
rect 7524 39312 7530 39364
rect 13357 39355 13415 39361
rect 13357 39352 13369 39355
rect 8404 39324 13369 39352
rect 8404 39293 8432 39324
rect 13357 39321 13369 39324
rect 13403 39321 13415 39355
rect 13357 39315 13415 39321
rect 13725 39355 13783 39361
rect 13725 39321 13737 39355
rect 13771 39352 13783 39355
rect 14826 39352 14832 39364
rect 13771 39324 14832 39352
rect 13771 39321 13783 39324
rect 13725 39315 13783 39321
rect 14826 39312 14832 39324
rect 14884 39312 14890 39364
rect 8389 39287 8447 39293
rect 8389 39253 8401 39287
rect 8435 39253 8447 39287
rect 8389 39247 8447 39253
rect 13081 39287 13139 39293
rect 13081 39253 13093 39287
rect 13127 39284 13139 39287
rect 14274 39284 14280 39296
rect 13127 39256 14280 39284
rect 13127 39253 13139 39256
rect 13081 39247 13139 39253
rect 14274 39244 14280 39256
rect 14332 39244 14338 39296
rect 1104 39194 14696 39216
rect 1104 39142 4308 39194
rect 4360 39142 4372 39194
rect 4424 39142 4436 39194
rect 4488 39142 4500 39194
rect 4552 39142 4564 39194
rect 4616 39142 7666 39194
rect 7718 39142 7730 39194
rect 7782 39142 7794 39194
rect 7846 39142 7858 39194
rect 7910 39142 7922 39194
rect 7974 39142 11024 39194
rect 11076 39142 11088 39194
rect 11140 39142 11152 39194
rect 11204 39142 11216 39194
rect 11268 39142 11280 39194
rect 11332 39142 14382 39194
rect 14434 39142 14446 39194
rect 14498 39142 14510 39194
rect 14562 39142 14574 39194
rect 14626 39142 14638 39194
rect 14690 39142 14696 39194
rect 1104 39120 14696 39142
rect 12437 39083 12495 39089
rect 12437 39049 12449 39083
rect 12483 39080 12495 39083
rect 12894 39080 12900 39092
rect 12483 39052 12900 39080
rect 12483 39049 12495 39052
rect 12437 39043 12495 39049
rect 12894 39040 12900 39052
rect 12952 39040 12958 39092
rect 13262 39040 13268 39092
rect 13320 39040 13326 39092
rect 13280 39012 13308 39040
rect 12636 38984 13308 39012
rect 12636 38953 12664 38984
rect 12621 38947 12679 38953
rect 12621 38913 12633 38947
rect 12667 38913 12679 38947
rect 12621 38907 12679 38913
rect 12897 38947 12955 38953
rect 12897 38913 12909 38947
rect 12943 38913 12955 38947
rect 12897 38907 12955 38913
rect 13081 38947 13139 38953
rect 13081 38913 13093 38947
rect 13127 38913 13139 38947
rect 13081 38907 13139 38913
rect 12250 38836 12256 38888
rect 12308 38876 12314 38888
rect 12912 38876 12940 38907
rect 12308 38848 12940 38876
rect 12308 38836 12314 38848
rect 12434 38768 12440 38820
rect 12492 38808 12498 38820
rect 13096 38808 13124 38907
rect 13630 38904 13636 38956
rect 13688 38904 13694 38956
rect 12492 38780 13124 38808
rect 12492 38768 12498 38780
rect 12713 38743 12771 38749
rect 12713 38709 12725 38743
rect 12759 38740 12771 38743
rect 13078 38740 13084 38752
rect 12759 38712 13084 38740
rect 12759 38709 12771 38712
rect 12713 38703 12771 38709
rect 13078 38700 13084 38712
rect 13136 38700 13142 38752
rect 13354 38700 13360 38752
rect 13412 38700 13418 38752
rect 13906 38700 13912 38752
rect 13964 38700 13970 38752
rect 1104 38650 14536 38672
rect 1104 38598 2629 38650
rect 2681 38598 2693 38650
rect 2745 38598 2757 38650
rect 2809 38598 2821 38650
rect 2873 38598 2885 38650
rect 2937 38598 5987 38650
rect 6039 38598 6051 38650
rect 6103 38598 6115 38650
rect 6167 38598 6179 38650
rect 6231 38598 6243 38650
rect 6295 38598 9345 38650
rect 9397 38598 9409 38650
rect 9461 38598 9473 38650
rect 9525 38598 9537 38650
rect 9589 38598 9601 38650
rect 9653 38598 12703 38650
rect 12755 38598 12767 38650
rect 12819 38598 12831 38650
rect 12883 38598 12895 38650
rect 12947 38598 12959 38650
rect 13011 38598 14536 38650
rect 1104 38576 14536 38598
rect 12345 38539 12403 38545
rect 12345 38505 12357 38539
rect 12391 38536 12403 38539
rect 13630 38536 13636 38548
rect 12391 38508 13636 38536
rect 12391 38505 12403 38508
rect 12345 38499 12403 38505
rect 13630 38496 13636 38508
rect 13688 38496 13694 38548
rect 12069 38471 12127 38477
rect 12069 38437 12081 38471
rect 12115 38437 12127 38471
rect 12069 38431 12127 38437
rect 12084 38400 12112 38431
rect 12158 38428 12164 38480
rect 12216 38468 12222 38480
rect 13446 38468 13452 38480
rect 12216 38440 13452 38468
rect 12216 38428 12222 38440
rect 13446 38428 13452 38440
rect 13504 38428 13510 38480
rect 12084 38372 12434 38400
rect 750 38292 756 38344
rect 808 38332 814 38344
rect 1397 38335 1455 38341
rect 1397 38332 1409 38335
rect 808 38304 1409 38332
rect 808 38292 814 38304
rect 1397 38301 1409 38304
rect 1443 38301 1455 38335
rect 11790 38332 11796 38344
rect 1397 38295 1455 38301
rect 2746 38304 11796 38332
rect 1581 38199 1639 38205
rect 1581 38165 1593 38199
rect 1627 38196 1639 38199
rect 2746 38196 2774 38304
rect 11790 38292 11796 38304
rect 11848 38332 11854 38344
rect 12253 38335 12311 38341
rect 12253 38332 12265 38335
rect 11848 38304 12265 38332
rect 11848 38292 11854 38304
rect 12253 38301 12265 38304
rect 12299 38301 12311 38335
rect 12406 38332 12434 38372
rect 12529 38335 12587 38341
rect 12529 38332 12541 38335
rect 12406 38304 12541 38332
rect 12253 38295 12311 38301
rect 12529 38301 12541 38304
rect 12575 38301 12587 38335
rect 12529 38295 12587 38301
rect 12618 38292 12624 38344
rect 12676 38332 12682 38344
rect 12805 38335 12863 38341
rect 12805 38332 12817 38335
rect 12676 38304 12817 38332
rect 12676 38292 12682 38304
rect 12805 38301 12817 38304
rect 12851 38301 12863 38335
rect 12805 38295 12863 38301
rect 12897 38335 12955 38341
rect 12897 38301 12909 38335
rect 12943 38301 12955 38335
rect 12897 38295 12955 38301
rect 11882 38224 11888 38276
rect 11940 38264 11946 38276
rect 12912 38264 12940 38295
rect 11940 38236 12940 38264
rect 11940 38224 11946 38236
rect 13354 38224 13360 38276
rect 13412 38224 13418 38276
rect 13725 38267 13783 38273
rect 13725 38233 13737 38267
rect 13771 38264 13783 38267
rect 14826 38264 14832 38276
rect 13771 38236 14832 38264
rect 13771 38233 13783 38236
rect 13725 38227 13783 38233
rect 14826 38224 14832 38236
rect 14884 38224 14890 38276
rect 1627 38168 2774 38196
rect 1627 38165 1639 38168
rect 1581 38159 1639 38165
rect 12618 38156 12624 38208
rect 12676 38156 12682 38208
rect 13081 38199 13139 38205
rect 13081 38165 13093 38199
rect 13127 38196 13139 38199
rect 14274 38196 14280 38208
rect 13127 38168 14280 38196
rect 13127 38165 13139 38168
rect 13081 38159 13139 38165
rect 14274 38156 14280 38168
rect 14332 38156 14338 38208
rect 1104 38106 14696 38128
rect 1104 38054 4308 38106
rect 4360 38054 4372 38106
rect 4424 38054 4436 38106
rect 4488 38054 4500 38106
rect 4552 38054 4564 38106
rect 4616 38054 7666 38106
rect 7718 38054 7730 38106
rect 7782 38054 7794 38106
rect 7846 38054 7858 38106
rect 7910 38054 7922 38106
rect 7974 38054 11024 38106
rect 11076 38054 11088 38106
rect 11140 38054 11152 38106
rect 11204 38054 11216 38106
rect 11268 38054 11280 38106
rect 11332 38054 14382 38106
rect 14434 38054 14446 38106
rect 14498 38054 14510 38106
rect 14562 38054 14574 38106
rect 14626 38054 14638 38106
rect 14690 38054 14696 38106
rect 1104 38032 14696 38054
rect 11517 37995 11575 38001
rect 11517 37961 11529 37995
rect 11563 37961 11575 37995
rect 11517 37955 11575 37961
rect 11532 37924 11560 37955
rect 11882 37952 11888 38004
rect 11940 37952 11946 38004
rect 12161 37995 12219 38001
rect 12161 37961 12173 37995
rect 12207 37992 12219 37995
rect 12342 37992 12348 38004
rect 12207 37964 12348 37992
rect 12207 37961 12219 37964
rect 12161 37955 12219 37961
rect 12342 37952 12348 37964
rect 12400 37952 12406 38004
rect 12437 37995 12495 38001
rect 12437 37961 12449 37995
rect 12483 37961 12495 37995
rect 12437 37955 12495 37961
rect 12452 37924 12480 37955
rect 12618 37952 12624 38004
rect 12676 37952 12682 38004
rect 13354 37952 13360 38004
rect 13412 37952 13418 38004
rect 13446 37952 13452 38004
rect 13504 37952 13510 38004
rect 11532 37896 12020 37924
rect 750 37816 756 37868
rect 808 37856 814 37868
rect 1397 37859 1455 37865
rect 1397 37856 1409 37859
rect 808 37828 1409 37856
rect 808 37816 814 37828
rect 1397 37825 1409 37828
rect 1443 37825 1455 37859
rect 1397 37819 1455 37825
rect 10318 37816 10324 37868
rect 10376 37856 10382 37868
rect 11149 37859 11207 37865
rect 11149 37856 11161 37859
rect 10376 37828 11161 37856
rect 10376 37816 10382 37828
rect 11149 37825 11161 37828
rect 11195 37825 11207 37859
rect 11701 37859 11759 37865
rect 11701 37856 11713 37859
rect 11149 37819 11207 37825
rect 11256 37828 11713 37856
rect 10410 37788 10416 37800
rect 2746 37760 10416 37788
rect 1581 37655 1639 37661
rect 1581 37621 1593 37655
rect 1627 37652 1639 37655
rect 2746 37652 2774 37760
rect 10410 37748 10416 37760
rect 10468 37788 10474 37800
rect 11256 37788 11284 37828
rect 11701 37825 11713 37828
rect 11747 37825 11759 37859
rect 11701 37819 11759 37825
rect 10468 37760 11284 37788
rect 11992 37788 12020 37896
rect 12084 37896 12480 37924
rect 12636 37924 12664 37952
rect 12636 37896 12756 37924
rect 12084 37865 12112 37896
rect 12069 37859 12127 37865
rect 12069 37825 12081 37859
rect 12115 37825 12127 37859
rect 12069 37819 12127 37825
rect 12345 37859 12403 37865
rect 12345 37825 12357 37859
rect 12391 37825 12403 37859
rect 12345 37819 12403 37825
rect 12360 37788 12388 37819
rect 12618 37816 12624 37868
rect 12676 37816 12682 37868
rect 12728 37865 12756 37896
rect 13078 37884 13084 37936
rect 13136 37924 13142 37936
rect 13173 37927 13231 37933
rect 13173 37924 13185 37927
rect 13136 37896 13185 37924
rect 13136 37884 13142 37896
rect 13173 37893 13185 37896
rect 13219 37893 13231 37927
rect 13173 37887 13231 37893
rect 12713 37859 12771 37865
rect 12713 37825 12725 37859
rect 12759 37825 12771 37859
rect 12713 37819 12771 37825
rect 13372 37788 13400 37952
rect 13464 37924 13492 37952
rect 13725 37927 13783 37933
rect 13725 37924 13737 37927
rect 13464 37896 13737 37924
rect 13725 37893 13737 37896
rect 13771 37893 13783 37927
rect 13725 37887 13783 37893
rect 13541 37859 13599 37865
rect 13541 37825 13553 37859
rect 13587 37825 13599 37859
rect 13541 37819 13599 37825
rect 11992 37760 12388 37788
rect 12820 37760 13400 37788
rect 13556 37788 13584 37819
rect 14366 37788 14372 37800
rect 13556 37760 14372 37788
rect 10468 37748 10474 37760
rect 10980 37692 12434 37720
rect 10980 37661 11008 37692
rect 1627 37624 2774 37652
rect 10965 37655 11023 37661
rect 1627 37621 1639 37624
rect 1581 37615 1639 37621
rect 10965 37621 10977 37655
rect 11011 37621 11023 37655
rect 12406 37652 12434 37692
rect 12820 37652 12848 37760
rect 14366 37748 14372 37760
rect 14424 37748 14430 37800
rect 14182 37720 14188 37732
rect 12912 37692 14188 37720
rect 12912 37661 12940 37692
rect 14182 37680 14188 37692
rect 14240 37680 14246 37732
rect 12406 37624 12848 37652
rect 12897 37655 12955 37661
rect 10965 37615 11023 37621
rect 12897 37621 12909 37655
rect 12943 37621 12955 37655
rect 12897 37615 12955 37621
rect 13722 37612 13728 37664
rect 13780 37652 13786 37664
rect 14001 37655 14059 37661
rect 14001 37652 14013 37655
rect 13780 37624 14013 37652
rect 13780 37612 13786 37624
rect 14001 37621 14013 37624
rect 14047 37621 14059 37655
rect 14001 37615 14059 37621
rect 1104 37562 14536 37584
rect 1104 37510 2629 37562
rect 2681 37510 2693 37562
rect 2745 37510 2757 37562
rect 2809 37510 2821 37562
rect 2873 37510 2885 37562
rect 2937 37510 5987 37562
rect 6039 37510 6051 37562
rect 6103 37510 6115 37562
rect 6167 37510 6179 37562
rect 6231 37510 6243 37562
rect 6295 37510 9345 37562
rect 9397 37510 9409 37562
rect 9461 37510 9473 37562
rect 9525 37510 9537 37562
rect 9589 37510 9601 37562
rect 9653 37510 12703 37562
rect 12755 37510 12767 37562
rect 12819 37510 12831 37562
rect 12883 37510 12895 37562
rect 12947 37510 12959 37562
rect 13011 37510 14536 37562
rect 1104 37488 14536 37510
rect 10318 37408 10324 37460
rect 10376 37408 10382 37460
rect 10502 37408 10508 37460
rect 10560 37448 10566 37460
rect 12618 37448 12624 37460
rect 10560 37420 12624 37448
rect 10560 37408 10566 37420
rect 12618 37408 12624 37420
rect 12676 37408 12682 37460
rect 12250 37340 12256 37392
rect 12308 37340 12314 37392
rect 12342 37272 12348 37324
rect 12400 37312 12406 37324
rect 12400 37284 13032 37312
rect 12400 37272 12406 37284
rect 8294 37204 8300 37256
rect 8352 37244 8358 37256
rect 10505 37247 10563 37253
rect 10505 37244 10517 37247
rect 8352 37216 10517 37244
rect 8352 37204 8358 37216
rect 10505 37213 10517 37216
rect 10551 37213 10563 37247
rect 10505 37207 10563 37213
rect 11882 37204 11888 37256
rect 11940 37204 11946 37256
rect 12161 37247 12219 37253
rect 12161 37220 12173 37247
rect 12084 37213 12173 37220
rect 12207 37213 12219 37247
rect 12084 37207 12219 37213
rect 12437 37247 12495 37253
rect 12437 37213 12449 37247
rect 12483 37244 12495 37247
rect 12618 37244 12624 37256
rect 12483 37216 12624 37244
rect 12483 37213 12495 37216
rect 12437 37207 12495 37213
rect 12084 37192 12204 37207
rect 12618 37204 12624 37216
rect 12676 37204 12682 37256
rect 12710 37204 12716 37256
rect 12768 37204 12774 37256
rect 13004 37253 13032 37284
rect 12989 37247 13047 37253
rect 12989 37213 13001 37247
rect 13035 37213 13047 37247
rect 12989 37207 13047 37213
rect 1578 37136 1584 37188
rect 1636 37176 1642 37188
rect 12084 37176 12112 37192
rect 1636 37148 12112 37176
rect 1636 37136 1642 37148
rect 13354 37136 13360 37188
rect 13412 37136 13418 37188
rect 13538 37136 13544 37188
rect 13596 37136 13602 37188
rect 11698 37068 11704 37120
rect 11756 37068 11762 37120
rect 11974 37068 11980 37120
rect 12032 37068 12038 37120
rect 12066 37068 12072 37120
rect 12124 37108 12130 37120
rect 12529 37111 12587 37117
rect 12529 37108 12541 37111
rect 12124 37080 12541 37108
rect 12124 37068 12130 37080
rect 12529 37077 12541 37080
rect 12575 37077 12587 37111
rect 12529 37071 12587 37077
rect 13630 37068 13636 37120
rect 13688 37068 13694 37120
rect 1104 37018 14696 37040
rect 1104 36966 4308 37018
rect 4360 36966 4372 37018
rect 4424 36966 4436 37018
rect 4488 36966 4500 37018
rect 4552 36966 4564 37018
rect 4616 36966 7666 37018
rect 7718 36966 7730 37018
rect 7782 36966 7794 37018
rect 7846 36966 7858 37018
rect 7910 36966 7922 37018
rect 7974 36966 11024 37018
rect 11076 36966 11088 37018
rect 11140 36966 11152 37018
rect 11204 36966 11216 37018
rect 11268 36966 11280 37018
rect 11332 36966 14382 37018
rect 14434 36966 14446 37018
rect 14498 36966 14510 37018
rect 14562 36966 14574 37018
rect 14626 36966 14638 37018
rect 14690 36966 14696 37018
rect 1104 36944 14696 36966
rect 1581 36907 1639 36913
rect 1581 36873 1593 36907
rect 1627 36904 1639 36907
rect 8294 36904 8300 36916
rect 1627 36876 8300 36904
rect 1627 36873 1639 36876
rect 1581 36867 1639 36873
rect 8294 36864 8300 36876
rect 8352 36864 8358 36916
rect 12253 36907 12311 36913
rect 12253 36873 12265 36907
rect 12299 36904 12311 36907
rect 13538 36904 13544 36916
rect 12299 36876 13544 36904
rect 12299 36873 12311 36876
rect 12253 36867 12311 36873
rect 13538 36864 13544 36876
rect 13596 36864 13602 36916
rect 10594 36796 10600 36848
rect 10652 36836 10658 36848
rect 13725 36839 13783 36845
rect 13725 36836 13737 36839
rect 10652 36808 13737 36836
rect 10652 36796 10658 36808
rect 13725 36805 13737 36808
rect 13771 36805 13783 36839
rect 13725 36799 13783 36805
rect 750 36728 756 36780
rect 808 36768 814 36780
rect 1397 36771 1455 36777
rect 1397 36768 1409 36771
rect 808 36740 1409 36768
rect 808 36728 814 36740
rect 1397 36737 1409 36740
rect 1443 36737 1455 36771
rect 1397 36731 1455 36737
rect 1946 36728 1952 36780
rect 2004 36728 2010 36780
rect 9766 36728 9772 36780
rect 9824 36768 9830 36780
rect 11885 36771 11943 36777
rect 11885 36768 11897 36771
rect 9824 36740 11897 36768
rect 9824 36728 9830 36740
rect 11885 36737 11897 36740
rect 11931 36737 11943 36771
rect 11885 36731 11943 36737
rect 11974 36728 11980 36780
rect 12032 36768 12038 36780
rect 12161 36771 12219 36777
rect 12161 36768 12173 36771
rect 12032 36740 12173 36768
rect 12032 36728 12038 36740
rect 12161 36737 12173 36740
rect 12207 36737 12219 36771
rect 12161 36731 12219 36737
rect 12434 36728 12440 36780
rect 12492 36728 12498 36780
rect 12526 36728 12532 36780
rect 12584 36768 12590 36780
rect 12713 36771 12771 36777
rect 12713 36768 12725 36771
rect 12584 36740 12725 36768
rect 12584 36728 12590 36740
rect 12713 36737 12725 36740
rect 12759 36737 12771 36771
rect 12713 36731 12771 36737
rect 13173 36771 13231 36777
rect 13173 36737 13185 36771
rect 13219 36737 13231 36771
rect 13173 36731 13231 36737
rect 13541 36771 13599 36777
rect 13541 36737 13553 36771
rect 13587 36768 13599 36771
rect 15010 36768 15016 36780
rect 13587 36740 15016 36768
rect 13587 36737 13599 36740
rect 13541 36731 13599 36737
rect 10226 36660 10232 36712
rect 10284 36700 10290 36712
rect 13188 36700 13216 36731
rect 15010 36728 15016 36740
rect 15068 36728 15074 36780
rect 10284 36672 13216 36700
rect 10284 36660 10290 36672
rect 1762 36592 1768 36644
rect 1820 36592 1826 36644
rect 11701 36635 11759 36641
rect 11701 36601 11713 36635
rect 11747 36632 11759 36635
rect 12802 36632 12808 36644
rect 11747 36604 12808 36632
rect 11747 36601 11759 36604
rect 11701 36595 11759 36601
rect 12802 36592 12808 36604
rect 12860 36592 12866 36644
rect 14182 36632 14188 36644
rect 12912 36604 14188 36632
rect 11977 36567 12035 36573
rect 11977 36533 11989 36567
rect 12023 36564 12035 36567
rect 12158 36564 12164 36576
rect 12023 36536 12164 36564
rect 12023 36533 12035 36536
rect 11977 36527 12035 36533
rect 12158 36524 12164 36536
rect 12216 36524 12222 36576
rect 12912 36573 12940 36604
rect 14182 36592 14188 36604
rect 14240 36592 14246 36644
rect 12897 36567 12955 36573
rect 12897 36533 12909 36567
rect 12943 36533 12955 36567
rect 12897 36527 12955 36533
rect 13538 36524 13544 36576
rect 13596 36564 13602 36576
rect 14001 36567 14059 36573
rect 14001 36564 14013 36567
rect 13596 36536 14013 36564
rect 13596 36524 13602 36536
rect 14001 36533 14013 36536
rect 14047 36533 14059 36567
rect 14001 36527 14059 36533
rect 1104 36474 14536 36496
rect 1104 36422 2629 36474
rect 2681 36422 2693 36474
rect 2745 36422 2757 36474
rect 2809 36422 2821 36474
rect 2873 36422 2885 36474
rect 2937 36422 5987 36474
rect 6039 36422 6051 36474
rect 6103 36422 6115 36474
rect 6167 36422 6179 36474
rect 6231 36422 6243 36474
rect 6295 36422 9345 36474
rect 9397 36422 9409 36474
rect 9461 36422 9473 36474
rect 9525 36422 9537 36474
rect 9589 36422 9601 36474
rect 9653 36422 12703 36474
rect 12755 36422 12767 36474
rect 12819 36422 12831 36474
rect 12883 36422 12895 36474
rect 12947 36422 12959 36474
rect 13011 36422 14536 36474
rect 1104 36400 14536 36422
rect 1946 36320 1952 36372
rect 2004 36320 2010 36372
rect 3694 36360 3700 36372
rect 2746 36332 3700 36360
rect 1765 36227 1823 36233
rect 1765 36193 1777 36227
rect 1811 36224 1823 36227
rect 2746 36224 2774 36332
rect 3694 36320 3700 36332
rect 3752 36360 3758 36372
rect 10502 36360 10508 36372
rect 3752 36332 10508 36360
rect 3752 36320 3758 36332
rect 10502 36320 10508 36332
rect 10560 36320 10566 36372
rect 11885 36363 11943 36369
rect 11885 36329 11897 36363
rect 11931 36360 11943 36363
rect 12434 36360 12440 36372
rect 11931 36332 12440 36360
rect 11931 36329 11943 36332
rect 11885 36323 11943 36329
rect 12434 36320 12440 36332
rect 12492 36320 12498 36372
rect 11333 36295 11391 36301
rect 11333 36261 11345 36295
rect 11379 36292 11391 36295
rect 11379 36264 12434 36292
rect 11379 36261 11391 36264
rect 11333 36255 11391 36261
rect 1811 36196 2774 36224
rect 1811 36193 1823 36196
rect 1765 36187 1823 36193
rect 10502 36184 10508 36236
rect 10560 36224 10566 36236
rect 10560 36196 12112 36224
rect 10560 36184 10566 36196
rect 2133 36159 2191 36165
rect 2133 36125 2145 36159
rect 2179 36156 2191 36159
rect 7374 36156 7380 36168
rect 2179 36128 7380 36156
rect 2179 36125 2191 36128
rect 2133 36119 2191 36125
rect 7374 36116 7380 36128
rect 7432 36116 7438 36168
rect 10870 36116 10876 36168
rect 10928 36156 10934 36168
rect 12084 36165 12112 36196
rect 11517 36159 11575 36165
rect 11517 36156 11529 36159
rect 10928 36128 11529 36156
rect 10928 36116 10934 36128
rect 11517 36125 11529 36128
rect 11563 36125 11575 36159
rect 11517 36119 11575 36125
rect 11793 36159 11851 36165
rect 11793 36125 11805 36159
rect 11839 36156 11851 36159
rect 12069 36159 12127 36165
rect 11839 36128 11928 36156
rect 11839 36125 11851 36128
rect 11793 36119 11851 36125
rect 1486 36048 1492 36100
rect 1544 36048 1550 36100
rect 11900 36032 11928 36128
rect 12069 36125 12081 36159
rect 12115 36125 12127 36159
rect 12406 36156 12434 36264
rect 12805 36159 12863 36165
rect 12805 36156 12817 36159
rect 12406 36128 12817 36156
rect 12069 36119 12127 36125
rect 12805 36125 12817 36128
rect 12851 36125 12863 36159
rect 12805 36119 12863 36125
rect 12250 36048 12256 36100
rect 12308 36048 12314 36100
rect 12618 36048 12624 36100
rect 12676 36048 12682 36100
rect 13170 36048 13176 36100
rect 13228 36048 13234 36100
rect 13354 36048 13360 36100
rect 13412 36048 13418 36100
rect 13722 36048 13728 36100
rect 13780 36048 13786 36100
rect 11609 36023 11667 36029
rect 11609 35989 11621 36023
rect 11655 36020 11667 36023
rect 11790 36020 11796 36032
rect 11655 35992 11796 36020
rect 11655 35989 11667 35992
rect 11609 35983 11667 35989
rect 11790 35980 11796 35992
rect 11848 35980 11854 36032
rect 11882 35980 11888 36032
rect 11940 35980 11946 36032
rect 1104 35930 14696 35952
rect 1104 35878 4308 35930
rect 4360 35878 4372 35930
rect 4424 35878 4436 35930
rect 4488 35878 4500 35930
rect 4552 35878 4564 35930
rect 4616 35878 7666 35930
rect 7718 35878 7730 35930
rect 7782 35878 7794 35930
rect 7846 35878 7858 35930
rect 7910 35878 7922 35930
rect 7974 35878 11024 35930
rect 11076 35878 11088 35930
rect 11140 35878 11152 35930
rect 11204 35878 11216 35930
rect 11268 35878 11280 35930
rect 11332 35878 14382 35930
rect 14434 35878 14446 35930
rect 14498 35878 14510 35930
rect 14562 35878 14574 35930
rect 14626 35878 14638 35930
rect 14690 35878 14696 35930
rect 1104 35856 14696 35878
rect 10226 35776 10232 35828
rect 10284 35776 10290 35828
rect 10594 35776 10600 35828
rect 10652 35776 10658 35828
rect 10870 35776 10876 35828
rect 10928 35776 10934 35828
rect 11149 35819 11207 35825
rect 11149 35785 11161 35819
rect 11195 35785 11207 35819
rect 11149 35779 11207 35785
rect 11164 35748 11192 35779
rect 11238 35776 11244 35828
rect 11296 35816 11302 35828
rect 11422 35816 11428 35828
rect 11296 35788 11428 35816
rect 11296 35776 11302 35788
rect 11422 35776 11428 35788
rect 11480 35776 11486 35828
rect 12158 35816 12164 35828
rect 11532 35788 12164 35816
rect 11532 35748 11560 35788
rect 12158 35776 12164 35788
rect 12216 35776 12222 35828
rect 10796 35720 11192 35748
rect 11256 35720 11560 35748
rect 8938 35640 8944 35692
rect 8996 35680 9002 35692
rect 9493 35683 9551 35689
rect 9493 35680 9505 35683
rect 8996 35652 9505 35680
rect 8996 35640 9002 35652
rect 9493 35649 9505 35652
rect 9539 35649 9551 35683
rect 9493 35643 9551 35649
rect 10410 35640 10416 35692
rect 10468 35640 10474 35692
rect 10796 35689 10824 35720
rect 10781 35683 10839 35689
rect 10781 35649 10793 35683
rect 10827 35649 10839 35683
rect 10781 35643 10839 35649
rect 11057 35683 11115 35689
rect 11057 35649 11069 35683
rect 11103 35680 11115 35683
rect 11256 35680 11284 35720
rect 11698 35708 11704 35760
rect 11756 35748 11762 35760
rect 11756 35720 12296 35748
rect 11756 35708 11762 35720
rect 11103 35652 11284 35680
rect 11333 35683 11391 35689
rect 11103 35649 11115 35652
rect 11057 35643 11115 35649
rect 11333 35649 11345 35683
rect 11379 35680 11391 35683
rect 11422 35680 11428 35692
rect 11379 35652 11428 35680
rect 11379 35649 11391 35652
rect 11333 35643 11391 35649
rect 11422 35640 11428 35652
rect 11480 35640 11486 35692
rect 11790 35640 11796 35692
rect 11848 35640 11854 35692
rect 12066 35640 12072 35692
rect 12124 35640 12130 35692
rect 12161 35683 12219 35689
rect 12161 35649 12173 35683
rect 12207 35649 12219 35683
rect 12268 35680 12296 35720
rect 12342 35708 12348 35760
rect 12400 35748 12406 35760
rect 13173 35751 13231 35757
rect 13173 35748 13185 35751
rect 12400 35720 13185 35748
rect 12400 35708 12406 35720
rect 13173 35717 13185 35720
rect 13219 35717 13231 35751
rect 13173 35711 13231 35717
rect 12434 35680 12440 35692
rect 12268 35652 12440 35680
rect 12161 35643 12219 35649
rect 10962 35572 10968 35624
rect 11020 35612 11026 35624
rect 12176 35612 12204 35643
rect 12434 35640 12440 35652
rect 12492 35640 12498 35692
rect 12526 35640 12532 35692
rect 12584 35680 12590 35692
rect 12621 35683 12679 35689
rect 12621 35680 12633 35683
rect 12584 35652 12633 35680
rect 12584 35640 12590 35652
rect 12621 35649 12633 35652
rect 12667 35649 12679 35683
rect 12621 35643 12679 35649
rect 13725 35683 13783 35689
rect 13725 35649 13737 35683
rect 13771 35680 13783 35683
rect 13814 35680 13820 35692
rect 13771 35652 13820 35680
rect 13771 35649 13783 35652
rect 13725 35643 13783 35649
rect 13814 35640 13820 35652
rect 13872 35640 13878 35692
rect 14090 35640 14096 35692
rect 14148 35640 14154 35692
rect 11020 35584 12204 35612
rect 11020 35572 11026 35584
rect 12250 35572 12256 35624
rect 12308 35572 12314 35624
rect 9309 35547 9367 35553
rect 9309 35513 9321 35547
rect 9355 35544 9367 35547
rect 11514 35544 11520 35556
rect 9355 35516 11520 35544
rect 9355 35513 9367 35516
rect 9309 35507 9367 35513
rect 11514 35504 11520 35516
rect 11572 35504 11578 35556
rect 11609 35547 11667 35553
rect 11609 35513 11621 35547
rect 11655 35544 11667 35547
rect 12268 35544 12296 35572
rect 11655 35516 12296 35544
rect 12345 35547 12403 35553
rect 11655 35513 11667 35516
rect 11609 35507 11667 35513
rect 12345 35513 12357 35547
rect 12391 35544 12403 35547
rect 13998 35544 14004 35556
rect 12391 35516 14004 35544
rect 12391 35513 12403 35516
rect 12345 35507 12403 35513
rect 13998 35504 14004 35516
rect 14056 35504 14062 35556
rect 10870 35436 10876 35488
rect 10928 35476 10934 35488
rect 11885 35479 11943 35485
rect 11885 35476 11897 35479
rect 10928 35448 11897 35476
rect 10928 35436 10934 35448
rect 11885 35445 11897 35448
rect 11931 35445 11943 35479
rect 11885 35439 11943 35445
rect 12897 35479 12955 35485
rect 12897 35445 12909 35479
rect 12943 35476 12955 35479
rect 13262 35476 13268 35488
rect 12943 35448 13268 35476
rect 12943 35445 12955 35448
rect 12897 35439 12955 35445
rect 13262 35436 13268 35448
rect 13320 35436 13326 35488
rect 13446 35436 13452 35488
rect 13504 35436 13510 35488
rect 1104 35386 14536 35408
rect 1104 35334 2629 35386
rect 2681 35334 2693 35386
rect 2745 35334 2757 35386
rect 2809 35334 2821 35386
rect 2873 35334 2885 35386
rect 2937 35334 5987 35386
rect 6039 35334 6051 35386
rect 6103 35334 6115 35386
rect 6167 35334 6179 35386
rect 6231 35334 6243 35386
rect 6295 35334 9345 35386
rect 9397 35334 9409 35386
rect 9461 35334 9473 35386
rect 9525 35334 9537 35386
rect 9589 35334 9601 35386
rect 9653 35334 12703 35386
rect 12755 35334 12767 35386
rect 12819 35334 12831 35386
rect 12883 35334 12895 35386
rect 12947 35334 12959 35386
rect 13011 35334 14536 35386
rect 1104 35312 14536 35334
rect 5534 35232 5540 35284
rect 5592 35232 5598 35284
rect 8938 35232 8944 35284
rect 8996 35232 9002 35284
rect 9493 35275 9551 35281
rect 9493 35241 9505 35275
rect 9539 35272 9551 35275
rect 10410 35272 10416 35284
rect 9539 35244 10416 35272
rect 9539 35241 9551 35244
rect 9493 35235 9551 35241
rect 10410 35232 10416 35244
rect 10468 35232 10474 35284
rect 10781 35275 10839 35281
rect 10781 35241 10793 35275
rect 10827 35272 10839 35275
rect 10962 35272 10968 35284
rect 10827 35244 10968 35272
rect 10827 35241 10839 35244
rect 10781 35235 10839 35241
rect 10962 35232 10968 35244
rect 11020 35232 11026 35284
rect 11057 35275 11115 35281
rect 11057 35241 11069 35275
rect 11103 35272 11115 35275
rect 13354 35272 13360 35284
rect 11103 35244 13360 35272
rect 11103 35241 11115 35244
rect 11057 35235 11115 35241
rect 13354 35232 13360 35244
rect 13412 35232 13418 35284
rect 9858 35164 9864 35216
rect 9916 35204 9922 35216
rect 11238 35204 11244 35216
rect 9916 35176 11244 35204
rect 9916 35164 9922 35176
rect 11238 35164 11244 35176
rect 11296 35164 11302 35216
rect 750 35028 756 35080
rect 808 35068 814 35080
rect 1397 35071 1455 35077
rect 1397 35068 1409 35071
rect 808 35040 1409 35068
rect 808 35028 814 35040
rect 1397 35037 1409 35040
rect 1443 35037 1455 35071
rect 1397 35031 1455 35037
rect 5718 35028 5724 35080
rect 5776 35028 5782 35080
rect 8110 35028 8116 35080
rect 8168 35068 8174 35080
rect 9125 35071 9183 35077
rect 9125 35068 9137 35071
rect 8168 35040 9137 35068
rect 8168 35028 8174 35040
rect 9125 35037 9137 35040
rect 9171 35037 9183 35071
rect 9125 35031 9183 35037
rect 9674 35028 9680 35080
rect 9732 35028 9738 35080
rect 10594 35028 10600 35080
rect 10652 35068 10658 35080
rect 10965 35071 11023 35077
rect 10965 35068 10977 35071
rect 10652 35040 10977 35068
rect 10652 35028 10658 35040
rect 10965 35037 10977 35040
rect 11011 35037 11023 35071
rect 10965 35031 11023 35037
rect 11241 35071 11299 35077
rect 11241 35037 11253 35071
rect 11287 35037 11299 35071
rect 11241 35031 11299 35037
rect 10410 34960 10416 35012
rect 10468 35000 10474 35012
rect 11256 35000 11284 35031
rect 11514 35028 11520 35080
rect 11572 35028 11578 35080
rect 11791 35061 11849 35067
rect 11791 35058 11803 35061
rect 10468 34972 11284 35000
rect 11790 35027 11803 35058
rect 11837 35027 11849 35061
rect 13078 35028 13084 35080
rect 13136 35028 13142 35080
rect 11790 35021 11849 35027
rect 10468 34960 10474 34972
rect 1581 34935 1639 34941
rect 1581 34901 1593 34935
rect 1627 34932 1639 34935
rect 6454 34932 6460 34944
rect 1627 34904 6460 34932
rect 1627 34901 1639 34904
rect 1581 34895 1639 34901
rect 6454 34892 6460 34904
rect 6512 34892 6518 34944
rect 11790 34932 11818 35021
rect 13170 34960 13176 35012
rect 13228 35000 13234 35012
rect 13357 35003 13415 35009
rect 13357 35000 13369 35003
rect 13228 34972 13369 35000
rect 13228 34960 13234 34972
rect 13357 34969 13369 34972
rect 13403 34969 13415 35003
rect 13357 34963 13415 34969
rect 11882 34932 11888 34944
rect 11790 34904 11888 34932
rect 11882 34892 11888 34904
rect 11940 34892 11946 34944
rect 12434 34892 12440 34944
rect 12492 34932 12498 34944
rect 12529 34935 12587 34941
rect 12529 34932 12541 34935
rect 12492 34904 12541 34932
rect 12492 34892 12498 34904
rect 12529 34901 12541 34904
rect 12575 34901 12587 34935
rect 12529 34895 12587 34901
rect 12618 34892 12624 34944
rect 12676 34932 12682 34944
rect 12897 34935 12955 34941
rect 12897 34932 12909 34935
rect 12676 34904 12909 34932
rect 12676 34892 12682 34904
rect 12897 34901 12909 34904
rect 12943 34901 12955 34935
rect 12897 34895 12955 34901
rect 13630 34892 13636 34944
rect 13688 34892 13694 34944
rect 1104 34842 14696 34864
rect 1104 34790 4308 34842
rect 4360 34790 4372 34842
rect 4424 34790 4436 34842
rect 4488 34790 4500 34842
rect 4552 34790 4564 34842
rect 4616 34790 7666 34842
rect 7718 34790 7730 34842
rect 7782 34790 7794 34842
rect 7846 34790 7858 34842
rect 7910 34790 7922 34842
rect 7974 34790 11024 34842
rect 11076 34790 11088 34842
rect 11140 34790 11152 34842
rect 11204 34790 11216 34842
rect 11268 34790 11280 34842
rect 11332 34790 14382 34842
rect 14434 34790 14446 34842
rect 14498 34790 14510 34842
rect 14562 34790 14574 34842
rect 14626 34790 14638 34842
rect 14690 34790 14696 34842
rect 1104 34768 14696 34790
rect 1581 34731 1639 34737
rect 1581 34697 1593 34731
rect 1627 34697 1639 34731
rect 1581 34691 1639 34697
rect 5537 34731 5595 34737
rect 5537 34697 5549 34731
rect 5583 34728 5595 34731
rect 5718 34728 5724 34740
rect 5583 34700 5724 34728
rect 5583 34697 5595 34700
rect 5537 34691 5595 34697
rect 1596 34660 1624 34691
rect 5718 34688 5724 34700
rect 5776 34688 5782 34740
rect 10594 34688 10600 34740
rect 10652 34688 10658 34740
rect 12713 34731 12771 34737
rect 12713 34697 12725 34731
rect 12759 34728 12771 34731
rect 12986 34728 12992 34740
rect 12759 34700 12992 34728
rect 12759 34697 12771 34700
rect 12713 34691 12771 34697
rect 12986 34688 12992 34700
rect 13044 34688 13050 34740
rect 13814 34688 13820 34740
rect 13872 34688 13878 34740
rect 5350 34660 5356 34672
rect 1596 34632 5356 34660
rect 5350 34620 5356 34632
rect 5408 34660 5414 34672
rect 9766 34660 9772 34672
rect 5408 34632 9772 34660
rect 5408 34620 5414 34632
rect 9766 34620 9772 34632
rect 9824 34620 9830 34672
rect 11238 34620 11244 34672
rect 11296 34660 11302 34672
rect 13832 34660 13860 34688
rect 11296 34632 13860 34660
rect 11296 34620 11302 34632
rect 1394 34552 1400 34604
rect 1452 34552 1458 34604
rect 5718 34552 5724 34604
rect 5776 34552 5782 34604
rect 8202 34552 8208 34604
rect 8260 34592 8266 34604
rect 10781 34595 10839 34601
rect 10781 34592 10793 34595
rect 8260 34564 10793 34592
rect 8260 34552 8266 34564
rect 10781 34561 10793 34564
rect 10827 34561 10839 34595
rect 10781 34555 10839 34561
rect 10962 34552 10968 34604
rect 11020 34552 11026 34604
rect 11330 34552 11336 34604
rect 11388 34552 11394 34604
rect 11422 34552 11428 34604
rect 11480 34592 11486 34604
rect 11943 34595 12001 34601
rect 11943 34592 11955 34595
rect 11480 34564 11955 34592
rect 11480 34552 11486 34564
rect 11943 34561 11955 34564
rect 11989 34561 12001 34595
rect 11943 34555 12001 34561
rect 13265 34595 13323 34601
rect 13265 34561 13277 34595
rect 13311 34592 13323 34595
rect 13311 34564 13584 34592
rect 13311 34561 13323 34564
rect 13265 34555 13323 34561
rect 11440 34524 11468 34552
rect 13556 34536 13584 34564
rect 13814 34552 13820 34604
rect 13872 34552 13878 34604
rect 14185 34595 14243 34601
rect 14185 34561 14197 34595
rect 14231 34592 14243 34595
rect 14918 34592 14924 34604
rect 14231 34564 14924 34592
rect 14231 34561 14243 34564
rect 14185 34555 14243 34561
rect 14918 34552 14924 34564
rect 14976 34552 14982 34604
rect 9784 34496 11468 34524
rect 9784 34400 9812 34496
rect 11514 34484 11520 34536
rect 11572 34524 11578 34536
rect 11701 34527 11759 34533
rect 11701 34524 11713 34527
rect 11572 34496 11713 34524
rect 11572 34484 11578 34496
rect 11701 34493 11713 34496
rect 11747 34493 11759 34527
rect 11701 34487 11759 34493
rect 13538 34484 13544 34536
rect 13596 34484 13602 34536
rect 9766 34348 9772 34400
rect 9824 34348 9830 34400
rect 13354 34348 13360 34400
rect 13412 34348 13418 34400
rect 1104 34298 14536 34320
rect 1104 34246 2629 34298
rect 2681 34246 2693 34298
rect 2745 34246 2757 34298
rect 2809 34246 2821 34298
rect 2873 34246 2885 34298
rect 2937 34246 5987 34298
rect 6039 34246 6051 34298
rect 6103 34246 6115 34298
rect 6167 34246 6179 34298
rect 6231 34246 6243 34298
rect 6295 34246 9345 34298
rect 9397 34246 9409 34298
rect 9461 34246 9473 34298
rect 9525 34246 9537 34298
rect 9589 34246 9601 34298
rect 9653 34246 12703 34298
rect 12755 34246 12767 34298
rect 12819 34246 12831 34298
rect 12883 34246 12895 34298
rect 12947 34246 12959 34298
rect 13011 34246 14536 34298
rect 1104 34224 14536 34246
rect 4982 34144 4988 34196
rect 5040 34184 5046 34196
rect 9858 34184 9864 34196
rect 5040 34156 9864 34184
rect 5040 34144 5046 34156
rect 9858 34144 9864 34156
rect 9916 34144 9922 34196
rect 10410 34144 10416 34196
rect 10468 34144 10474 34196
rect 10962 34144 10968 34196
rect 11020 34144 11026 34196
rect 11238 34144 11244 34196
rect 11296 34144 11302 34196
rect 11517 34187 11575 34193
rect 11517 34153 11529 34187
rect 11563 34184 11575 34187
rect 12342 34184 12348 34196
rect 11563 34156 12348 34184
rect 11563 34153 11575 34156
rect 11517 34147 11575 34153
rect 12342 34144 12348 34156
rect 12400 34144 12406 34196
rect 10689 34119 10747 34125
rect 10689 34085 10701 34119
rect 10735 34116 10747 34119
rect 12526 34116 12532 34128
rect 10735 34088 12532 34116
rect 10735 34085 10747 34088
rect 10689 34079 10747 34085
rect 12526 34076 12532 34088
rect 12584 34076 12590 34128
rect 9950 34008 9956 34060
rect 10008 34048 10014 34060
rect 12618 34048 12624 34060
rect 10008 34020 10640 34048
rect 10008 34008 10014 34020
rect 9858 33940 9864 33992
rect 9916 33980 9922 33992
rect 10045 33983 10103 33989
rect 10045 33980 10057 33983
rect 9916 33952 10057 33980
rect 9916 33940 9922 33952
rect 10045 33949 10057 33952
rect 10091 33949 10103 33983
rect 10045 33943 10103 33949
rect 10134 33940 10140 33992
rect 10192 33980 10198 33992
rect 10612 33989 10640 34020
rect 11440 34020 12624 34048
rect 10321 33983 10379 33989
rect 10321 33980 10333 33983
rect 10192 33952 10333 33980
rect 10192 33940 10198 33952
rect 10321 33949 10333 33952
rect 10367 33949 10379 33983
rect 10321 33943 10379 33949
rect 10597 33983 10655 33989
rect 10597 33949 10609 33983
rect 10643 33949 10655 33983
rect 10597 33943 10655 33949
rect 10870 33940 10876 33992
rect 10928 33976 10934 33992
rect 11440 33989 11468 34020
rect 12618 34008 12624 34020
rect 12676 34008 12682 34060
rect 13265 34051 13323 34057
rect 13265 34017 13277 34051
rect 13311 34048 13323 34051
rect 13906 34048 13912 34060
rect 13311 34020 13912 34048
rect 13311 34017 13323 34020
rect 13265 34011 13323 34017
rect 13906 34008 13912 34020
rect 13964 34008 13970 34060
rect 11149 33983 11207 33989
rect 10928 33948 10969 33976
rect 11149 33949 11161 33983
rect 11195 33949 11207 33983
rect 10928 33940 10934 33948
rect 11149 33943 11207 33949
rect 11425 33983 11483 33989
rect 11425 33949 11437 33983
rect 11471 33949 11483 33983
rect 11425 33943 11483 33949
rect 11701 33983 11759 33989
rect 11701 33949 11713 33983
rect 11747 33949 11759 33983
rect 11701 33943 11759 33949
rect 10873 33939 10931 33940
rect 9858 33804 9864 33856
rect 9916 33804 9922 33856
rect 10137 33847 10195 33853
rect 10137 33813 10149 33847
rect 10183 33844 10195 33847
rect 11164 33844 11192 33943
rect 11716 33912 11744 33943
rect 11440 33884 11744 33912
rect 11440 33856 11468 33884
rect 11790 33872 11796 33924
rect 11848 33912 11854 33924
rect 11885 33915 11943 33921
rect 11885 33912 11897 33915
rect 11848 33884 11897 33912
rect 11848 33872 11854 33884
rect 11885 33881 11897 33884
rect 11931 33881 11943 33915
rect 11885 33875 11943 33881
rect 12250 33872 12256 33924
rect 12308 33872 12314 33924
rect 12437 33915 12495 33921
rect 12437 33881 12449 33915
rect 12483 33881 12495 33915
rect 12437 33875 12495 33881
rect 12989 33915 13047 33921
rect 12989 33881 13001 33915
rect 13035 33912 13047 33915
rect 13262 33912 13268 33924
rect 13035 33884 13268 33912
rect 13035 33881 13047 33884
rect 12989 33875 13047 33881
rect 10183 33816 11192 33844
rect 10183 33813 10195 33816
rect 10137 33807 10195 33813
rect 11422 33804 11428 33856
rect 11480 33804 11486 33856
rect 11606 33804 11612 33856
rect 11664 33844 11670 33856
rect 12452 33844 12480 33875
rect 13262 33872 13268 33884
rect 13320 33872 13326 33924
rect 13538 33872 13544 33924
rect 13596 33872 13602 33924
rect 11664 33816 12480 33844
rect 11664 33804 11670 33816
rect 12526 33804 12532 33856
rect 12584 33844 12590 33856
rect 12713 33847 12771 33853
rect 12713 33844 12725 33847
rect 12584 33816 12725 33844
rect 12584 33804 12590 33816
rect 12713 33813 12725 33816
rect 12759 33813 12771 33847
rect 12713 33807 12771 33813
rect 13722 33804 13728 33856
rect 13780 33844 13786 33856
rect 13817 33847 13875 33853
rect 13817 33844 13829 33847
rect 13780 33816 13829 33844
rect 13780 33804 13786 33816
rect 13817 33813 13829 33816
rect 13863 33813 13875 33847
rect 13817 33807 13875 33813
rect 1104 33754 14696 33776
rect 1104 33702 4308 33754
rect 4360 33702 4372 33754
rect 4424 33702 4436 33754
rect 4488 33702 4500 33754
rect 4552 33702 4564 33754
rect 4616 33702 7666 33754
rect 7718 33702 7730 33754
rect 7782 33702 7794 33754
rect 7846 33702 7858 33754
rect 7910 33702 7922 33754
rect 7974 33702 11024 33754
rect 11076 33702 11088 33754
rect 11140 33702 11152 33754
rect 11204 33702 11216 33754
rect 11268 33702 11280 33754
rect 11332 33702 14382 33754
rect 14434 33702 14446 33754
rect 14498 33702 14510 33754
rect 14562 33702 14574 33754
rect 14626 33702 14638 33754
rect 14690 33702 14696 33754
rect 1104 33680 14696 33702
rect 9858 33600 9864 33652
rect 9916 33600 9922 33652
rect 10413 33643 10471 33649
rect 10413 33609 10425 33643
rect 10459 33640 10471 33643
rect 10459 33612 12434 33640
rect 10459 33609 10471 33612
rect 10413 33603 10471 33609
rect 750 33464 756 33516
rect 808 33504 814 33516
rect 1397 33507 1455 33513
rect 1397 33504 1409 33507
rect 808 33476 1409 33504
rect 808 33464 814 33476
rect 1397 33473 1409 33476
rect 1443 33473 1455 33507
rect 9876 33504 9904 33600
rect 11606 33572 11612 33584
rect 11256 33544 11612 33572
rect 10597 33507 10655 33513
rect 10597 33504 10609 33507
rect 9876 33476 10609 33504
rect 1397 33467 1455 33473
rect 10597 33473 10609 33476
rect 10643 33473 10655 33507
rect 10597 33467 10655 33473
rect 10686 33464 10692 33516
rect 10744 33504 10750 33516
rect 10873 33507 10931 33513
rect 10873 33504 10885 33507
rect 10744 33476 10885 33504
rect 10744 33464 10750 33476
rect 10873 33473 10885 33476
rect 10919 33473 10931 33507
rect 10873 33467 10931 33473
rect 5534 33396 5540 33448
rect 5592 33436 5598 33448
rect 9674 33436 9680 33448
rect 5592 33408 9680 33436
rect 5592 33396 5598 33408
rect 9674 33396 9680 33408
rect 9732 33396 9738 33448
rect 11149 33371 11207 33377
rect 11149 33337 11161 33371
rect 11195 33368 11207 33371
rect 11256 33368 11284 33544
rect 11606 33532 11612 33544
rect 11664 33532 11670 33584
rect 12406 33572 12434 33612
rect 13170 33600 13176 33652
rect 13228 33600 13234 33652
rect 13722 33600 13728 33652
rect 13780 33600 13786 33652
rect 13188 33572 13216 33600
rect 13740 33572 13768 33600
rect 12406 33544 13216 33572
rect 13648 33544 13768 33572
rect 11791 33517 11849 33523
rect 11330 33464 11336 33516
rect 11388 33464 11394 33516
rect 11422 33464 11428 33516
rect 11480 33464 11486 33516
rect 11791 33483 11803 33517
rect 11837 33514 11849 33517
rect 11837 33504 11928 33514
rect 12158 33504 12164 33516
rect 11837 33486 12164 33504
rect 11837 33483 11849 33486
rect 11791 33477 11849 33483
rect 11900 33476 12164 33486
rect 12158 33464 12164 33476
rect 12216 33464 12222 33516
rect 13170 33464 13176 33516
rect 13228 33464 13234 33516
rect 11195 33340 11284 33368
rect 11195 33337 11207 33340
rect 11149 33331 11207 33337
rect 1581 33303 1639 33309
rect 1581 33269 1593 33303
rect 1627 33300 1639 33303
rect 4982 33300 4988 33312
rect 1627 33272 4988 33300
rect 1627 33269 1639 33272
rect 1581 33263 1639 33269
rect 4982 33260 4988 33272
rect 5040 33260 5046 33312
rect 10689 33303 10747 33309
rect 10689 33269 10701 33303
rect 10735 33300 10747 33303
rect 11440 33300 11468 33464
rect 13648 33448 13676 33544
rect 13722 33464 13728 33516
rect 13780 33464 13786 33516
rect 11514 33396 11520 33448
rect 11572 33396 11578 33448
rect 13630 33396 13636 33448
rect 13688 33396 13694 33448
rect 13538 33368 13544 33380
rect 12406 33340 13544 33368
rect 10735 33272 11468 33300
rect 10735 33269 10747 33272
rect 10689 33263 10747 33269
rect 11974 33260 11980 33312
rect 12032 33300 12038 33312
rect 12406 33300 12434 33340
rect 13538 33328 13544 33340
rect 13596 33328 13602 33380
rect 14182 33368 14188 33380
rect 13924 33340 14188 33368
rect 12032 33272 12434 33300
rect 12032 33260 12038 33272
rect 12526 33260 12532 33312
rect 12584 33260 12590 33312
rect 13449 33303 13507 33309
rect 13449 33269 13461 33303
rect 13495 33300 13507 33303
rect 13924 33300 13952 33340
rect 14182 33328 14188 33340
rect 14240 33328 14246 33380
rect 13495 33272 13952 33300
rect 14001 33303 14059 33309
rect 13495 33269 13507 33272
rect 13449 33263 13507 33269
rect 14001 33269 14013 33303
rect 14047 33300 14059 33303
rect 15010 33300 15016 33312
rect 14047 33272 15016 33300
rect 14047 33269 14059 33272
rect 14001 33263 14059 33269
rect 15010 33260 15016 33272
rect 15068 33260 15074 33312
rect 1104 33210 14536 33232
rect 1104 33158 2629 33210
rect 2681 33158 2693 33210
rect 2745 33158 2757 33210
rect 2809 33158 2821 33210
rect 2873 33158 2885 33210
rect 2937 33158 5987 33210
rect 6039 33158 6051 33210
rect 6103 33158 6115 33210
rect 6167 33158 6179 33210
rect 6231 33158 6243 33210
rect 6295 33158 9345 33210
rect 9397 33158 9409 33210
rect 9461 33158 9473 33210
rect 9525 33158 9537 33210
rect 9589 33158 9601 33210
rect 9653 33158 12703 33210
rect 12755 33158 12767 33210
rect 12819 33158 12831 33210
rect 12883 33158 12895 33210
rect 12947 33158 12959 33210
rect 13011 33158 14536 33210
rect 1104 33136 14536 33158
rect 10413 33099 10471 33105
rect 10413 33065 10425 33099
rect 10459 33096 10471 33099
rect 13538 33096 13544 33108
rect 10459 33068 13544 33096
rect 10459 33065 10471 33068
rect 10413 33059 10471 33065
rect 13538 33056 13544 33068
rect 13596 33056 13602 33108
rect 8754 32988 8760 33040
rect 8812 33028 8818 33040
rect 11146 33028 11152 33040
rect 8812 33000 11152 33028
rect 8812 32988 8818 33000
rect 11146 32988 11152 33000
rect 11204 32988 11210 33040
rect 12434 32988 12440 33040
rect 12492 33028 12498 33040
rect 12894 33028 12900 33040
rect 12492 33000 12900 33028
rect 12492 32988 12498 33000
rect 12894 32988 12900 33000
rect 12952 32988 12958 33040
rect 9416 32932 10916 32960
rect 9416 32904 9444 32932
rect 750 32852 756 32904
rect 808 32892 814 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 808 32864 1409 32892
rect 808 32852 814 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 9398 32852 9404 32904
rect 9456 32852 9462 32904
rect 10318 32852 10324 32904
rect 10376 32852 10382 32904
rect 10888 32901 10916 32932
rect 11514 32920 11520 32972
rect 11572 32920 11578 32972
rect 13265 32963 13323 32969
rect 13265 32929 13277 32963
rect 13311 32960 13323 32963
rect 13538 32960 13544 32972
rect 13311 32932 13544 32960
rect 13311 32929 13323 32932
rect 13265 32923 13323 32929
rect 13538 32920 13544 32932
rect 13596 32920 13602 32972
rect 10597 32895 10655 32901
rect 10597 32861 10609 32895
rect 10643 32861 10655 32895
rect 10597 32855 10655 32861
rect 10873 32895 10931 32901
rect 10873 32861 10885 32895
rect 10919 32861 10931 32895
rect 10873 32855 10931 32861
rect 6914 32784 6920 32836
rect 6972 32824 6978 32836
rect 10502 32824 10508 32836
rect 6972 32796 10508 32824
rect 6972 32784 6978 32796
rect 10502 32784 10508 32796
rect 10560 32784 10566 32836
rect 1578 32716 1584 32768
rect 1636 32756 1642 32768
rect 1854 32756 1860 32768
rect 1636 32728 1860 32756
rect 1636 32716 1642 32728
rect 1854 32716 1860 32728
rect 1912 32716 1918 32768
rect 10134 32716 10140 32768
rect 10192 32716 10198 32768
rect 10612 32756 10640 32855
rect 10962 32852 10968 32904
rect 11020 32892 11026 32904
rect 11759 32895 11817 32901
rect 11759 32892 11771 32895
rect 11020 32864 11771 32892
rect 11020 32852 11026 32864
rect 11759 32861 11771 32864
rect 11805 32861 11817 32895
rect 11759 32855 11817 32861
rect 10778 32784 10784 32836
rect 10836 32824 10842 32836
rect 11057 32827 11115 32833
rect 11057 32824 11069 32827
rect 10836 32796 11069 32824
rect 10836 32784 10842 32796
rect 11057 32793 11069 32796
rect 11103 32793 11115 32827
rect 11057 32787 11115 32793
rect 11146 32784 11152 32836
rect 11204 32824 11210 32836
rect 12989 32827 13047 32833
rect 11204 32796 12940 32824
rect 11204 32784 11210 32796
rect 10689 32759 10747 32765
rect 10689 32756 10701 32759
rect 10612 32728 10701 32756
rect 10689 32725 10701 32728
rect 10735 32725 10747 32759
rect 10689 32719 10747 32725
rect 11238 32716 11244 32768
rect 11296 32756 11302 32768
rect 11333 32759 11391 32765
rect 11333 32756 11345 32759
rect 11296 32728 11345 32756
rect 11296 32716 11302 32728
rect 11333 32725 11345 32728
rect 11379 32725 11391 32759
rect 11333 32719 11391 32725
rect 12529 32759 12587 32765
rect 12529 32725 12541 32759
rect 12575 32756 12587 32759
rect 12802 32756 12808 32768
rect 12575 32728 12808 32756
rect 12575 32725 12587 32728
rect 12529 32719 12587 32725
rect 12802 32716 12808 32728
rect 12860 32716 12866 32768
rect 12912 32756 12940 32796
rect 12989 32793 13001 32827
rect 13035 32824 13047 32827
rect 13354 32824 13360 32836
rect 13035 32796 13360 32824
rect 13035 32793 13047 32796
rect 12989 32787 13047 32793
rect 13354 32784 13360 32796
rect 13412 32784 13418 32836
rect 13541 32827 13599 32833
rect 13541 32793 13553 32827
rect 13587 32793 13599 32827
rect 13541 32787 13599 32793
rect 13909 32827 13967 32833
rect 13909 32793 13921 32827
rect 13955 32824 13967 32827
rect 14274 32824 14280 32836
rect 13955 32796 14280 32824
rect 13955 32793 13967 32796
rect 13909 32787 13967 32793
rect 13556 32756 13584 32787
rect 14274 32784 14280 32796
rect 14332 32784 14338 32836
rect 12912 32728 13584 32756
rect 1104 32666 14696 32688
rect 1104 32614 4308 32666
rect 4360 32614 4372 32666
rect 4424 32614 4436 32666
rect 4488 32614 4500 32666
rect 4552 32614 4564 32666
rect 4616 32614 7666 32666
rect 7718 32614 7730 32666
rect 7782 32614 7794 32666
rect 7846 32614 7858 32666
rect 7910 32614 7922 32666
rect 7974 32614 11024 32666
rect 11076 32614 11088 32666
rect 11140 32614 11152 32666
rect 11204 32614 11216 32666
rect 11268 32614 11280 32666
rect 11332 32614 14382 32666
rect 14434 32614 14446 32666
rect 14498 32614 14510 32666
rect 14562 32614 14574 32666
rect 14626 32614 14638 32666
rect 14690 32614 14696 32666
rect 1104 32592 14696 32614
rect 10134 32512 10140 32564
rect 10192 32512 10198 32564
rect 10505 32555 10563 32561
rect 10505 32521 10517 32555
rect 10551 32552 10563 32555
rect 10551 32524 13124 32552
rect 10551 32521 10563 32524
rect 10505 32515 10563 32521
rect 10152 32484 10180 32512
rect 12989 32487 13047 32493
rect 12989 32484 13001 32487
rect 10152 32456 13001 32484
rect 12989 32453 13001 32456
rect 13035 32453 13047 32487
rect 13096 32484 13124 32524
rect 13170 32512 13176 32564
rect 13228 32552 13234 32564
rect 13449 32555 13507 32561
rect 13449 32552 13461 32555
rect 13228 32524 13461 32552
rect 13228 32512 13234 32524
rect 13449 32521 13461 32524
rect 13495 32521 13507 32555
rect 13449 32515 13507 32521
rect 13262 32484 13268 32496
rect 13096 32456 13268 32484
rect 12989 32447 13047 32453
rect 13262 32444 13268 32456
rect 13320 32444 13326 32496
rect 8570 32376 8576 32428
rect 8628 32416 8634 32428
rect 9398 32425 9404 32428
rect 9367 32419 9404 32425
rect 9367 32416 9379 32419
rect 8628 32388 9379 32416
rect 8628 32376 8634 32388
rect 9367 32385 9379 32388
rect 9367 32379 9404 32385
rect 9398 32376 9404 32379
rect 9456 32376 9462 32428
rect 10686 32376 10692 32428
rect 10744 32376 10750 32428
rect 10965 32419 11023 32425
rect 10965 32385 10977 32419
rect 11011 32385 11023 32419
rect 10965 32379 11023 32385
rect 7374 32308 7380 32360
rect 7432 32348 7438 32360
rect 9125 32351 9183 32357
rect 9125 32348 9137 32351
rect 7432 32320 9137 32348
rect 7432 32308 7438 32320
rect 9125 32317 9137 32320
rect 9171 32317 9183 32351
rect 9125 32311 9183 32317
rect 9858 32308 9864 32360
rect 9916 32348 9922 32360
rect 10980 32348 11008 32379
rect 11146 32376 11152 32428
rect 11204 32416 11210 32428
rect 11759 32419 11817 32425
rect 11759 32416 11771 32419
rect 11204 32388 11771 32416
rect 11204 32376 11210 32388
rect 11759 32385 11771 32388
rect 11805 32416 11817 32419
rect 12342 32416 12348 32428
rect 11805 32388 12348 32416
rect 11805 32385 11817 32388
rect 11759 32379 11817 32385
rect 12342 32376 12348 32388
rect 12400 32376 12406 32428
rect 13633 32419 13691 32425
rect 13633 32385 13645 32419
rect 13679 32385 13691 32419
rect 13633 32379 13691 32385
rect 13817 32419 13875 32425
rect 13817 32385 13829 32419
rect 13863 32416 13875 32419
rect 15102 32416 15108 32428
rect 13863 32388 15108 32416
rect 13863 32385 13875 32388
rect 13817 32379 13875 32385
rect 9916 32320 11008 32348
rect 9916 32308 9922 32320
rect 11054 32308 11060 32360
rect 11112 32348 11118 32360
rect 11514 32348 11520 32360
rect 11112 32320 11520 32348
rect 11112 32308 11118 32320
rect 11514 32308 11520 32320
rect 11572 32308 11578 32360
rect 13648 32348 13676 32379
rect 15102 32376 15108 32388
rect 15160 32376 15166 32428
rect 13906 32348 13912 32360
rect 13648 32320 13912 32348
rect 13906 32308 13912 32320
rect 13964 32308 13970 32360
rect 4798 32240 4804 32292
rect 4856 32240 4862 32292
rect 11146 32280 11152 32292
rect 10060 32252 11152 32280
rect 4816 32212 4844 32240
rect 10060 32212 10088 32252
rect 11146 32240 11152 32252
rect 11204 32240 11210 32292
rect 4816 32184 10088 32212
rect 10134 32172 10140 32224
rect 10192 32172 10198 32224
rect 11241 32215 11299 32221
rect 11241 32181 11253 32215
rect 11287 32212 11299 32215
rect 12250 32212 12256 32224
rect 11287 32184 12256 32212
rect 11287 32181 11299 32184
rect 11241 32175 11299 32181
rect 12250 32172 12256 32184
rect 12308 32172 12314 32224
rect 12526 32172 12532 32224
rect 12584 32172 12590 32224
rect 13262 32172 13268 32224
rect 13320 32172 13326 32224
rect 14093 32215 14151 32221
rect 14093 32181 14105 32215
rect 14139 32212 14151 32215
rect 15194 32212 15200 32224
rect 14139 32184 15200 32212
rect 14139 32181 14151 32184
rect 14093 32175 14151 32181
rect 15194 32172 15200 32184
rect 15252 32172 15258 32224
rect 1104 32122 14536 32144
rect 1104 32070 2629 32122
rect 2681 32070 2693 32122
rect 2745 32070 2757 32122
rect 2809 32070 2821 32122
rect 2873 32070 2885 32122
rect 2937 32070 5987 32122
rect 6039 32070 6051 32122
rect 6103 32070 6115 32122
rect 6167 32070 6179 32122
rect 6231 32070 6243 32122
rect 6295 32070 9345 32122
rect 9397 32070 9409 32122
rect 9461 32070 9473 32122
rect 9525 32070 9537 32122
rect 9589 32070 9601 32122
rect 9653 32070 12703 32122
rect 12755 32070 12767 32122
rect 12819 32070 12831 32122
rect 12883 32070 12895 32122
rect 12947 32070 12959 32122
rect 13011 32070 14536 32122
rect 1104 32048 14536 32070
rect 9493 32011 9551 32017
rect 9493 31977 9505 32011
rect 9539 32008 9551 32011
rect 10686 32008 10692 32020
rect 9539 31980 10692 32008
rect 9539 31977 9551 31980
rect 9493 31971 9551 31977
rect 10686 31968 10692 31980
rect 10744 31968 10750 32020
rect 10778 31968 10784 32020
rect 10836 31968 10842 32020
rect 11149 32011 11207 32017
rect 11149 31977 11161 32011
rect 11195 32008 11207 32011
rect 11974 32008 11980 32020
rect 11195 31980 11980 32008
rect 11195 31977 11207 31980
rect 11149 31971 11207 31977
rect 11974 31968 11980 31980
rect 12032 31968 12038 32020
rect 12250 31968 12256 32020
rect 12308 31968 12314 32020
rect 12621 32011 12679 32017
rect 12621 31977 12633 32011
rect 12667 32008 12679 32011
rect 15378 32008 15384 32020
rect 12667 31980 15384 32008
rect 12667 31977 12679 31980
rect 12621 31971 12679 31977
rect 15378 31968 15384 31980
rect 15436 31968 15442 32020
rect 9953 31943 10011 31949
rect 9953 31909 9965 31943
rect 9999 31909 10011 31943
rect 9953 31903 10011 31909
rect 10229 31943 10287 31949
rect 10229 31909 10241 31943
rect 10275 31940 10287 31943
rect 11238 31940 11244 31952
rect 10275 31912 11244 31940
rect 10275 31909 10287 31912
rect 10229 31903 10287 31909
rect 7374 31832 7380 31884
rect 7432 31872 7438 31884
rect 7469 31875 7527 31881
rect 7469 31872 7481 31875
rect 7432 31844 7481 31872
rect 7432 31832 7438 31844
rect 7469 31841 7481 31844
rect 7515 31841 7527 31875
rect 9968 31872 9996 31903
rect 11238 31900 11244 31912
rect 11296 31900 11302 31952
rect 11790 31900 11796 31952
rect 11848 31900 11854 31952
rect 11808 31872 11836 31900
rect 9968 31844 10732 31872
rect 7469 31835 7527 31841
rect 1394 31764 1400 31816
rect 1452 31764 1458 31816
rect 7190 31764 7196 31816
rect 7248 31804 7254 31816
rect 7743 31807 7801 31813
rect 7743 31804 7755 31807
rect 7248 31776 7755 31804
rect 7248 31764 7254 31776
rect 7743 31773 7755 31776
rect 7789 31804 7801 31807
rect 8202 31804 8208 31816
rect 7789 31776 8208 31804
rect 7789 31773 7801 31776
rect 7743 31767 7801 31773
rect 8202 31764 8208 31776
rect 8260 31764 8266 31816
rect 8846 31764 8852 31816
rect 8904 31764 8910 31816
rect 9677 31807 9735 31813
rect 9677 31804 9689 31807
rect 9600 31776 9689 31804
rect 8864 31736 8892 31764
rect 9600 31736 9628 31776
rect 9677 31773 9689 31776
rect 9723 31773 9735 31807
rect 9677 31767 9735 31773
rect 10134 31764 10140 31816
rect 10192 31764 10198 31816
rect 10413 31807 10471 31813
rect 10413 31773 10425 31807
rect 10459 31804 10471 31807
rect 10502 31804 10508 31816
rect 10459 31776 10508 31804
rect 10459 31773 10471 31776
rect 10413 31767 10471 31773
rect 10502 31764 10508 31776
rect 10560 31764 10566 31816
rect 10704 31813 10732 31844
rect 11072 31844 11836 31872
rect 10689 31807 10747 31813
rect 10689 31773 10701 31807
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 10778 31764 10784 31816
rect 10836 31804 10842 31816
rect 10965 31807 11023 31813
rect 10965 31804 10977 31807
rect 10836 31776 10977 31804
rect 10836 31764 10842 31776
rect 10965 31773 10977 31776
rect 11011 31773 11023 31807
rect 10965 31767 11023 31773
rect 10870 31736 10876 31748
rect 8864 31708 9628 31736
rect 9692 31708 10876 31736
rect 9692 31680 9720 31708
rect 10870 31696 10876 31708
rect 10928 31696 10934 31748
rect 1581 31671 1639 31677
rect 1581 31637 1593 31671
rect 1627 31668 1639 31671
rect 1762 31668 1768 31680
rect 1627 31640 1768 31668
rect 1627 31637 1639 31640
rect 1581 31631 1639 31637
rect 1762 31628 1768 31640
rect 1820 31628 1826 31680
rect 8481 31671 8539 31677
rect 8481 31637 8493 31671
rect 8527 31668 8539 31671
rect 9214 31668 9220 31680
rect 8527 31640 9220 31668
rect 8527 31637 8539 31640
rect 8481 31631 8539 31637
rect 9214 31628 9220 31640
rect 9272 31628 9278 31680
rect 9674 31628 9680 31680
rect 9732 31628 9738 31680
rect 10505 31671 10563 31677
rect 10505 31637 10517 31671
rect 10551 31668 10563 31671
rect 11072 31668 11100 31844
rect 12066 31832 12072 31884
rect 12124 31872 12130 31884
rect 12124 31844 12204 31872
rect 12124 31832 12130 31844
rect 11330 31764 11336 31816
rect 11388 31764 11394 31816
rect 11698 31764 11704 31816
rect 11756 31764 11762 31816
rect 11790 31696 11796 31748
rect 11848 31736 11854 31748
rect 12069 31739 12127 31745
rect 12069 31736 12081 31739
rect 11848 31708 12081 31736
rect 11848 31696 11854 31708
rect 12069 31705 12081 31708
rect 12115 31705 12127 31739
rect 12176 31736 12204 31844
rect 12268 31816 12296 31968
rect 13998 31872 14004 31884
rect 12912 31844 14004 31872
rect 12250 31764 12256 31816
rect 12308 31764 12314 31816
rect 12912 31745 12940 31844
rect 13998 31832 14004 31844
rect 14056 31832 14062 31884
rect 13265 31807 13323 31813
rect 13265 31773 13277 31807
rect 13311 31804 13323 31807
rect 13630 31804 13636 31816
rect 13311 31776 13636 31804
rect 13311 31773 13323 31776
rect 13265 31767 13323 31773
rect 13630 31764 13636 31776
rect 13688 31764 13694 31816
rect 15286 31804 15292 31816
rect 13740 31776 15292 31804
rect 12345 31739 12403 31745
rect 12345 31736 12357 31739
rect 12176 31708 12357 31736
rect 12069 31699 12127 31705
rect 12345 31705 12357 31708
rect 12391 31705 12403 31739
rect 12345 31699 12403 31705
rect 12897 31739 12955 31745
rect 12897 31705 12909 31739
rect 12943 31705 12955 31739
rect 12897 31699 12955 31705
rect 13449 31739 13507 31745
rect 13449 31705 13461 31739
rect 13495 31736 13507 31739
rect 13740 31736 13768 31776
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 13495 31708 13768 31736
rect 13817 31739 13875 31745
rect 13495 31705 13507 31708
rect 13449 31699 13507 31705
rect 13817 31705 13829 31739
rect 13863 31705 13875 31739
rect 13817 31699 13875 31705
rect 10551 31640 11100 31668
rect 10551 31637 10563 31640
rect 10505 31631 10563 31637
rect 12986 31628 12992 31680
rect 13044 31668 13050 31680
rect 13538 31668 13544 31680
rect 13044 31640 13544 31668
rect 13044 31628 13050 31640
rect 13538 31628 13544 31640
rect 13596 31628 13602 31680
rect 13832 31668 13860 31699
rect 15562 31696 15568 31748
rect 15620 31736 15626 31748
rect 15620 31708 15700 31736
rect 15620 31696 15626 31708
rect 14274 31668 14280 31680
rect 13832 31640 14280 31668
rect 14274 31628 14280 31640
rect 14332 31628 14338 31680
rect 1104 31578 14696 31600
rect 1104 31526 4308 31578
rect 4360 31526 4372 31578
rect 4424 31526 4436 31578
rect 4488 31526 4500 31578
rect 4552 31526 4564 31578
rect 4616 31526 7666 31578
rect 7718 31526 7730 31578
rect 7782 31526 7794 31578
rect 7846 31526 7858 31578
rect 7910 31526 7922 31578
rect 7974 31526 11024 31578
rect 11076 31526 11088 31578
rect 11140 31526 11152 31578
rect 11204 31526 11216 31578
rect 11268 31526 11280 31578
rect 11332 31526 14382 31578
rect 14434 31526 14446 31578
rect 14498 31526 14510 31578
rect 14562 31526 14574 31578
rect 14626 31526 14638 31578
rect 14690 31526 14696 31578
rect 1104 31504 14696 31526
rect 7006 31424 7012 31476
rect 7064 31464 7070 31476
rect 7064 31436 9720 31464
rect 7064 31424 7070 31436
rect 9692 31396 9720 31436
rect 9858 31424 9864 31476
rect 9916 31424 9922 31476
rect 9953 31467 10011 31473
rect 9953 31433 9965 31467
rect 9999 31464 10011 31467
rect 10778 31464 10784 31476
rect 9999 31436 10784 31464
rect 9999 31433 10011 31436
rect 9953 31427 10011 31433
rect 10778 31424 10784 31436
rect 10836 31424 10842 31476
rect 12710 31464 12716 31476
rect 10980 31436 12716 31464
rect 10980 31405 11008 31436
rect 12710 31424 12716 31436
rect 12768 31424 12774 31476
rect 13354 31424 13360 31476
rect 13412 31464 13418 31476
rect 13541 31467 13599 31473
rect 13541 31464 13553 31467
rect 13412 31436 13553 31464
rect 13412 31424 13418 31436
rect 13541 31433 13553 31436
rect 13587 31433 13599 31467
rect 13541 31427 13599 31433
rect 10965 31399 11023 31405
rect 9692 31368 10180 31396
rect 750 31288 756 31340
rect 808 31328 814 31340
rect 1397 31331 1455 31337
rect 1397 31328 1409 31331
rect 808 31300 1409 31328
rect 808 31288 814 31300
rect 1397 31297 1409 31300
rect 1443 31297 1455 31331
rect 1397 31291 1455 31297
rect 6546 31288 6552 31340
rect 6604 31328 6610 31340
rect 6604 31300 8340 31328
rect 6604 31288 6610 31300
rect 8018 31220 8024 31272
rect 8076 31220 8082 31272
rect 8205 31263 8263 31269
rect 8205 31229 8217 31263
rect 8251 31229 8263 31263
rect 8312 31260 8340 31300
rect 8938 31288 8944 31340
rect 8996 31288 9002 31340
rect 9214 31288 9220 31340
rect 9272 31288 9278 31340
rect 10152 31337 10180 31368
rect 10965 31365 10977 31399
rect 11011 31365 11023 31399
rect 10965 31359 11023 31365
rect 10137 31331 10195 31337
rect 10137 31297 10149 31331
rect 10183 31297 10195 31331
rect 10137 31291 10195 31297
rect 10686 31288 10692 31340
rect 10744 31288 10750 31340
rect 12894 31288 12900 31340
rect 12952 31288 12958 31340
rect 13725 31331 13783 31337
rect 13725 31297 13737 31331
rect 13771 31328 13783 31331
rect 14182 31328 14188 31340
rect 13771 31300 14188 31328
rect 13771 31297 13783 31300
rect 13725 31291 13783 31297
rect 14182 31288 14188 31300
rect 14240 31288 14246 31340
rect 9058 31263 9116 31269
rect 9058 31260 9070 31263
rect 8312 31232 9070 31260
rect 8205 31223 8263 31229
rect 9058 31229 9070 31232
rect 9104 31229 9116 31263
rect 9058 31223 9116 31229
rect 1581 31127 1639 31133
rect 1581 31093 1593 31127
rect 1627 31124 1639 31127
rect 3786 31124 3792 31136
rect 1627 31096 3792 31124
rect 1627 31093 1639 31096
rect 1581 31087 1639 31093
rect 3786 31084 3792 31096
rect 3844 31084 3850 31136
rect 8220 31124 8248 31223
rect 9766 31220 9772 31272
rect 9824 31260 9830 31272
rect 10410 31260 10416 31272
rect 9824 31232 10416 31260
rect 9824 31220 9830 31232
rect 10410 31220 10416 31232
rect 10468 31220 10474 31272
rect 11514 31220 11520 31272
rect 11572 31260 11578 31272
rect 11701 31263 11759 31269
rect 11701 31260 11713 31263
rect 11572 31232 11713 31260
rect 11572 31220 11578 31232
rect 11701 31229 11713 31232
rect 11747 31229 11759 31263
rect 11701 31223 11759 31229
rect 11882 31220 11888 31272
rect 11940 31220 11946 31272
rect 12342 31220 12348 31272
rect 12400 31220 12406 31272
rect 12618 31220 12624 31272
rect 12676 31220 12682 31272
rect 12738 31263 12796 31269
rect 12738 31229 12750 31263
rect 12784 31260 12796 31263
rect 12784 31232 13676 31260
rect 12784 31229 12796 31232
rect 12738 31223 12796 31229
rect 8662 31152 8668 31204
rect 8720 31152 8726 31204
rect 10505 31195 10563 31201
rect 10505 31161 10517 31195
rect 10551 31192 10563 31195
rect 11422 31192 11428 31204
rect 10551 31164 11428 31192
rect 10551 31161 10563 31164
rect 10505 31155 10563 31161
rect 11422 31152 11428 31164
rect 11480 31152 11486 31204
rect 13648 31136 13676 31232
rect 9122 31124 9128 31136
rect 8220 31096 9128 31124
rect 9122 31084 9128 31096
rect 9180 31084 9186 31136
rect 9214 31084 9220 31136
rect 9272 31124 9278 31136
rect 11146 31124 11152 31136
rect 9272 31096 11152 31124
rect 9272 31084 9278 31096
rect 11146 31084 11152 31096
rect 11204 31084 11210 31136
rect 11241 31127 11299 31133
rect 11241 31093 11253 31127
rect 11287 31124 11299 31127
rect 11606 31124 11612 31136
rect 11287 31096 11612 31124
rect 11287 31093 11299 31096
rect 11241 31087 11299 31093
rect 11606 31084 11612 31096
rect 11664 31084 11670 31136
rect 12710 31084 12716 31136
rect 12768 31124 12774 31136
rect 13262 31124 13268 31136
rect 12768 31096 13268 31124
rect 12768 31084 12774 31096
rect 13262 31084 13268 31096
rect 13320 31084 13326 31136
rect 13630 31084 13636 31136
rect 13688 31084 13694 31136
rect 14001 31127 14059 31133
rect 14001 31093 14013 31127
rect 14047 31124 14059 31127
rect 14274 31124 14280 31136
rect 14047 31096 14280 31124
rect 14047 31093 14059 31096
rect 14001 31087 14059 31093
rect 14274 31084 14280 31096
rect 14332 31084 14338 31136
rect 15562 31084 15568 31136
rect 15620 31124 15626 31136
rect 15672 31124 15700 31708
rect 15620 31096 15700 31124
rect 15620 31084 15626 31096
rect 1104 31034 14536 31056
rect 1104 30982 2629 31034
rect 2681 30982 2693 31034
rect 2745 30982 2757 31034
rect 2809 30982 2821 31034
rect 2873 30982 2885 31034
rect 2937 30982 5987 31034
rect 6039 30982 6051 31034
rect 6103 30982 6115 31034
rect 6167 30982 6179 31034
rect 6231 30982 6243 31034
rect 6295 30982 9345 31034
rect 9397 30982 9409 31034
rect 9461 30982 9473 31034
rect 9525 30982 9537 31034
rect 9589 30982 9601 31034
rect 9653 30982 12703 31034
rect 12755 30982 12767 31034
rect 12819 30982 12831 31034
rect 12883 30982 12895 31034
rect 12947 30982 12959 31034
rect 13011 30982 14536 31034
rect 1104 30960 14536 30982
rect 7374 30880 7380 30932
rect 7432 30920 7438 30932
rect 8297 30923 8355 30929
rect 7432 30892 7972 30920
rect 7432 30880 7438 30892
rect 7392 30852 7420 30880
rect 7300 30824 7420 30852
rect 7300 30793 7328 30824
rect 7285 30787 7343 30793
rect 7285 30753 7297 30787
rect 7331 30753 7343 30787
rect 7285 30747 7343 30753
rect 7527 30719 7585 30725
rect 7527 30716 7539 30719
rect 7392 30688 7539 30716
rect 7392 30592 7420 30688
rect 7527 30685 7539 30688
rect 7573 30685 7585 30719
rect 7944 30716 7972 30892
rect 8297 30889 8309 30923
rect 8343 30920 8355 30923
rect 8662 30920 8668 30932
rect 8343 30892 8668 30920
rect 8343 30889 8355 30892
rect 8297 30883 8355 30889
rect 8662 30880 8668 30892
rect 8720 30880 8726 30932
rect 9030 30880 9036 30932
rect 9088 30920 9094 30932
rect 9950 30920 9956 30932
rect 9088 30892 9956 30920
rect 9088 30880 9094 30892
rect 9950 30880 9956 30892
rect 10008 30880 10014 30932
rect 10318 30880 10324 30932
rect 10376 30920 10382 30932
rect 10376 30892 11100 30920
rect 10376 30880 10382 30892
rect 8941 30787 8999 30793
rect 8941 30784 8953 30787
rect 8864 30756 8953 30784
rect 8864 30750 8892 30756
rect 8772 30722 8892 30750
rect 8941 30753 8953 30756
rect 8987 30753 8999 30787
rect 10413 30787 10471 30793
rect 10413 30784 10425 30787
rect 8941 30747 8999 30753
rect 9692 30756 10425 30784
rect 9692 30728 9720 30756
rect 10413 30753 10425 30756
rect 10459 30753 10471 30787
rect 11072 30784 11100 30892
rect 11146 30880 11152 30932
rect 11204 30920 11210 30932
rect 11204 30892 13952 30920
rect 11204 30880 11210 30892
rect 12434 30812 12440 30864
rect 12492 30812 12498 30864
rect 13633 30855 13691 30861
rect 13633 30821 13645 30855
rect 13679 30852 13691 30855
rect 13722 30852 13728 30864
rect 13679 30824 13728 30852
rect 13679 30821 13691 30824
rect 13633 30815 13691 30821
rect 13722 30812 13728 30824
rect 13780 30812 13786 30864
rect 11072 30756 13768 30784
rect 10413 30747 10471 30753
rect 8772 30716 8800 30722
rect 9199 30719 9257 30725
rect 9199 30716 9211 30719
rect 7944 30688 8800 30716
rect 9140 30688 9211 30716
rect 7527 30679 7585 30685
rect 8846 30608 8852 30660
rect 8904 30648 8910 30660
rect 9140 30648 9168 30688
rect 9199 30685 9211 30688
rect 9245 30685 9257 30719
rect 9199 30679 9257 30685
rect 9674 30676 9680 30728
rect 9732 30676 9738 30728
rect 10594 30716 10600 30728
rect 10428 30706 10600 30716
rect 10336 30688 10600 30706
rect 10336 30678 10456 30688
rect 10336 30648 10364 30678
rect 10594 30676 10600 30688
rect 10652 30716 10658 30728
rect 10687 30719 10745 30725
rect 10687 30716 10699 30719
rect 10652 30688 10699 30716
rect 10652 30676 10658 30688
rect 10687 30685 10699 30688
rect 10733 30685 10745 30719
rect 10687 30679 10745 30685
rect 11790 30676 11796 30728
rect 11848 30676 11854 30728
rect 11882 30676 11888 30728
rect 11940 30716 11946 30728
rect 11977 30719 12035 30725
rect 11977 30716 11989 30719
rect 11940 30688 11989 30716
rect 11940 30676 11946 30688
rect 11977 30685 11989 30688
rect 12023 30685 12035 30719
rect 11977 30679 12035 30685
rect 12710 30676 12716 30728
rect 12768 30676 12774 30728
rect 12802 30676 12808 30728
rect 12860 30725 12866 30728
rect 12860 30719 12888 30725
rect 12876 30685 12888 30719
rect 12860 30679 12888 30685
rect 12860 30676 12866 30679
rect 12986 30676 12992 30728
rect 13044 30676 13050 30728
rect 8904 30620 9168 30648
rect 9324 30620 10364 30648
rect 8904 30608 8910 30620
rect 7374 30540 7380 30592
rect 7432 30580 7438 30592
rect 9030 30580 9036 30592
rect 7432 30552 9036 30580
rect 7432 30540 7438 30552
rect 9030 30540 9036 30552
rect 9088 30540 9094 30592
rect 9214 30540 9220 30592
rect 9272 30580 9278 30592
rect 9324 30580 9352 30620
rect 9272 30552 9352 30580
rect 9272 30540 9278 30552
rect 9582 30540 9588 30592
rect 9640 30580 9646 30592
rect 9953 30583 10011 30589
rect 9953 30580 9965 30583
rect 9640 30552 9965 30580
rect 9640 30540 9646 30552
rect 9953 30549 9965 30552
rect 9999 30549 10011 30583
rect 9953 30543 10011 30549
rect 11425 30583 11483 30589
rect 11425 30549 11437 30583
rect 11471 30580 11483 30583
rect 12250 30580 12256 30592
rect 11471 30552 12256 30580
rect 11471 30549 11483 30552
rect 11425 30543 11483 30549
rect 12250 30540 12256 30552
rect 12308 30540 12314 30592
rect 13740 30589 13768 30756
rect 13924 30725 13952 30892
rect 13909 30719 13967 30725
rect 13909 30685 13921 30719
rect 13955 30685 13967 30719
rect 13909 30679 13967 30685
rect 14366 30608 14372 30660
rect 14424 30648 14430 30660
rect 15470 30648 15476 30660
rect 14424 30620 15476 30648
rect 14424 30608 14430 30620
rect 15470 30608 15476 30620
rect 15528 30608 15534 30660
rect 13725 30583 13783 30589
rect 13725 30549 13737 30583
rect 13771 30549 13783 30583
rect 13725 30543 13783 30549
rect 1104 30490 14696 30512
rect 1104 30438 4308 30490
rect 4360 30438 4372 30490
rect 4424 30438 4436 30490
rect 4488 30438 4500 30490
rect 4552 30438 4564 30490
rect 4616 30438 7666 30490
rect 7718 30438 7730 30490
rect 7782 30438 7794 30490
rect 7846 30438 7858 30490
rect 7910 30438 7922 30490
rect 7974 30438 11024 30490
rect 11076 30438 11088 30490
rect 11140 30438 11152 30490
rect 11204 30438 11216 30490
rect 11268 30438 11280 30490
rect 11332 30438 14382 30490
rect 14434 30438 14446 30490
rect 14498 30438 14510 30490
rect 14562 30438 14574 30490
rect 14626 30438 14638 30490
rect 14690 30438 14696 30490
rect 1104 30416 14696 30438
rect 8202 30336 8208 30388
rect 8260 30376 8266 30388
rect 10686 30376 10692 30388
rect 8260 30348 10692 30376
rect 8260 30336 8266 30348
rect 10686 30336 10692 30348
rect 10744 30336 10750 30388
rect 12434 30336 12440 30388
rect 12492 30376 12498 30388
rect 12802 30376 12808 30388
rect 12492 30348 12808 30376
rect 12492 30336 12498 30348
rect 12802 30336 12808 30348
rect 12860 30336 12866 30388
rect 10873 30311 10931 30317
rect 10873 30277 10885 30311
rect 10919 30308 10931 30311
rect 11698 30308 11704 30320
rect 10919 30280 11704 30308
rect 10919 30277 10931 30280
rect 10873 30271 10931 30277
rect 11698 30268 11704 30280
rect 11756 30268 11762 30320
rect 13814 30268 13820 30320
rect 13872 30268 13878 30320
rect 750 30200 756 30252
rect 808 30240 814 30252
rect 1397 30243 1455 30249
rect 1397 30240 1409 30243
rect 808 30212 1409 30240
rect 808 30200 814 30212
rect 1397 30209 1409 30212
rect 1443 30209 1455 30243
rect 1397 30203 1455 30209
rect 10226 30200 10232 30252
rect 10284 30200 10290 30252
rect 13170 30200 13176 30252
rect 13228 30200 13234 30252
rect 14093 30243 14151 30249
rect 14093 30209 14105 30243
rect 14139 30209 14151 30243
rect 14093 30203 14151 30209
rect 9030 30132 9036 30184
rect 9088 30132 9094 30184
rect 9122 30132 9128 30184
rect 9180 30172 9186 30184
rect 9217 30175 9275 30181
rect 9217 30172 9229 30175
rect 9180 30144 9229 30172
rect 9180 30132 9186 30144
rect 9217 30141 9229 30144
rect 9263 30141 9275 30175
rect 9217 30135 9275 30141
rect 9582 30132 9588 30184
rect 9640 30172 9646 30184
rect 9677 30175 9735 30181
rect 9677 30172 9689 30175
rect 9640 30144 9689 30172
rect 9640 30132 9646 30144
rect 9677 30141 9689 30144
rect 9723 30141 9735 30175
rect 9953 30175 10011 30181
rect 9953 30172 9965 30175
rect 9677 30135 9735 30141
rect 9784 30144 9965 30172
rect 8662 30064 8668 30116
rect 8720 30104 8726 30116
rect 9306 30104 9312 30116
rect 8720 30076 9312 30104
rect 8720 30064 8726 30076
rect 9306 30064 9312 30076
rect 9364 30064 9370 30116
rect 1581 30039 1639 30045
rect 1581 30005 1593 30039
rect 1627 30036 1639 30039
rect 5534 30036 5540 30048
rect 1627 30008 5540 30036
rect 1627 30005 1639 30008
rect 1581 29999 1639 30005
rect 5534 29996 5540 30008
rect 5592 29996 5598 30048
rect 8478 29996 8484 30048
rect 8536 30036 8542 30048
rect 8938 30036 8944 30048
rect 8536 30008 8944 30036
rect 8536 29996 8542 30008
rect 8938 29996 8944 30008
rect 8996 30036 9002 30048
rect 9784 30036 9812 30144
rect 9953 30141 9965 30144
rect 9999 30141 10011 30175
rect 9953 30135 10011 30141
rect 10042 30132 10048 30184
rect 10100 30181 10106 30184
rect 10100 30175 10128 30181
rect 10116 30141 10128 30175
rect 10100 30135 10128 30141
rect 10100 30132 10106 30135
rect 11974 30132 11980 30184
rect 12032 30132 12038 30184
rect 12158 30132 12164 30184
rect 12216 30132 12222 30184
rect 12250 30132 12256 30184
rect 12308 30172 12314 30184
rect 12621 30175 12679 30181
rect 12621 30172 12633 30175
rect 12308 30144 12633 30172
rect 12308 30132 12314 30144
rect 12621 30141 12633 30144
rect 12667 30141 12679 30175
rect 12621 30135 12679 30141
rect 12710 30132 12716 30184
rect 12768 30172 12774 30184
rect 12897 30175 12955 30181
rect 12897 30172 12909 30175
rect 12768 30144 12909 30172
rect 12768 30132 12774 30144
rect 12897 30141 12909 30144
rect 12943 30141 12955 30175
rect 12897 30135 12955 30141
rect 12986 30132 12992 30184
rect 13044 30181 13050 30184
rect 13044 30175 13072 30181
rect 13060 30141 13072 30175
rect 13044 30135 13072 30141
rect 13044 30132 13050 30135
rect 10686 30064 10692 30116
rect 10744 30104 10750 30116
rect 10744 30076 12756 30104
rect 10744 30064 10750 30076
rect 8996 30008 9812 30036
rect 12728 30036 12756 30076
rect 13906 30064 13912 30116
rect 13964 30064 13970 30116
rect 14108 30036 14136 30203
rect 12728 30008 14136 30036
rect 8996 29996 9002 30008
rect 1104 29946 14536 29968
rect 1104 29894 2629 29946
rect 2681 29894 2693 29946
rect 2745 29894 2757 29946
rect 2809 29894 2821 29946
rect 2873 29894 2885 29946
rect 2937 29894 5987 29946
rect 6039 29894 6051 29946
rect 6103 29894 6115 29946
rect 6167 29894 6179 29946
rect 6231 29894 6243 29946
rect 6295 29894 9345 29946
rect 9397 29894 9409 29946
rect 9461 29894 9473 29946
rect 9525 29894 9537 29946
rect 9589 29894 9601 29946
rect 9653 29894 12703 29946
rect 12755 29894 12767 29946
rect 12819 29894 12831 29946
rect 12883 29894 12895 29946
rect 12947 29894 12959 29946
rect 13011 29894 14536 29946
rect 1104 29872 14536 29894
rect 2130 29792 2136 29844
rect 2188 29792 2194 29844
rect 7098 29832 7104 29844
rect 6104 29804 7104 29832
rect 6104 29705 6132 29804
rect 7098 29792 7104 29804
rect 7156 29792 7162 29844
rect 7282 29792 7288 29844
rect 7340 29832 7346 29844
rect 7340 29804 11008 29832
rect 7340 29792 7346 29804
rect 6089 29699 6147 29705
rect 6089 29696 6101 29699
rect 2746 29668 6101 29696
rect 750 29588 756 29640
rect 808 29628 814 29640
rect 1397 29631 1455 29637
rect 1397 29628 1409 29631
rect 808 29600 1409 29628
rect 808 29588 814 29600
rect 1397 29597 1409 29600
rect 1443 29597 1455 29631
rect 1397 29591 1455 29597
rect 1949 29631 2007 29637
rect 1949 29597 1961 29631
rect 1995 29628 2007 29631
rect 2746 29628 2774 29668
rect 6089 29665 6101 29668
rect 6135 29665 6147 29699
rect 8110 29696 8116 29708
rect 6089 29659 6147 29665
rect 7024 29668 8116 29696
rect 1995 29600 2774 29628
rect 1995 29597 2007 29600
rect 1949 29591 2007 29597
rect 3786 29588 3792 29640
rect 3844 29628 3850 29640
rect 7024 29628 7052 29668
rect 8110 29656 8116 29668
rect 8168 29656 8174 29708
rect 3844 29601 7052 29628
rect 3844 29600 6359 29601
rect 3844 29588 3850 29600
rect 6347 29567 6359 29600
rect 6393 29600 7052 29601
rect 6393 29570 6408 29600
rect 7282 29588 7288 29640
rect 7340 29628 7346 29640
rect 7466 29628 7472 29640
rect 7340 29600 7472 29628
rect 7340 29588 7346 29600
rect 7466 29588 7472 29600
rect 7524 29628 7530 29640
rect 7524 29600 8892 29628
rect 7524 29588 7530 29600
rect 6393 29567 6405 29570
rect 6347 29561 6405 29567
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 2038 29492 2044 29504
rect 1627 29464 2044 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 2038 29452 2044 29464
rect 2096 29492 2102 29504
rect 6822 29492 6828 29504
rect 2096 29464 6828 29492
rect 2096 29452 2102 29464
rect 6822 29452 6828 29464
rect 6880 29452 6886 29504
rect 7101 29495 7159 29501
rect 7101 29461 7113 29495
rect 7147 29492 7159 29495
rect 7466 29492 7472 29504
rect 7147 29464 7472 29492
rect 7147 29461 7159 29464
rect 7101 29455 7159 29461
rect 7466 29452 7472 29464
rect 7524 29452 7530 29504
rect 8864 29492 8892 29600
rect 9674 29588 9680 29640
rect 9732 29628 9738 29640
rect 10321 29631 10379 29637
rect 10321 29628 10333 29631
rect 9732 29600 10333 29628
rect 9732 29588 9738 29600
rect 10321 29597 10333 29600
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 10502 29588 10508 29640
rect 10560 29628 10566 29640
rect 10595 29631 10653 29637
rect 10595 29628 10607 29631
rect 10560 29600 10607 29628
rect 10560 29588 10566 29600
rect 10595 29597 10607 29600
rect 10641 29597 10653 29631
rect 10980 29628 11008 29804
rect 12066 29792 12072 29844
rect 12124 29832 12130 29844
rect 14918 29832 14924 29844
rect 12124 29804 14924 29832
rect 12124 29792 12130 29804
rect 14918 29792 14924 29804
rect 14976 29792 14982 29844
rect 11790 29656 11796 29708
rect 11848 29696 11854 29708
rect 12621 29699 12679 29705
rect 12621 29696 12633 29699
rect 11848 29668 12633 29696
rect 11848 29656 11854 29668
rect 12621 29665 12633 29668
rect 12667 29665 12679 29699
rect 12621 29659 12679 29665
rect 12863 29631 12921 29637
rect 12863 29628 12875 29631
rect 10980 29600 12875 29628
rect 10595 29591 10653 29597
rect 12863 29597 12875 29600
rect 12909 29628 12921 29631
rect 12909 29600 13216 29628
rect 12909 29597 12921 29600
rect 12863 29591 12921 29597
rect 13188 29572 13216 29600
rect 8938 29520 8944 29572
rect 8996 29560 9002 29572
rect 9861 29563 9919 29569
rect 9861 29560 9873 29563
rect 8996 29532 9873 29560
rect 8996 29520 9002 29532
rect 9861 29529 9873 29532
rect 9907 29529 9919 29563
rect 9861 29523 9919 29529
rect 10229 29563 10287 29569
rect 10229 29529 10241 29563
rect 10275 29560 10287 29563
rect 11422 29560 11428 29572
rect 10275 29532 11428 29560
rect 10275 29529 10287 29532
rect 10229 29523 10287 29529
rect 11422 29520 11428 29532
rect 11480 29520 11486 29572
rect 11698 29520 11704 29572
rect 11756 29560 11762 29572
rect 12161 29563 12219 29569
rect 12161 29560 12173 29563
rect 11756 29532 12173 29560
rect 11756 29520 11762 29532
rect 12161 29529 12173 29532
rect 12207 29529 12219 29563
rect 12161 29523 12219 29529
rect 13170 29520 13176 29572
rect 13228 29520 13234 29572
rect 9674 29492 9680 29504
rect 8864 29464 9680 29492
rect 9674 29452 9680 29464
rect 9732 29452 9738 29504
rect 9766 29452 9772 29504
rect 9824 29492 9830 29504
rect 10686 29492 10692 29504
rect 9824 29464 10692 29492
rect 9824 29452 9830 29464
rect 10686 29452 10692 29464
rect 10744 29452 10750 29504
rect 11333 29495 11391 29501
rect 11333 29461 11345 29495
rect 11379 29492 11391 29495
rect 12066 29492 12072 29504
rect 11379 29464 12072 29492
rect 11379 29461 11391 29464
rect 11333 29455 11391 29461
rect 12066 29452 12072 29464
rect 12124 29452 12130 29504
rect 12250 29452 12256 29504
rect 12308 29452 12314 29504
rect 12342 29452 12348 29504
rect 12400 29492 12406 29504
rect 12526 29492 12532 29504
rect 12400 29464 12532 29492
rect 12400 29452 12406 29464
rect 12526 29452 12532 29464
rect 12584 29452 12590 29504
rect 13538 29452 13544 29504
rect 13596 29492 13602 29504
rect 13633 29495 13691 29501
rect 13633 29492 13645 29495
rect 13596 29464 13645 29492
rect 13596 29452 13602 29464
rect 13633 29461 13645 29464
rect 13679 29461 13691 29495
rect 13633 29455 13691 29461
rect 1104 29402 14696 29424
rect 1104 29350 4308 29402
rect 4360 29350 4372 29402
rect 4424 29350 4436 29402
rect 4488 29350 4500 29402
rect 4552 29350 4564 29402
rect 4616 29350 7666 29402
rect 7718 29350 7730 29402
rect 7782 29350 7794 29402
rect 7846 29350 7858 29402
rect 7910 29350 7922 29402
rect 7974 29350 11024 29402
rect 11076 29350 11088 29402
rect 11140 29350 11152 29402
rect 11204 29350 11216 29402
rect 11268 29350 11280 29402
rect 11332 29350 14382 29402
rect 14434 29350 14446 29402
rect 14498 29350 14510 29402
rect 14562 29350 14574 29402
rect 14626 29350 14638 29402
rect 14690 29350 14696 29402
rect 1104 29328 14696 29350
rect 6822 29248 6828 29300
rect 6880 29288 6886 29300
rect 11882 29288 11888 29300
rect 6880 29260 11888 29288
rect 6880 29248 6886 29260
rect 11882 29248 11888 29260
rect 11940 29288 11946 29300
rect 13354 29288 13360 29300
rect 11940 29260 13360 29288
rect 11940 29248 11946 29260
rect 13354 29248 13360 29260
rect 13412 29248 13418 29300
rect 5552 29192 9996 29220
rect 5552 28960 5580 29192
rect 7098 29112 7104 29164
rect 7156 29112 7162 29164
rect 7375 29155 7433 29161
rect 7375 29121 7387 29155
rect 7421 29152 7433 29155
rect 8386 29152 8392 29164
rect 7421 29124 8392 29152
rect 7421 29121 7433 29124
rect 7375 29115 7433 29121
rect 8386 29112 8392 29124
rect 8444 29152 8450 29164
rect 8662 29152 8668 29164
rect 8444 29124 8668 29152
rect 8444 29112 8450 29124
rect 8662 29112 8668 29124
rect 8720 29112 8726 29164
rect 8755 29155 8813 29161
rect 8755 29121 8767 29155
rect 8801 29152 8813 29155
rect 9766 29152 9772 29164
rect 8801 29124 9772 29152
rect 8801 29121 8813 29124
rect 8755 29115 8813 29121
rect 9766 29112 9772 29124
rect 9824 29112 9830 29164
rect 9968 29152 9996 29192
rect 10226 29180 10232 29232
rect 10284 29220 10290 29232
rect 10502 29220 10508 29232
rect 10284 29192 10508 29220
rect 10284 29180 10290 29192
rect 10502 29180 10508 29192
rect 10560 29180 10566 29232
rect 10778 29180 10784 29232
rect 10836 29220 10842 29232
rect 12618 29220 12624 29232
rect 10836 29192 12624 29220
rect 10836 29180 10842 29192
rect 12618 29180 12624 29192
rect 12676 29180 12682 29232
rect 10134 29152 10140 29164
rect 9968 29124 10140 29152
rect 10134 29112 10140 29124
rect 10192 29112 10198 29164
rect 11054 29112 11060 29164
rect 11112 29152 11118 29164
rect 12035 29155 12093 29161
rect 12035 29152 12047 29155
rect 11112 29124 12047 29152
rect 11112 29112 11118 29124
rect 12035 29121 12047 29124
rect 12081 29121 12093 29155
rect 12035 29115 12093 29121
rect 13541 29155 13599 29161
rect 13541 29121 13553 29155
rect 13587 29152 13599 29155
rect 13630 29152 13636 29164
rect 13587 29124 13636 29152
rect 13587 29121 13599 29124
rect 13541 29115 13599 29121
rect 13630 29112 13636 29124
rect 13688 29112 13694 29164
rect 5534 28908 5540 28960
rect 5592 28908 5598 28960
rect 7116 28948 7144 29112
rect 8481 29087 8539 29093
rect 8481 29084 8493 29087
rect 8036 29056 8493 29084
rect 8036 28948 8064 29056
rect 8481 29053 8493 29056
rect 8527 29053 8539 29087
rect 8481 29047 8539 29053
rect 9674 29044 9680 29096
rect 9732 29084 9738 29096
rect 9861 29087 9919 29093
rect 9861 29084 9873 29087
rect 9732 29056 9873 29084
rect 9732 29044 9738 29056
rect 9861 29053 9873 29056
rect 9907 29053 9919 29087
rect 9861 29047 9919 29053
rect 11606 29044 11612 29096
rect 11664 29084 11670 29096
rect 11790 29084 11796 29096
rect 11664 29056 11796 29084
rect 11664 29044 11670 29056
rect 11790 29044 11796 29056
rect 11848 29044 11854 29096
rect 9493 29019 9551 29025
rect 9493 28985 9505 29019
rect 9539 29016 9551 29019
rect 9539 28988 9996 29016
rect 9539 28985 9551 28988
rect 9493 28979 9551 28985
rect 7116 28920 8064 28948
rect 8110 28908 8116 28960
rect 8168 28908 8174 28960
rect 9968 28948 9996 28988
rect 11330 28976 11336 29028
rect 11388 29016 11394 29028
rect 11698 29016 11704 29028
rect 11388 28988 11704 29016
rect 11388 28976 11394 28988
rect 11698 28976 11704 28988
rect 11756 28976 11762 29028
rect 13814 28976 13820 29028
rect 13872 28976 13878 29028
rect 10134 28948 10140 28960
rect 9968 28920 10140 28948
rect 10134 28908 10140 28920
rect 10192 28908 10198 28960
rect 10870 28908 10876 28960
rect 10928 28908 10934 28960
rect 12250 28908 12256 28960
rect 12308 28948 12314 28960
rect 12710 28948 12716 28960
rect 12308 28920 12716 28948
rect 12308 28908 12314 28920
rect 12710 28908 12716 28920
rect 12768 28908 12774 28960
rect 12805 28951 12863 28957
rect 12805 28917 12817 28951
rect 12851 28948 12863 28951
rect 13078 28948 13084 28960
rect 12851 28920 13084 28948
rect 12851 28917 12863 28920
rect 12805 28911 12863 28917
rect 13078 28908 13084 28920
rect 13136 28908 13142 28960
rect 1104 28858 14536 28880
rect 1104 28806 2629 28858
rect 2681 28806 2693 28858
rect 2745 28806 2757 28858
rect 2809 28806 2821 28858
rect 2873 28806 2885 28858
rect 2937 28806 5987 28858
rect 6039 28806 6051 28858
rect 6103 28806 6115 28858
rect 6167 28806 6179 28858
rect 6231 28806 6243 28858
rect 6295 28806 9345 28858
rect 9397 28806 9409 28858
rect 9461 28806 9473 28858
rect 9525 28806 9537 28858
rect 9589 28806 9601 28858
rect 9653 28806 12703 28858
rect 12755 28806 12767 28858
rect 12819 28806 12831 28858
rect 12883 28806 12895 28858
rect 12947 28806 12959 28858
rect 13011 28806 14536 28858
rect 1104 28784 14536 28806
rect 1581 28747 1639 28753
rect 1581 28713 1593 28747
rect 1627 28744 1639 28747
rect 1946 28744 1952 28756
rect 1627 28716 1952 28744
rect 1627 28713 1639 28716
rect 1581 28707 1639 28713
rect 1946 28704 1952 28716
rect 2004 28744 2010 28756
rect 12250 28744 12256 28756
rect 2004 28716 12256 28744
rect 2004 28704 2010 28716
rect 12250 28704 12256 28716
rect 12308 28704 12314 28756
rect 13262 28704 13268 28756
rect 13320 28704 13326 28756
rect 10870 28636 10876 28688
rect 10928 28676 10934 28688
rect 11517 28679 11575 28685
rect 11517 28676 11529 28679
rect 10928 28648 11529 28676
rect 10928 28636 10934 28648
rect 11517 28645 11529 28648
rect 11563 28645 11575 28679
rect 11517 28639 11575 28645
rect 12713 28679 12771 28685
rect 12713 28645 12725 28679
rect 12759 28676 12771 28679
rect 13280 28676 13308 28704
rect 12759 28648 13308 28676
rect 12759 28645 12771 28648
rect 12713 28639 12771 28645
rect 7098 28608 7104 28620
rect 6472 28580 7104 28608
rect 6472 28552 6500 28580
rect 7098 28568 7104 28580
rect 7156 28568 7162 28620
rect 11790 28568 11796 28620
rect 11848 28568 11854 28620
rect 13173 28611 13231 28617
rect 13173 28577 13185 28611
rect 13219 28608 13231 28611
rect 15010 28608 15016 28620
rect 13219 28580 15016 28608
rect 13219 28577 13231 28580
rect 13173 28571 13231 28577
rect 15010 28568 15016 28580
rect 15068 28568 15074 28620
rect 750 28500 756 28552
rect 808 28540 814 28552
rect 1397 28543 1455 28549
rect 1397 28540 1409 28543
rect 808 28512 1409 28540
rect 808 28500 814 28512
rect 1397 28509 1409 28512
rect 1443 28509 1455 28543
rect 1397 28503 1455 28509
rect 6454 28500 6460 28552
rect 6512 28500 6518 28552
rect 6914 28500 6920 28552
rect 6972 28540 6978 28552
rect 7343 28543 7401 28549
rect 7343 28540 7355 28543
rect 6972 28512 7355 28540
rect 6972 28500 6978 28512
rect 7343 28509 7355 28512
rect 7389 28509 7401 28543
rect 7343 28503 7401 28509
rect 8938 28500 8944 28552
rect 8996 28540 9002 28552
rect 9214 28540 9220 28552
rect 8996 28512 9220 28540
rect 8996 28500 9002 28512
rect 9214 28500 9220 28512
rect 9272 28500 9278 28552
rect 10873 28543 10931 28549
rect 10873 28509 10885 28543
rect 10919 28509 10931 28543
rect 10873 28503 10931 28509
rect 11057 28543 11115 28549
rect 11057 28509 11069 28543
rect 11103 28509 11115 28543
rect 11057 28503 11115 28509
rect 10888 28472 10916 28503
rect 7300 28444 8984 28472
rect 7098 28364 7104 28416
rect 7156 28404 7162 28416
rect 7300 28404 7328 28444
rect 8956 28416 8984 28444
rect 10520 28444 10916 28472
rect 7156 28376 7328 28404
rect 7156 28364 7162 28376
rect 7558 28364 7564 28416
rect 7616 28404 7622 28416
rect 8113 28407 8171 28413
rect 8113 28404 8125 28407
rect 7616 28376 8125 28404
rect 7616 28364 7622 28376
rect 8113 28373 8125 28376
rect 8159 28373 8171 28407
rect 8113 28367 8171 28373
rect 8294 28364 8300 28416
rect 8352 28404 8358 28416
rect 8662 28404 8668 28416
rect 8352 28376 8668 28404
rect 8352 28364 8358 28376
rect 8662 28364 8668 28376
rect 8720 28364 8726 28416
rect 8938 28364 8944 28416
rect 8996 28364 9002 28416
rect 9674 28364 9680 28416
rect 9732 28404 9738 28416
rect 10520 28413 10548 28444
rect 10505 28407 10563 28413
rect 10505 28404 10517 28407
rect 9732 28376 10517 28404
rect 9732 28364 9738 28376
rect 10505 28373 10517 28376
rect 10551 28373 10563 28407
rect 11072 28404 11100 28503
rect 11882 28500 11888 28552
rect 11940 28549 11946 28552
rect 11940 28543 11968 28549
rect 11956 28509 11968 28543
rect 11940 28503 11968 28509
rect 11940 28500 11946 28503
rect 12066 28500 12072 28552
rect 12124 28500 12130 28552
rect 12710 28500 12716 28552
rect 12768 28540 12774 28552
rect 12768 28512 13492 28540
rect 12768 28500 12774 28512
rect 12802 28432 12808 28484
rect 12860 28472 12866 28484
rect 13464 28481 13492 28512
rect 12897 28475 12955 28481
rect 12897 28472 12909 28475
rect 12860 28444 12909 28472
rect 12860 28432 12866 28444
rect 12897 28441 12909 28444
rect 12943 28441 12955 28475
rect 12897 28435 12955 28441
rect 13449 28475 13507 28481
rect 13449 28441 13461 28475
rect 13495 28441 13507 28475
rect 13449 28435 13507 28441
rect 11882 28404 11888 28416
rect 11072 28376 11888 28404
rect 10505 28367 10563 28373
rect 11882 28364 11888 28376
rect 11940 28364 11946 28416
rect 12710 28364 12716 28416
rect 12768 28404 12774 28416
rect 13078 28404 13084 28416
rect 12768 28376 13084 28404
rect 12768 28364 12774 28376
rect 13078 28364 13084 28376
rect 13136 28364 13142 28416
rect 13722 28364 13728 28416
rect 13780 28364 13786 28416
rect 1104 28314 14696 28336
rect 1104 28262 4308 28314
rect 4360 28262 4372 28314
rect 4424 28262 4436 28314
rect 4488 28262 4500 28314
rect 4552 28262 4564 28314
rect 4616 28262 7666 28314
rect 7718 28262 7730 28314
rect 7782 28262 7794 28314
rect 7846 28262 7858 28314
rect 7910 28262 7922 28314
rect 7974 28262 11024 28314
rect 11076 28262 11088 28314
rect 11140 28262 11152 28314
rect 11204 28262 11216 28314
rect 11268 28262 11280 28314
rect 11332 28262 14382 28314
rect 14434 28262 14446 28314
rect 14498 28262 14510 28314
rect 14562 28262 14574 28314
rect 14626 28262 14638 28314
rect 14690 28262 14696 28314
rect 1104 28240 14696 28262
rect 7098 28160 7104 28212
rect 7156 28160 7162 28212
rect 8849 28203 8907 28209
rect 7208 28172 8800 28200
rect 1394 28024 1400 28076
rect 1452 28024 1458 28076
rect 7009 28067 7067 28073
rect 7009 28033 7021 28067
rect 7055 28064 7067 28067
rect 7116 28064 7144 28160
rect 7055 28036 7144 28064
rect 7055 28033 7067 28036
rect 7009 28027 7067 28033
rect 7208 28005 7236 28172
rect 8772 28132 8800 28172
rect 8849 28169 8861 28203
rect 8895 28200 8907 28203
rect 8895 28172 11652 28200
rect 8895 28169 8907 28172
rect 8849 28163 8907 28169
rect 11624 28141 11652 28172
rect 11882 28160 11888 28212
rect 11940 28200 11946 28212
rect 13446 28200 13452 28212
rect 11940 28172 13452 28200
rect 11940 28160 11946 28172
rect 11609 28135 11667 28141
rect 8772 28104 9168 28132
rect 8202 28024 8208 28076
rect 8260 28024 8266 28076
rect 9140 28073 9168 28104
rect 11609 28101 11621 28135
rect 11655 28101 11667 28135
rect 11609 28095 11667 28101
rect 9125 28067 9183 28073
rect 8864 28036 9076 28064
rect 7193 27999 7251 28005
rect 7193 27965 7205 27999
rect 7239 27996 7251 27999
rect 7282 27996 7288 28008
rect 7239 27968 7288 27996
rect 7239 27965 7251 27968
rect 7193 27959 7251 27965
rect 7282 27956 7288 27968
rect 7340 27956 7346 28008
rect 7558 27956 7564 28008
rect 7616 27996 7622 28008
rect 7653 27999 7711 28005
rect 7653 27996 7665 27999
rect 7616 27968 7665 27996
rect 7616 27956 7622 27968
rect 7653 27965 7665 27968
rect 7699 27965 7711 27999
rect 7653 27959 7711 27965
rect 7926 27956 7932 28008
rect 7984 27956 7990 28008
rect 8067 27999 8125 28005
rect 8067 27965 8079 27999
rect 8113 27996 8125 27999
rect 8864 27996 8892 28036
rect 8113 27968 8892 27996
rect 8113 27965 8125 27968
rect 8067 27959 8125 27965
rect 8938 27956 8944 28008
rect 8996 27956 9002 28008
rect 9048 27996 9076 28036
rect 9125 28033 9137 28067
rect 9171 28033 9183 28067
rect 9125 28027 9183 28033
rect 9950 28024 9956 28076
rect 10008 28073 10014 28076
rect 10008 28067 10036 28073
rect 10024 28033 10036 28067
rect 10008 28027 10036 28033
rect 10008 28024 10014 28027
rect 10134 28024 10140 28076
rect 10192 28024 10198 28076
rect 10962 28024 10968 28076
rect 11020 28024 11026 28076
rect 11974 28024 11980 28076
rect 12032 28064 12038 28076
rect 12406 28064 12434 28172
rect 13446 28160 13452 28172
rect 13504 28160 13510 28212
rect 14182 28160 14188 28212
rect 14240 28160 14246 28212
rect 12529 28067 12587 28073
rect 12529 28064 12541 28067
rect 12032 28036 12296 28064
rect 12406 28036 12541 28064
rect 12032 28024 12038 28036
rect 9306 27996 9312 28008
rect 9048 27968 9312 27996
rect 9306 27956 9312 27968
rect 9364 27956 9370 28008
rect 9861 27999 9919 28005
rect 9861 27996 9873 27999
rect 9692 27968 9873 27996
rect 9585 27931 9643 27937
rect 9585 27928 9597 27931
rect 8864 27900 9597 27928
rect 1578 27820 1584 27872
rect 1636 27820 1642 27872
rect 8110 27820 8116 27872
rect 8168 27860 8174 27872
rect 8864 27860 8892 27900
rect 9585 27897 9597 27900
rect 9631 27897 9643 27931
rect 9585 27891 9643 27897
rect 8168 27832 8892 27860
rect 8168 27820 8174 27832
rect 8938 27820 8944 27872
rect 8996 27860 9002 27872
rect 9692 27860 9720 27968
rect 9861 27965 9873 27968
rect 9907 27996 9919 27999
rect 10778 27996 10784 28008
rect 9907 27968 10784 27996
rect 9907 27965 9919 27968
rect 9861 27959 9919 27965
rect 10778 27956 10784 27968
rect 10836 27956 10842 28008
rect 8996 27832 9720 27860
rect 8996 27820 9002 27832
rect 10042 27820 10048 27872
rect 10100 27860 10106 27872
rect 10686 27860 10692 27872
rect 10100 27832 10692 27860
rect 10100 27820 10106 27832
rect 10686 27820 10692 27832
rect 10744 27820 10750 27872
rect 10778 27820 10784 27872
rect 10836 27820 10842 27872
rect 11241 27863 11299 27869
rect 11241 27829 11253 27863
rect 11287 27860 11299 27863
rect 11606 27860 11612 27872
rect 11287 27832 11612 27860
rect 11287 27829 11299 27832
rect 11241 27823 11299 27829
rect 11606 27820 11612 27832
rect 11664 27820 11670 27872
rect 11885 27863 11943 27869
rect 11885 27829 11897 27863
rect 11931 27860 11943 27863
rect 12066 27860 12072 27872
rect 11931 27832 12072 27860
rect 11931 27829 11943 27832
rect 11885 27823 11943 27829
rect 12066 27820 12072 27832
rect 12124 27820 12130 27872
rect 12268 27860 12296 28036
rect 12529 28033 12541 28036
rect 12575 28033 12587 28067
rect 12529 28027 12587 28033
rect 13538 28024 13544 28076
rect 13596 28024 13602 28076
rect 12342 27956 12348 28008
rect 12400 27956 12406 28008
rect 12710 27956 12716 28008
rect 12768 27996 12774 28008
rect 12989 27999 13047 28005
rect 12989 27996 13001 27999
rect 12768 27968 13001 27996
rect 12768 27956 12774 27968
rect 12989 27965 13001 27968
rect 13035 27965 13047 27999
rect 13265 27999 13323 28005
rect 13265 27996 13277 27999
rect 12989 27959 13047 27965
rect 13096 27968 13277 27996
rect 13096 27872 13124 27968
rect 13265 27965 13277 27968
rect 13311 27965 13323 27999
rect 13265 27959 13323 27965
rect 13354 27956 13360 28008
rect 13412 28005 13418 28008
rect 13412 27999 13440 28005
rect 13428 27965 13440 27999
rect 13412 27959 13440 27965
rect 13412 27956 13418 27959
rect 13078 27860 13084 27872
rect 12268 27832 13084 27860
rect 13078 27820 13084 27832
rect 13136 27820 13142 27872
rect 1104 27770 14536 27792
rect 1104 27718 2629 27770
rect 2681 27718 2693 27770
rect 2745 27718 2757 27770
rect 2809 27718 2821 27770
rect 2873 27718 2885 27770
rect 2937 27718 5987 27770
rect 6039 27718 6051 27770
rect 6103 27718 6115 27770
rect 6167 27718 6179 27770
rect 6231 27718 6243 27770
rect 6295 27718 9345 27770
rect 9397 27718 9409 27770
rect 9461 27718 9473 27770
rect 9525 27718 9537 27770
rect 9589 27718 9601 27770
rect 9653 27718 12703 27770
rect 12755 27718 12767 27770
rect 12819 27718 12831 27770
rect 12883 27718 12895 27770
rect 12947 27718 12959 27770
rect 13011 27718 14536 27770
rect 1104 27696 14536 27718
rect 6822 27616 6828 27668
rect 6880 27656 6886 27668
rect 6880 27628 8156 27656
rect 6880 27616 6886 27628
rect 2869 27591 2927 27597
rect 2869 27557 2881 27591
rect 2915 27588 2927 27591
rect 3050 27588 3056 27600
rect 2915 27560 3056 27588
rect 2915 27557 2927 27560
rect 2869 27551 2927 27557
rect 3050 27548 3056 27560
rect 3108 27548 3114 27600
rect 3878 27548 3884 27600
rect 3936 27588 3942 27600
rect 7466 27588 7472 27600
rect 3936 27560 7472 27588
rect 3936 27548 3942 27560
rect 7466 27548 7472 27560
rect 7524 27548 7530 27600
rect 1670 27480 1676 27532
rect 1728 27520 1734 27532
rect 7374 27520 7380 27532
rect 1728 27492 7380 27520
rect 1728 27480 1734 27492
rect 7374 27480 7380 27492
rect 7432 27480 7438 27532
rect 1854 27412 1860 27464
rect 1912 27412 1918 27464
rect 2682 27412 2688 27464
rect 2740 27412 2746 27464
rect 6454 27412 6460 27464
rect 6512 27452 6518 27464
rect 7469 27455 7527 27461
rect 7469 27452 7481 27455
rect 6512 27424 7481 27452
rect 6512 27412 6518 27424
rect 7469 27421 7481 27424
rect 7515 27421 7527 27455
rect 7711 27455 7769 27461
rect 7711 27452 7723 27455
rect 7469 27415 7527 27421
rect 7576 27424 7723 27452
rect 1872 27384 1900 27412
rect 7576 27384 7604 27424
rect 7711 27421 7723 27424
rect 7757 27421 7769 27455
rect 7711 27415 7769 27421
rect 1872 27356 7604 27384
rect 8128 27384 8156 27628
rect 8202 27616 8208 27668
rect 8260 27616 8266 27668
rect 10962 27656 10968 27668
rect 8588 27628 10968 27656
rect 8220 27588 8248 27616
rect 8481 27591 8539 27597
rect 8481 27588 8493 27591
rect 8220 27560 8493 27588
rect 8481 27557 8493 27560
rect 8527 27557 8539 27591
rect 8481 27551 8539 27557
rect 8202 27412 8208 27464
rect 8260 27452 8266 27464
rect 8588 27452 8616 27628
rect 10962 27616 10968 27628
rect 11020 27616 11026 27668
rect 11698 27616 11704 27668
rect 11756 27616 11762 27668
rect 9674 27548 9680 27600
rect 9732 27588 9738 27600
rect 9950 27588 9956 27600
rect 9732 27560 9956 27588
rect 9732 27548 9738 27560
rect 9950 27548 9956 27560
rect 10008 27548 10014 27600
rect 11716 27588 11744 27616
rect 11624 27560 11744 27588
rect 11624 27529 11652 27560
rect 11609 27523 11667 27529
rect 11609 27489 11621 27523
rect 11655 27489 11667 27523
rect 11609 27483 11667 27489
rect 8260 27424 8616 27452
rect 8260 27412 8266 27424
rect 10226 27412 10232 27464
rect 10284 27412 10290 27464
rect 11624 27452 11652 27483
rect 10487 27425 10545 27431
rect 10487 27422 10499 27425
rect 10428 27394 10499 27422
rect 10428 27384 10456 27394
rect 10487 27391 10499 27394
rect 10533 27391 10545 27425
rect 10487 27385 10545 27391
rect 10704 27424 11652 27452
rect 11882 27431 11888 27464
rect 11867 27425 11888 27431
rect 8128 27356 10456 27384
rect 7190 27276 7196 27328
rect 7248 27316 7254 27328
rect 8754 27316 8760 27328
rect 7248 27288 8760 27316
rect 7248 27276 7254 27288
rect 8754 27276 8760 27288
rect 8812 27276 8818 27328
rect 9674 27276 9680 27328
rect 9732 27316 9738 27328
rect 10226 27316 10232 27328
rect 9732 27288 10232 27316
rect 9732 27276 9738 27288
rect 10226 27276 10232 27288
rect 10284 27316 10290 27328
rect 10704 27316 10732 27424
rect 11867 27391 11879 27425
rect 11940 27412 11946 27464
rect 11913 27394 11928 27412
rect 11913 27391 11925 27394
rect 11867 27385 11925 27391
rect 12342 27344 12348 27396
rect 12400 27384 12406 27396
rect 13081 27387 13139 27393
rect 13081 27384 13093 27387
rect 12400 27356 13093 27384
rect 12400 27344 12406 27356
rect 13081 27353 13093 27356
rect 13127 27353 13139 27387
rect 13081 27347 13139 27353
rect 13446 27344 13452 27396
rect 13504 27344 13510 27396
rect 10284 27288 10732 27316
rect 11241 27319 11299 27325
rect 10284 27276 10290 27288
rect 11241 27285 11253 27319
rect 11287 27316 11299 27319
rect 11698 27316 11704 27328
rect 11287 27288 11704 27316
rect 11287 27285 11299 27288
rect 11241 27279 11299 27285
rect 11698 27276 11704 27288
rect 11756 27276 11762 27328
rect 12621 27319 12679 27325
rect 12621 27285 12633 27319
rect 12667 27316 12679 27319
rect 12710 27316 12716 27328
rect 12667 27288 12716 27316
rect 12667 27285 12679 27288
rect 12621 27279 12679 27285
rect 12710 27276 12716 27288
rect 12768 27276 12774 27328
rect 1104 27226 14696 27248
rect 1104 27174 4308 27226
rect 4360 27174 4372 27226
rect 4424 27174 4436 27226
rect 4488 27174 4500 27226
rect 4552 27174 4564 27226
rect 4616 27174 7666 27226
rect 7718 27174 7730 27226
rect 7782 27174 7794 27226
rect 7846 27174 7858 27226
rect 7910 27174 7922 27226
rect 7974 27174 11024 27226
rect 11076 27174 11088 27226
rect 11140 27174 11152 27226
rect 11204 27174 11216 27226
rect 11268 27174 11280 27226
rect 11332 27174 14382 27226
rect 14434 27174 14446 27226
rect 14498 27174 14510 27226
rect 14562 27174 14574 27226
rect 14626 27174 14638 27226
rect 14690 27174 14696 27226
rect 1104 27152 14696 27174
rect 1581 27115 1639 27121
rect 1581 27081 1593 27115
rect 1627 27112 1639 27115
rect 1670 27112 1676 27124
rect 1627 27084 1676 27112
rect 1627 27081 1639 27084
rect 1581 27075 1639 27081
rect 1670 27072 1676 27084
rect 1728 27072 1734 27124
rect 2682 27072 2688 27124
rect 2740 27112 2746 27124
rect 2777 27115 2835 27121
rect 2777 27112 2789 27115
rect 2740 27084 2789 27112
rect 2740 27072 2746 27084
rect 2777 27081 2789 27084
rect 2823 27081 2835 27115
rect 2777 27075 2835 27081
rect 4908 27084 6500 27112
rect 4908 26988 4936 27084
rect 6472 27056 6500 27084
rect 7374 27072 7380 27124
rect 7432 27112 7438 27124
rect 7432 27084 8156 27112
rect 7432 27072 7438 27084
rect 5442 27044 5448 27056
rect 5184 27016 5448 27044
rect 5184 26988 5212 27016
rect 5442 27004 5448 27016
rect 5500 27004 5506 27056
rect 6454 27004 6460 27056
rect 6512 27004 6518 27056
rect 8128 27044 8156 27084
rect 8202 27072 8208 27124
rect 8260 27072 8266 27124
rect 10594 27072 10600 27124
rect 10652 27112 10658 27124
rect 11790 27112 11796 27124
rect 10652 27084 11796 27112
rect 10652 27072 10658 27084
rect 11790 27072 11796 27084
rect 11848 27072 11854 27124
rect 14185 27115 14243 27121
rect 14185 27112 14197 27115
rect 12406 27084 14197 27112
rect 11609 27047 11667 27053
rect 8128 27016 9812 27044
rect 750 26936 756 26988
rect 808 26976 814 26988
rect 1489 26979 1547 26985
rect 1489 26976 1501 26979
rect 808 26948 1501 26976
rect 808 26936 814 26948
rect 1489 26945 1501 26948
rect 1535 26945 1547 26979
rect 1489 26939 1547 26945
rect 2961 26979 3019 26985
rect 2961 26945 2973 26979
rect 3007 26976 3019 26979
rect 4154 26976 4160 26988
rect 3007 26948 4160 26976
rect 3007 26945 3019 26948
rect 2961 26939 3019 26945
rect 4154 26936 4160 26948
rect 4212 26936 4218 26988
rect 4890 26936 4896 26988
rect 4948 26936 4954 26988
rect 5166 26976 5172 26988
rect 5127 26948 5172 26976
rect 5166 26936 5172 26948
rect 5224 26936 5230 26988
rect 5902 26936 5908 26988
rect 5960 26976 5966 26988
rect 6365 26979 6423 26985
rect 6365 26976 6377 26979
rect 5960 26948 6377 26976
rect 5960 26936 5966 26948
rect 6365 26945 6377 26948
rect 6411 26945 6423 26979
rect 6365 26939 6423 26945
rect 7558 26936 7564 26988
rect 7616 26936 7622 26988
rect 9674 26936 9680 26988
rect 9732 26936 9738 26988
rect 9784 26986 9812 27016
rect 11609 27013 11621 27047
rect 11655 27044 11667 27047
rect 12406 27044 12434 27084
rect 14185 27081 14197 27084
rect 14231 27081 14243 27115
rect 14185 27075 14243 27081
rect 11655 27016 12434 27044
rect 11655 27013 11667 27016
rect 11609 27007 11667 27013
rect 10103 26989 10161 26995
rect 9784 26976 9994 26986
rect 10103 26976 10115 26989
rect 9784 26958 10115 26976
rect 9966 26955 10115 26958
rect 10149 26986 10161 26989
rect 10149 26955 10162 26986
rect 12345 26979 12403 26985
rect 12345 26976 12357 26979
rect 9966 26948 10162 26955
rect 12268 26948 12357 26976
rect 6546 26868 6552 26920
rect 6604 26868 6610 26920
rect 7285 26911 7343 26917
rect 7285 26908 7297 26911
rect 7116 26880 7297 26908
rect 5905 26843 5963 26849
rect 5905 26809 5917 26843
rect 5951 26840 5963 26843
rect 7009 26843 7067 26849
rect 7009 26840 7021 26843
rect 5951 26812 7021 26840
rect 5951 26809 5963 26812
rect 5905 26803 5963 26809
rect 7009 26809 7021 26812
rect 7055 26809 7067 26843
rect 7009 26803 7067 26809
rect 5810 26732 5816 26784
rect 5868 26772 5874 26784
rect 7116 26772 7144 26880
rect 7285 26877 7297 26880
rect 7331 26877 7343 26911
rect 7285 26871 7343 26877
rect 7374 26868 7380 26920
rect 7432 26917 7438 26920
rect 7432 26911 7460 26917
rect 7448 26877 7460 26911
rect 7432 26871 7460 26877
rect 7432 26868 7438 26871
rect 7742 26868 7748 26920
rect 7800 26908 7806 26920
rect 9692 26908 9720 26936
rect 12268 26920 12296 26948
rect 12345 26945 12357 26948
rect 12391 26945 12403 26979
rect 12345 26939 12403 26945
rect 12710 26936 12716 26988
rect 12768 26936 12774 26988
rect 9861 26911 9919 26917
rect 9861 26908 9873 26911
rect 7800 26880 8616 26908
rect 9692 26880 9873 26908
rect 7800 26868 7806 26880
rect 8478 26772 8484 26784
rect 5868 26744 8484 26772
rect 5868 26732 5874 26744
rect 8478 26732 8484 26744
rect 8536 26732 8542 26784
rect 8588 26772 8616 26880
rect 9861 26877 9873 26880
rect 9907 26877 9919 26911
rect 9861 26871 9919 26877
rect 10870 26868 10876 26920
rect 10928 26908 10934 26920
rect 11790 26908 11796 26920
rect 10928 26880 11796 26908
rect 10928 26868 10934 26880
rect 11790 26868 11796 26880
rect 11848 26868 11854 26920
rect 12250 26868 12256 26920
rect 12308 26868 12314 26920
rect 12526 26868 12532 26920
rect 12584 26868 12590 26920
rect 12728 26908 12756 26936
rect 12989 26911 13047 26917
rect 12989 26908 13001 26911
rect 12728 26880 13001 26908
rect 12989 26877 13001 26880
rect 13035 26877 13047 26911
rect 12989 26871 13047 26877
rect 13078 26868 13084 26920
rect 13136 26908 13142 26920
rect 13265 26911 13323 26917
rect 13265 26908 13277 26911
rect 13136 26880 13277 26908
rect 13136 26868 13142 26880
rect 13265 26877 13277 26880
rect 13311 26877 13323 26911
rect 13265 26871 13323 26877
rect 13354 26868 13360 26920
rect 13412 26917 13418 26920
rect 13412 26911 13440 26917
rect 13428 26877 13440 26911
rect 13412 26871 13440 26877
rect 13412 26868 13418 26871
rect 13538 26868 13544 26920
rect 13596 26868 13602 26920
rect 12342 26840 12348 26852
rect 10520 26812 12348 26840
rect 10520 26772 10548 26812
rect 12342 26800 12348 26812
rect 12400 26800 12406 26852
rect 8588 26744 10548 26772
rect 10870 26732 10876 26784
rect 10928 26732 10934 26784
rect 11885 26775 11943 26781
rect 11885 26741 11897 26775
rect 11931 26772 11943 26775
rect 13998 26772 14004 26784
rect 11931 26744 14004 26772
rect 11931 26741 11943 26744
rect 11885 26735 11943 26741
rect 13998 26732 14004 26744
rect 14056 26732 14062 26784
rect 1104 26682 14536 26704
rect 1104 26630 2629 26682
rect 2681 26630 2693 26682
rect 2745 26630 2757 26682
rect 2809 26630 2821 26682
rect 2873 26630 2885 26682
rect 2937 26630 5987 26682
rect 6039 26630 6051 26682
rect 6103 26630 6115 26682
rect 6167 26630 6179 26682
rect 6231 26630 6243 26682
rect 6295 26630 9345 26682
rect 9397 26630 9409 26682
rect 9461 26630 9473 26682
rect 9525 26630 9537 26682
rect 9589 26630 9601 26682
rect 9653 26630 12703 26682
rect 12755 26630 12767 26682
rect 12819 26630 12831 26682
rect 12883 26630 12895 26682
rect 12947 26630 12959 26682
rect 13011 26630 14536 26682
rect 1104 26608 14536 26630
rect 8205 26571 8263 26577
rect 5828 26540 7972 26568
rect 4890 26460 4896 26512
rect 4948 26460 4954 26512
rect 4908 26432 4936 26460
rect 4985 26435 5043 26441
rect 4985 26432 4997 26435
rect 4908 26404 4997 26432
rect 4985 26401 4997 26404
rect 5031 26401 5043 26435
rect 4985 26395 5043 26401
rect 4890 26324 4896 26376
rect 4948 26364 4954 26376
rect 5259 26367 5317 26373
rect 5259 26364 5271 26367
rect 4948 26336 5271 26364
rect 4948 26324 4954 26336
rect 5259 26333 5271 26336
rect 5305 26364 5317 26367
rect 5828 26364 5856 26540
rect 5997 26503 6055 26509
rect 5997 26469 6009 26503
rect 6043 26500 6055 26503
rect 7009 26503 7067 26509
rect 7009 26500 7021 26503
rect 6043 26472 7021 26500
rect 6043 26469 6055 26472
rect 5997 26463 6055 26469
rect 7009 26469 7021 26472
rect 7055 26469 7067 26503
rect 7944 26500 7972 26540
rect 8205 26537 8217 26571
rect 8251 26568 8263 26571
rect 10042 26568 10048 26580
rect 8251 26540 10048 26568
rect 8251 26537 8263 26540
rect 8205 26531 8263 26537
rect 10042 26528 10048 26540
rect 10100 26528 10106 26580
rect 10870 26528 10876 26580
rect 10928 26528 10934 26580
rect 12345 26571 12403 26577
rect 12345 26537 12357 26571
rect 12391 26568 12403 26571
rect 12618 26568 12624 26580
rect 12391 26540 12624 26568
rect 12391 26537 12403 26540
rect 12345 26531 12403 26537
rect 12618 26528 12624 26540
rect 12676 26528 12682 26580
rect 13538 26528 13544 26580
rect 13596 26568 13602 26580
rect 13633 26571 13691 26577
rect 13633 26568 13645 26571
rect 13596 26540 13645 26568
rect 13596 26528 13602 26540
rect 13633 26537 13645 26540
rect 13679 26537 13691 26571
rect 13633 26531 13691 26537
rect 9122 26500 9128 26512
rect 7944 26472 9128 26500
rect 7009 26463 7067 26469
rect 9122 26460 9128 26472
rect 9180 26460 9186 26512
rect 10502 26460 10508 26512
rect 10560 26500 10566 26512
rect 10888 26500 10916 26528
rect 11149 26503 11207 26509
rect 11149 26500 11161 26503
rect 10560 26472 10732 26500
rect 10888 26472 11161 26500
rect 10560 26460 10566 26472
rect 10704 26444 10732 26472
rect 11149 26469 11161 26472
rect 11195 26469 11207 26503
rect 11149 26463 11207 26469
rect 7374 26392 7380 26444
rect 7432 26441 7438 26444
rect 7432 26435 7460 26441
rect 7448 26401 7460 26435
rect 7432 26395 7460 26401
rect 7432 26392 7438 26395
rect 10686 26392 10692 26444
rect 10744 26392 10750 26444
rect 10870 26432 10876 26444
rect 10778 26404 10876 26432
rect 5305 26336 5856 26364
rect 5305 26333 5317 26336
rect 5259 26327 5317 26333
rect 5902 26324 5908 26376
rect 5960 26364 5966 26376
rect 6365 26367 6423 26373
rect 6365 26364 6377 26367
rect 5960 26336 6377 26364
rect 5960 26324 5966 26336
rect 6365 26333 6377 26336
rect 6411 26333 6423 26367
rect 6365 26327 6423 26333
rect 6546 26324 6552 26376
rect 6604 26324 6610 26376
rect 7282 26324 7288 26376
rect 7340 26324 7346 26376
rect 7558 26324 7564 26376
rect 7616 26324 7622 26376
rect 10505 26367 10563 26373
rect 10505 26333 10517 26367
rect 10551 26364 10563 26367
rect 10594 26364 10600 26376
rect 10551 26336 10600 26364
rect 10551 26333 10563 26336
rect 10505 26327 10563 26333
rect 10594 26324 10600 26336
rect 10652 26324 10658 26376
rect 10778 26364 10806 26404
rect 10870 26392 10876 26404
rect 10928 26432 10934 26444
rect 11425 26435 11483 26441
rect 11425 26432 11437 26435
rect 10928 26404 11437 26432
rect 10928 26392 10934 26404
rect 11425 26401 11437 26404
rect 11471 26401 11483 26435
rect 11425 26395 11483 26401
rect 11563 26435 11621 26441
rect 11563 26401 11575 26435
rect 11609 26432 11621 26435
rect 12066 26432 12072 26444
rect 11609 26404 12072 26432
rect 11609 26401 11621 26404
rect 11563 26395 11621 26401
rect 12066 26392 12072 26404
rect 12124 26392 12130 26444
rect 10704 26336 10806 26364
rect 1486 26256 1492 26308
rect 1544 26256 1550 26308
rect 1673 26299 1731 26305
rect 1673 26265 1685 26299
rect 1719 26296 1731 26299
rect 5718 26296 5724 26308
rect 1719 26268 5724 26296
rect 1719 26265 1731 26268
rect 1673 26259 1731 26265
rect 5718 26256 5724 26268
rect 5776 26256 5782 26308
rect 6270 26256 6276 26308
rect 6328 26296 6334 26308
rect 6564 26296 6592 26324
rect 6328 26268 6592 26296
rect 6328 26256 6334 26268
rect 9858 26256 9864 26308
rect 9916 26296 9922 26308
rect 10704 26296 10732 26336
rect 11698 26324 11704 26376
rect 11756 26324 11762 26376
rect 12621 26367 12679 26373
rect 12621 26364 12633 26367
rect 12268 26336 12633 26364
rect 9916 26268 10732 26296
rect 9916 26256 9922 26268
rect 5166 26188 5172 26240
rect 5224 26228 5230 26240
rect 6546 26228 6552 26240
rect 5224 26200 6552 26228
rect 5224 26188 5230 26200
rect 6546 26188 6552 26200
rect 6604 26188 6610 26240
rect 6822 26188 6828 26240
rect 6880 26228 6886 26240
rect 7374 26228 7380 26240
rect 6880 26200 7380 26228
rect 6880 26188 6886 26200
rect 7374 26188 7380 26200
rect 7432 26188 7438 26240
rect 9582 26188 9588 26240
rect 9640 26228 9646 26240
rect 12268 26228 12296 26336
rect 12621 26333 12633 26336
rect 12667 26333 12679 26367
rect 13262 26364 13268 26376
rect 12912 26343 13268 26364
rect 12879 26337 13268 26343
rect 12879 26334 12891 26337
rect 12621 26327 12679 26333
rect 12526 26256 12532 26308
rect 12584 26296 12590 26308
rect 12820 26306 12891 26334
rect 12820 26296 12848 26306
rect 12879 26303 12891 26306
rect 12925 26336 13268 26337
rect 12925 26306 12940 26336
rect 13262 26324 13268 26336
rect 13320 26324 13326 26376
rect 12925 26303 12937 26306
rect 12879 26297 12937 26303
rect 12584 26268 12848 26296
rect 12584 26256 12590 26268
rect 9640 26200 12296 26228
rect 9640 26188 9646 26200
rect 1104 26138 14696 26160
rect 1104 26086 4308 26138
rect 4360 26086 4372 26138
rect 4424 26086 4436 26138
rect 4488 26086 4500 26138
rect 4552 26086 4564 26138
rect 4616 26086 7666 26138
rect 7718 26086 7730 26138
rect 7782 26086 7794 26138
rect 7846 26086 7858 26138
rect 7910 26086 7922 26138
rect 7974 26086 11024 26138
rect 11076 26086 11088 26138
rect 11140 26086 11152 26138
rect 11204 26086 11216 26138
rect 11268 26086 11280 26138
rect 11332 26086 14382 26138
rect 14434 26086 14446 26138
rect 14498 26086 14510 26138
rect 14562 26086 14574 26138
rect 14626 26086 14638 26138
rect 14690 26086 14696 26138
rect 1104 26064 14696 26086
rect 8662 26024 8668 26036
rect 8128 25996 8668 26024
rect 6914 25916 6920 25968
rect 6972 25956 6978 25968
rect 6972 25928 7052 25956
rect 6972 25916 6978 25928
rect 7024 25888 7052 25928
rect 7175 25921 7233 25927
rect 7175 25888 7187 25921
rect 7024 25887 7187 25888
rect 7221 25918 7233 25921
rect 7221 25888 7236 25918
rect 8128 25888 8156 25996
rect 8662 25984 8668 25996
rect 8720 25984 8726 26036
rect 10042 26024 10048 26036
rect 8772 25996 10048 26024
rect 8772 25956 8800 25996
rect 10042 25984 10048 25996
rect 10100 25984 10106 26036
rect 10410 25984 10416 26036
rect 10468 25984 10474 26036
rect 13630 25984 13636 26036
rect 13688 26024 13694 26036
rect 14185 26027 14243 26033
rect 14185 26024 14197 26027
rect 13688 25996 14197 26024
rect 13688 25984 13694 25996
rect 14185 25993 14197 25996
rect 14231 25993 14243 26027
rect 14185 25987 14243 25993
rect 10226 25956 10232 25968
rect 8588 25928 8800 25956
rect 9692 25928 10232 25956
rect 8588 25927 8616 25928
rect 7221 25887 8156 25888
rect 7024 25860 8156 25887
rect 8555 25921 8616 25927
rect 8555 25887 8567 25921
rect 8601 25890 8616 25921
rect 9692 25897 9720 25928
rect 10226 25916 10232 25928
rect 10284 25916 10290 25968
rect 9677 25891 9735 25897
rect 8601 25887 8613 25890
rect 8555 25881 8613 25887
rect 9677 25857 9689 25891
rect 9723 25857 9735 25891
rect 9677 25851 9735 25857
rect 9951 25891 10009 25897
rect 9951 25857 9963 25891
rect 9997 25888 10009 25891
rect 10428 25888 10456 25984
rect 12250 25916 12256 25968
rect 12308 25956 12314 25968
rect 12308 25928 12572 25956
rect 12308 25916 12314 25928
rect 9997 25860 10456 25888
rect 9997 25857 10009 25860
rect 9951 25851 10009 25857
rect 11606 25848 11612 25900
rect 11664 25848 11670 25900
rect 12066 25848 12072 25900
rect 12124 25888 12130 25900
rect 12434 25888 12440 25900
rect 12124 25860 12440 25888
rect 12124 25848 12130 25860
rect 12434 25848 12440 25860
rect 12492 25848 12498 25900
rect 12544 25888 12572 25928
rect 12544 25860 12652 25888
rect 6917 25823 6975 25829
rect 6917 25789 6929 25823
rect 6963 25789 6975 25823
rect 8297 25823 8355 25829
rect 8297 25820 8309 25823
rect 6917 25783 6975 25789
rect 8220 25792 8309 25820
rect 6454 25644 6460 25696
rect 6512 25684 6518 25696
rect 6932 25684 6960 25783
rect 8220 25764 8248 25792
rect 8297 25789 8309 25792
rect 8343 25789 8355 25823
rect 8297 25783 8355 25789
rect 12342 25780 12348 25832
rect 12400 25780 12406 25832
rect 12452 25820 12480 25848
rect 12529 25823 12587 25829
rect 12529 25820 12541 25823
rect 12452 25792 12541 25820
rect 12529 25789 12541 25792
rect 12575 25789 12587 25823
rect 12624 25820 12652 25860
rect 13262 25848 13268 25900
rect 13320 25848 13326 25900
rect 13382 25823 13440 25829
rect 13382 25820 13394 25823
rect 12624 25792 13394 25820
rect 12529 25783 12587 25789
rect 13382 25789 13394 25792
rect 13428 25789 13440 25823
rect 13382 25783 13440 25789
rect 13538 25780 13544 25832
rect 13596 25780 13602 25832
rect 8202 25752 8208 25764
rect 7576 25724 8208 25752
rect 7576 25684 7604 25724
rect 8202 25712 8208 25724
rect 8260 25712 8266 25764
rect 9582 25752 9588 25764
rect 8956 25724 9588 25752
rect 6512 25656 7604 25684
rect 6512 25644 6518 25656
rect 7926 25644 7932 25696
rect 7984 25644 7990 25696
rect 8220 25684 8248 25712
rect 8956 25684 8984 25724
rect 9582 25712 9588 25724
rect 9640 25752 9646 25764
rect 11146 25752 11152 25764
rect 9640 25724 9812 25752
rect 9640 25712 9646 25724
rect 8220 25656 8984 25684
rect 9309 25687 9367 25693
rect 9309 25653 9321 25687
rect 9355 25684 9367 25687
rect 9674 25684 9680 25696
rect 9355 25656 9680 25684
rect 9355 25653 9367 25656
rect 9309 25647 9367 25653
rect 9674 25644 9680 25656
rect 9732 25644 9738 25696
rect 9784 25684 9812 25724
rect 10612 25724 11152 25752
rect 10612 25684 10640 25724
rect 11146 25712 11152 25724
rect 11204 25712 11210 25764
rect 12618 25712 12624 25764
rect 12676 25752 12682 25764
rect 12969 25755 13027 25761
rect 12969 25752 12981 25755
rect 12676 25724 12981 25752
rect 12676 25712 12682 25724
rect 12969 25721 12981 25724
rect 13015 25721 13027 25755
rect 12969 25715 13027 25721
rect 9784 25656 10640 25684
rect 10686 25644 10692 25696
rect 10744 25644 10750 25696
rect 11882 25644 11888 25696
rect 11940 25644 11946 25696
rect 12802 25644 12808 25696
rect 12860 25684 12866 25696
rect 13262 25684 13268 25696
rect 12860 25656 13268 25684
rect 12860 25644 12866 25656
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 1104 25594 14536 25616
rect 1104 25542 2629 25594
rect 2681 25542 2693 25594
rect 2745 25542 2757 25594
rect 2809 25542 2821 25594
rect 2873 25542 2885 25594
rect 2937 25542 5987 25594
rect 6039 25542 6051 25594
rect 6103 25542 6115 25594
rect 6167 25542 6179 25594
rect 6231 25542 6243 25594
rect 6295 25542 9345 25594
rect 9397 25542 9409 25594
rect 9461 25542 9473 25594
rect 9525 25542 9537 25594
rect 9589 25542 9601 25594
rect 9653 25542 12703 25594
rect 12755 25542 12767 25594
rect 12819 25542 12831 25594
rect 12883 25542 12895 25594
rect 12947 25542 12959 25594
rect 13011 25542 14536 25594
rect 1104 25520 14536 25542
rect 7469 25483 7527 25489
rect 7469 25449 7481 25483
rect 7515 25480 7527 25483
rect 7558 25480 7564 25492
rect 7515 25452 7564 25480
rect 7515 25449 7527 25452
rect 7469 25443 7527 25449
rect 7558 25440 7564 25452
rect 7616 25440 7622 25492
rect 7926 25440 7932 25492
rect 7984 25440 7990 25492
rect 10781 25483 10839 25489
rect 10781 25449 10793 25483
rect 10827 25480 10839 25483
rect 11422 25480 11428 25492
rect 10827 25452 11428 25480
rect 10827 25449 10839 25452
rect 10781 25443 10839 25449
rect 11422 25440 11428 25452
rect 11480 25440 11486 25492
rect 11606 25440 11612 25492
rect 11664 25480 11670 25492
rect 12345 25483 12403 25489
rect 11664 25452 12020 25480
rect 11664 25440 11670 25452
rect 7944 25412 7972 25440
rect 9585 25415 9643 25421
rect 9585 25412 9597 25415
rect 7944 25384 9597 25412
rect 9585 25381 9597 25384
rect 9631 25381 9643 25415
rect 11992 25412 12020 25452
rect 12345 25449 12357 25483
rect 12391 25480 12403 25483
rect 12618 25480 12624 25492
rect 12391 25452 12624 25480
rect 12391 25449 12403 25452
rect 12345 25443 12403 25449
rect 12618 25440 12624 25452
rect 12676 25440 12682 25492
rect 14090 25412 14096 25424
rect 11992 25384 14096 25412
rect 9585 25375 9643 25381
rect 14090 25372 14096 25384
rect 14148 25372 14154 25424
rect 1673 25347 1731 25353
rect 1673 25313 1685 25347
rect 1719 25344 1731 25347
rect 4890 25344 4896 25356
rect 1719 25316 4896 25344
rect 1719 25313 1731 25316
rect 1673 25307 1731 25313
rect 4890 25304 4896 25316
rect 4948 25304 4954 25356
rect 6454 25304 6460 25356
rect 6512 25304 6518 25356
rect 7558 25304 7564 25356
rect 7616 25344 7622 25356
rect 9125 25347 9183 25353
rect 9125 25344 9137 25347
rect 7616 25316 9137 25344
rect 7616 25304 7622 25316
rect 9125 25313 9137 25316
rect 9171 25313 9183 25347
rect 9125 25307 9183 25313
rect 9858 25304 9864 25356
rect 9916 25304 9922 25356
rect 10962 25344 10968 25356
rect 10152 25316 10968 25344
rect 750 25236 756 25288
rect 808 25276 814 25288
rect 1397 25279 1455 25285
rect 1397 25276 1409 25279
rect 808 25248 1409 25276
rect 808 25236 814 25248
rect 1397 25245 1409 25248
rect 1443 25245 1455 25279
rect 1397 25239 1455 25245
rect 5718 25236 5724 25288
rect 5776 25276 5782 25288
rect 6699 25279 6757 25285
rect 6699 25276 6711 25279
rect 5776 25248 6711 25276
rect 5776 25236 5782 25248
rect 6699 25245 6711 25248
rect 6745 25276 6757 25279
rect 6745 25248 6868 25276
rect 6745 25245 6757 25248
rect 6699 25239 6757 25245
rect 6840 25140 6868 25248
rect 8938 25236 8944 25288
rect 8996 25236 9002 25288
rect 9950 25236 9956 25288
rect 10008 25285 10014 25288
rect 10152 25285 10180 25316
rect 10962 25304 10968 25316
rect 11020 25304 11026 25356
rect 11146 25304 11152 25356
rect 11204 25344 11210 25356
rect 11333 25347 11391 25353
rect 11333 25344 11345 25347
rect 11204 25316 11345 25344
rect 11204 25304 11210 25316
rect 11333 25313 11345 25316
rect 11379 25313 11391 25347
rect 11333 25307 11391 25313
rect 13081 25347 13139 25353
rect 13081 25313 13093 25347
rect 13127 25344 13139 25347
rect 14182 25344 14188 25356
rect 13127 25316 14188 25344
rect 13127 25313 13139 25316
rect 13081 25307 13139 25313
rect 10008 25279 10036 25285
rect 10024 25245 10036 25279
rect 10008 25239 10036 25245
rect 10137 25279 10195 25285
rect 10137 25245 10149 25279
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 10008 25238 10021 25239
rect 10008 25236 10014 25238
rect 10410 25140 10416 25152
rect 6840 25112 10416 25140
rect 10410 25100 10416 25112
rect 10468 25100 10474 25152
rect 11348 25140 11376 25307
rect 14182 25304 14188 25316
rect 14240 25304 14246 25356
rect 11575 25279 11633 25285
rect 11575 25276 11587 25279
rect 11440 25248 11587 25276
rect 11440 25220 11468 25248
rect 11575 25245 11587 25248
rect 11621 25276 11633 25279
rect 11621 25248 11928 25276
rect 11621 25245 11633 25248
rect 11575 25239 11633 25245
rect 11900 25220 11928 25248
rect 11422 25168 11428 25220
rect 11480 25168 11486 25220
rect 11882 25168 11888 25220
rect 11940 25168 11946 25220
rect 12802 25168 12808 25220
rect 12860 25168 12866 25220
rect 13078 25168 13084 25220
rect 13136 25208 13142 25220
rect 13541 25211 13599 25217
rect 13541 25208 13553 25211
rect 13136 25180 13553 25208
rect 13136 25168 13142 25180
rect 13541 25177 13553 25180
rect 13587 25177 13599 25211
rect 13541 25171 13599 25177
rect 11606 25140 11612 25152
rect 11348 25112 11612 25140
rect 11606 25100 11612 25112
rect 11664 25100 11670 25152
rect 13814 25100 13820 25152
rect 13872 25100 13878 25152
rect 1104 25050 14696 25072
rect 1104 24998 4308 25050
rect 4360 24998 4372 25050
rect 4424 24998 4436 25050
rect 4488 24998 4500 25050
rect 4552 24998 4564 25050
rect 4616 24998 7666 25050
rect 7718 24998 7730 25050
rect 7782 24998 7794 25050
rect 7846 24998 7858 25050
rect 7910 24998 7922 25050
rect 7974 24998 11024 25050
rect 11076 24998 11088 25050
rect 11140 24998 11152 25050
rect 11204 24998 11216 25050
rect 11268 24998 11280 25050
rect 11332 24998 14382 25050
rect 14434 24998 14446 25050
rect 14498 24998 14510 25050
rect 14562 24998 14574 25050
rect 14626 24998 14638 25050
rect 14690 24998 14696 25050
rect 1104 24976 14696 24998
rect 7650 24896 7656 24948
rect 7708 24936 7714 24948
rect 8202 24936 8208 24948
rect 7708 24908 8208 24936
rect 7708 24896 7714 24908
rect 8202 24896 8208 24908
rect 8260 24896 8266 24948
rect 8662 24896 8668 24948
rect 8720 24936 8726 24948
rect 9582 24936 9588 24948
rect 8720 24908 9588 24936
rect 8720 24896 8726 24908
rect 9582 24896 9588 24908
rect 9640 24896 9646 24948
rect 13449 24939 13507 24945
rect 13449 24905 13461 24939
rect 13495 24936 13507 24939
rect 13538 24936 13544 24948
rect 13495 24908 13544 24936
rect 13495 24905 13507 24908
rect 13449 24899 13507 24905
rect 13538 24896 13544 24908
rect 13596 24896 13602 24948
rect 6730 24868 6736 24880
rect 6654 24840 6736 24868
rect 6654 24839 6682 24840
rect 6623 24833 6682 24839
rect 750 24760 756 24812
rect 808 24800 814 24812
rect 1489 24803 1547 24809
rect 1489 24800 1501 24803
rect 808 24772 1501 24800
rect 808 24760 814 24772
rect 1489 24769 1501 24772
rect 1535 24769 1547 24803
rect 6623 24799 6635 24833
rect 6669 24802 6682 24833
rect 6730 24828 6736 24840
rect 6788 24868 6794 24880
rect 7006 24868 7012 24880
rect 6788 24840 7012 24868
rect 6788 24828 6794 24840
rect 7006 24828 7012 24840
rect 7064 24828 7070 24880
rect 12406 24840 12848 24868
rect 6669 24799 6681 24802
rect 6623 24793 6681 24799
rect 1489 24763 1547 24769
rect 10410 24760 10416 24812
rect 10468 24760 10474 24812
rect 10962 24760 10968 24812
rect 11020 24760 11026 24812
rect 11333 24803 11391 24809
rect 11333 24769 11345 24803
rect 11379 24769 11391 24803
rect 11333 24763 11391 24769
rect 11977 24803 12035 24809
rect 11977 24769 11989 24803
rect 12023 24800 12035 24803
rect 12158 24800 12164 24812
rect 12023 24772 12164 24800
rect 12023 24769 12035 24772
rect 11977 24763 12035 24769
rect 4154 24692 4160 24744
rect 4212 24732 4218 24744
rect 6365 24735 6423 24741
rect 6365 24732 6377 24735
rect 4212 24704 6377 24732
rect 4212 24692 4218 24704
rect 6365 24701 6377 24704
rect 6411 24701 6423 24735
rect 11348 24732 11376 24763
rect 12158 24760 12164 24772
rect 12216 24760 12222 24812
rect 12406 24800 12434 24840
rect 12710 24800 12716 24812
rect 12268 24772 12434 24800
rect 12671 24772 12716 24800
rect 12268 24732 12296 24772
rect 12710 24760 12716 24772
rect 12768 24760 12774 24812
rect 12820 24800 12848 24840
rect 14090 24828 14096 24880
rect 14148 24868 14154 24880
rect 15010 24868 15016 24880
rect 14148 24840 15016 24868
rect 14148 24828 14154 24840
rect 15010 24828 15016 24840
rect 15068 24828 15074 24880
rect 14274 24800 14280 24812
rect 12820 24772 14280 24800
rect 14274 24760 14280 24772
rect 14332 24760 14338 24812
rect 15194 24760 15200 24812
rect 15252 24800 15258 24812
rect 15562 24800 15568 24812
rect 15252 24772 15568 24800
rect 15252 24760 15258 24772
rect 15562 24760 15568 24772
rect 15620 24760 15626 24812
rect 11348 24704 12296 24732
rect 12440 24735 12498 24741
rect 6365 24695 6423 24701
rect 12440 24701 12452 24735
rect 12486 24701 12498 24735
rect 12440 24695 12498 24701
rect 1673 24667 1731 24673
rect 1673 24633 1685 24667
rect 1719 24664 1731 24667
rect 5718 24664 5724 24676
rect 1719 24636 5724 24664
rect 1719 24633 1731 24636
rect 1673 24627 1731 24633
rect 5718 24624 5724 24636
rect 5776 24624 5782 24676
rect 6380 24596 6408 24695
rect 7466 24664 7472 24676
rect 7300 24636 7472 24664
rect 7300 24596 7328 24636
rect 7466 24624 7472 24636
rect 7524 24624 7530 24676
rect 11606 24624 11612 24676
rect 11664 24664 11670 24676
rect 12452 24664 12480 24695
rect 11664 24636 12480 24664
rect 11664 24624 11670 24636
rect 6380 24568 7328 24596
rect 7374 24556 7380 24608
rect 7432 24556 7438 24608
rect 7558 24556 7564 24608
rect 7616 24596 7622 24608
rect 7742 24596 7748 24608
rect 7616 24568 7748 24596
rect 7616 24556 7622 24568
rect 7742 24556 7748 24568
rect 7800 24556 7806 24608
rect 10689 24599 10747 24605
rect 10689 24565 10701 24599
rect 10735 24596 10747 24599
rect 11422 24596 11428 24608
rect 10735 24568 11428 24596
rect 10735 24565 10747 24568
rect 10689 24559 10747 24565
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 12253 24599 12311 24605
rect 12253 24565 12265 24599
rect 12299 24596 12311 24599
rect 13998 24596 14004 24608
rect 12299 24568 14004 24596
rect 12299 24565 12311 24568
rect 12253 24559 12311 24565
rect 13998 24556 14004 24568
rect 14056 24556 14062 24608
rect 1104 24506 14536 24528
rect 1104 24454 2629 24506
rect 2681 24454 2693 24506
rect 2745 24454 2757 24506
rect 2809 24454 2821 24506
rect 2873 24454 2885 24506
rect 2937 24454 5987 24506
rect 6039 24454 6051 24506
rect 6103 24454 6115 24506
rect 6167 24454 6179 24506
rect 6231 24454 6243 24506
rect 6295 24454 9345 24506
rect 9397 24454 9409 24506
rect 9461 24454 9473 24506
rect 9525 24454 9537 24506
rect 9589 24454 9601 24506
rect 9653 24454 12703 24506
rect 12755 24454 12767 24506
rect 12819 24454 12831 24506
rect 12883 24454 12895 24506
rect 12947 24454 12959 24506
rect 13011 24454 14536 24506
rect 1104 24432 14536 24454
rect 5810 24352 5816 24404
rect 5868 24392 5874 24404
rect 6270 24392 6276 24404
rect 5868 24364 6276 24392
rect 5868 24352 5874 24364
rect 6270 24352 6276 24364
rect 6328 24392 6334 24404
rect 6328 24364 6592 24392
rect 6328 24352 6334 24364
rect 5445 24327 5503 24333
rect 5445 24293 5457 24327
rect 5491 24324 5503 24327
rect 6457 24327 6515 24333
rect 6457 24324 6469 24327
rect 5491 24296 6469 24324
rect 5491 24293 5503 24296
rect 5445 24287 5503 24293
rect 6457 24293 6469 24296
rect 6503 24293 6515 24327
rect 6457 24287 6515 24293
rect 4154 24216 4160 24268
rect 4212 24256 4218 24268
rect 4433 24259 4491 24265
rect 4433 24256 4445 24259
rect 4212 24228 4445 24256
rect 4212 24216 4218 24228
rect 4433 24225 4445 24228
rect 4479 24225 4491 24259
rect 4433 24219 4491 24225
rect 5994 24216 6000 24268
rect 6052 24216 6058 24268
rect 6564 24256 6592 24364
rect 7374 24352 7380 24404
rect 7432 24352 7438 24404
rect 7466 24352 7472 24404
rect 7524 24352 7530 24404
rect 7653 24395 7711 24401
rect 7653 24361 7665 24395
rect 7699 24392 7711 24395
rect 10410 24392 10416 24404
rect 7699 24364 10416 24392
rect 7699 24361 7711 24364
rect 7653 24355 7711 24361
rect 10410 24352 10416 24364
rect 10468 24352 10474 24404
rect 10520 24364 11192 24392
rect 6733 24259 6791 24265
rect 6733 24256 6745 24259
rect 6564 24228 6745 24256
rect 6733 24225 6745 24228
rect 6779 24225 6791 24259
rect 6733 24219 6791 24225
rect 7009 24259 7067 24265
rect 7009 24225 7021 24259
rect 7055 24256 7067 24259
rect 7392 24256 7420 24352
rect 7055 24228 7420 24256
rect 7484 24256 7512 24352
rect 9950 24284 9956 24336
rect 10008 24284 10014 24336
rect 10520 24265 10548 24364
rect 8941 24259 8999 24265
rect 8941 24256 8953 24259
rect 7484 24228 8953 24256
rect 7055 24225 7067 24228
rect 7009 24219 7067 24225
rect 8941 24225 8953 24228
rect 8987 24225 8999 24259
rect 10505 24259 10563 24265
rect 10505 24256 10517 24259
rect 8941 24219 8999 24225
rect 9968 24228 10517 24256
rect 4706 24188 4712 24200
rect 4667 24160 4712 24188
rect 4706 24148 4712 24160
rect 4764 24188 4770 24200
rect 5442 24188 5448 24200
rect 4764 24160 5448 24188
rect 4764 24148 4770 24160
rect 5442 24148 5448 24160
rect 5500 24148 5506 24200
rect 5813 24191 5871 24197
rect 5813 24157 5825 24191
rect 5859 24188 5871 24191
rect 5902 24188 5908 24200
rect 5859 24160 5908 24188
rect 5859 24157 5871 24160
rect 5813 24151 5871 24157
rect 5902 24148 5908 24160
rect 5960 24188 5966 24200
rect 6178 24188 6184 24200
rect 5960 24160 6184 24188
rect 5960 24148 5966 24160
rect 6178 24148 6184 24160
rect 6236 24148 6242 24200
rect 6822 24148 6828 24200
rect 6880 24197 6886 24200
rect 6880 24191 6908 24197
rect 6896 24157 6908 24191
rect 6880 24151 6908 24157
rect 6880 24148 6886 24151
rect 8956 24120 8984 24219
rect 9122 24148 9128 24200
rect 9180 24188 9186 24200
rect 9215 24191 9273 24197
rect 9215 24188 9227 24191
rect 9180 24160 9227 24188
rect 9180 24148 9186 24160
rect 9215 24157 9227 24160
rect 9261 24157 9273 24191
rect 9215 24151 9273 24157
rect 9968 24120 9996 24228
rect 10505 24225 10517 24228
rect 10551 24225 10563 24259
rect 11164 24256 11192 24364
rect 12158 24352 12164 24404
rect 12216 24392 12222 24404
rect 15470 24392 15476 24404
rect 12216 24364 15476 24392
rect 12216 24352 12222 24364
rect 15470 24352 15476 24364
rect 15528 24352 15534 24404
rect 11885 24259 11943 24265
rect 11885 24256 11897 24259
rect 11164 24228 11897 24256
rect 10505 24219 10563 24225
rect 11885 24225 11897 24228
rect 11931 24225 11943 24259
rect 11885 24219 11943 24225
rect 10042 24148 10048 24200
rect 10100 24188 10106 24200
rect 11790 24188 11796 24200
rect 10100 24161 10824 24188
rect 10100 24160 10775 24161
rect 10100 24148 10106 24160
rect 10226 24120 10232 24132
rect 8956 24092 10232 24120
rect 10226 24080 10232 24092
rect 10284 24080 10290 24132
rect 10763 24127 10775 24160
rect 10809 24130 10824 24161
rect 10888 24160 11796 24188
rect 10809 24127 10821 24130
rect 10763 24121 10821 24127
rect 5534 24012 5540 24064
rect 5592 24052 5598 24064
rect 5902 24052 5908 24064
rect 5592 24024 5908 24052
rect 5592 24012 5598 24024
rect 5902 24012 5908 24024
rect 5960 24012 5966 24064
rect 5994 24012 6000 24064
rect 6052 24052 6058 24064
rect 6362 24052 6368 24064
rect 6052 24024 6368 24052
rect 6052 24012 6058 24024
rect 6362 24012 6368 24024
rect 6420 24052 6426 24064
rect 6730 24052 6736 24064
rect 6420 24024 6736 24052
rect 6420 24012 6426 24024
rect 6730 24012 6736 24024
rect 6788 24012 6794 24064
rect 7466 24012 7472 24064
rect 7524 24052 7530 24064
rect 10888 24052 10916 24160
rect 11790 24148 11796 24160
rect 11848 24188 11854 24200
rect 12127 24191 12185 24197
rect 12127 24188 12139 24191
rect 11848 24160 12139 24188
rect 11848 24148 11854 24160
rect 12127 24157 12139 24160
rect 12173 24157 12185 24191
rect 14090 24188 14096 24200
rect 12127 24151 12185 24157
rect 13372 24160 14096 24188
rect 10962 24080 10968 24132
rect 11020 24120 11026 24132
rect 13372 24129 13400 24160
rect 14090 24148 14096 24160
rect 14148 24148 14154 24200
rect 13357 24123 13415 24129
rect 11020 24092 13308 24120
rect 11020 24080 11026 24092
rect 7524 24024 10916 24052
rect 11517 24055 11575 24061
rect 7524 24012 7530 24024
rect 11517 24021 11529 24055
rect 11563 24052 11575 24055
rect 11790 24052 11796 24064
rect 11563 24024 11796 24052
rect 11563 24021 11575 24024
rect 11517 24015 11575 24021
rect 11790 24012 11796 24024
rect 11848 24012 11854 24064
rect 12894 24012 12900 24064
rect 12952 24012 12958 24064
rect 13280 24052 13308 24092
rect 13357 24089 13369 24123
rect 13403 24089 13415 24123
rect 13357 24083 13415 24089
rect 13722 24080 13728 24132
rect 13780 24080 13786 24132
rect 14182 24052 14188 24064
rect 13280 24024 14188 24052
rect 14182 24012 14188 24024
rect 14240 24012 14246 24064
rect 1104 23962 14696 23984
rect 1104 23910 4308 23962
rect 4360 23910 4372 23962
rect 4424 23910 4436 23962
rect 4488 23910 4500 23962
rect 4552 23910 4564 23962
rect 4616 23910 7666 23962
rect 7718 23910 7730 23962
rect 7782 23910 7794 23962
rect 7846 23910 7858 23962
rect 7910 23910 7922 23962
rect 7974 23910 11024 23962
rect 11076 23910 11088 23962
rect 11140 23910 11152 23962
rect 11204 23910 11216 23962
rect 11268 23910 11280 23962
rect 11332 23910 14382 23962
rect 14434 23910 14446 23962
rect 14498 23910 14510 23962
rect 14562 23910 14574 23962
rect 14626 23910 14638 23962
rect 14690 23910 14696 23962
rect 1104 23888 14696 23910
rect 3510 23808 3516 23860
rect 3568 23848 3574 23860
rect 7466 23848 7472 23860
rect 3568 23820 7472 23848
rect 3568 23808 3574 23820
rect 7466 23808 7472 23820
rect 7524 23808 7530 23860
rect 9214 23808 9220 23860
rect 9272 23808 9278 23860
rect 9674 23808 9680 23860
rect 9732 23848 9738 23860
rect 12161 23851 12219 23857
rect 9732 23820 10166 23848
rect 9732 23808 9738 23820
rect 10138 23731 10166 23820
rect 12161 23817 12173 23851
rect 12207 23848 12219 23851
rect 13998 23848 14004 23860
rect 12207 23820 14004 23848
rect 12207 23817 12219 23820
rect 12161 23811 12219 23817
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 14182 23808 14188 23860
rect 14240 23808 14246 23860
rect 10410 23740 10416 23792
rect 10468 23740 10474 23792
rect 10778 23740 10784 23792
rect 10836 23780 10842 23792
rect 11885 23783 11943 23789
rect 11885 23780 11897 23783
rect 10836 23752 11897 23780
rect 10836 23740 10842 23752
rect 11885 23749 11897 23752
rect 11931 23749 11943 23783
rect 11885 23743 11943 23749
rect 10103 23725 10166 23731
rect 750 23672 756 23724
rect 808 23712 814 23724
rect 1489 23715 1547 23721
rect 1489 23712 1501 23715
rect 808 23684 1501 23712
rect 808 23672 814 23684
rect 1489 23681 1501 23684
rect 1535 23681 1547 23715
rect 1489 23675 1547 23681
rect 7558 23672 7564 23724
rect 7616 23672 7622 23724
rect 10103 23691 10115 23725
rect 10149 23694 10166 23725
rect 10428 23712 10456 23740
rect 12250 23712 12256 23724
rect 10149 23691 10161 23694
rect 10103 23685 10161 23691
rect 10428 23684 12256 23712
rect 12250 23672 12256 23684
rect 12308 23712 12314 23724
rect 13446 23721 13452 23724
rect 12345 23715 12403 23721
rect 12345 23712 12357 23715
rect 12308 23684 12357 23712
rect 12308 23672 12314 23684
rect 12345 23681 12357 23684
rect 12391 23681 12403 23715
rect 12345 23675 12403 23681
rect 13403 23715 13452 23721
rect 13403 23681 13415 23715
rect 13449 23681 13452 23715
rect 13403 23675 13452 23681
rect 13446 23672 13452 23675
rect 13504 23672 13510 23724
rect 5166 23604 5172 23656
rect 5224 23644 5230 23656
rect 7377 23647 7435 23653
rect 7377 23644 7389 23647
rect 5224 23616 7389 23644
rect 5224 23604 5230 23616
rect 7377 23613 7389 23616
rect 7423 23613 7435 23647
rect 7377 23607 7435 23613
rect 8294 23604 8300 23656
rect 8352 23604 8358 23656
rect 8478 23653 8484 23656
rect 8435 23647 8484 23653
rect 8435 23613 8447 23647
rect 8481 23613 8484 23647
rect 8435 23607 8484 23613
rect 8478 23604 8484 23607
rect 8536 23604 8542 23656
rect 8573 23647 8631 23653
rect 8573 23613 8585 23647
rect 8619 23644 8631 23647
rect 8754 23644 8760 23656
rect 8619 23616 8760 23644
rect 8619 23613 8631 23616
rect 8573 23607 8631 23613
rect 8754 23604 8760 23616
rect 8812 23604 8818 23656
rect 9674 23604 9680 23656
rect 9732 23644 9738 23656
rect 9861 23647 9919 23653
rect 9861 23644 9873 23647
rect 9732 23616 9873 23644
rect 9732 23604 9738 23616
rect 9861 23613 9873 23616
rect 9907 23613 9919 23647
rect 12529 23647 12587 23653
rect 12529 23644 12541 23647
rect 9861 23607 9919 23613
rect 12406 23616 12541 23644
rect 1673 23579 1731 23585
rect 1673 23545 1685 23579
rect 1719 23576 1731 23579
rect 5074 23576 5080 23588
rect 1719 23548 5080 23576
rect 1719 23545 1731 23548
rect 1673 23539 1731 23545
rect 5074 23536 5080 23548
rect 5132 23536 5138 23588
rect 7834 23536 7840 23588
rect 7892 23576 7898 23588
rect 8021 23579 8079 23585
rect 8021 23576 8033 23579
rect 7892 23548 8033 23576
rect 7892 23536 7898 23548
rect 8021 23545 8033 23548
rect 8067 23545 8079 23579
rect 8021 23539 8079 23545
rect 12406 23520 12434 23616
rect 12529 23613 12541 23616
rect 12575 23613 12587 23647
rect 12529 23607 12587 23613
rect 12894 23604 12900 23656
rect 12952 23644 12958 23656
rect 12989 23647 13047 23653
rect 12989 23644 13001 23647
rect 12952 23616 13001 23644
rect 12952 23604 12958 23616
rect 12989 23613 13001 23616
rect 13035 23613 13047 23647
rect 12989 23607 13047 23613
rect 13262 23604 13268 23656
rect 13320 23604 13326 23656
rect 13538 23604 13544 23656
rect 13596 23604 13602 23656
rect 6178 23468 6184 23520
rect 6236 23508 6242 23520
rect 8478 23508 8484 23520
rect 6236 23480 8484 23508
rect 6236 23468 6242 23480
rect 8478 23468 8484 23480
rect 8536 23508 8542 23520
rect 10226 23508 10232 23520
rect 8536 23480 10232 23508
rect 8536 23468 8542 23480
rect 10226 23468 10232 23480
rect 10284 23468 10290 23520
rect 10873 23511 10931 23517
rect 10873 23477 10885 23511
rect 10919 23508 10931 23511
rect 11054 23508 11060 23520
rect 10919 23480 11060 23508
rect 10919 23477 10931 23480
rect 10873 23471 10931 23477
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 12158 23468 12164 23520
rect 12216 23508 12222 23520
rect 12342 23508 12348 23520
rect 12216 23480 12348 23508
rect 12216 23468 12222 23480
rect 12342 23468 12348 23480
rect 12400 23480 12434 23520
rect 12400 23468 12406 23480
rect 1104 23418 14536 23440
rect 1104 23366 2629 23418
rect 2681 23366 2693 23418
rect 2745 23366 2757 23418
rect 2809 23366 2821 23418
rect 2873 23366 2885 23418
rect 2937 23366 5987 23418
rect 6039 23366 6051 23418
rect 6103 23366 6115 23418
rect 6167 23366 6179 23418
rect 6231 23366 6243 23418
rect 6295 23366 9345 23418
rect 9397 23366 9409 23418
rect 9461 23366 9473 23418
rect 9525 23366 9537 23418
rect 9589 23366 9601 23418
rect 9653 23366 12703 23418
rect 12755 23366 12767 23418
rect 12819 23366 12831 23418
rect 12883 23366 12895 23418
rect 12947 23366 12959 23418
rect 13011 23366 14536 23418
rect 1104 23344 14536 23366
rect 2498 23264 2504 23316
rect 2556 23304 2562 23316
rect 11606 23304 11612 23316
rect 2556 23276 11612 23304
rect 2556 23264 2562 23276
rect 11606 23264 11612 23276
rect 11664 23264 11670 23316
rect 12437 23307 12495 23313
rect 12437 23273 12449 23307
rect 12483 23304 12495 23307
rect 13078 23304 13084 23316
rect 12483 23276 13084 23304
rect 12483 23273 12495 23276
rect 12437 23267 12495 23273
rect 13078 23264 13084 23276
rect 13136 23264 13142 23316
rect 13538 23264 13544 23316
rect 13596 23304 13602 23316
rect 13633 23307 13691 23313
rect 13633 23304 13645 23307
rect 13596 23276 13645 23304
rect 13596 23264 13602 23276
rect 13633 23273 13645 23276
rect 13679 23273 13691 23307
rect 13633 23267 13691 23273
rect 8389 23239 8447 23245
rect 8389 23205 8401 23239
rect 8435 23236 8447 23239
rect 8754 23236 8760 23248
rect 8435 23208 8760 23236
rect 8435 23205 8447 23208
rect 8389 23199 8447 23205
rect 8754 23196 8760 23208
rect 8812 23196 8818 23248
rect 10318 23196 10324 23248
rect 10376 23236 10382 23248
rect 10778 23236 10784 23248
rect 10376 23208 10784 23236
rect 10376 23196 10382 23208
rect 10778 23196 10784 23208
rect 10836 23196 10842 23248
rect 11054 23196 11060 23248
rect 11112 23236 11118 23248
rect 11241 23239 11299 23245
rect 11241 23236 11253 23239
rect 11112 23208 11253 23236
rect 11112 23196 11118 23208
rect 11241 23205 11253 23208
rect 11287 23205 11299 23239
rect 11241 23199 11299 23205
rect 7190 23128 7196 23180
rect 7248 23168 7254 23180
rect 7377 23171 7435 23177
rect 7377 23168 7389 23171
rect 7248 23140 7389 23168
rect 7248 23128 7254 23140
rect 7377 23137 7389 23140
rect 7423 23137 7435 23171
rect 7377 23131 7435 23137
rect 8294 23128 8300 23180
rect 8352 23168 8358 23180
rect 10870 23168 10876 23180
rect 8352 23140 10876 23168
rect 8352 23128 8358 23140
rect 10870 23128 10876 23140
rect 10928 23168 10934 23180
rect 11517 23171 11575 23177
rect 11517 23168 11529 23171
rect 10928 23140 11529 23168
rect 10928 23128 10934 23140
rect 11517 23137 11529 23140
rect 11563 23137 11575 23171
rect 11517 23131 11575 23137
rect 11655 23171 11713 23177
rect 11655 23137 11667 23171
rect 11701 23168 11713 23171
rect 12434 23168 12440 23180
rect 11701 23140 12440 23168
rect 11701 23137 11713 23140
rect 11655 23131 11713 23137
rect 12434 23128 12440 23140
rect 12492 23128 12498 23180
rect 7651 23103 7709 23109
rect 7651 23069 7663 23103
rect 7697 23100 7709 23103
rect 8202 23100 8208 23112
rect 7697 23072 8208 23100
rect 7697 23069 7709 23072
rect 7651 23063 7709 23069
rect 750 22992 756 23044
rect 808 23032 814 23044
rect 1489 23035 1547 23041
rect 1489 23032 1501 23035
rect 808 23004 1501 23032
rect 808 22992 814 23004
rect 1489 23001 1501 23004
rect 1535 23001 1547 23035
rect 1489 22995 1547 23001
rect 1673 23035 1731 23041
rect 1673 23001 1685 23035
rect 1719 23032 1731 23035
rect 1719 23004 2774 23032
rect 1719 23001 1731 23004
rect 1673 22995 1731 23001
rect 2746 22964 2774 23004
rect 7466 22992 7472 23044
rect 7524 23032 7530 23044
rect 7666 23032 7694 23063
rect 8202 23060 8208 23072
rect 8260 23060 8266 23112
rect 10502 23060 10508 23112
rect 10560 23060 10566 23112
rect 10594 23060 10600 23112
rect 10652 23060 10658 23112
rect 10781 23103 10839 23109
rect 10781 23069 10793 23103
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 7524 23004 7694 23032
rect 7524 22992 7530 23004
rect 10318 22992 10324 23044
rect 10376 23032 10382 23044
rect 10520 23032 10548 23060
rect 10796 23032 10824 23063
rect 11790 23060 11796 23112
rect 11848 23060 11854 23112
rect 12609 23103 12667 23109
rect 12609 23069 12621 23103
rect 12655 23069 12667 23103
rect 12609 23063 12667 23069
rect 12879 23073 12937 23079
rect 10376 23004 10824 23032
rect 10376 22992 10382 23004
rect 12342 22992 12348 23044
rect 12400 23032 12406 23044
rect 12624 23032 12652 23063
rect 12879 23039 12891 23073
rect 12925 23070 12937 23073
rect 12925 23039 12940 23070
rect 12879 23033 12940 23039
rect 12400 23004 12652 23032
rect 12912 23032 12940 23033
rect 13170 23032 13176 23044
rect 12912 23004 13176 23032
rect 12400 22992 12406 23004
rect 13170 22992 13176 23004
rect 13228 22992 13234 23044
rect 8386 22964 8392 22976
rect 2746 22936 8392 22964
rect 8386 22924 8392 22936
rect 8444 22924 8450 22976
rect 9030 22924 9036 22976
rect 9088 22964 9094 22976
rect 15194 22964 15200 22976
rect 9088 22936 15200 22964
rect 9088 22924 9094 22936
rect 15194 22924 15200 22936
rect 15252 22924 15258 22976
rect 1104 22874 14696 22896
rect 1104 22822 4308 22874
rect 4360 22822 4372 22874
rect 4424 22822 4436 22874
rect 4488 22822 4500 22874
rect 4552 22822 4564 22874
rect 4616 22822 7666 22874
rect 7718 22822 7730 22874
rect 7782 22822 7794 22874
rect 7846 22822 7858 22874
rect 7910 22822 7922 22874
rect 7974 22822 11024 22874
rect 11076 22822 11088 22874
rect 11140 22822 11152 22874
rect 11204 22822 11216 22874
rect 11268 22822 11280 22874
rect 11332 22822 14382 22874
rect 14434 22822 14446 22874
rect 14498 22822 14510 22874
rect 14562 22822 14574 22874
rect 14626 22822 14638 22874
rect 14690 22822 14696 22874
rect 1104 22800 14696 22822
rect 7190 22720 7196 22772
rect 7248 22720 7254 22772
rect 7837 22763 7895 22769
rect 7837 22729 7849 22763
rect 7883 22760 7895 22763
rect 8018 22760 8024 22772
rect 7883 22732 8024 22760
rect 7883 22729 7895 22732
rect 7837 22723 7895 22729
rect 8018 22720 8024 22732
rect 8076 22720 8082 22772
rect 8386 22720 8392 22772
rect 8444 22760 8450 22772
rect 10778 22760 10784 22772
rect 8444 22732 10784 22760
rect 8444 22720 8450 22732
rect 10778 22720 10784 22732
rect 10836 22760 10842 22772
rect 13354 22760 13360 22772
rect 10836 22732 13360 22760
rect 10836 22720 10842 22732
rect 13354 22720 13360 22732
rect 13412 22720 13418 22772
rect 14093 22763 14151 22769
rect 14093 22729 14105 22763
rect 14139 22760 14151 22763
rect 14918 22760 14924 22772
rect 14139 22732 14924 22760
rect 14139 22729 14151 22732
rect 14093 22723 14151 22729
rect 14918 22720 14924 22732
rect 14976 22720 14982 22772
rect 7208 22692 7236 22720
rect 9674 22692 9680 22704
rect 6840 22664 7326 22692
rect 5534 22584 5540 22636
rect 5592 22624 5598 22636
rect 6840 22633 6868 22664
rect 6825 22627 6883 22633
rect 6825 22624 6837 22627
rect 5592 22596 6837 22624
rect 5592 22584 5598 22596
rect 6825 22593 6837 22596
rect 6871 22593 6883 22627
rect 6825 22587 6883 22593
rect 7099 22627 7157 22633
rect 7099 22593 7111 22627
rect 7145 22624 7157 22627
rect 7190 22624 7196 22636
rect 7145 22596 7196 22624
rect 7145 22593 7157 22596
rect 7099 22587 7157 22593
rect 7190 22584 7196 22596
rect 7248 22584 7254 22636
rect 7298 22624 7326 22664
rect 8588 22664 9680 22692
rect 7298 22596 7445 22624
rect 7417 22556 7445 22596
rect 8588 22556 8616 22664
rect 9674 22652 9680 22664
rect 9732 22652 9738 22704
rect 11977 22695 12035 22701
rect 11977 22661 11989 22695
rect 12023 22692 12035 22695
rect 13998 22692 14004 22704
rect 12023 22664 14004 22692
rect 12023 22661 12035 22664
rect 11977 22655 12035 22661
rect 13998 22652 14004 22664
rect 14056 22652 14062 22704
rect 8662 22584 8668 22636
rect 8720 22624 8726 22636
rect 8999 22627 9057 22633
rect 8999 22624 9011 22627
rect 8720 22596 9011 22624
rect 8720 22584 8726 22596
rect 8999 22593 9011 22596
rect 9045 22593 9057 22627
rect 12618 22624 12624 22636
rect 8999 22587 9057 22593
rect 9416 22596 12624 22624
rect 8757 22559 8815 22565
rect 8757 22556 8769 22559
rect 7417 22528 8769 22556
rect 8757 22525 8769 22528
rect 8803 22525 8815 22559
rect 8757 22519 8815 22525
rect 5810 22380 5816 22432
rect 5868 22420 5874 22432
rect 9416 22420 9444 22596
rect 12618 22584 12624 22596
rect 12676 22633 12682 22636
rect 12676 22627 12737 22633
rect 12676 22593 12691 22627
rect 12725 22624 12737 22627
rect 13909 22627 13967 22633
rect 12725 22596 12769 22624
rect 12725 22593 12737 22596
rect 12676 22587 12737 22593
rect 13909 22593 13921 22627
rect 13955 22624 13967 22627
rect 15378 22624 15384 22636
rect 13955 22596 15384 22624
rect 13955 22593 13967 22596
rect 13909 22587 13967 22593
rect 12676 22584 12682 22587
rect 15378 22584 15384 22596
rect 15436 22584 15442 22636
rect 12250 22516 12256 22568
rect 12308 22556 12314 22568
rect 12437 22559 12495 22565
rect 12437 22556 12449 22559
rect 12308 22528 12449 22556
rect 12308 22516 12314 22528
rect 12437 22525 12449 22528
rect 12483 22525 12495 22559
rect 12437 22519 12495 22525
rect 14918 22516 14924 22568
rect 14976 22556 14982 22568
rect 15286 22556 15292 22568
rect 14976 22528 15292 22556
rect 14976 22516 14982 22528
rect 15286 22516 15292 22528
rect 15344 22516 15350 22568
rect 13814 22488 13820 22500
rect 13372 22460 13820 22488
rect 5868 22392 9444 22420
rect 5868 22380 5874 22392
rect 9766 22380 9772 22432
rect 9824 22380 9830 22432
rect 10226 22380 10232 22432
rect 10284 22420 10290 22432
rect 10594 22420 10600 22432
rect 10284 22392 10600 22420
rect 10284 22380 10290 22392
rect 10594 22380 10600 22392
rect 10652 22380 10658 22432
rect 12253 22423 12311 22429
rect 12253 22389 12265 22423
rect 12299 22420 12311 22423
rect 13372 22420 13400 22460
rect 13814 22448 13820 22460
rect 13872 22448 13878 22500
rect 12299 22392 13400 22420
rect 12299 22389 12311 22392
rect 12253 22383 12311 22389
rect 13446 22380 13452 22432
rect 13504 22380 13510 22432
rect 1104 22330 14536 22352
rect 1104 22278 2629 22330
rect 2681 22278 2693 22330
rect 2745 22278 2757 22330
rect 2809 22278 2821 22330
rect 2873 22278 2885 22330
rect 2937 22278 5987 22330
rect 6039 22278 6051 22330
rect 6103 22278 6115 22330
rect 6167 22278 6179 22330
rect 6231 22278 6243 22330
rect 6295 22278 9345 22330
rect 9397 22278 9409 22330
rect 9461 22278 9473 22330
rect 9525 22278 9537 22330
rect 9589 22278 9601 22330
rect 9653 22278 12703 22330
rect 12755 22278 12767 22330
rect 12819 22278 12831 22330
rect 12883 22278 12895 22330
rect 12947 22278 12959 22330
rect 13011 22278 14536 22330
rect 1104 22256 14536 22278
rect 9858 22176 9864 22228
rect 9916 22216 9922 22228
rect 9916 22188 12388 22216
rect 9916 22176 9922 22188
rect 9766 22108 9772 22160
rect 9824 22148 9830 22160
rect 10413 22151 10471 22157
rect 10413 22148 10425 22151
rect 9824 22120 10425 22148
rect 9824 22108 9830 22120
rect 10413 22117 10425 22120
rect 10459 22117 10471 22151
rect 10413 22111 10471 22117
rect 9953 22083 10011 22089
rect 9953 22080 9965 22083
rect 9324 22052 9965 22080
rect 9324 22024 9352 22052
rect 9953 22049 9965 22052
rect 9999 22049 10011 22083
rect 10134 22080 10140 22092
rect 9953 22043 10011 22049
rect 10060 22052 10140 22080
rect 4890 21972 4896 22024
rect 4948 22012 4954 22024
rect 5534 22012 5540 22024
rect 4948 21984 5540 22012
rect 4948 21972 4954 21984
rect 5534 21972 5540 21984
rect 5592 21972 5598 22024
rect 5810 22021 5816 22024
rect 5779 22015 5816 22021
rect 5779 21981 5791 22015
rect 5779 21975 5816 21981
rect 5810 21972 5816 21975
rect 5868 21972 5874 22024
rect 7006 21972 7012 22024
rect 7064 21972 7070 22024
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7374 22012 7380 22024
rect 7156 21984 7380 22012
rect 7156 21972 7162 21984
rect 7374 21972 7380 21984
rect 7432 22012 7438 22024
rect 7469 22015 7527 22021
rect 7469 22012 7481 22015
rect 7432 21984 7481 22012
rect 7432 21972 7438 21984
rect 7469 21981 7481 21984
rect 7515 21981 7527 22015
rect 7711 22015 7769 22021
rect 7711 22012 7723 22015
rect 7469 21975 7527 21981
rect 7576 21984 7723 22012
rect 750 21904 756 21956
rect 808 21944 814 21956
rect 1489 21947 1547 21953
rect 1489 21944 1501 21947
rect 808 21916 1501 21944
rect 808 21904 814 21916
rect 1489 21913 1501 21916
rect 1535 21913 1547 21947
rect 7024 21944 7052 21972
rect 7576 21956 7604 21984
rect 7711 21981 7723 21984
rect 7757 21981 7769 22015
rect 7711 21975 7769 21981
rect 8294 21972 8300 22024
rect 8352 22012 8358 22024
rect 8662 22012 8668 22024
rect 8352 21984 8668 22012
rect 8352 21972 8358 21984
rect 8662 21972 8668 21984
rect 8720 21972 8726 22024
rect 9306 21972 9312 22024
rect 9364 21972 9370 22024
rect 9766 21972 9772 22024
rect 9824 21972 9830 22024
rect 10060 22012 10088 22052
rect 10134 22040 10140 22052
rect 10192 22040 10198 22092
rect 10520 22080 10548 22188
rect 12360 22148 12388 22188
rect 12434 22176 12440 22228
rect 12492 22216 12498 22228
rect 13170 22216 13176 22228
rect 12492 22188 13176 22216
rect 12492 22176 12498 22188
rect 13170 22176 13176 22188
rect 13228 22176 13234 22228
rect 13262 22148 13268 22160
rect 12360 22120 13268 22148
rect 13262 22108 13268 22120
rect 13320 22108 13326 22160
rect 10689 22083 10747 22089
rect 10689 22080 10701 22083
rect 10520 22052 10701 22080
rect 10689 22049 10701 22052
rect 10735 22049 10747 22083
rect 10689 22043 10747 22049
rect 11606 22040 11612 22092
rect 11664 22040 11670 22092
rect 13633 22083 13691 22089
rect 13633 22049 13645 22083
rect 13679 22080 13691 22083
rect 13722 22080 13728 22092
rect 13679 22052 13728 22080
rect 13679 22049 13691 22052
rect 13633 22043 13691 22049
rect 13722 22040 13728 22052
rect 13780 22040 13786 22092
rect 9876 21984 10088 22012
rect 7558 21944 7564 21956
rect 7024 21916 7564 21944
rect 1489 21907 1547 21913
rect 7558 21904 7564 21916
rect 7616 21904 7622 21956
rect 9122 21904 9128 21956
rect 9180 21944 9186 21956
rect 9876 21944 9904 21984
rect 10778 21972 10784 22024
rect 10836 22021 10842 22024
rect 10836 22015 10864 22021
rect 10852 21981 10864 22015
rect 10836 21975 10864 21981
rect 10836 21972 10842 21975
rect 10962 21972 10968 22024
rect 11020 21972 11026 22024
rect 11701 22015 11759 22021
rect 11701 22012 11713 22015
rect 11624 21984 11713 22012
rect 11624 21956 11652 21984
rect 11701 21981 11713 21984
rect 11747 21981 11759 22015
rect 11701 21975 11759 21981
rect 11882 21972 11888 22024
rect 11940 22012 11946 22024
rect 11975 22015 12033 22021
rect 11975 22012 11987 22015
rect 11940 21984 11987 22012
rect 11940 21972 11946 21984
rect 11975 21981 11987 21984
rect 12021 21981 12033 22015
rect 11975 21975 12033 21981
rect 9180 21916 9904 21944
rect 9180 21904 9186 21916
rect 11606 21904 11612 21956
rect 11664 21944 11670 21956
rect 12250 21944 12256 21956
rect 11664 21916 12256 21944
rect 11664 21904 11670 21916
rect 12250 21904 12256 21916
rect 12308 21904 12314 21956
rect 13357 21947 13415 21953
rect 13357 21913 13369 21947
rect 13403 21944 13415 21947
rect 13814 21944 13820 21956
rect 13403 21916 13820 21944
rect 13403 21913 13415 21916
rect 13357 21907 13415 21913
rect 13814 21904 13820 21916
rect 13872 21904 13878 21956
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 2314 21876 2320 21888
rect 1627 21848 2320 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 2314 21836 2320 21848
rect 2372 21876 2378 21888
rect 4798 21876 4804 21888
rect 2372 21848 4804 21876
rect 2372 21836 2378 21848
rect 4798 21836 4804 21848
rect 4856 21836 4862 21888
rect 6362 21836 6368 21888
rect 6420 21876 6426 21888
rect 6549 21879 6607 21885
rect 6549 21876 6561 21879
rect 6420 21848 6561 21876
rect 6420 21836 6426 21848
rect 6549 21845 6561 21848
rect 6595 21845 6607 21879
rect 6549 21839 6607 21845
rect 8481 21879 8539 21885
rect 8481 21845 8493 21879
rect 8527 21876 8539 21879
rect 8754 21876 8760 21888
rect 8527 21848 8760 21876
rect 8527 21845 8539 21848
rect 8481 21839 8539 21845
rect 8754 21836 8760 21848
rect 8812 21836 8818 21888
rect 9766 21836 9772 21888
rect 9824 21876 9830 21888
rect 10226 21876 10232 21888
rect 9824 21848 10232 21876
rect 9824 21836 9830 21848
rect 10226 21836 10232 21848
rect 10284 21836 10290 21888
rect 10778 21836 10784 21888
rect 10836 21876 10842 21888
rect 12158 21876 12164 21888
rect 10836 21848 12164 21876
rect 10836 21836 10842 21848
rect 12158 21836 12164 21848
rect 12216 21836 12222 21888
rect 12713 21879 12771 21885
rect 12713 21845 12725 21879
rect 12759 21876 12771 21879
rect 12986 21876 12992 21888
rect 12759 21848 12992 21876
rect 12759 21845 12771 21848
rect 12713 21839 12771 21845
rect 12986 21836 12992 21848
rect 13044 21836 13050 21888
rect 13630 21836 13636 21888
rect 13688 21876 13694 21888
rect 15378 21876 15384 21888
rect 13688 21848 15384 21876
rect 13688 21836 13694 21848
rect 15378 21836 15384 21848
rect 15436 21836 15442 21888
rect 1104 21786 14696 21808
rect 1104 21734 4308 21786
rect 4360 21734 4372 21786
rect 4424 21734 4436 21786
rect 4488 21734 4500 21786
rect 4552 21734 4564 21786
rect 4616 21734 7666 21786
rect 7718 21734 7730 21786
rect 7782 21734 7794 21786
rect 7846 21734 7858 21786
rect 7910 21734 7922 21786
rect 7974 21734 11024 21786
rect 11076 21734 11088 21786
rect 11140 21734 11152 21786
rect 11204 21734 11216 21786
rect 11268 21734 11280 21786
rect 11332 21734 14382 21786
rect 14434 21734 14446 21786
rect 14498 21734 14510 21786
rect 14562 21734 14574 21786
rect 14626 21734 14638 21786
rect 14690 21734 14696 21786
rect 1104 21712 14696 21734
rect 5074 21632 5080 21684
rect 5132 21672 5138 21684
rect 5132 21644 9258 21672
rect 5132 21632 5138 21644
rect 1673 21607 1731 21613
rect 1673 21573 1685 21607
rect 1719 21604 1731 21607
rect 4522 21604 4528 21616
rect 1719 21576 4528 21604
rect 1719 21573 1731 21576
rect 1673 21567 1731 21573
rect 4522 21564 4528 21576
rect 4580 21564 4586 21616
rect 750 21496 756 21548
rect 808 21536 814 21548
rect 1489 21539 1547 21545
rect 1489 21536 1501 21539
rect 808 21508 1501 21536
rect 808 21496 814 21508
rect 1489 21505 1501 21508
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 4890 21496 4896 21548
rect 4948 21496 4954 21548
rect 5092 21536 5120 21632
rect 5534 21564 5540 21616
rect 5592 21604 5598 21616
rect 6822 21604 6828 21616
rect 5592 21576 6828 21604
rect 5592 21564 5598 21576
rect 6822 21564 6828 21576
rect 6880 21564 6886 21616
rect 9230 21604 9258 21644
rect 9398 21632 9404 21684
rect 9456 21632 9462 21684
rect 13630 21672 13636 21684
rect 9646 21644 11836 21672
rect 9646 21604 9674 21644
rect 11808 21616 11836 21644
rect 12406 21644 13636 21672
rect 9230 21576 9674 21604
rect 11790 21564 11796 21616
rect 11848 21564 11854 21616
rect 11885 21607 11943 21613
rect 11885 21573 11897 21607
rect 11931 21604 11943 21607
rect 12406 21604 12434 21644
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 15470 21632 15476 21684
rect 15528 21632 15534 21684
rect 11931 21576 12434 21604
rect 11931 21573 11943 21576
rect 11885 21567 11943 21573
rect 5151 21539 5209 21545
rect 5151 21536 5163 21539
rect 5092 21508 5163 21536
rect 5151 21505 5163 21508
rect 5197 21505 5209 21539
rect 5151 21499 5209 21505
rect 5258 21496 5264 21548
rect 5316 21536 5322 21548
rect 7561 21539 7619 21545
rect 5316 21508 7512 21536
rect 5316 21496 5322 21508
rect 7484 21468 7512 21508
rect 7561 21505 7573 21539
rect 7607 21536 7619 21539
rect 7607 21508 7972 21536
rect 7607 21505 7619 21508
rect 7561 21499 7619 21505
rect 7944 21480 7972 21508
rect 8478 21496 8484 21548
rect 8536 21496 8542 21548
rect 8754 21496 8760 21548
rect 8812 21496 8818 21548
rect 10686 21496 10692 21548
rect 10744 21496 10750 21548
rect 11698 21496 11704 21548
rect 11756 21496 11762 21548
rect 12345 21539 12403 21545
rect 12345 21505 12357 21539
rect 12391 21505 12403 21539
rect 12345 21499 12403 21505
rect 7742 21468 7748 21480
rect 7484 21440 7748 21468
rect 7742 21428 7748 21440
rect 7800 21428 7806 21480
rect 7926 21428 7932 21480
rect 7984 21428 7990 21480
rect 8598 21471 8656 21477
rect 8598 21468 8610 21471
rect 8036 21440 8610 21468
rect 5902 21292 5908 21344
rect 5960 21292 5966 21344
rect 7374 21292 7380 21344
rect 7432 21332 7438 21344
rect 8036 21332 8064 21440
rect 8598 21437 8610 21440
rect 8644 21468 8656 21471
rect 8644 21440 9168 21468
rect 8644 21437 8656 21440
rect 8598 21431 8656 21437
rect 8202 21360 8208 21412
rect 8260 21360 8266 21412
rect 7432 21304 8064 21332
rect 7432 21292 7438 21304
rect 8662 21292 8668 21344
rect 8720 21332 8726 21344
rect 8938 21332 8944 21344
rect 8720 21304 8944 21332
rect 8720 21292 8726 21304
rect 8938 21292 8944 21304
rect 8996 21292 9002 21344
rect 9140 21332 9168 21440
rect 9306 21428 9312 21480
rect 9364 21468 9370 21480
rect 9493 21471 9551 21477
rect 9493 21468 9505 21471
rect 9364 21440 9505 21468
rect 9364 21428 9370 21440
rect 9493 21437 9505 21440
rect 9539 21437 9551 21471
rect 9493 21431 9551 21437
rect 9677 21471 9735 21477
rect 9677 21437 9689 21471
rect 9723 21468 9735 21471
rect 9766 21468 9772 21480
rect 9723 21440 9772 21468
rect 9723 21437 9735 21440
rect 9677 21431 9735 21437
rect 9766 21428 9772 21440
rect 9824 21428 9830 21480
rect 10134 21428 10140 21480
rect 10192 21428 10198 21480
rect 10413 21471 10471 21477
rect 10413 21468 10425 21471
rect 10244 21440 10425 21468
rect 10244 21400 10272 21440
rect 10413 21437 10425 21440
rect 10459 21437 10471 21471
rect 10413 21431 10471 21437
rect 10551 21471 10609 21477
rect 10551 21437 10563 21471
rect 10597 21468 10609 21471
rect 11054 21468 11060 21480
rect 10597 21440 11060 21468
rect 10597 21437 10609 21440
rect 10551 21431 10609 21437
rect 11054 21428 11060 21440
rect 11112 21428 11118 21480
rect 11238 21428 11244 21480
rect 11296 21468 11302 21480
rect 12360 21468 12388 21499
rect 13538 21496 13544 21548
rect 13596 21496 13602 21548
rect 15488 21480 15516 21632
rect 11296 21440 12388 21468
rect 12529 21471 12587 21477
rect 11296 21428 11302 21440
rect 12529 21437 12541 21471
rect 12575 21437 12587 21471
rect 12529 21431 12587 21437
rect 11517 21403 11575 21409
rect 11517 21400 11529 21403
rect 10152 21372 10272 21400
rect 11072 21372 11529 21400
rect 10152 21344 10180 21372
rect 10042 21332 10048 21344
rect 9140 21304 10048 21332
rect 10042 21292 10048 21304
rect 10100 21292 10106 21344
rect 10134 21292 10140 21344
rect 10192 21332 10198 21344
rect 10594 21332 10600 21344
rect 10192 21304 10600 21332
rect 10192 21292 10198 21304
rect 10594 21292 10600 21304
rect 10652 21292 10658 21344
rect 10686 21292 10692 21344
rect 10744 21332 10750 21344
rect 11072 21332 11100 21372
rect 11517 21369 11529 21372
rect 11563 21369 11575 21403
rect 11517 21363 11575 21369
rect 11606 21360 11612 21412
rect 11664 21400 11670 21412
rect 11790 21400 11796 21412
rect 11664 21372 11796 21400
rect 11664 21360 11670 21372
rect 11790 21360 11796 21372
rect 11848 21360 11854 21412
rect 12544 21400 12572 21431
rect 12986 21428 12992 21480
rect 13044 21428 13050 21480
rect 13262 21428 13268 21480
rect 13320 21428 13326 21480
rect 13354 21428 13360 21480
rect 13412 21477 13418 21480
rect 13412 21471 13440 21477
rect 13428 21437 13440 21471
rect 13412 21431 13440 21437
rect 13412 21428 13418 21431
rect 15470 21428 15476 21480
rect 15528 21428 15534 21480
rect 13078 21400 13084 21412
rect 12544 21372 13084 21400
rect 13078 21360 13084 21372
rect 13136 21360 13142 21412
rect 10744 21304 11100 21332
rect 11333 21335 11391 21341
rect 10744 21292 10750 21304
rect 11333 21301 11345 21335
rect 11379 21332 11391 21335
rect 11882 21332 11888 21344
rect 11379 21304 11888 21332
rect 11379 21301 11391 21304
rect 11333 21295 11391 21301
rect 11882 21292 11888 21304
rect 11940 21292 11946 21344
rect 12161 21335 12219 21341
rect 12161 21301 12173 21335
rect 12207 21332 12219 21335
rect 14090 21332 14096 21344
rect 12207 21304 14096 21332
rect 12207 21301 12219 21304
rect 12161 21295 12219 21301
rect 14090 21292 14096 21304
rect 14148 21292 14154 21344
rect 14185 21335 14243 21341
rect 14185 21301 14197 21335
rect 14231 21332 14243 21335
rect 14231 21304 14596 21332
rect 14231 21301 14243 21304
rect 14185 21295 14243 21301
rect 1104 21242 14536 21264
rect 1104 21190 2629 21242
rect 2681 21190 2693 21242
rect 2745 21190 2757 21242
rect 2809 21190 2821 21242
rect 2873 21190 2885 21242
rect 2937 21190 5987 21242
rect 6039 21190 6051 21242
rect 6103 21190 6115 21242
rect 6167 21190 6179 21242
rect 6231 21190 6243 21242
rect 6295 21190 9345 21242
rect 9397 21190 9409 21242
rect 9461 21190 9473 21242
rect 9525 21190 9537 21242
rect 9589 21190 9601 21242
rect 9653 21190 12703 21242
rect 12755 21190 12767 21242
rect 12819 21190 12831 21242
rect 12883 21190 12895 21242
rect 12947 21190 12959 21242
rect 13011 21190 14536 21242
rect 1104 21168 14536 21190
rect 3234 21088 3240 21140
rect 3292 21088 3298 21140
rect 7282 21088 7288 21140
rect 7340 21088 7346 21140
rect 8478 21088 8484 21140
rect 8536 21128 8542 21140
rect 8938 21128 8944 21140
rect 8536 21100 8944 21128
rect 8536 21088 8542 21100
rect 8938 21088 8944 21100
rect 8996 21088 9002 21140
rect 9766 21128 9772 21140
rect 9048 21100 9772 21128
rect 9048 21060 9076 21100
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 10781 21131 10839 21137
rect 9876 21100 10732 21128
rect 9876 21060 9904 21100
rect 7114 21032 9076 21060
rect 9784 21032 9904 21060
rect 10704 21060 10732 21100
rect 10781 21097 10793 21131
rect 10827 21128 10839 21131
rect 10870 21128 10876 21140
rect 10827 21100 10876 21128
rect 10827 21097 10839 21100
rect 10781 21091 10839 21097
rect 10870 21088 10876 21100
rect 10928 21088 10934 21140
rect 11609 21131 11667 21137
rect 11609 21097 11621 21131
rect 11655 21128 11667 21131
rect 13998 21128 14004 21140
rect 11655 21100 14004 21128
rect 11655 21097 11667 21100
rect 11609 21091 11667 21097
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 11238 21060 11244 21072
rect 10704 21032 11244 21060
rect 5902 20952 5908 21004
rect 5960 20952 5966 21004
rect 3050 20884 3056 20936
rect 3108 20884 3114 20936
rect 6362 20884 6368 20936
rect 6420 20884 6426 20936
rect 6454 20884 6460 20936
rect 6512 20884 6518 20936
rect 7114 20924 7142 21032
rect 7742 20952 7748 21004
rect 7800 20992 7806 21004
rect 9784 20992 9812 21032
rect 11238 21020 11244 21032
rect 11296 21020 11302 21072
rect 14568 21060 14596 21304
rect 15010 21088 15016 21140
rect 15068 21128 15074 21140
rect 15194 21128 15200 21140
rect 15068 21100 15200 21128
rect 15068 21088 15074 21100
rect 15194 21088 15200 21100
rect 15252 21088 15258 21140
rect 11348 21032 14596 21060
rect 7800 20964 9812 20992
rect 7800 20952 7806 20964
rect 6564 20896 7142 20924
rect 5718 20816 5724 20868
rect 5776 20856 5782 20868
rect 6273 20859 6331 20865
rect 5776 20828 6132 20856
rect 5776 20816 5782 20828
rect 5534 20748 5540 20800
rect 5592 20788 5598 20800
rect 5902 20788 5908 20800
rect 5592 20760 5908 20788
rect 5592 20748 5598 20760
rect 5902 20748 5908 20760
rect 5960 20788 5966 20800
rect 5997 20791 6055 20797
rect 5997 20788 6009 20791
rect 5960 20760 6009 20788
rect 5960 20748 5966 20760
rect 5997 20757 6009 20760
rect 6043 20757 6055 20791
rect 6104 20788 6132 20828
rect 6273 20825 6285 20859
rect 6319 20856 6331 20859
rect 6472 20856 6500 20884
rect 6319 20828 6500 20856
rect 6319 20825 6331 20828
rect 6273 20819 6331 20825
rect 6564 20788 6592 20896
rect 8110 20884 8116 20936
rect 8168 20924 8174 20936
rect 8846 20924 8852 20936
rect 8168 20896 8852 20924
rect 8168 20884 8174 20896
rect 8846 20884 8852 20896
rect 8904 20884 8910 20936
rect 9582 20884 9588 20936
rect 9640 20924 9646 20936
rect 9640 20884 9674 20924
rect 9766 20884 9772 20936
rect 9824 20884 9830 20936
rect 11348 20933 11376 21032
rect 12710 20952 12716 21004
rect 12768 20952 12774 21004
rect 13265 20995 13323 21001
rect 13265 20961 13277 20995
rect 13311 20992 13323 20995
rect 15010 20992 15016 21004
rect 13311 20964 15016 20992
rect 13311 20961 13323 20964
rect 13265 20955 13323 20961
rect 15010 20952 15016 20964
rect 15068 20952 15074 21004
rect 10011 20927 10069 20933
rect 10011 20924 10023 20927
rect 9876 20896 10023 20924
rect 6730 20816 6736 20868
rect 6788 20816 6794 20868
rect 9646 20856 9674 20884
rect 9876 20856 9904 20896
rect 10011 20893 10023 20896
rect 10057 20893 10069 20927
rect 10011 20887 10069 20893
rect 11333 20927 11391 20933
rect 11333 20893 11345 20927
rect 11379 20893 11391 20927
rect 11333 20887 11391 20893
rect 12437 20927 12495 20933
rect 12437 20893 12449 20927
rect 12483 20924 12495 20927
rect 13354 20924 13360 20936
rect 12483 20896 13360 20924
rect 12483 20893 12495 20896
rect 12437 20887 12495 20893
rect 13354 20884 13360 20896
rect 13412 20884 13418 20936
rect 13909 20927 13967 20933
rect 13909 20893 13921 20927
rect 13955 20924 13967 20927
rect 14274 20924 14280 20936
rect 13955 20896 14280 20924
rect 13955 20893 13967 20896
rect 13909 20887 13967 20893
rect 14274 20884 14280 20896
rect 14332 20884 14338 20936
rect 11885 20859 11943 20865
rect 11885 20856 11897 20859
rect 9646 20828 9904 20856
rect 10152 20828 11897 20856
rect 6104 20760 6592 20788
rect 7101 20791 7159 20797
rect 5997 20751 6055 20757
rect 7101 20757 7113 20791
rect 7147 20788 7159 20791
rect 8110 20788 8116 20800
rect 7147 20760 8116 20788
rect 7147 20757 7159 20760
rect 7101 20751 7159 20757
rect 8110 20748 8116 20760
rect 8168 20748 8174 20800
rect 8478 20748 8484 20800
rect 8536 20788 8542 20800
rect 10152 20788 10180 20828
rect 11885 20825 11897 20828
rect 11931 20825 11943 20859
rect 11885 20819 11943 20825
rect 12253 20859 12311 20865
rect 12253 20825 12265 20859
rect 12299 20856 12311 20859
rect 12299 20828 12434 20856
rect 12299 20825 12311 20828
rect 12253 20819 12311 20825
rect 8536 20760 10180 20788
rect 8536 20748 8542 20760
rect 10226 20748 10232 20800
rect 10284 20788 10290 20800
rect 10870 20788 10876 20800
rect 10284 20760 10876 20788
rect 10284 20748 10290 20760
rect 10870 20748 10876 20760
rect 10928 20748 10934 20800
rect 12406 20788 12434 20828
rect 12526 20816 12532 20868
rect 12584 20856 12590 20868
rect 12989 20859 13047 20865
rect 12989 20856 13001 20859
rect 12584 20828 13001 20856
rect 12584 20816 12590 20828
rect 12989 20825 13001 20828
rect 13035 20825 13047 20859
rect 12989 20819 13047 20825
rect 13541 20859 13599 20865
rect 13541 20825 13553 20859
rect 13587 20856 13599 20859
rect 13998 20856 14004 20868
rect 13587 20828 14004 20856
rect 13587 20825 13599 20828
rect 13541 20819 13599 20825
rect 13998 20816 14004 20828
rect 14056 20816 14062 20868
rect 15286 20788 15292 20800
rect 12406 20760 15292 20788
rect 15286 20748 15292 20760
rect 15344 20748 15350 20800
rect 1104 20698 14696 20720
rect 1104 20646 4308 20698
rect 4360 20646 4372 20698
rect 4424 20646 4436 20698
rect 4488 20646 4500 20698
rect 4552 20646 4564 20698
rect 4616 20646 7666 20698
rect 7718 20646 7730 20698
rect 7782 20646 7794 20698
rect 7846 20646 7858 20698
rect 7910 20646 7922 20698
rect 7974 20646 11024 20698
rect 11076 20646 11088 20698
rect 11140 20646 11152 20698
rect 11204 20646 11216 20698
rect 11268 20646 11280 20698
rect 11332 20646 14382 20698
rect 14434 20646 14446 20698
rect 14498 20646 14510 20698
rect 14562 20646 14574 20698
rect 14626 20646 14638 20698
rect 14690 20646 14696 20698
rect 1104 20624 14696 20646
rect 8021 20587 8079 20593
rect 5184 20556 7972 20584
rect 1670 20476 1676 20528
rect 1728 20516 1734 20528
rect 1728 20488 2774 20516
rect 1728 20476 1734 20488
rect 2746 20448 2774 20488
rect 5184 20460 5212 20556
rect 5442 20476 5448 20528
rect 5500 20516 5506 20528
rect 7098 20516 7104 20528
rect 5500 20488 7104 20516
rect 5500 20476 5506 20488
rect 7098 20476 7104 20488
rect 7156 20516 7162 20528
rect 7944 20516 7972 20556
rect 8021 20553 8033 20587
rect 8067 20584 8079 20587
rect 8202 20584 8208 20596
rect 8067 20556 8208 20584
rect 8067 20553 8079 20556
rect 8021 20547 8079 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 9122 20544 9128 20596
rect 9180 20584 9186 20596
rect 9766 20584 9772 20596
rect 9180 20556 9772 20584
rect 9180 20544 9186 20556
rect 9766 20544 9772 20556
rect 9824 20544 9830 20596
rect 11149 20587 11207 20593
rect 11149 20553 11161 20587
rect 11195 20553 11207 20587
rect 11149 20547 11207 20553
rect 11164 20516 11192 20547
rect 11882 20544 11888 20596
rect 11940 20584 11946 20596
rect 13633 20587 13691 20593
rect 11940 20556 12296 20584
rect 11940 20544 11946 20556
rect 7156 20488 7236 20516
rect 7944 20488 10042 20516
rect 11164 20488 11744 20516
rect 7156 20476 7162 20488
rect 7208 20478 7236 20488
rect 10014 20487 10042 20488
rect 7267 20481 7325 20487
rect 7267 20478 7279 20481
rect 2746 20420 5120 20448
rect 750 20340 756 20392
rect 808 20380 814 20392
rect 1397 20383 1455 20389
rect 1397 20380 1409 20383
rect 808 20352 1409 20380
rect 808 20340 814 20352
rect 1397 20349 1409 20352
rect 1443 20349 1455 20383
rect 1397 20343 1455 20349
rect 1673 20383 1731 20389
rect 1673 20349 1685 20383
rect 1719 20349 1731 20383
rect 5092 20380 5120 20420
rect 5166 20408 5172 20460
rect 5224 20408 5230 20460
rect 7208 20450 7279 20478
rect 7267 20447 7279 20450
rect 7313 20447 7325 20481
rect 10014 20481 10085 20487
rect 7267 20441 7325 20447
rect 7926 20408 7932 20460
rect 7984 20448 7990 20460
rect 9122 20448 9128 20460
rect 7984 20420 9128 20448
rect 7984 20408 7990 20420
rect 9122 20408 9128 20420
rect 9180 20408 9186 20460
rect 10014 20450 10039 20481
rect 10027 20447 10039 20450
rect 10073 20447 10085 20481
rect 11716 20457 11744 20488
rect 12158 20487 12164 20528
rect 12143 20481 12164 20487
rect 10027 20441 10085 20447
rect 11333 20451 11391 20457
rect 11333 20417 11345 20451
rect 11379 20417 11391 20451
rect 11333 20411 11391 20417
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20417 11759 20451
rect 12143 20447 12155 20481
rect 12216 20476 12222 20528
rect 12189 20450 12204 20476
rect 12189 20447 12201 20450
rect 12143 20441 12201 20447
rect 12268 20448 12296 20556
rect 13633 20553 13645 20587
rect 13679 20584 13691 20587
rect 13722 20584 13728 20596
rect 13679 20556 13728 20584
rect 13679 20553 13691 20556
rect 13633 20547 13691 20553
rect 13722 20544 13728 20556
rect 13780 20544 13786 20596
rect 13357 20451 13415 20457
rect 13357 20448 13369 20451
rect 12268 20420 13369 20448
rect 11701 20411 11759 20417
rect 13357 20417 13369 20420
rect 13403 20417 13415 20451
rect 13357 20411 13415 20417
rect 6914 20380 6920 20392
rect 5092 20352 6920 20380
rect 1673 20343 1731 20349
rect 1688 20312 1716 20343
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7006 20340 7012 20392
rect 7064 20340 7070 20392
rect 8754 20340 8760 20392
rect 8812 20340 8818 20392
rect 9674 20340 9680 20392
rect 9732 20380 9738 20392
rect 9769 20383 9827 20389
rect 9769 20380 9781 20383
rect 9732 20352 9781 20380
rect 9732 20340 9738 20352
rect 9769 20349 9781 20352
rect 9815 20349 9827 20383
rect 11348 20380 11376 20411
rect 9769 20343 9827 20349
rect 10486 20352 11376 20380
rect 8772 20312 8800 20340
rect 9122 20312 9128 20324
rect 1688 20284 6893 20312
rect 6865 20244 6893 20284
rect 7666 20284 9128 20312
rect 7666 20244 7694 20284
rect 9122 20272 9128 20284
rect 9180 20272 9186 20324
rect 6865 20216 7694 20244
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 9030 20244 9036 20256
rect 8352 20216 9036 20244
rect 8352 20204 8358 20216
rect 9030 20204 9036 20216
rect 9088 20244 9094 20256
rect 10486 20244 10514 20352
rect 10781 20315 10839 20321
rect 10781 20281 10793 20315
rect 10827 20312 10839 20315
rect 10962 20312 10968 20324
rect 10827 20284 10968 20312
rect 10827 20281 10839 20284
rect 10781 20275 10839 20281
rect 10962 20272 10968 20284
rect 11020 20312 11026 20324
rect 11532 20312 11560 20411
rect 14182 20408 14188 20460
rect 14240 20408 14246 20460
rect 11882 20340 11888 20392
rect 11940 20340 11946 20392
rect 13262 20340 13268 20392
rect 13320 20380 13326 20392
rect 13722 20380 13728 20392
rect 13320 20352 13728 20380
rect 13320 20340 13326 20352
rect 13722 20340 13728 20352
rect 13780 20340 13786 20392
rect 11020 20284 11560 20312
rect 11020 20272 11026 20284
rect 14200 20256 14228 20408
rect 9088 20216 10514 20244
rect 9088 20204 9094 20216
rect 11606 20204 11612 20256
rect 11664 20204 11670 20256
rect 12618 20204 12624 20256
rect 12676 20244 12682 20256
rect 12897 20247 12955 20253
rect 12897 20244 12909 20247
rect 12676 20216 12909 20244
rect 12676 20204 12682 20216
rect 12897 20213 12909 20216
rect 12943 20213 12955 20247
rect 12897 20207 12955 20213
rect 14182 20204 14188 20256
rect 14240 20204 14246 20256
rect 1104 20154 14536 20176
rect 1104 20102 2629 20154
rect 2681 20102 2693 20154
rect 2745 20102 2757 20154
rect 2809 20102 2821 20154
rect 2873 20102 2885 20154
rect 2937 20102 5987 20154
rect 6039 20102 6051 20154
rect 6103 20102 6115 20154
rect 6167 20102 6179 20154
rect 6231 20102 6243 20154
rect 6295 20102 9345 20154
rect 9397 20102 9409 20154
rect 9461 20102 9473 20154
rect 9525 20102 9537 20154
rect 9589 20102 9601 20154
rect 9653 20102 12703 20154
rect 12755 20102 12767 20154
rect 12819 20102 12831 20154
rect 12883 20102 12895 20154
rect 12947 20102 12959 20154
rect 13011 20102 14536 20154
rect 1104 20080 14536 20102
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 1670 20040 1676 20052
rect 1627 20012 1676 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 1670 20000 1676 20012
rect 1728 20000 1734 20052
rect 9858 20040 9864 20052
rect 7024 20012 9864 20040
rect 6365 19975 6423 19981
rect 6365 19941 6377 19975
rect 6411 19972 6423 19975
rect 7024 19972 7052 20012
rect 9858 20000 9864 20012
rect 9916 20000 9922 20052
rect 11606 20000 11612 20052
rect 11664 20000 11670 20052
rect 11974 20000 11980 20052
rect 12032 20040 12038 20052
rect 12032 20012 12848 20040
rect 12032 20000 12038 20012
rect 6411 19944 7052 19972
rect 6411 19941 6423 19944
rect 6365 19935 6423 19941
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 7024 19845 7052 19944
rect 7282 19932 7288 19984
rect 7340 19972 7346 19984
rect 7466 19972 7472 19984
rect 7340 19944 7472 19972
rect 7340 19932 7346 19944
rect 7466 19932 7472 19944
rect 7524 19932 7530 19984
rect 8938 19864 8944 19916
rect 8996 19864 9002 19916
rect 10781 19907 10839 19913
rect 10781 19873 10793 19907
rect 10827 19904 10839 19907
rect 11057 19907 11115 19913
rect 11057 19904 11069 19907
rect 10827 19876 11069 19904
rect 10827 19873 10839 19876
rect 10781 19867 10839 19873
rect 11057 19873 11069 19876
rect 11103 19873 11115 19907
rect 11057 19867 11115 19873
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19904 11299 19907
rect 11624 19904 11652 20000
rect 12618 19904 12624 19916
rect 11287 19876 11652 19904
rect 11808 19876 12624 19904
rect 11287 19873 11299 19876
rect 11241 19867 11299 19873
rect 4617 19839 4675 19845
rect 4617 19836 4629 19839
rect 4212 19808 4629 19836
rect 4212 19796 4218 19808
rect 4617 19805 4629 19808
rect 4663 19805 4675 19839
rect 4617 19799 4675 19805
rect 7009 19839 7067 19845
rect 7009 19805 7021 19839
rect 7055 19805 7067 19839
rect 7009 19799 7067 19805
rect 7466 19796 7472 19848
rect 7524 19796 7530 19848
rect 7743 19839 7801 19845
rect 7743 19805 7755 19839
rect 7789 19805 7801 19839
rect 8956 19836 8984 19864
rect 8956 19808 9042 19836
rect 7743 19799 7801 19805
rect 750 19728 756 19780
rect 808 19768 814 19780
rect 4890 19777 4896 19780
rect 1489 19771 1547 19777
rect 1489 19768 1501 19771
rect 808 19740 1501 19768
rect 808 19728 814 19740
rect 1489 19737 1501 19740
rect 1535 19737 1547 19771
rect 4884 19768 4896 19777
rect 4851 19740 4896 19768
rect 1489 19731 1547 19737
rect 4884 19731 4896 19740
rect 4948 19768 4954 19780
rect 6181 19771 6239 19777
rect 6181 19768 6193 19771
rect 4948 19740 6193 19768
rect 4890 19728 4896 19731
rect 4948 19728 4954 19740
rect 6181 19737 6193 19740
rect 6227 19737 6239 19771
rect 7758 19768 7786 19799
rect 8754 19768 8760 19780
rect 6181 19731 6239 19737
rect 6748 19740 7696 19768
rect 7758 19740 8760 19768
rect 5997 19703 6055 19709
rect 5997 19669 6009 19703
rect 6043 19700 6055 19703
rect 6748 19700 6776 19740
rect 6043 19672 6776 19700
rect 6043 19669 6055 19672
rect 5997 19663 6055 19669
rect 6822 19660 6828 19712
rect 6880 19660 6886 19712
rect 7668 19700 7696 19740
rect 8754 19728 8760 19740
rect 8812 19728 8818 19780
rect 8294 19700 8300 19712
rect 7668 19672 8300 19700
rect 8294 19660 8300 19672
rect 8352 19660 8358 19712
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8846 19700 8852 19712
rect 8527 19672 8852 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9014 19700 9042 19808
rect 9122 19796 9128 19848
rect 9180 19836 9186 19848
rect 9215 19839 9273 19845
rect 9215 19836 9227 19839
rect 9180 19808 9227 19836
rect 9180 19796 9186 19808
rect 9215 19805 9227 19808
rect 9261 19805 9273 19839
rect 9215 19799 9273 19805
rect 10686 19796 10692 19848
rect 10744 19796 10750 19848
rect 10962 19796 10968 19848
rect 11020 19796 11026 19848
rect 11808 19845 11836 19876
rect 12618 19864 12624 19876
rect 12676 19864 12682 19916
rect 12710 19864 12716 19916
rect 12768 19864 12774 19916
rect 12820 19904 12848 20012
rect 13906 20000 13912 20052
rect 13964 20000 13970 20052
rect 13106 19907 13164 19913
rect 13106 19904 13118 19907
rect 12820 19876 13118 19904
rect 13106 19873 13118 19876
rect 13152 19904 13164 19907
rect 13630 19904 13636 19916
rect 13152 19876 13636 19904
rect 13152 19873 13164 19876
rect 13106 19867 13164 19873
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 11793 19839 11851 19845
rect 11793 19805 11805 19839
rect 11839 19805 11851 19839
rect 11793 19799 11851 19805
rect 12066 19796 12072 19848
rect 12124 19796 12130 19848
rect 12250 19796 12256 19848
rect 12308 19796 12314 19848
rect 12986 19796 12992 19848
rect 13044 19796 13050 19848
rect 13262 19796 13268 19848
rect 13320 19796 13326 19848
rect 11241 19771 11299 19777
rect 11241 19737 11253 19771
rect 11287 19768 11299 19771
rect 11330 19768 11336 19780
rect 11287 19740 11336 19768
rect 11287 19737 11299 19740
rect 11241 19731 11299 19737
rect 11330 19728 11336 19740
rect 11388 19728 11394 19780
rect 11425 19771 11483 19777
rect 11425 19737 11437 19771
rect 11471 19768 11483 19771
rect 11471 19740 11928 19768
rect 11471 19737 11483 19740
rect 11425 19731 11483 19737
rect 9858 19700 9864 19712
rect 9014 19672 9864 19700
rect 9858 19660 9864 19672
rect 9916 19660 9922 19712
rect 9950 19660 9956 19712
rect 10008 19660 10014 19712
rect 11900 19700 11928 19740
rect 13814 19700 13820 19712
rect 11900 19672 13820 19700
rect 13814 19660 13820 19672
rect 13872 19660 13878 19712
rect 1104 19610 14696 19632
rect 1104 19558 4308 19610
rect 4360 19558 4372 19610
rect 4424 19558 4436 19610
rect 4488 19558 4500 19610
rect 4552 19558 4564 19610
rect 4616 19558 7666 19610
rect 7718 19558 7730 19610
rect 7782 19558 7794 19610
rect 7846 19558 7858 19610
rect 7910 19558 7922 19610
rect 7974 19558 11024 19610
rect 11076 19558 11088 19610
rect 11140 19558 11152 19610
rect 11204 19558 11216 19610
rect 11268 19558 11280 19610
rect 11332 19558 14382 19610
rect 14434 19558 14446 19610
rect 14498 19558 14510 19610
rect 14562 19558 14574 19610
rect 14626 19558 14638 19610
rect 14690 19558 14696 19610
rect 1104 19536 14696 19558
rect 6822 19456 6828 19508
rect 6880 19456 6886 19508
rect 7466 19456 7472 19508
rect 7524 19496 7530 19508
rect 11882 19496 11888 19508
rect 7524 19468 11888 19496
rect 7524 19456 7530 19468
rect 11882 19456 11888 19468
rect 11940 19496 11946 19508
rect 11940 19468 12204 19496
rect 11940 19456 11946 19468
rect 6840 19428 6868 19456
rect 6840 19400 7972 19428
rect 3694 19320 3700 19372
rect 3752 19360 3758 19372
rect 5166 19360 5172 19372
rect 3752 19332 5172 19360
rect 3752 19320 3758 19332
rect 5166 19320 5172 19332
rect 5224 19320 5230 19372
rect 6362 19320 6368 19372
rect 6420 19320 6426 19372
rect 6638 19360 6644 19372
rect 6599 19332 6644 19360
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 7006 19320 7012 19372
rect 7064 19360 7070 19372
rect 7064 19332 7236 19360
rect 7064 19320 7070 19332
rect 7116 19306 7236 19332
rect 7282 19320 7288 19372
rect 7340 19334 7346 19372
rect 7340 19320 7420 19334
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 7944 19369 7972 19400
rect 10318 19388 10324 19440
rect 10376 19428 10382 19440
rect 11793 19431 11851 19437
rect 11793 19428 11805 19431
rect 10376 19400 11805 19428
rect 10376 19388 10382 19400
rect 11793 19397 11805 19400
rect 11839 19397 11851 19431
rect 11793 19391 11851 19397
rect 7745 19363 7803 19369
rect 7745 19360 7757 19363
rect 7524 19332 7757 19360
rect 7524 19320 7530 19332
rect 7745 19329 7757 19332
rect 7791 19329 7803 19363
rect 7745 19323 7803 19329
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 8573 19363 8631 19369
rect 8573 19329 8585 19363
rect 8619 19360 8631 19363
rect 8938 19360 8944 19372
rect 8619 19332 8944 19360
rect 8619 19329 8631 19332
rect 8573 19323 8631 19329
rect 8938 19320 8944 19332
rect 8996 19320 9002 19372
rect 10965 19363 11023 19369
rect 10965 19329 10977 19363
rect 11011 19360 11023 19363
rect 11606 19360 11612 19372
rect 11011 19332 11612 19360
rect 11011 19329 11023 19332
rect 10965 19323 11023 19329
rect 11606 19320 11612 19332
rect 11664 19320 11670 19372
rect 12176 19360 12204 19468
rect 12250 19456 12256 19508
rect 12308 19496 12314 19508
rect 12308 19468 13216 19496
rect 12308 19456 12314 19468
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 13188 19428 13216 19468
rect 13262 19456 13268 19508
rect 13320 19496 13326 19508
rect 13541 19499 13599 19505
rect 13541 19496 13553 19499
rect 13320 19468 13553 19496
rect 13320 19456 13326 19468
rect 13541 19465 13553 19468
rect 13587 19465 13599 19499
rect 13541 19459 13599 19465
rect 14090 19456 14096 19508
rect 14148 19456 14154 19508
rect 12492 19400 12756 19428
rect 13188 19400 13676 19428
rect 12492 19388 12498 19400
rect 12728 19390 12756 19400
rect 12787 19393 12845 19399
rect 12787 19390 12799 19393
rect 12728 19362 12799 19390
rect 12176 19332 12480 19360
rect 12787 19359 12799 19362
rect 12833 19359 12845 19393
rect 13648 19372 13676 19400
rect 12787 19353 12845 19359
rect 7300 19306 7420 19320
rect 7116 19292 7144 19306
rect 7022 19264 7144 19292
rect 7392 19292 7420 19306
rect 12452 19304 12480 19332
rect 13262 19320 13268 19372
rect 13320 19360 13326 19372
rect 13538 19360 13544 19372
rect 13320 19332 13544 19360
rect 13320 19320 13326 19332
rect 13538 19320 13544 19332
rect 13596 19320 13602 19372
rect 13630 19320 13636 19372
rect 13688 19320 13694 19372
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19360 13967 19363
rect 14090 19360 14096 19372
rect 13955 19332 14096 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 14090 19320 14096 19332
rect 14148 19320 14154 19372
rect 7650 19292 7656 19304
rect 7392 19264 7656 19292
rect 6822 19116 6828 19168
rect 6880 19156 6886 19168
rect 7022 19156 7050 19264
rect 7650 19252 7656 19264
rect 7708 19252 7714 19304
rect 8754 19252 8760 19304
rect 8812 19252 8818 19304
rect 8846 19252 8852 19304
rect 8904 19292 8910 19304
rect 9217 19295 9275 19301
rect 9217 19292 9229 19295
rect 8904 19264 9229 19292
rect 8904 19252 8910 19264
rect 9217 19261 9229 19264
rect 9263 19261 9275 19295
rect 9493 19295 9551 19301
rect 9493 19292 9505 19295
rect 9217 19255 9275 19261
rect 9324 19264 9505 19292
rect 7377 19227 7435 19233
rect 7377 19193 7389 19227
rect 7423 19224 7435 19227
rect 7466 19224 7472 19236
rect 7423 19196 7472 19224
rect 7423 19193 7435 19196
rect 7377 19187 7435 19193
rect 7466 19184 7472 19196
rect 7524 19184 7530 19236
rect 6880 19128 7050 19156
rect 6880 19116 6886 19128
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 7742 19156 7748 19168
rect 7616 19128 7748 19156
rect 7616 19116 7622 19128
rect 7742 19116 7748 19128
rect 7800 19116 7806 19168
rect 7834 19116 7840 19168
rect 7892 19116 7898 19168
rect 8846 19116 8852 19168
rect 8904 19156 8910 19168
rect 9324 19156 9352 19264
rect 9493 19261 9505 19264
rect 9539 19261 9551 19295
rect 9493 19255 9551 19261
rect 9582 19252 9588 19304
rect 9640 19301 9646 19304
rect 9640 19295 9668 19301
rect 9656 19261 9668 19295
rect 9640 19255 9668 19261
rect 9640 19252 9646 19255
rect 9766 19252 9772 19304
rect 9824 19252 9830 19304
rect 10778 19292 10784 19304
rect 10336 19264 10784 19292
rect 10336 19156 10364 19264
rect 10778 19252 10784 19264
rect 10836 19252 10842 19304
rect 11238 19252 11244 19304
rect 11296 19252 11302 19304
rect 12069 19295 12127 19301
rect 12069 19261 12081 19295
rect 12115 19292 12127 19295
rect 12158 19292 12164 19304
rect 12115 19264 12164 19292
rect 12115 19261 12127 19264
rect 12069 19255 12127 19261
rect 12158 19252 12164 19264
rect 12216 19252 12222 19304
rect 12434 19252 12440 19304
rect 12492 19292 12498 19304
rect 12529 19295 12587 19301
rect 12529 19292 12541 19295
rect 12492 19264 12541 19292
rect 12492 19252 12498 19264
rect 12529 19261 12541 19264
rect 12575 19261 12587 19295
rect 12529 19255 12587 19261
rect 10428 19196 12434 19224
rect 10428 19165 10456 19196
rect 8904 19128 10364 19156
rect 10413 19159 10471 19165
rect 8904 19116 8910 19128
rect 10413 19125 10425 19159
rect 10459 19125 10471 19159
rect 12406 19156 12434 19196
rect 12526 19156 12532 19168
rect 12406 19128 12532 19156
rect 10413 19119 10471 19125
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 1104 19066 14536 19088
rect 1104 19014 2629 19066
rect 2681 19014 2693 19066
rect 2745 19014 2757 19066
rect 2809 19014 2821 19066
rect 2873 19014 2885 19066
rect 2937 19014 5987 19066
rect 6039 19014 6051 19066
rect 6103 19014 6115 19066
rect 6167 19014 6179 19066
rect 6231 19014 6243 19066
rect 6295 19014 9345 19066
rect 9397 19014 9409 19066
rect 9461 19014 9473 19066
rect 9525 19014 9537 19066
rect 9589 19014 9601 19066
rect 9653 19014 12703 19066
rect 12755 19014 12767 19066
rect 12819 19014 12831 19066
rect 12883 19014 12895 19066
rect 12947 19014 12959 19066
rect 13011 19014 14536 19066
rect 1104 18992 14536 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 5810 18952 5816 18964
rect 1627 18924 5816 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 6454 18912 6460 18964
rect 6512 18912 6518 18964
rect 7834 18952 7840 18964
rect 7300 18924 7840 18952
rect 6472 18816 6500 18912
rect 6380 18788 6500 18816
rect 5902 18708 5908 18760
rect 5960 18748 5966 18760
rect 6380 18757 6408 18788
rect 6730 18776 6736 18828
rect 6788 18776 6794 18828
rect 7300 18825 7328 18924
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 8294 18912 8300 18964
rect 8352 18912 8358 18964
rect 8570 18912 8576 18964
rect 8628 18912 8634 18964
rect 9766 18912 9772 18964
rect 9824 18952 9830 18964
rect 9953 18955 10011 18961
rect 9953 18952 9965 18955
rect 9824 18924 9965 18952
rect 9824 18912 9830 18924
rect 9953 18921 9965 18924
rect 9999 18921 10011 18955
rect 9953 18915 10011 18921
rect 10226 18912 10232 18964
rect 10284 18952 10290 18964
rect 12161 18955 12219 18961
rect 10284 18924 11008 18952
rect 10284 18912 10290 18924
rect 7466 18844 7472 18896
rect 7524 18884 7530 18896
rect 7929 18887 7987 18893
rect 7929 18884 7941 18887
rect 7524 18856 7941 18884
rect 7524 18844 7530 18856
rect 7929 18853 7941 18856
rect 7975 18853 7987 18887
rect 7929 18847 7987 18853
rect 7285 18819 7343 18825
rect 7285 18785 7297 18819
rect 7331 18785 7343 18819
rect 8312 18816 8340 18912
rect 7285 18779 7343 18785
rect 7852 18788 8340 18816
rect 6365 18751 6423 18757
rect 6365 18748 6377 18751
rect 5960 18720 6377 18748
rect 5960 18708 5966 18720
rect 6365 18717 6377 18720
rect 6411 18717 6423 18751
rect 6365 18711 6423 18717
rect 6457 18751 6515 18757
rect 6457 18717 6469 18751
rect 6503 18717 6515 18751
rect 6457 18711 6515 18717
rect 6549 18751 6607 18757
rect 6549 18717 6561 18751
rect 6595 18748 6607 18751
rect 6914 18748 6920 18760
rect 6595 18720 6920 18748
rect 6595 18717 6607 18720
rect 6549 18711 6607 18717
rect 750 18640 756 18692
rect 808 18680 814 18692
rect 1489 18683 1547 18689
rect 1489 18680 1501 18683
rect 808 18652 1501 18680
rect 808 18640 814 18652
rect 1489 18649 1501 18652
rect 1535 18649 1547 18683
rect 1489 18643 1547 18649
rect 5169 18683 5227 18689
rect 5169 18649 5181 18683
rect 5215 18649 5227 18683
rect 6472 18680 6500 18711
rect 6914 18708 6920 18720
rect 6972 18708 6978 18760
rect 7006 18708 7012 18760
rect 7064 18708 7070 18760
rect 7852 18757 7880 18788
rect 7101 18751 7159 18757
rect 7101 18717 7113 18751
rect 7147 18717 7159 18751
rect 7101 18711 7159 18717
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18748 7435 18751
rect 7837 18751 7895 18757
rect 7423 18720 7696 18748
rect 7423 18717 7435 18720
rect 7377 18711 7435 18717
rect 5169 18643 5227 18649
rect 6380 18652 6500 18680
rect 7116 18680 7144 18711
rect 7469 18683 7527 18689
rect 7469 18680 7481 18683
rect 7116 18652 7481 18680
rect 4798 18572 4804 18624
rect 4856 18612 4862 18624
rect 5184 18612 5212 18643
rect 6380 18624 6408 18652
rect 7469 18649 7481 18652
rect 7515 18649 7527 18683
rect 7469 18643 7527 18649
rect 4856 18584 5212 18612
rect 5261 18615 5319 18621
rect 4856 18572 4862 18584
rect 5261 18581 5273 18615
rect 5307 18612 5319 18615
rect 6086 18612 6092 18624
rect 5307 18584 6092 18612
rect 5307 18581 5319 18584
rect 5261 18575 5319 18581
rect 6086 18572 6092 18584
rect 6144 18572 6150 18624
rect 6178 18572 6184 18624
rect 6236 18572 6242 18624
rect 6362 18572 6368 18624
rect 6420 18572 6426 18624
rect 6733 18615 6791 18621
rect 6733 18581 6745 18615
rect 6779 18612 6791 18615
rect 7006 18612 7012 18624
rect 6779 18584 7012 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 7282 18572 7288 18624
rect 7340 18572 7346 18624
rect 7668 18621 7696 18720
rect 7837 18717 7849 18751
rect 7883 18717 7895 18751
rect 7837 18711 7895 18717
rect 8113 18751 8171 18757
rect 8113 18717 8125 18751
rect 8159 18748 8171 18751
rect 8159 18720 8248 18748
rect 8159 18717 8171 18720
rect 8113 18711 8171 18717
rect 8220 18624 8248 18720
rect 8312 18624 8340 18788
rect 8588 18748 8616 18912
rect 10980 18884 11008 18924
rect 12161 18921 12173 18955
rect 12207 18952 12219 18955
rect 13998 18952 14004 18964
rect 12207 18924 14004 18952
rect 12207 18921 12219 18924
rect 12161 18915 12219 18921
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 12342 18884 12348 18896
rect 10980 18856 12348 18884
rect 12342 18844 12348 18856
rect 12400 18844 12406 18896
rect 8846 18776 8852 18828
rect 8904 18816 8910 18828
rect 8941 18819 8999 18825
rect 8941 18816 8953 18819
rect 8904 18788 8953 18816
rect 8904 18776 8910 18788
rect 8941 18785 8953 18788
rect 8987 18785 8999 18819
rect 8941 18779 8999 18785
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 10321 18819 10379 18825
rect 10321 18816 10333 18819
rect 9916 18788 10333 18816
rect 9916 18776 9922 18788
rect 10321 18785 10333 18788
rect 10367 18785 10379 18819
rect 10321 18779 10379 18785
rect 9183 18751 9241 18757
rect 9183 18748 9195 18751
rect 8588 18720 9195 18748
rect 9183 18717 9195 18720
rect 9229 18748 9241 18751
rect 10563 18751 10621 18757
rect 10563 18748 10575 18751
rect 9229 18720 10575 18748
rect 9229 18717 9241 18720
rect 9183 18711 9241 18717
rect 10563 18717 10575 18720
rect 10609 18717 10621 18751
rect 10563 18711 10621 18717
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 12711 18751 12769 18757
rect 12492 18720 12572 18748
rect 12492 18708 12498 18720
rect 11885 18683 11943 18689
rect 11885 18680 11897 18683
rect 8772 18652 11897 18680
rect 7653 18615 7711 18621
rect 7653 18581 7665 18615
rect 7699 18581 7711 18615
rect 7653 18575 7711 18581
rect 8202 18572 8208 18624
rect 8260 18572 8266 18624
rect 8294 18572 8300 18624
rect 8352 18572 8358 18624
rect 8662 18572 8668 18624
rect 8720 18612 8726 18624
rect 8772 18612 8800 18652
rect 11885 18649 11897 18652
rect 11931 18649 11943 18683
rect 11885 18643 11943 18649
rect 12544 18624 12572 18720
rect 12711 18717 12723 18751
rect 12757 18748 12769 18751
rect 13446 18748 13452 18760
rect 12757 18720 13452 18748
rect 12757 18717 12769 18720
rect 12711 18711 12769 18717
rect 13446 18708 13452 18720
rect 13504 18708 13510 18760
rect 14366 18708 14372 18760
rect 14424 18748 14430 18760
rect 15562 18748 15568 18760
rect 14424 18720 15568 18748
rect 14424 18708 14430 18720
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 8720 18584 8800 18612
rect 8720 18572 8726 18584
rect 10226 18572 10232 18624
rect 10284 18612 10290 18624
rect 10502 18612 10508 18624
rect 10284 18584 10508 18612
rect 10284 18572 10290 18584
rect 10502 18572 10508 18584
rect 10560 18572 10566 18624
rect 11333 18615 11391 18621
rect 11333 18581 11345 18615
rect 11379 18612 11391 18615
rect 11514 18612 11520 18624
rect 11379 18584 11520 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11514 18572 11520 18584
rect 11572 18572 11578 18624
rect 12526 18572 12532 18624
rect 12584 18572 12590 18624
rect 13449 18615 13507 18621
rect 13449 18581 13461 18615
rect 13495 18612 13507 18615
rect 13538 18612 13544 18624
rect 13495 18584 13544 18612
rect 13495 18581 13507 18584
rect 13449 18575 13507 18581
rect 13538 18572 13544 18584
rect 13596 18572 13602 18624
rect 1104 18522 14696 18544
rect 1104 18470 4308 18522
rect 4360 18470 4372 18522
rect 4424 18470 4436 18522
rect 4488 18470 4500 18522
rect 4552 18470 4564 18522
rect 4616 18470 7666 18522
rect 7718 18470 7730 18522
rect 7782 18470 7794 18522
rect 7846 18470 7858 18522
rect 7910 18470 7922 18522
rect 7974 18470 11024 18522
rect 11076 18470 11088 18522
rect 11140 18470 11152 18522
rect 11204 18470 11216 18522
rect 11268 18470 11280 18522
rect 11332 18470 14382 18522
rect 14434 18470 14446 18522
rect 14498 18470 14510 18522
rect 14562 18470 14574 18522
rect 14626 18470 14638 18522
rect 14690 18470 14696 18522
rect 1104 18448 14696 18470
rect 5902 18368 5908 18420
rect 5960 18368 5966 18420
rect 6641 18411 6699 18417
rect 6641 18377 6653 18411
rect 6687 18408 6699 18411
rect 6730 18408 6736 18420
rect 6687 18380 6736 18408
rect 6687 18377 6699 18380
rect 6641 18371 6699 18377
rect 6730 18368 6736 18380
rect 6788 18368 6794 18420
rect 6914 18368 6920 18420
rect 6972 18368 6978 18420
rect 7006 18368 7012 18420
rect 7064 18368 7070 18420
rect 11974 18408 11980 18420
rect 8128 18380 11980 18408
rect 1673 18343 1731 18349
rect 1673 18309 1685 18343
rect 1719 18340 1731 18343
rect 3694 18340 3700 18352
rect 1719 18312 3700 18340
rect 1719 18309 1731 18312
rect 1673 18303 1731 18309
rect 3694 18300 3700 18312
rect 3752 18300 3758 18352
rect 4982 18300 4988 18352
rect 5040 18300 5046 18352
rect 6178 18300 6184 18352
rect 6236 18340 6242 18352
rect 7024 18340 7052 18368
rect 8128 18340 8156 18380
rect 11974 18368 11980 18380
rect 12032 18368 12038 18420
rect 12069 18411 12127 18417
rect 12069 18377 12081 18411
rect 12115 18408 12127 18411
rect 15010 18408 15016 18420
rect 12115 18380 15016 18408
rect 12115 18377 12127 18380
rect 12069 18371 12127 18377
rect 15010 18368 15016 18380
rect 15068 18368 15074 18420
rect 11793 18343 11851 18349
rect 11793 18340 11805 18343
rect 6236 18312 6592 18340
rect 7024 18312 8156 18340
rect 8220 18312 11805 18340
rect 6236 18300 6242 18312
rect 1486 18232 1492 18284
rect 1544 18232 1550 18284
rect 2958 18232 2964 18284
rect 3016 18272 3022 18284
rect 4798 18281 4804 18284
rect 4781 18275 4804 18281
rect 4781 18272 4793 18275
rect 3016 18244 4793 18272
rect 3016 18232 3022 18244
rect 4781 18241 4793 18244
rect 4781 18235 4804 18241
rect 4798 18232 4804 18235
rect 4856 18232 4862 18284
rect 5000 18272 5028 18300
rect 5000 18244 6316 18272
rect 474 18164 480 18216
rect 532 18204 538 18216
rect 4154 18204 4160 18216
rect 532 18176 4160 18204
rect 532 18164 538 18176
rect 4154 18164 4160 18176
rect 4212 18204 4218 18216
rect 4525 18207 4583 18213
rect 4525 18204 4537 18207
rect 4212 18176 4537 18204
rect 4212 18164 4218 18176
rect 4525 18173 4537 18176
rect 4571 18173 4583 18207
rect 4525 18167 4583 18173
rect 6288 18136 6316 18244
rect 6362 18232 6368 18284
rect 6420 18272 6426 18284
rect 6457 18275 6515 18281
rect 6457 18272 6469 18275
rect 6420 18244 6469 18272
rect 6420 18232 6426 18244
rect 6457 18241 6469 18244
rect 6503 18241 6515 18275
rect 6564 18272 6592 18312
rect 6641 18275 6699 18281
rect 6641 18272 6653 18275
rect 6564 18244 6653 18272
rect 6457 18235 6515 18241
rect 6641 18241 6653 18244
rect 6687 18241 6699 18275
rect 6641 18235 6699 18241
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18272 6883 18275
rect 7466 18272 7472 18284
rect 6871 18244 7472 18272
rect 6871 18241 6883 18244
rect 6825 18235 6883 18241
rect 7466 18232 7472 18244
rect 7524 18232 7530 18284
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 8220 18204 8248 18312
rect 11793 18309 11805 18312
rect 11839 18309 11851 18343
rect 11793 18303 11851 18309
rect 8294 18232 8300 18284
rect 8352 18232 8358 18284
rect 10043 18275 10101 18281
rect 10043 18241 10055 18275
rect 10089 18272 10101 18275
rect 10686 18272 10692 18284
rect 10089 18244 10692 18272
rect 10089 18241 10101 18244
rect 10043 18235 10101 18241
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 11333 18275 11391 18281
rect 11333 18241 11345 18275
rect 11379 18241 11391 18275
rect 11333 18235 11391 18241
rect 7340 18176 8248 18204
rect 7340 18164 7346 18176
rect 8312 18136 8340 18232
rect 9674 18164 9680 18216
rect 9732 18204 9738 18216
rect 9769 18207 9827 18213
rect 9769 18204 9781 18207
rect 9732 18176 9781 18204
rect 9732 18164 9738 18176
rect 9769 18173 9781 18176
rect 9815 18173 9827 18207
rect 9769 18167 9827 18173
rect 11348 18136 11376 18235
rect 11698 18232 11704 18284
rect 11756 18272 11762 18284
rect 12342 18272 12348 18284
rect 11756 18244 12348 18272
rect 11756 18232 11762 18244
rect 12342 18232 12348 18244
rect 12400 18232 12406 18284
rect 13446 18281 13452 18284
rect 13403 18275 13452 18281
rect 13403 18241 13415 18275
rect 13449 18241 13452 18275
rect 13403 18235 13452 18241
rect 13446 18232 13452 18235
rect 13504 18232 13510 18284
rect 13538 18232 13544 18284
rect 13596 18232 13602 18284
rect 11790 18164 11796 18216
rect 11848 18204 11854 18216
rect 12529 18207 12587 18213
rect 12529 18204 12541 18207
rect 11848 18176 12541 18204
rect 11848 18164 11854 18176
rect 12529 18173 12541 18176
rect 12575 18173 12587 18207
rect 12529 18167 12587 18173
rect 12618 18164 12624 18216
rect 12676 18204 12682 18216
rect 12989 18207 13047 18213
rect 12989 18204 13001 18207
rect 12676 18176 13001 18204
rect 12676 18164 12682 18176
rect 12989 18173 13001 18176
rect 13035 18173 13047 18207
rect 13265 18207 13323 18213
rect 13265 18204 13277 18207
rect 12989 18167 13047 18173
rect 13121 18176 13277 18204
rect 13121 18136 13149 18176
rect 13265 18173 13277 18176
rect 13311 18173 13323 18207
rect 13265 18167 13323 18173
rect 13906 18164 13912 18216
rect 13964 18204 13970 18216
rect 14185 18207 14243 18213
rect 14185 18204 14197 18207
rect 13964 18176 14197 18204
rect 13964 18164 13970 18176
rect 14185 18173 14197 18176
rect 14231 18173 14243 18207
rect 14185 18167 14243 18173
rect 6288 18108 8340 18136
rect 10428 18108 11376 18136
rect 13004 18108 13149 18136
rect 4154 18028 4160 18080
rect 4212 18068 4218 18080
rect 5626 18068 5632 18080
rect 4212 18040 5632 18068
rect 4212 18028 4218 18040
rect 5626 18028 5632 18040
rect 5684 18028 5690 18080
rect 6086 18028 6092 18080
rect 6144 18068 6150 18080
rect 9030 18068 9036 18080
rect 6144 18040 9036 18068
rect 6144 18028 6150 18040
rect 9030 18028 9036 18040
rect 9088 18068 9094 18080
rect 10428 18068 10456 18108
rect 9088 18040 10456 18068
rect 9088 18028 9094 18040
rect 10778 18028 10784 18080
rect 10836 18028 10842 18080
rect 11146 18028 11152 18080
rect 11204 18028 11210 18080
rect 12434 18028 12440 18080
rect 12492 18068 12498 18080
rect 13004 18068 13032 18108
rect 12492 18040 13032 18068
rect 12492 18028 12498 18040
rect 1104 17978 14536 18000
rect 1104 17926 2629 17978
rect 2681 17926 2693 17978
rect 2745 17926 2757 17978
rect 2809 17926 2821 17978
rect 2873 17926 2885 17978
rect 2937 17926 5987 17978
rect 6039 17926 6051 17978
rect 6103 17926 6115 17978
rect 6167 17926 6179 17978
rect 6231 17926 6243 17978
rect 6295 17926 9345 17978
rect 9397 17926 9409 17978
rect 9461 17926 9473 17978
rect 9525 17926 9537 17978
rect 9589 17926 9601 17978
rect 9653 17926 12703 17978
rect 12755 17926 12767 17978
rect 12819 17926 12831 17978
rect 12883 17926 12895 17978
rect 12947 17926 12959 17978
rect 13011 17926 14536 17978
rect 1104 17904 14536 17926
rect 6089 17867 6147 17873
rect 6089 17833 6101 17867
rect 6135 17864 6147 17867
rect 6362 17864 6368 17876
rect 6135 17836 6368 17864
rect 6135 17833 6147 17836
rect 6089 17827 6147 17833
rect 6362 17824 6368 17836
rect 6420 17824 6426 17876
rect 8846 17824 8852 17876
rect 8904 17864 8910 17876
rect 11517 17867 11575 17873
rect 8904 17836 11468 17864
rect 8904 17824 8910 17836
rect 11146 17796 11152 17808
rect 10704 17768 11152 17796
rect 1394 17620 1400 17672
rect 1452 17660 1458 17672
rect 1671 17663 1729 17669
rect 1452 17632 1624 17660
rect 1452 17620 1458 17632
rect 1596 17592 1624 17632
rect 1671 17629 1683 17663
rect 1717 17660 1729 17663
rect 2038 17660 2044 17672
rect 1717 17632 2044 17660
rect 1717 17629 1729 17632
rect 1671 17623 1729 17629
rect 2038 17620 2044 17632
rect 2096 17620 2102 17672
rect 5077 17663 5135 17669
rect 5077 17629 5089 17663
rect 5123 17629 5135 17663
rect 5350 17660 5356 17672
rect 5311 17632 5356 17660
rect 5077 17623 5135 17629
rect 3050 17592 3056 17604
rect 1596 17564 3056 17592
rect 3050 17552 3056 17564
rect 3108 17592 3114 17604
rect 5092 17592 5120 17623
rect 5350 17620 5356 17632
rect 5408 17620 5414 17672
rect 6454 17620 6460 17672
rect 6512 17620 6518 17672
rect 10704 17669 10732 17768
rect 11146 17756 11152 17768
rect 11204 17756 11210 17808
rect 11440 17796 11468 17836
rect 11517 17833 11529 17867
rect 11563 17864 11575 17867
rect 12066 17864 12072 17876
rect 11563 17836 12072 17864
rect 11563 17833 11575 17836
rect 11517 17827 11575 17833
rect 12066 17824 12072 17836
rect 12124 17824 12130 17876
rect 12618 17824 12624 17876
rect 12676 17864 12682 17876
rect 12713 17867 12771 17873
rect 12713 17864 12725 17867
rect 12676 17836 12725 17864
rect 12676 17824 12682 17836
rect 12713 17833 12725 17836
rect 12759 17833 12771 17867
rect 12713 17827 12771 17833
rect 11440 17768 11744 17796
rect 11716 17672 11744 17768
rect 13078 17756 13084 17808
rect 13136 17756 13142 17808
rect 12618 17688 12624 17740
rect 12676 17728 12682 17740
rect 13096 17728 13124 17756
rect 12676 17700 13124 17728
rect 12676 17688 12682 17700
rect 6731 17663 6789 17669
rect 6731 17629 6743 17663
rect 6777 17660 6789 17663
rect 10505 17663 10563 17669
rect 6777 17632 6960 17660
rect 6777 17629 6789 17632
rect 6731 17623 6789 17629
rect 6472 17592 6500 17620
rect 6932 17604 6960 17632
rect 10505 17629 10517 17663
rect 10551 17629 10563 17663
rect 10505 17623 10563 17629
rect 10689 17663 10747 17669
rect 10689 17629 10701 17663
rect 10735 17629 10747 17663
rect 10689 17623 10747 17629
rect 10781 17663 10839 17669
rect 10781 17629 10793 17663
rect 10827 17660 10839 17663
rect 10870 17660 10876 17672
rect 10827 17632 10876 17660
rect 10827 17629 10839 17632
rect 10781 17623 10839 17629
rect 3108 17564 6500 17592
rect 3108 17552 3114 17564
rect 6914 17552 6920 17604
rect 6972 17552 6978 17604
rect 10520 17592 10548 17623
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17660 11299 17663
rect 11422 17660 11428 17672
rect 11287 17632 11428 17660
rect 11287 17629 11299 17632
rect 11241 17623 11299 17629
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 11698 17620 11704 17672
rect 11756 17620 11762 17672
rect 11943 17663 12001 17669
rect 11943 17660 11955 17663
rect 11806 17632 11955 17660
rect 11806 17592 11834 17632
rect 11943 17629 11955 17632
rect 11989 17629 12001 17663
rect 11943 17623 12001 17629
rect 13078 17620 13084 17672
rect 13136 17620 13142 17672
rect 13170 17620 13176 17672
rect 13228 17660 13234 17672
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 13228 17632 13369 17660
rect 13228 17620 13234 17632
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 13357 17623 13415 17629
rect 10520 17564 11468 17592
rect 10796 17536 10824 17564
rect 11440 17536 11468 17564
rect 11716 17564 11834 17592
rect 11716 17536 11744 17564
rect 2406 17484 2412 17536
rect 2464 17484 2470 17536
rect 7466 17484 7472 17536
rect 7524 17484 7530 17536
rect 7926 17484 7932 17536
rect 7984 17524 7990 17536
rect 8478 17524 8484 17536
rect 7984 17496 8484 17524
rect 7984 17484 7990 17496
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 9674 17484 9680 17536
rect 9732 17524 9738 17536
rect 10597 17527 10655 17533
rect 10597 17524 10609 17527
rect 9732 17496 10609 17524
rect 9732 17484 9738 17496
rect 10597 17493 10609 17496
rect 10643 17493 10655 17527
rect 10597 17487 10655 17493
rect 10778 17484 10784 17536
rect 10836 17484 10842 17536
rect 10870 17484 10876 17536
rect 10928 17484 10934 17536
rect 11422 17484 11428 17536
rect 11480 17484 11486 17536
rect 11698 17484 11704 17536
rect 11756 17484 11762 17536
rect 1104 17434 14696 17456
rect 1104 17382 4308 17434
rect 4360 17382 4372 17434
rect 4424 17382 4436 17434
rect 4488 17382 4500 17434
rect 4552 17382 4564 17434
rect 4616 17382 7666 17434
rect 7718 17382 7730 17434
rect 7782 17382 7794 17434
rect 7846 17382 7858 17434
rect 7910 17382 7922 17434
rect 7974 17382 11024 17434
rect 11076 17382 11088 17434
rect 11140 17382 11152 17434
rect 11204 17382 11216 17434
rect 11268 17382 11280 17434
rect 11332 17382 14382 17434
rect 14434 17382 14446 17434
rect 14498 17382 14510 17434
rect 14562 17382 14574 17434
rect 14626 17382 14638 17434
rect 14690 17382 14696 17434
rect 1104 17360 14696 17382
rect 2406 17280 2412 17332
rect 2464 17280 2470 17332
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 8478 17320 8484 17332
rect 7892 17292 8484 17320
rect 7892 17280 7898 17292
rect 8478 17280 8484 17292
rect 8536 17280 8542 17332
rect 8662 17280 8668 17332
rect 8720 17280 8726 17332
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 9766 17320 9772 17332
rect 8904 17292 9772 17320
rect 8904 17280 8910 17292
rect 9766 17280 9772 17292
rect 9824 17320 9830 17332
rect 9824 17292 10806 17320
rect 9824 17280 9830 17292
rect 750 17144 756 17196
rect 808 17184 814 17196
rect 1489 17187 1547 17193
rect 1489 17184 1501 17187
rect 808 17156 1501 17184
rect 808 17144 814 17156
rect 1489 17153 1501 17156
rect 1535 17153 1547 17187
rect 1489 17147 1547 17153
rect 1949 17187 2007 17193
rect 1949 17153 1961 17187
rect 1995 17184 2007 17187
rect 2424 17184 2452 17280
rect 9582 17252 9588 17264
rect 8588 17224 9588 17252
rect 7190 17184 7196 17196
rect 1995 17156 2452 17184
rect 5184 17156 7196 17184
rect 1995 17153 2007 17156
rect 1949 17147 2007 17153
rect 1673 17119 1731 17125
rect 1673 17085 1685 17119
rect 1719 17085 1731 17119
rect 1673 17079 1731 17085
rect 1688 17048 1716 17079
rect 1854 17076 1860 17128
rect 1912 17116 1918 17128
rect 2130 17116 2136 17128
rect 1912 17088 2136 17116
rect 1912 17076 1918 17088
rect 2130 17076 2136 17088
rect 2188 17076 2194 17128
rect 5184 17048 5212 17156
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 7834 17144 7840 17196
rect 7892 17193 7898 17196
rect 7892 17187 7920 17193
rect 7908 17153 7920 17187
rect 7892 17147 7920 17153
rect 7892 17144 7898 17147
rect 5258 17076 5264 17128
rect 5316 17116 5322 17128
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 5316 17088 6837 17116
rect 5316 17076 5322 17088
rect 6825 17085 6837 17088
rect 6871 17116 6883 17119
rect 7009 17119 7067 17125
rect 6871 17088 6960 17116
rect 6871 17085 6883 17088
rect 6825 17079 6883 17085
rect 1688 17020 5212 17048
rect 1486 16940 1492 16992
rect 1544 16980 1550 16992
rect 1765 16983 1823 16989
rect 1765 16980 1777 16983
rect 1544 16952 1777 16980
rect 1544 16940 1550 16952
rect 1765 16949 1777 16952
rect 1811 16949 1823 16983
rect 6932 16980 6960 17088
rect 7009 17085 7021 17119
rect 7055 17116 7067 17119
rect 7098 17116 7104 17128
rect 7055 17088 7104 17116
rect 7055 17085 7067 17088
rect 7009 17079 7067 17085
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 7466 17076 7472 17128
rect 7524 17076 7530 17128
rect 7745 17119 7803 17125
rect 7745 17116 7757 17119
rect 7576 17088 7757 17116
rect 7374 17008 7380 17060
rect 7432 17048 7438 17060
rect 7576 17048 7604 17088
rect 7745 17085 7757 17088
rect 7791 17085 7803 17119
rect 7745 17079 7803 17085
rect 8018 17076 8024 17128
rect 8076 17076 8082 17128
rect 8386 17076 8392 17128
rect 8444 17116 8450 17128
rect 8588 17116 8616 17224
rect 9582 17212 9588 17224
rect 9640 17212 9646 17264
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 10778 17252 10806 17292
rect 11330 17280 11336 17332
rect 11388 17320 11394 17332
rect 11388 17292 13584 17320
rect 11388 17280 11394 17292
rect 13556 17264 13584 17292
rect 13722 17280 13728 17332
rect 13780 17320 13786 17332
rect 14093 17323 14151 17329
rect 14093 17320 14105 17323
rect 13780 17292 14105 17320
rect 13780 17280 13786 17292
rect 14093 17289 14105 17292
rect 14139 17289 14151 17323
rect 14093 17283 14151 17289
rect 11793 17255 11851 17261
rect 9732 17224 10732 17252
rect 10778 17224 11652 17252
rect 9732 17212 9738 17224
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 8999 17187 9057 17193
rect 8999 17184 9011 17187
rect 8720 17156 9011 17184
rect 8720 17144 8726 17156
rect 8999 17153 9011 17156
rect 9045 17153 9057 17187
rect 8999 17147 9057 17153
rect 10410 17144 10416 17196
rect 10468 17144 10474 17196
rect 10502 17144 10508 17196
rect 10560 17144 10566 17196
rect 8757 17119 8815 17125
rect 8757 17116 8769 17119
rect 8444 17088 8769 17116
rect 8444 17076 8450 17088
rect 8757 17085 8769 17088
rect 8803 17085 8815 17119
rect 8757 17079 8815 17085
rect 10042 17076 10048 17128
rect 10100 17076 10106 17128
rect 7432 17020 7604 17048
rect 7432 17008 7438 17020
rect 9674 16980 9680 16992
rect 6932 16952 9680 16980
rect 1765 16943 1823 16949
rect 9674 16940 9680 16952
rect 9732 16940 9738 16992
rect 9766 16940 9772 16992
rect 9824 16940 9830 16992
rect 10060 16980 10088 17076
rect 10428 17048 10456 17144
rect 10704 17116 10732 17224
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17184 10839 17187
rect 11146 17184 11152 17196
rect 10827 17156 11152 17184
rect 10827 17153 10839 17156
rect 10781 17147 10839 17153
rect 11146 17144 11152 17156
rect 11204 17144 11210 17196
rect 11241 17187 11299 17193
rect 11241 17153 11253 17187
rect 11287 17184 11299 17187
rect 11330 17184 11336 17196
rect 11287 17156 11336 17184
rect 11287 17153 11299 17156
rect 11241 17147 11299 17153
rect 11330 17144 11336 17156
rect 11388 17144 11394 17196
rect 11422 17144 11428 17196
rect 11480 17184 11486 17196
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11480 17156 11529 17184
rect 11480 17144 11486 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11624 17184 11652 17224
rect 11793 17221 11805 17255
rect 11839 17252 11851 17255
rect 12069 17255 12127 17261
rect 12069 17252 12081 17255
rect 11839 17224 12081 17252
rect 11839 17221 11851 17224
rect 11793 17215 11851 17221
rect 12069 17221 12081 17224
rect 12115 17221 12127 17255
rect 12069 17215 12127 17221
rect 13538 17212 13544 17264
rect 13596 17212 13602 17264
rect 12771 17187 12829 17193
rect 12771 17184 12783 17187
rect 11624 17156 12783 17184
rect 11517 17147 11575 17153
rect 12771 17153 12783 17156
rect 12817 17153 12829 17187
rect 12771 17147 12829 17153
rect 13998 17144 14004 17196
rect 14056 17144 14062 17196
rect 10704 17088 10916 17116
rect 10888 17048 10916 17088
rect 10962 17076 10968 17128
rect 11020 17116 11026 17128
rect 11609 17119 11667 17125
rect 11609 17116 11621 17119
rect 11020 17088 11621 17116
rect 11020 17076 11026 17088
rect 11609 17085 11621 17088
rect 11655 17085 11667 17119
rect 11609 17079 11667 17085
rect 11793 17119 11851 17125
rect 11793 17085 11805 17119
rect 11839 17085 11851 17119
rect 11793 17079 11851 17085
rect 11808 17048 11836 17079
rect 12066 17076 12072 17128
rect 12124 17076 12130 17128
rect 12342 17076 12348 17128
rect 12400 17076 12406 17128
rect 12526 17076 12532 17128
rect 12584 17076 12590 17128
rect 13906 17076 13912 17128
rect 13964 17116 13970 17128
rect 15562 17116 15568 17128
rect 13964 17088 15568 17116
rect 13964 17076 13970 17088
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 10428 17020 10806 17048
rect 10888 17020 11836 17048
rect 12084 17048 12112 17076
rect 12544 17048 12572 17076
rect 12084 17020 12572 17048
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10060 16952 10701 16980
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10778 16980 10806 17020
rect 10965 16983 11023 16989
rect 10965 16980 10977 16983
rect 10778 16952 10977 16980
rect 10689 16943 10747 16949
rect 10965 16949 10977 16952
rect 11011 16949 11023 16983
rect 10965 16943 11023 16949
rect 11054 16940 11060 16992
rect 11112 16940 11118 16992
rect 11238 16940 11244 16992
rect 11296 16980 11302 16992
rect 12250 16980 12256 16992
rect 11296 16952 12256 16980
rect 11296 16940 11302 16952
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 12526 16940 12532 16992
rect 12584 16980 12590 16992
rect 12986 16980 12992 16992
rect 12584 16952 12992 16980
rect 12584 16940 12590 16952
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 13446 16940 13452 16992
rect 13504 16980 13510 16992
rect 13541 16983 13599 16989
rect 13541 16980 13553 16983
rect 13504 16952 13553 16980
rect 13504 16940 13510 16952
rect 13541 16949 13553 16952
rect 13587 16949 13599 16983
rect 13541 16943 13599 16949
rect 1104 16890 14536 16912
rect 1104 16838 2629 16890
rect 2681 16838 2693 16890
rect 2745 16838 2757 16890
rect 2809 16838 2821 16890
rect 2873 16838 2885 16890
rect 2937 16838 5987 16890
rect 6039 16838 6051 16890
rect 6103 16838 6115 16890
rect 6167 16838 6179 16890
rect 6231 16838 6243 16890
rect 6295 16838 9345 16890
rect 9397 16838 9409 16890
rect 9461 16838 9473 16890
rect 9525 16838 9537 16890
rect 9589 16838 9601 16890
rect 9653 16838 12703 16890
rect 12755 16838 12767 16890
rect 12819 16838 12831 16890
rect 12883 16838 12895 16890
rect 12947 16838 12959 16890
rect 13011 16838 14536 16890
rect 1104 16816 14536 16838
rect 1581 16779 1639 16785
rect 1581 16745 1593 16779
rect 1627 16776 1639 16779
rect 7745 16779 7803 16785
rect 1627 16748 7696 16776
rect 1627 16745 1639 16748
rect 1581 16739 1639 16745
rect 6454 16600 6460 16652
rect 6512 16640 6518 16652
rect 6733 16643 6791 16649
rect 6733 16640 6745 16643
rect 6512 16612 6745 16640
rect 6512 16600 6518 16612
rect 6733 16609 6745 16612
rect 6779 16609 6791 16643
rect 7668 16640 7696 16748
rect 7745 16745 7757 16779
rect 7791 16776 7803 16779
rect 8018 16776 8024 16788
rect 7791 16748 8024 16776
rect 7791 16745 7803 16748
rect 7745 16739 7803 16745
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 8478 16736 8484 16788
rect 8536 16776 8542 16788
rect 8536 16748 9674 16776
rect 8536 16736 8542 16748
rect 8846 16640 8852 16652
rect 7668 16612 8852 16640
rect 6733 16603 6791 16609
rect 3418 16532 3424 16584
rect 3476 16572 3482 16584
rect 4890 16572 4896 16584
rect 3476 16544 4896 16572
rect 3476 16532 3482 16544
rect 4890 16532 4896 16544
rect 4948 16532 4954 16584
rect 750 16464 756 16516
rect 808 16504 814 16516
rect 1489 16507 1547 16513
rect 1489 16504 1501 16507
rect 808 16476 1501 16504
rect 808 16464 814 16476
rect 1489 16473 1501 16476
rect 1535 16473 1547 16507
rect 1489 16467 1547 16473
rect 3510 16464 3516 16516
rect 3568 16464 3574 16516
rect 6748 16504 6776 16603
rect 8846 16600 8852 16612
rect 8904 16600 8910 16652
rect 9214 16600 9220 16652
rect 9272 16600 9278 16652
rect 9401 16643 9459 16649
rect 9401 16609 9413 16643
rect 9447 16640 9459 16643
rect 9490 16640 9496 16652
rect 9447 16612 9496 16640
rect 9447 16609 9459 16612
rect 9401 16603 9459 16609
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 9646 16640 9674 16748
rect 9766 16736 9772 16788
rect 9824 16776 9830 16788
rect 11057 16779 11115 16785
rect 9824 16748 9904 16776
rect 9824 16736 9830 16748
rect 9876 16717 9904 16748
rect 9968 16748 11008 16776
rect 9861 16711 9919 16717
rect 9861 16677 9873 16711
rect 9907 16677 9919 16711
rect 9861 16671 9919 16677
rect 9968 16640 9996 16748
rect 10870 16668 10876 16720
rect 10928 16668 10934 16720
rect 10980 16708 11008 16748
rect 11057 16745 11069 16779
rect 11103 16776 11115 16779
rect 11606 16776 11612 16788
rect 11103 16748 11612 16776
rect 11103 16745 11115 16748
rect 11057 16739 11115 16745
rect 11606 16736 11612 16748
rect 11664 16736 11670 16788
rect 11974 16736 11980 16788
rect 12032 16776 12038 16788
rect 12710 16776 12716 16788
rect 12032 16748 12716 16776
rect 12032 16736 12038 16748
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 13170 16776 13176 16788
rect 12820 16748 13176 16776
rect 11238 16708 11244 16720
rect 10980 16680 11244 16708
rect 11238 16668 11244 16680
rect 11296 16668 11302 16720
rect 11333 16711 11391 16717
rect 11333 16677 11345 16711
rect 11379 16708 11391 16711
rect 12526 16708 12532 16720
rect 11379 16680 12532 16708
rect 11379 16677 11391 16680
rect 11333 16671 11391 16677
rect 12526 16668 12532 16680
rect 12584 16668 12590 16720
rect 9646 16612 9996 16640
rect 10275 16643 10333 16649
rect 10275 16609 10287 16643
rect 10321 16640 10333 16643
rect 10594 16640 10600 16652
rect 10321 16612 10600 16640
rect 10321 16609 10333 16612
rect 10275 16603 10333 16609
rect 10594 16600 10600 16612
rect 10652 16640 10658 16652
rect 10888 16640 10916 16668
rect 10652 16612 10916 16640
rect 12069 16643 12127 16649
rect 10652 16600 10658 16612
rect 12069 16609 12081 16643
rect 12115 16640 12127 16643
rect 12158 16640 12164 16652
rect 12115 16612 12164 16640
rect 12115 16609 12127 16612
rect 12069 16603 12127 16609
rect 12158 16600 12164 16612
rect 12216 16600 12222 16652
rect 12710 16600 12716 16652
rect 12768 16600 12774 16652
rect 12820 16640 12848 16748
rect 13170 16736 13176 16748
rect 13228 16736 13234 16788
rect 13814 16736 13820 16788
rect 13872 16776 13878 16788
rect 13909 16779 13967 16785
rect 13909 16776 13921 16779
rect 13872 16748 13921 16776
rect 13872 16736 13878 16748
rect 13909 16745 13921 16748
rect 13955 16745 13967 16779
rect 13909 16739 13967 16745
rect 12989 16643 13047 16649
rect 12989 16640 13001 16643
rect 12820 16612 13001 16640
rect 12989 16609 13001 16612
rect 13035 16609 13047 16643
rect 12989 16603 13047 16609
rect 13265 16643 13323 16649
rect 13265 16609 13277 16643
rect 13311 16640 13323 16643
rect 13446 16640 13452 16652
rect 13311 16612 13452 16640
rect 13311 16609 13323 16612
rect 13265 16603 13323 16609
rect 13446 16600 13452 16612
rect 13504 16600 13510 16652
rect 7007 16575 7065 16581
rect 7007 16541 7019 16575
rect 7053 16572 7065 16575
rect 9582 16572 9588 16584
rect 7053 16544 9588 16572
rect 7053 16541 7065 16544
rect 7007 16535 7065 16541
rect 9582 16532 9588 16544
rect 9640 16532 9646 16584
rect 10134 16532 10140 16584
rect 10192 16532 10198 16584
rect 10410 16532 10416 16584
rect 10468 16532 10474 16584
rect 11146 16532 11152 16584
rect 11204 16532 11210 16584
rect 11425 16575 11483 16581
rect 11425 16541 11437 16575
rect 11471 16572 11483 16575
rect 11882 16572 11888 16584
rect 11471 16544 11888 16572
rect 11471 16541 11483 16544
rect 11425 16535 11483 16541
rect 11882 16532 11888 16544
rect 11940 16532 11946 16584
rect 13170 16581 13176 16584
rect 12253 16575 12311 16581
rect 12253 16541 12265 16575
rect 12299 16541 12311 16575
rect 12253 16535 12311 16541
rect 13127 16575 13176 16581
rect 13127 16541 13139 16575
rect 13173 16541 13176 16575
rect 13127 16535 13176 16541
rect 8386 16504 8392 16516
rect 6748 16476 8392 16504
rect 8386 16464 8392 16476
rect 8444 16464 8450 16516
rect 11793 16507 11851 16513
rect 11440 16476 11744 16504
rect 3528 16436 3556 16464
rect 11440 16448 11468 16476
rect 8662 16436 8668 16448
rect 3528 16408 8668 16436
rect 8662 16396 8668 16408
rect 8720 16396 8726 16448
rect 10226 16396 10232 16448
rect 10284 16436 10290 16448
rect 11422 16436 11428 16448
rect 10284 16408 11428 16436
rect 10284 16396 10290 16408
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 11606 16396 11612 16448
rect 11664 16396 11670 16448
rect 11716 16436 11744 16476
rect 11793 16473 11805 16507
rect 11839 16504 11851 16507
rect 11839 16476 12112 16504
rect 11839 16473 11851 16476
rect 11793 16467 11851 16473
rect 11885 16439 11943 16445
rect 11885 16436 11897 16439
rect 11716 16408 11897 16436
rect 11885 16405 11897 16408
rect 11931 16405 11943 16439
rect 12084 16436 12112 16476
rect 12158 16464 12164 16516
rect 12216 16504 12222 16516
rect 12268 16504 12296 16535
rect 13170 16532 13176 16535
rect 13228 16532 13234 16584
rect 12216 16476 12296 16504
rect 12216 16464 12222 16476
rect 13814 16436 13820 16448
rect 12084 16408 13820 16436
rect 11885 16399 11943 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 1104 16346 14696 16368
rect 1104 16294 4308 16346
rect 4360 16294 4372 16346
rect 4424 16294 4436 16346
rect 4488 16294 4500 16346
rect 4552 16294 4564 16346
rect 4616 16294 7666 16346
rect 7718 16294 7730 16346
rect 7782 16294 7794 16346
rect 7846 16294 7858 16346
rect 7910 16294 7922 16346
rect 7974 16294 11024 16346
rect 11076 16294 11088 16346
rect 11140 16294 11152 16346
rect 11204 16294 11216 16346
rect 11268 16294 11280 16346
rect 11332 16294 14382 16346
rect 14434 16294 14446 16346
rect 14498 16294 14510 16346
rect 14562 16294 14574 16346
rect 14626 16294 14638 16346
rect 14690 16294 14696 16346
rect 1104 16272 14696 16294
rect 1946 16232 1952 16244
rect 1688 16204 1952 16232
rect 1688 16135 1716 16204
rect 1946 16192 1952 16204
rect 2004 16192 2010 16244
rect 10045 16235 10103 16241
rect 10045 16201 10057 16235
rect 10091 16232 10103 16235
rect 10410 16232 10416 16244
rect 10091 16204 10416 16232
rect 10091 16201 10103 16204
rect 10045 16195 10103 16201
rect 10410 16192 10416 16204
rect 10468 16192 10474 16244
rect 12710 16192 12716 16244
rect 12768 16232 12774 16244
rect 12805 16235 12863 16241
rect 12805 16232 12817 16235
rect 12768 16204 12817 16232
rect 12768 16192 12774 16204
rect 12805 16201 12817 16204
rect 12851 16201 12863 16235
rect 12805 16195 12863 16201
rect 14093 16235 14151 16241
rect 14093 16201 14105 16235
rect 14139 16232 14151 16235
rect 15286 16232 15292 16244
rect 14139 16204 15292 16232
rect 14139 16201 14151 16204
rect 14093 16195 14151 16201
rect 15286 16192 15292 16204
rect 15344 16192 15350 16244
rect 1655 16129 1716 16135
rect 1394 16056 1400 16108
rect 1452 16056 1458 16108
rect 1655 16095 1667 16129
rect 1701 16098 1716 16129
rect 7374 16124 7380 16176
rect 7432 16164 7438 16176
rect 8294 16164 8300 16176
rect 7432 16136 8300 16164
rect 7432 16124 7438 16136
rect 8294 16124 8300 16136
rect 8352 16164 8358 16176
rect 8352 16136 10548 16164
rect 8352 16124 8358 16136
rect 1701 16095 1713 16098
rect 1655 16089 1713 16095
rect 6454 16056 6460 16108
rect 6512 16096 6518 16108
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 6512 16068 6837 16096
rect 6512 16056 6518 16068
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7099 16099 7157 16105
rect 7099 16096 7111 16099
rect 7064 16068 7111 16096
rect 7064 16056 7070 16068
rect 7099 16065 7111 16068
rect 7145 16065 7157 16099
rect 9275 16099 9333 16105
rect 9275 16096 9287 16099
rect 7099 16059 7157 16065
rect 7484 16068 9287 16096
rect 2406 15852 2412 15904
rect 2464 15852 2470 15904
rect 2498 15852 2504 15904
rect 2556 15892 2562 15904
rect 5534 15892 5540 15904
rect 2556 15864 5540 15892
rect 2556 15852 2562 15864
rect 5534 15852 5540 15864
rect 5592 15892 5598 15904
rect 7484 15892 7512 16068
rect 9275 16065 9287 16068
rect 9321 16065 9333 16099
rect 9275 16059 9333 16065
rect 9766 16056 9772 16108
rect 9824 16096 9830 16108
rect 10410 16096 10416 16108
rect 9824 16068 10416 16096
rect 9824 16056 9830 16068
rect 10410 16056 10416 16068
rect 10468 16056 10474 16108
rect 10520 16096 10548 16136
rect 11054 16124 11060 16176
rect 11112 16164 11118 16176
rect 11790 16164 11796 16176
rect 11112 16136 11796 16164
rect 11112 16124 11118 16136
rect 11790 16124 11796 16136
rect 11848 16124 11854 16176
rect 13449 16167 13507 16173
rect 13449 16133 13461 16167
rect 13495 16164 13507 16167
rect 15010 16164 15016 16176
rect 13495 16136 15016 16164
rect 13495 16133 13507 16136
rect 13449 16127 13507 16133
rect 15010 16124 15016 16136
rect 15068 16124 15074 16176
rect 15470 16124 15476 16176
rect 15528 16124 15534 16176
rect 15562 16124 15568 16176
rect 15620 16124 15626 16176
rect 12035 16099 12093 16105
rect 12035 16096 12047 16099
rect 10520 16068 12047 16096
rect 12035 16065 12047 16068
rect 12081 16065 12093 16099
rect 12035 16059 12093 16065
rect 12802 16056 12808 16108
rect 12860 16096 12866 16108
rect 13817 16099 13875 16105
rect 13817 16096 13829 16099
rect 12860 16068 13829 16096
rect 12860 16056 12866 16068
rect 13817 16065 13829 16068
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 9033 16031 9091 16037
rect 9033 16028 9045 16031
rect 8444 16000 9045 16028
rect 8444 15988 8450 16000
rect 9033 15997 9045 16000
rect 9079 15997 9091 16031
rect 9033 15991 9091 15997
rect 11606 15988 11612 16040
rect 11664 16028 11670 16040
rect 11790 16028 11796 16040
rect 11664 16000 11796 16028
rect 11664 15988 11670 16000
rect 11790 15988 11796 16000
rect 11848 15988 11854 16040
rect 15378 15988 15384 16040
rect 15436 16028 15442 16040
rect 15488 16028 15516 16124
rect 15436 16000 15516 16028
rect 15436 15988 15442 16000
rect 15580 15972 15608 16124
rect 15562 15920 15568 15972
rect 15620 15920 15626 15972
rect 5592 15864 7512 15892
rect 7837 15895 7895 15901
rect 5592 15852 5598 15864
rect 7837 15861 7849 15895
rect 7883 15892 7895 15895
rect 8386 15892 8392 15904
rect 7883 15864 8392 15892
rect 7883 15861 7895 15864
rect 7837 15855 7895 15861
rect 8386 15852 8392 15864
rect 8444 15852 8450 15904
rect 10134 15852 10140 15904
rect 10192 15892 10198 15904
rect 13541 15895 13599 15901
rect 13541 15892 13553 15895
rect 10192 15864 13553 15892
rect 10192 15852 10198 15864
rect 13541 15861 13553 15864
rect 13587 15861 13599 15895
rect 13541 15855 13599 15861
rect 1104 15802 14536 15824
rect 1104 15750 2629 15802
rect 2681 15750 2693 15802
rect 2745 15750 2757 15802
rect 2809 15750 2821 15802
rect 2873 15750 2885 15802
rect 2937 15750 5987 15802
rect 6039 15750 6051 15802
rect 6103 15750 6115 15802
rect 6167 15750 6179 15802
rect 6231 15750 6243 15802
rect 6295 15750 9345 15802
rect 9397 15750 9409 15802
rect 9461 15750 9473 15802
rect 9525 15750 9537 15802
rect 9589 15750 9601 15802
rect 9653 15750 12703 15802
rect 12755 15750 12767 15802
rect 12819 15750 12831 15802
rect 12883 15750 12895 15802
rect 12947 15750 12959 15802
rect 13011 15750 14536 15802
rect 1104 15728 14536 15750
rect 6914 15648 6920 15700
rect 6972 15688 6978 15700
rect 7190 15688 7196 15700
rect 6972 15660 7196 15688
rect 6972 15648 6978 15660
rect 7190 15648 7196 15660
rect 7248 15648 7254 15700
rect 11054 15688 11060 15700
rect 10888 15660 11060 15688
rect 1673 15623 1731 15629
rect 1673 15589 1685 15623
rect 1719 15620 1731 15623
rect 7374 15620 7380 15632
rect 1719 15592 7380 15620
rect 1719 15589 1731 15592
rect 1673 15583 1731 15589
rect 7374 15580 7380 15592
rect 7432 15580 7438 15632
rect 9950 15580 9956 15632
rect 10008 15620 10014 15632
rect 10781 15623 10839 15629
rect 10781 15620 10793 15623
rect 10008 15592 10793 15620
rect 10008 15580 10014 15592
rect 10781 15589 10793 15592
rect 10827 15589 10839 15623
rect 10781 15583 10839 15589
rect 6454 15512 6460 15564
rect 6512 15552 6518 15564
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 6512 15524 7481 15552
rect 6512 15512 6518 15524
rect 7469 15521 7481 15524
rect 7515 15521 7527 15555
rect 10321 15555 10379 15561
rect 10321 15552 10333 15555
rect 7469 15515 7527 15521
rect 8864 15524 10333 15552
rect 8864 15496 8892 15524
rect 10321 15521 10333 15524
rect 10367 15552 10379 15555
rect 10888 15552 10916 15660
rect 11054 15648 11060 15660
rect 11112 15648 11118 15700
rect 11698 15648 11704 15700
rect 11756 15648 11762 15700
rect 11977 15691 12035 15697
rect 11977 15657 11989 15691
rect 12023 15688 12035 15691
rect 13906 15688 13912 15700
rect 12023 15660 13912 15688
rect 12023 15657 12035 15660
rect 11977 15651 12035 15657
rect 13906 15648 13912 15660
rect 13964 15648 13970 15700
rect 10367 15524 10916 15552
rect 10367 15521 10379 15524
rect 10321 15515 10379 15521
rect 11054 15512 11060 15564
rect 11112 15512 11118 15564
rect 11333 15555 11391 15561
rect 11333 15521 11345 15555
rect 11379 15552 11391 15555
rect 11514 15552 11520 15564
rect 11379 15524 11520 15552
rect 11379 15521 11391 15524
rect 11333 15515 11391 15521
rect 11514 15512 11520 15524
rect 11572 15512 11578 15564
rect 11716 15552 11744 15648
rect 11882 15580 11888 15632
rect 11940 15620 11946 15632
rect 11940 15592 12112 15620
rect 11940 15580 11946 15592
rect 12084 15564 12112 15592
rect 11716 15524 11928 15552
rect 7374 15484 7380 15496
rect 5644 15456 7380 15484
rect 5644 15428 5672 15456
rect 7374 15444 7380 15456
rect 7432 15484 7438 15496
rect 7711 15487 7769 15493
rect 7711 15484 7723 15487
rect 7432 15456 7723 15484
rect 7432 15444 7438 15456
rect 7711 15453 7723 15456
rect 7757 15453 7769 15487
rect 7711 15447 7769 15453
rect 8846 15444 8852 15496
rect 8904 15444 8910 15496
rect 10134 15444 10140 15496
rect 10192 15444 10198 15496
rect 11146 15444 11152 15496
rect 11204 15493 11210 15496
rect 11204 15487 11232 15493
rect 11220 15453 11232 15487
rect 11900 15484 11928 15524
rect 12066 15512 12072 15564
rect 12124 15512 12130 15564
rect 12311 15487 12369 15493
rect 12311 15484 12323 15487
rect 11900 15456 12323 15484
rect 11204 15447 11232 15453
rect 12311 15453 12323 15456
rect 12357 15453 12369 15487
rect 12311 15447 12369 15453
rect 13725 15487 13783 15493
rect 13725 15453 13737 15487
rect 13771 15484 13783 15487
rect 14642 15484 14648 15496
rect 13771 15456 14648 15484
rect 13771 15453 13783 15456
rect 13725 15447 13783 15453
rect 11204 15444 11210 15447
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 750 15376 756 15428
rect 808 15416 814 15428
rect 1489 15419 1547 15425
rect 1489 15416 1501 15419
rect 808 15388 1501 15416
rect 808 15376 814 15388
rect 1489 15385 1501 15388
rect 1535 15385 1547 15419
rect 1489 15379 1547 15385
rect 5626 15376 5632 15428
rect 5684 15376 5690 15428
rect 8481 15351 8539 15357
rect 8481 15317 8493 15351
rect 8527 15348 8539 15351
rect 9306 15348 9312 15360
rect 8527 15320 9312 15348
rect 8527 15317 8539 15320
rect 8481 15311 8539 15317
rect 9306 15308 9312 15320
rect 9364 15308 9370 15360
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 11146 15348 11152 15360
rect 10284 15320 11152 15348
rect 10284 15308 10290 15320
rect 11146 15308 11152 15320
rect 11204 15348 11210 15360
rect 12158 15348 12164 15360
rect 11204 15320 12164 15348
rect 11204 15308 11210 15320
rect 12158 15308 12164 15320
rect 12216 15308 12222 15360
rect 12986 15308 12992 15360
rect 13044 15348 13050 15360
rect 13081 15351 13139 15357
rect 13081 15348 13093 15351
rect 13044 15320 13093 15348
rect 13044 15308 13050 15320
rect 13081 15317 13093 15320
rect 13127 15317 13139 15351
rect 13081 15311 13139 15317
rect 13814 15308 13820 15360
rect 13872 15308 13878 15360
rect 1104 15258 14696 15280
rect 1104 15206 4308 15258
rect 4360 15206 4372 15258
rect 4424 15206 4436 15258
rect 4488 15206 4500 15258
rect 4552 15206 4564 15258
rect 4616 15206 7666 15258
rect 7718 15206 7730 15258
rect 7782 15206 7794 15258
rect 7846 15206 7858 15258
rect 7910 15206 7922 15258
rect 7974 15206 11024 15258
rect 11076 15206 11088 15258
rect 11140 15206 11152 15258
rect 11204 15206 11216 15258
rect 11268 15206 11280 15258
rect 11332 15206 14382 15258
rect 14434 15206 14446 15258
rect 14498 15206 14510 15258
rect 14562 15206 14574 15258
rect 14626 15206 14638 15258
rect 14690 15206 14696 15258
rect 1104 15184 14696 15206
rect 1302 15104 1308 15156
rect 1360 15144 1366 15156
rect 1360 15116 5304 15144
rect 1360 15104 1366 15116
rect 1486 15036 1492 15088
rect 1544 15036 1550 15088
rect 2406 15036 2412 15088
rect 2464 15036 2470 15088
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 15008 2191 15011
rect 2424 15008 2452 15036
rect 5135 15011 5193 15017
rect 5135 15008 5147 15011
rect 2179 14980 2452 15008
rect 2746 14980 5147 15008
rect 2179 14977 2191 14980
rect 2133 14971 2191 14977
rect 1578 14900 1584 14952
rect 1636 14940 1642 14952
rect 2746 14940 2774 14980
rect 5135 14977 5147 14980
rect 5181 14977 5193 15011
rect 5276 15008 5304 15116
rect 5902 15104 5908 15156
rect 5960 15144 5966 15156
rect 6730 15144 6736 15156
rect 5960 15116 6736 15144
rect 5960 15104 5966 15116
rect 6730 15104 6736 15116
rect 6788 15104 6794 15156
rect 7098 15104 7104 15156
rect 7156 15144 7162 15156
rect 9953 15147 10011 15153
rect 7156 15116 9904 15144
rect 7156 15104 7162 15116
rect 9876 15076 9904 15116
rect 9953 15113 9965 15147
rect 9999 15144 10011 15147
rect 10318 15144 10324 15156
rect 9999 15116 10324 15144
rect 9999 15113 10011 15116
rect 9953 15107 10011 15113
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 11885 15147 11943 15153
rect 11885 15113 11897 15147
rect 11931 15113 11943 15147
rect 11885 15107 11943 15113
rect 14185 15147 14243 15153
rect 14185 15113 14197 15147
rect 14231 15144 14243 15147
rect 15194 15144 15200 15156
rect 14231 15116 15200 15144
rect 14231 15113 14243 15116
rect 14185 15107 14243 15113
rect 10042 15076 10048 15088
rect 9876 15048 10048 15076
rect 10042 15036 10048 15048
rect 10100 15076 10106 15088
rect 11900 15076 11928 15107
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 12342 15076 12348 15088
rect 10100 15048 10732 15076
rect 11900 15048 12348 15076
rect 10100 15036 10106 15048
rect 6607 15011 6665 15017
rect 6607 15008 6619 15011
rect 5276 14980 6619 15008
rect 5135 14971 5193 14977
rect 6607 14977 6619 14980
rect 6653 14977 6665 15011
rect 6607 14971 6665 14977
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 8110 15008 8116 15020
rect 7156 14980 8116 15008
rect 7156 14968 7162 14980
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 9030 14968 9036 15020
rect 9088 14968 9094 15020
rect 9306 14968 9312 15020
rect 9364 14968 9370 15020
rect 10318 15017 10324 15020
rect 10287 15011 10324 15017
rect 10287 14977 10299 15011
rect 10287 14971 10324 14977
rect 10318 14968 10324 14971
rect 10376 14968 10382 15020
rect 1636 14912 2774 14940
rect 4893 14943 4951 14949
rect 1636 14900 1642 14912
rect 4893 14909 4905 14943
rect 4939 14909 4951 14943
rect 6362 14940 6368 14952
rect 4893 14903 4951 14909
rect 5828 14912 6368 14940
rect 842 14764 848 14816
rect 900 14804 906 14816
rect 1581 14807 1639 14813
rect 1581 14804 1593 14807
rect 900 14776 1593 14804
rect 900 14764 906 14776
rect 1581 14773 1593 14776
rect 1627 14773 1639 14807
rect 1581 14767 1639 14773
rect 1946 14764 1952 14816
rect 2004 14764 2010 14816
rect 4908 14804 4936 14903
rect 5828 14804 5856 14912
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 8294 14900 8300 14952
rect 8352 14900 8358 14952
rect 8386 14900 8392 14952
rect 8444 14940 8450 14952
rect 8757 14943 8815 14949
rect 8757 14940 8769 14943
rect 8444 14912 8769 14940
rect 8444 14900 8450 14912
rect 8757 14909 8769 14912
rect 8803 14909 8815 14943
rect 9150 14943 9208 14949
rect 9150 14940 9162 14943
rect 8757 14903 8815 14909
rect 8864 14912 9162 14940
rect 8662 14872 8668 14884
rect 7300 14844 8668 14872
rect 4908 14776 5856 14804
rect 5902 14764 5908 14816
rect 5960 14764 5966 14816
rect 6822 14764 6828 14816
rect 6880 14804 6886 14816
rect 7300 14804 7328 14844
rect 8662 14832 8668 14844
rect 8720 14872 8726 14884
rect 8864 14872 8892 14912
rect 9150 14909 9162 14912
rect 9196 14909 9208 14943
rect 9150 14903 9208 14909
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 10045 14943 10103 14949
rect 10045 14940 10057 14943
rect 9732 14912 10057 14940
rect 9732 14900 9738 14912
rect 10045 14909 10057 14912
rect 10091 14909 10103 14943
rect 10045 14903 10103 14909
rect 8720 14844 8892 14872
rect 10704 14872 10732 15048
rect 12342 15036 12348 15048
rect 12400 15036 12406 15088
rect 11698 14968 11704 15020
rect 11756 14968 11762 15020
rect 12066 14968 12072 15020
rect 12124 14968 12130 15020
rect 12253 15011 12311 15017
rect 12253 14977 12265 15011
rect 12299 15008 12311 15011
rect 12299 14980 12480 15008
rect 12299 14977 12311 14980
rect 12253 14971 12311 14977
rect 12452 14952 12480 14980
rect 12526 14968 12532 15020
rect 12584 14968 12590 15020
rect 13265 15011 13323 15017
rect 13265 14977 13277 15011
rect 13311 14977 13323 15011
rect 13265 14971 13323 14977
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 12345 14943 12403 14949
rect 12345 14940 12357 14943
rect 11112 14912 12357 14940
rect 11112 14900 11118 14912
rect 12345 14909 12357 14912
rect 12391 14909 12403 14943
rect 12345 14903 12403 14909
rect 12434 14900 12440 14952
rect 12492 14900 12498 14952
rect 12986 14900 12992 14952
rect 13044 14900 13050 14952
rect 13280 14940 13308 14971
rect 13096 14912 13308 14940
rect 13096 14872 13124 14912
rect 13354 14900 13360 14952
rect 13412 14949 13418 14952
rect 13412 14943 13440 14949
rect 13428 14909 13440 14943
rect 13412 14903 13440 14909
rect 13412 14900 13418 14903
rect 13538 14900 13544 14952
rect 13596 14900 13602 14952
rect 10704 14844 13124 14872
rect 8720 14832 8726 14844
rect 6880 14776 7328 14804
rect 6880 14764 6886 14776
rect 7374 14764 7380 14816
rect 7432 14764 7438 14816
rect 11057 14807 11115 14813
rect 11057 14773 11069 14807
rect 11103 14804 11115 14807
rect 11330 14804 11336 14816
rect 11103 14776 11336 14804
rect 11103 14773 11115 14776
rect 11057 14767 11115 14773
rect 11330 14764 11336 14776
rect 11388 14764 11394 14816
rect 12066 14764 12072 14816
rect 12124 14804 12130 14816
rect 14366 14804 14372 14816
rect 12124 14776 14372 14804
rect 12124 14764 12130 14776
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 1104 14714 14536 14736
rect 1104 14662 2629 14714
rect 2681 14662 2693 14714
rect 2745 14662 2757 14714
rect 2809 14662 2821 14714
rect 2873 14662 2885 14714
rect 2937 14662 5987 14714
rect 6039 14662 6051 14714
rect 6103 14662 6115 14714
rect 6167 14662 6179 14714
rect 6231 14662 6243 14714
rect 6295 14662 9345 14714
rect 9397 14662 9409 14714
rect 9461 14662 9473 14714
rect 9525 14662 9537 14714
rect 9589 14662 9601 14714
rect 9653 14662 12703 14714
rect 12755 14662 12767 14714
rect 12819 14662 12831 14714
rect 12883 14662 12895 14714
rect 12947 14662 12959 14714
rect 13011 14662 14536 14714
rect 1104 14640 14536 14662
rect 5902 14560 5908 14612
rect 5960 14560 5966 14612
rect 7098 14600 7104 14612
rect 6564 14572 7104 14600
rect 5920 14532 5948 14560
rect 6457 14535 6515 14541
rect 6457 14532 6469 14535
rect 5920 14504 6469 14532
rect 6457 14501 6469 14504
rect 6503 14501 6515 14535
rect 6457 14495 6515 14501
rect 1394 14424 1400 14476
rect 1452 14424 1458 14476
rect 5813 14467 5871 14473
rect 5813 14433 5825 14467
rect 5859 14464 5871 14467
rect 6564 14464 6592 14572
rect 7098 14560 7104 14572
rect 7156 14560 7162 14612
rect 7374 14560 7380 14612
rect 7432 14560 7438 14612
rect 7653 14603 7711 14609
rect 7653 14569 7665 14603
rect 7699 14600 7711 14603
rect 8018 14600 8024 14612
rect 7699 14572 8024 14600
rect 7699 14569 7711 14572
rect 7653 14563 7711 14569
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 8570 14560 8576 14612
rect 8628 14600 8634 14612
rect 10502 14600 10508 14612
rect 8628 14572 10508 14600
rect 8628 14560 8634 14572
rect 10502 14560 10508 14572
rect 10560 14560 10566 14612
rect 10612 14572 13216 14600
rect 5859 14436 6592 14464
rect 5859 14433 5871 14436
rect 5813 14427 5871 14433
rect 6822 14424 6828 14476
rect 6880 14473 6886 14476
rect 6880 14467 6908 14473
rect 6896 14433 6908 14467
rect 6880 14427 6908 14433
rect 7009 14467 7067 14473
rect 7009 14433 7021 14467
rect 7055 14464 7067 14467
rect 7392 14464 7420 14560
rect 7558 14492 7564 14544
rect 7616 14532 7622 14544
rect 7926 14532 7932 14544
rect 7616 14504 7932 14532
rect 7616 14492 7622 14504
rect 7926 14492 7932 14504
rect 7984 14532 7990 14544
rect 9766 14532 9772 14544
rect 7984 14504 9772 14532
rect 7984 14492 7990 14504
rect 9766 14492 9772 14504
rect 9824 14492 9830 14544
rect 10612 14532 10640 14572
rect 10244 14504 10640 14532
rect 11977 14535 12035 14541
rect 9030 14464 9036 14476
rect 7055 14436 7420 14464
rect 7668 14436 9036 14464
rect 7055 14433 7067 14436
rect 7009 14427 7067 14433
rect 6880 14424 6886 14427
rect 1302 14356 1308 14408
rect 1360 14396 1366 14408
rect 1639 14399 1697 14405
rect 1639 14396 1651 14399
rect 1360 14368 1651 14396
rect 1360 14356 1366 14368
rect 1639 14365 1651 14368
rect 1685 14365 1697 14399
rect 1639 14359 1697 14365
rect 5994 14356 6000 14408
rect 6052 14356 6058 14408
rect 6730 14356 6736 14408
rect 6788 14356 6794 14408
rect 7668 14328 7696 14436
rect 9030 14424 9036 14436
rect 9088 14464 9094 14476
rect 10244 14464 10272 14504
rect 11977 14501 11989 14535
rect 12023 14532 12035 14535
rect 12158 14532 12164 14544
rect 12023 14504 12164 14532
rect 12023 14501 12035 14504
rect 11977 14495 12035 14501
rect 12158 14492 12164 14504
rect 12216 14492 12222 14544
rect 13188 14532 13216 14572
rect 13538 14560 13544 14612
rect 13596 14560 13602 14612
rect 13188 14504 13860 14532
rect 13832 14476 13860 14504
rect 9088 14436 10272 14464
rect 9088 14424 9094 14436
rect 10318 14424 10324 14476
rect 10376 14424 10382 14476
rect 10778 14424 10784 14476
rect 10836 14424 10842 14476
rect 11054 14424 11060 14476
rect 11112 14473 11118 14476
rect 11112 14467 11133 14473
rect 11121 14433 11133 14467
rect 11112 14427 11133 14433
rect 11112 14424 11118 14427
rect 12434 14424 12440 14476
rect 12492 14464 12498 14476
rect 12529 14467 12587 14473
rect 12529 14464 12541 14467
rect 12492 14436 12541 14464
rect 12492 14424 12498 14436
rect 12529 14433 12541 14436
rect 12575 14433 12587 14467
rect 12529 14427 12587 14433
rect 13814 14424 13820 14476
rect 13872 14424 13878 14476
rect 10137 14399 10195 14405
rect 10137 14396 10149 14399
rect 7576 14300 7696 14328
rect 8312 14368 10149 14396
rect 2406 14220 2412 14272
rect 2464 14220 2470 14272
rect 6730 14220 6736 14272
rect 6788 14260 6794 14272
rect 7576 14260 7604 14300
rect 6788 14232 7604 14260
rect 6788 14220 6794 14232
rect 7650 14220 7656 14272
rect 7708 14260 7714 14272
rect 8312 14260 8340 14368
rect 10137 14365 10149 14368
rect 10183 14396 10195 14399
rect 10502 14396 10508 14408
rect 10183 14368 10508 14396
rect 10183 14365 10195 14368
rect 10137 14359 10195 14365
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 11238 14405 11244 14408
rect 11195 14399 11244 14405
rect 11195 14365 11207 14399
rect 11241 14365 11244 14399
rect 11195 14359 11244 14365
rect 11238 14356 11244 14359
rect 11296 14356 11302 14408
rect 11330 14356 11336 14408
rect 11388 14356 11394 14408
rect 12279 14399 12337 14405
rect 12279 14365 12291 14399
rect 12325 14396 12337 14399
rect 12803 14399 12861 14405
rect 12325 14368 12756 14396
rect 12325 14365 12337 14368
rect 12279 14359 12337 14365
rect 8386 14288 8392 14340
rect 8444 14328 8450 14340
rect 8570 14328 8576 14340
rect 8444 14300 8576 14328
rect 8444 14288 8450 14300
rect 8570 14288 8576 14300
rect 8628 14328 8634 14340
rect 9858 14328 9864 14340
rect 8628 14300 9864 14328
rect 8628 14288 8634 14300
rect 9858 14288 9864 14300
rect 9916 14288 9922 14340
rect 11882 14288 11888 14340
rect 11940 14328 11946 14340
rect 12158 14328 12164 14340
rect 11940 14300 12164 14328
rect 11940 14288 11946 14300
rect 12158 14288 12164 14300
rect 12216 14288 12222 14340
rect 12728 14328 12756 14368
rect 12803 14365 12815 14399
rect 12849 14396 12861 14399
rect 12894 14396 12900 14408
rect 12849 14368 12900 14396
rect 12849 14365 12861 14368
rect 12803 14359 12861 14365
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 15010 14328 15016 14340
rect 12728 14300 15016 14328
rect 15010 14288 15016 14300
rect 15068 14288 15074 14340
rect 7708 14232 8340 14260
rect 7708 14220 7714 14232
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 12437 14263 12495 14269
rect 12437 14260 12449 14263
rect 11020 14232 12449 14260
rect 11020 14220 11026 14232
rect 12437 14229 12449 14232
rect 12483 14229 12495 14263
rect 12437 14223 12495 14229
rect 1104 14170 14696 14192
rect 1104 14118 4308 14170
rect 4360 14118 4372 14170
rect 4424 14118 4436 14170
rect 4488 14118 4500 14170
rect 4552 14118 4564 14170
rect 4616 14118 7666 14170
rect 7718 14118 7730 14170
rect 7782 14118 7794 14170
rect 7846 14118 7858 14170
rect 7910 14118 7922 14170
rect 7974 14118 11024 14170
rect 11076 14118 11088 14170
rect 11140 14118 11152 14170
rect 11204 14118 11216 14170
rect 11268 14118 11280 14170
rect 11332 14118 14382 14170
rect 14434 14118 14446 14170
rect 14498 14118 14510 14170
rect 14562 14118 14574 14170
rect 14626 14118 14638 14170
rect 14690 14118 14696 14170
rect 1104 14096 14696 14118
rect 1946 14056 1952 14068
rect 1504 14028 1952 14056
rect 1504 13997 1532 14028
rect 1946 14016 1952 14028
rect 2004 14016 2010 14068
rect 7282 14016 7288 14068
rect 7340 14056 7346 14068
rect 7340 14028 9812 14056
rect 7340 14016 7346 14028
rect 1489 13991 1547 13997
rect 1489 13957 1501 13991
rect 1535 13957 1547 13991
rect 9674 13988 9680 14000
rect 1489 13951 1547 13957
rect 9646 13948 9680 13988
rect 9732 13948 9738 14000
rect 1670 13880 1676 13932
rect 1728 13920 1734 13932
rect 1854 13920 1860 13932
rect 1728 13892 1860 13920
rect 1728 13880 1734 13892
rect 1854 13880 1860 13892
rect 1912 13880 1918 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 7193 13923 7251 13929
rect 7193 13920 7205 13923
rect 5132 13892 7205 13920
rect 5132 13880 5138 13892
rect 7193 13889 7205 13892
rect 7239 13920 7251 13923
rect 7558 13920 7564 13932
rect 7239 13892 7564 13920
rect 7239 13889 7251 13892
rect 7193 13883 7251 13889
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 8113 13923 8171 13929
rect 8113 13889 8125 13923
rect 8159 13889 8171 13923
rect 8113 13883 8171 13889
rect 8251 13923 8309 13929
rect 8251 13889 8263 13923
rect 8297 13889 8309 13923
rect 8251 13886 8309 13889
rect 8251 13883 8340 13886
rect 7377 13855 7435 13861
rect 7377 13821 7389 13855
rect 7423 13821 7435 13855
rect 7377 13815 7435 13821
rect 5074 13744 5080 13796
rect 5132 13784 5138 13796
rect 5442 13784 5448 13796
rect 5132 13756 5448 13784
rect 5132 13744 5138 13756
rect 5442 13744 5448 13756
rect 5500 13744 5506 13796
rect 1578 13676 1584 13728
rect 1636 13676 1642 13728
rect 7392 13716 7420 13815
rect 7834 13812 7840 13864
rect 7892 13812 7898 13864
rect 8128 13852 8156 13883
rect 8266 13864 8340 13883
rect 8386 13880 8392 13932
rect 8444 13880 8450 13932
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9646 13920 9674 13948
rect 9784 13939 9812 14028
rect 9858 14016 9864 14068
rect 9916 14016 9922 14068
rect 10505 14059 10563 14065
rect 10505 14025 10517 14059
rect 10551 14056 10563 14059
rect 10778 14056 10784 14068
rect 10551 14028 10784 14056
rect 10551 14025 10563 14028
rect 10505 14019 10563 14025
rect 10778 14016 10784 14028
rect 10836 14016 10842 14068
rect 13354 14056 13360 14068
rect 10888 14028 13360 14056
rect 9876 13988 9904 14016
rect 10888 13988 10916 14028
rect 13354 14016 13360 14028
rect 13412 14016 13418 14068
rect 9876 13960 10916 13988
rect 11189 13960 11974 13988
rect 9079 13892 9674 13920
rect 9767 13933 9825 13939
rect 9767 13899 9779 13933
rect 9813 13899 9825 13933
rect 9767 13893 9825 13899
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9858 13880 9864 13932
rect 9916 13920 9922 13932
rect 10686 13920 10692 13932
rect 9916 13892 10692 13920
rect 9916 13880 9922 13892
rect 10686 13880 10692 13892
rect 10744 13920 10750 13932
rect 11189 13920 11217 13960
rect 10744 13892 11217 13920
rect 10744 13880 10750 13892
rect 11790 13880 11796 13932
rect 11848 13920 11854 13932
rect 11946 13920 11974 13960
rect 12342 13948 12348 14000
rect 12400 13988 12406 14000
rect 12434 13988 12440 14000
rect 12400 13960 12440 13988
rect 12400 13948 12406 13960
rect 12434 13948 12440 13960
rect 12492 13988 12498 14000
rect 12492 13960 13400 13988
rect 12492 13948 12498 13960
rect 13372 13932 13400 13960
rect 13906 13948 13912 14000
rect 13964 13948 13970 14000
rect 11848 13892 11891 13920
rect 11946 13892 13308 13920
rect 11848 13880 11854 13892
rect 8266 13858 8300 13864
rect 7926 13824 8156 13852
rect 7650 13744 7656 13796
rect 7708 13784 7714 13796
rect 7926 13784 7954 13824
rect 8294 13812 8300 13858
rect 8352 13812 8358 13864
rect 9490 13812 9496 13864
rect 9548 13812 9554 13864
rect 11514 13812 11520 13864
rect 11572 13812 11578 13864
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 13078 13852 13084 13864
rect 12943 13824 13084 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 13173 13855 13231 13861
rect 13173 13821 13185 13855
rect 13219 13821 13231 13855
rect 13280 13852 13308 13892
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 14093 13855 14151 13861
rect 14093 13852 14105 13855
rect 13280 13824 14105 13852
rect 13173 13815 13231 13821
rect 14093 13821 14105 13824
rect 14139 13821 14151 13855
rect 14093 13815 14151 13821
rect 7708 13756 7954 13784
rect 13188 13784 13216 13815
rect 13188 13756 13400 13784
rect 7708 13744 7714 13756
rect 13372 13728 13400 13756
rect 11790 13716 11796 13728
rect 7392 13688 11796 13716
rect 11790 13676 11796 13688
rect 11848 13676 11854 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12529 13719 12587 13725
rect 12529 13716 12541 13719
rect 12492 13688 12541 13716
rect 12492 13676 12498 13688
rect 12529 13685 12541 13688
rect 12575 13685 12587 13719
rect 12529 13679 12587 13685
rect 13354 13676 13360 13728
rect 13412 13676 13418 13728
rect 1104 13626 14536 13648
rect 1104 13574 2629 13626
rect 2681 13574 2693 13626
rect 2745 13574 2757 13626
rect 2809 13574 2821 13626
rect 2873 13574 2885 13626
rect 2937 13574 5987 13626
rect 6039 13574 6051 13626
rect 6103 13574 6115 13626
rect 6167 13574 6179 13626
rect 6231 13574 6243 13626
rect 6295 13574 9345 13626
rect 9397 13574 9409 13626
rect 9461 13574 9473 13626
rect 9525 13574 9537 13626
rect 9589 13574 9601 13626
rect 9653 13574 12703 13626
rect 12755 13574 12767 13626
rect 12819 13574 12831 13626
rect 12883 13574 12895 13626
rect 12947 13574 12959 13626
rect 13011 13574 14536 13626
rect 1104 13552 14536 13574
rect 6362 13512 6368 13524
rect 6196 13484 6368 13512
rect 6196 13444 6224 13484
rect 6362 13472 6368 13484
rect 6420 13512 6426 13524
rect 7101 13515 7159 13521
rect 6420 13484 7052 13512
rect 6420 13472 6426 13484
rect 6104 13416 6224 13444
rect 6104 13385 6132 13416
rect 6089 13379 6147 13385
rect 6089 13345 6101 13379
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 2406 13308 2412 13320
rect 2179 13280 2412 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 2406 13268 2412 13280
rect 2464 13268 2470 13320
rect 7024 13308 7052 13484
rect 7101 13481 7113 13515
rect 7147 13512 7159 13515
rect 7834 13512 7840 13524
rect 7147 13484 7840 13512
rect 7147 13481 7159 13484
rect 7101 13475 7159 13481
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8846 13512 8852 13524
rect 8352 13484 8852 13512
rect 8352 13472 8358 13484
rect 8846 13472 8852 13484
rect 8904 13472 8910 13524
rect 9398 13472 9404 13524
rect 9456 13512 9462 13524
rect 9456 13484 9720 13512
rect 9456 13472 9462 13484
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 9585 13447 9643 13453
rect 9585 13444 9597 13447
rect 8527 13416 9597 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9585 13413 9597 13416
rect 9631 13413 9643 13447
rect 9585 13407 9643 13413
rect 8938 13336 8944 13388
rect 8996 13336 9002 13388
rect 9692 13376 9720 13484
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10318 13512 10324 13524
rect 10192 13484 10324 13512
rect 10192 13472 10198 13484
rect 10318 13472 10324 13484
rect 10376 13512 10382 13524
rect 10781 13515 10839 13521
rect 10376 13484 10732 13512
rect 10376 13472 10382 13484
rect 10704 13444 10732 13484
rect 10781 13481 10793 13515
rect 10827 13512 10839 13515
rect 10870 13512 10876 13524
rect 10827 13484 10876 13512
rect 10827 13481 10839 13484
rect 10781 13475 10839 13481
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 13081 13515 13139 13521
rect 11992 13484 13032 13512
rect 10704 13416 11468 13444
rect 11440 13385 11468 13416
rect 9978 13379 10036 13385
rect 9978 13376 9990 13379
rect 9692 13348 9990 13376
rect 9978 13345 9990 13348
rect 10024 13376 10036 13379
rect 11425 13379 11483 13385
rect 10024 13348 10732 13376
rect 10024 13345 10036 13348
rect 9978 13339 10036 13345
rect 7098 13308 7104 13320
rect 6347 13281 6405 13287
rect 1489 13243 1547 13249
rect 1489 13209 1501 13243
rect 1535 13240 1547 13243
rect 6347 13247 6359 13281
rect 6393 13278 6405 13281
rect 7024 13280 7104 13308
rect 6393 13247 6408 13278
rect 7098 13268 7104 13280
rect 7156 13308 7162 13320
rect 7469 13311 7527 13317
rect 7156 13304 7420 13308
rect 7469 13304 7481 13311
rect 7156 13280 7481 13304
rect 7156 13268 7162 13280
rect 7392 13277 7481 13280
rect 7515 13277 7527 13311
rect 7392 13276 7527 13277
rect 7469 13271 7527 13276
rect 7650 13268 7656 13320
rect 7708 13308 7714 13320
rect 7743 13311 7801 13317
rect 7743 13308 7755 13311
rect 7708 13280 7755 13308
rect 7708 13268 7714 13280
rect 7743 13277 7755 13280
rect 7789 13277 7801 13311
rect 7743 13271 7801 13277
rect 8202 13268 8208 13320
rect 8260 13308 8266 13320
rect 8478 13308 8484 13320
rect 8260 13280 8484 13308
rect 8260 13268 8266 13280
rect 8478 13268 8484 13280
rect 8536 13268 8542 13320
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 6347 13241 6408 13247
rect 6380 13240 6408 13241
rect 6546 13240 6552 13252
rect 1535 13212 1992 13240
rect 6380 13212 6552 13240
rect 1535 13209 1547 13212
rect 1489 13203 1547 13209
rect 842 13132 848 13184
rect 900 13172 906 13184
rect 1964 13181 1992 13212
rect 6546 13200 6552 13212
rect 6604 13240 6610 13252
rect 6822 13240 6828 13252
rect 6604 13212 6828 13240
rect 6604 13200 6610 13212
rect 6822 13200 6828 13212
rect 6880 13200 6886 13252
rect 8938 13200 8944 13252
rect 8996 13240 9002 13252
rect 9140 13240 9168 13271
rect 9858 13268 9864 13320
rect 9916 13268 9922 13320
rect 10134 13268 10140 13320
rect 10192 13268 10198 13320
rect 10704 13252 10732 13348
rect 11425 13345 11437 13379
rect 11471 13345 11483 13379
rect 11425 13339 11483 13345
rect 11882 13336 11888 13388
rect 11940 13336 11946 13388
rect 11992 13376 12020 13484
rect 13004 13444 13032 13484
rect 13081 13481 13093 13515
rect 13127 13512 13139 13515
rect 13446 13512 13452 13524
rect 13127 13484 13452 13512
rect 13127 13481 13139 13484
rect 13081 13475 13139 13481
rect 13446 13472 13452 13484
rect 13504 13472 13510 13524
rect 13817 13515 13875 13521
rect 13817 13481 13829 13515
rect 13863 13512 13875 13515
rect 15286 13512 15292 13524
rect 13863 13484 15292 13512
rect 13863 13481 13875 13484
rect 13817 13475 13875 13481
rect 13170 13444 13176 13456
rect 13004 13416 13176 13444
rect 12342 13385 12348 13388
rect 12161 13379 12219 13385
rect 12161 13376 12173 13379
rect 11992 13348 12173 13376
rect 12161 13345 12173 13348
rect 12207 13345 12219 13379
rect 12161 13339 12219 13345
rect 12299 13379 12348 13385
rect 12299 13345 12311 13379
rect 12345 13345 12348 13379
rect 12299 13339 12348 13345
rect 12342 13336 12348 13339
rect 12400 13336 12406 13388
rect 12434 13336 12440 13388
rect 12492 13336 12498 13388
rect 13004 13376 13032 13416
rect 13170 13404 13176 13416
rect 13228 13404 13234 13456
rect 13262 13404 13268 13456
rect 13320 13444 13326 13456
rect 13357 13447 13415 13453
rect 13357 13444 13369 13447
rect 13320 13416 13369 13444
rect 13320 13404 13326 13416
rect 13357 13413 13369 13416
rect 13403 13413 13415 13447
rect 13357 13407 13415 13413
rect 13832 13376 13860 13475
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 13004 13348 13860 13376
rect 11238 13308 11244 13320
rect 10796 13280 11244 13308
rect 10796 13252 10824 13280
rect 11238 13268 11244 13280
rect 11296 13268 11302 13320
rect 13173 13311 13231 13317
rect 13173 13277 13185 13311
rect 13219 13308 13231 13311
rect 14366 13308 14372 13320
rect 13219 13280 14372 13308
rect 13219 13277 13231 13280
rect 13173 13271 13231 13277
rect 14366 13268 14372 13280
rect 14424 13268 14430 13320
rect 8996 13212 9168 13240
rect 8996 13200 9002 13212
rect 10686 13200 10692 13252
rect 10744 13200 10750 13252
rect 10778 13200 10784 13252
rect 10836 13200 10842 13252
rect 13722 13200 13728 13252
rect 13780 13200 13786 13252
rect 1581 13175 1639 13181
rect 1581 13172 1593 13175
rect 900 13144 1593 13172
rect 900 13132 906 13144
rect 1581 13141 1593 13144
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 1949 13175 2007 13181
rect 1949 13141 1961 13175
rect 1995 13141 2007 13175
rect 1949 13135 2007 13141
rect 4062 13132 4068 13184
rect 4120 13172 4126 13184
rect 8570 13172 8576 13184
rect 4120 13144 8576 13172
rect 4120 13132 4126 13144
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 8662 13132 8668 13184
rect 8720 13172 8726 13184
rect 11422 13172 11428 13184
rect 8720 13144 11428 13172
rect 8720 13132 8726 13144
rect 11422 13132 11428 13144
rect 11480 13132 11486 13184
rect 1104 13082 14696 13104
rect 1104 13030 4308 13082
rect 4360 13030 4372 13082
rect 4424 13030 4436 13082
rect 4488 13030 4500 13082
rect 4552 13030 4564 13082
rect 4616 13030 7666 13082
rect 7718 13030 7730 13082
rect 7782 13030 7794 13082
rect 7846 13030 7858 13082
rect 7910 13030 7922 13082
rect 7974 13030 11024 13082
rect 11076 13030 11088 13082
rect 11140 13030 11152 13082
rect 11204 13030 11216 13082
rect 11268 13030 11280 13082
rect 11332 13030 14382 13082
rect 14434 13030 14446 13082
rect 14498 13030 14510 13082
rect 14562 13030 14574 13082
rect 14626 13030 14638 13082
rect 14690 13030 14696 13082
rect 1104 13008 14696 13030
rect 1670 12928 1676 12980
rect 1728 12928 1734 12980
rect 3786 12928 3792 12980
rect 3844 12968 3850 12980
rect 6914 12968 6920 12980
rect 3844 12940 6920 12968
rect 3844 12928 3850 12940
rect 6914 12928 6920 12940
rect 6972 12968 6978 12980
rect 7282 12968 7288 12980
rect 6972 12940 7288 12968
rect 6972 12928 6978 12940
rect 7282 12928 7288 12940
rect 7340 12928 7346 12980
rect 8021 12971 8079 12977
rect 8021 12937 8033 12971
rect 8067 12968 8079 12971
rect 8386 12968 8392 12980
rect 8067 12940 8392 12968
rect 8067 12937 8079 12940
rect 8021 12931 8079 12937
rect 8386 12928 8392 12940
rect 8444 12928 8450 12980
rect 8570 12928 8576 12980
rect 8628 12968 8634 12980
rect 9861 12971 9919 12977
rect 8628 12940 9812 12968
rect 8628 12928 8634 12940
rect 1688 12871 1716 12928
rect 7098 12900 7104 12912
rect 1655 12865 1716 12871
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 1655 12831 1667 12865
rect 1701 12834 1716 12865
rect 7024 12872 7104 12900
rect 7024 12841 7052 12872
rect 7098 12860 7104 12872
rect 7156 12900 7162 12912
rect 8846 12900 8852 12912
rect 7156 12872 8852 12900
rect 7156 12860 7162 12872
rect 8846 12860 8852 12872
rect 8904 12900 8910 12912
rect 9674 12900 9680 12912
rect 8904 12872 9680 12900
rect 8904 12860 8910 12872
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 9784 12900 9812 12940
rect 9861 12937 9873 12971
rect 9907 12968 9919 12971
rect 10134 12968 10140 12980
rect 9907 12940 10140 12968
rect 9907 12937 9919 12940
rect 9861 12931 9919 12937
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10778 12928 10784 12980
rect 10836 12928 10842 12980
rect 13998 12968 14004 12980
rect 12084 12940 14004 12968
rect 10796 12900 10824 12928
rect 9784 12872 10824 12900
rect 7009 12835 7067 12841
rect 1701 12831 1713 12834
rect 1655 12825 1713 12831
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7282 12832 7288 12844
rect 7243 12804 7288 12832
rect 7009 12795 7067 12801
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 8662 12792 8668 12844
rect 8720 12836 8726 12844
rect 8720 12832 8800 12836
rect 9091 12835 9149 12841
rect 9091 12832 9103 12835
rect 8720 12808 9103 12832
rect 8720 12792 8726 12808
rect 8772 12804 9103 12808
rect 9091 12801 9103 12804
rect 9137 12801 9149 12835
rect 9091 12795 9149 12801
rect 10410 12792 10416 12844
rect 10468 12832 10474 12844
rect 12084 12841 12112 12940
rect 13998 12928 14004 12940
rect 14056 12928 14062 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 15470 12968 15476 12980
rect 14231 12940 15476 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 10781 12835 10839 12841
rect 10781 12832 10793 12835
rect 10468 12804 10793 12832
rect 10468 12792 10474 12804
rect 10781 12801 10793 12804
rect 10827 12801 10839 12835
rect 10781 12795 10839 12801
rect 12069 12835 12127 12841
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12529 12835 12587 12841
rect 12529 12801 12541 12835
rect 12575 12832 12587 12835
rect 12710 12832 12716 12844
rect 12575 12804 12716 12832
rect 12575 12801 12587 12804
rect 12529 12795 12587 12801
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 8846 12724 8852 12776
rect 8904 12724 8910 12776
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 9858 12656 9864 12708
rect 9916 12696 9922 12708
rect 10042 12696 10048 12708
rect 9916 12668 10048 12696
rect 9916 12656 9922 12668
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 10520 12696 10548 12727
rect 11974 12724 11980 12776
rect 12032 12764 12038 12776
rect 12345 12767 12403 12773
rect 12032 12736 12296 12764
rect 12032 12724 12038 12736
rect 12158 12696 12164 12708
rect 10520 12668 12164 12696
rect 12158 12656 12164 12668
rect 12216 12656 12222 12708
rect 12268 12705 12296 12736
rect 12345 12733 12357 12767
rect 12391 12733 12403 12767
rect 12345 12727 12403 12733
rect 12253 12699 12311 12705
rect 12253 12665 12265 12699
rect 12299 12665 12311 12699
rect 12253 12659 12311 12665
rect 2406 12588 2412 12640
rect 2464 12588 2470 12640
rect 5350 12588 5356 12640
rect 5408 12628 5414 12640
rect 8662 12628 8668 12640
rect 5408 12600 8668 12628
rect 5408 12588 5414 12600
rect 8662 12588 8668 12600
rect 8720 12628 8726 12640
rect 8846 12628 8852 12640
rect 8720 12600 8852 12628
rect 8720 12588 8726 12600
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 11330 12628 11336 12640
rect 8996 12600 11336 12628
rect 8996 12588 9002 12600
rect 11330 12588 11336 12600
rect 11388 12588 11394 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 12360 12628 12388 12727
rect 12618 12724 12624 12776
rect 12676 12764 12682 12776
rect 13446 12773 13452 12776
rect 13265 12767 13323 12773
rect 13265 12764 13277 12767
rect 12676 12736 13277 12764
rect 12676 12724 12682 12736
rect 13265 12733 13277 12736
rect 13311 12733 13323 12767
rect 13265 12727 13323 12733
rect 13403 12767 13452 12773
rect 13403 12733 13415 12767
rect 13449 12733 13452 12767
rect 13403 12727 13452 12733
rect 13446 12724 13452 12727
rect 13504 12724 13510 12776
rect 13538 12724 13544 12776
rect 13596 12724 13602 12776
rect 12986 12656 12992 12708
rect 13044 12656 13050 12708
rect 11848 12600 12388 12628
rect 11848 12588 11854 12600
rect 12434 12588 12440 12640
rect 12492 12628 12498 12640
rect 12618 12628 12624 12640
rect 12492 12600 12624 12628
rect 12492 12588 12498 12600
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 1104 12538 14536 12560
rect 1104 12486 2629 12538
rect 2681 12486 2693 12538
rect 2745 12486 2757 12538
rect 2809 12486 2821 12538
rect 2873 12486 2885 12538
rect 2937 12486 5987 12538
rect 6039 12486 6051 12538
rect 6103 12486 6115 12538
rect 6167 12486 6179 12538
rect 6231 12486 6243 12538
rect 6295 12486 9345 12538
rect 9397 12486 9409 12538
rect 9461 12486 9473 12538
rect 9525 12486 9537 12538
rect 9589 12486 9601 12538
rect 9653 12486 12703 12538
rect 12755 12486 12767 12538
rect 12819 12486 12831 12538
rect 12883 12486 12895 12538
rect 12947 12486 12959 12538
rect 13011 12486 14536 12538
rect 1104 12464 14536 12486
rect 4706 12424 4712 12436
rect 4356 12396 4712 12424
rect 4356 12297 4384 12396
rect 4706 12384 4712 12396
rect 4764 12384 4770 12436
rect 7190 12384 7196 12436
rect 7248 12384 7254 12436
rect 11517 12427 11575 12433
rect 11517 12393 11529 12427
rect 11563 12424 11575 12427
rect 11882 12424 11888 12436
rect 11563 12396 11888 12424
rect 11563 12393 11575 12396
rect 11517 12387 11575 12393
rect 11882 12384 11888 12396
rect 11940 12384 11946 12436
rect 13078 12384 13084 12436
rect 13136 12424 13142 12436
rect 13173 12427 13231 12433
rect 13173 12424 13185 12427
rect 13136 12396 13185 12424
rect 13136 12384 13142 12396
rect 13173 12393 13185 12396
rect 13219 12393 13231 12427
rect 13173 12387 13231 12393
rect 6822 12316 6828 12368
rect 6880 12356 6886 12368
rect 7208 12356 7236 12384
rect 6880 12328 7236 12356
rect 6880 12316 6886 12328
rect 4341 12291 4399 12297
rect 4341 12257 4353 12291
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 7098 12248 7104 12300
rect 7156 12248 7162 12300
rect 9674 12248 9680 12300
rect 9732 12288 9738 12300
rect 10502 12288 10508 12300
rect 9732 12260 10508 12288
rect 9732 12248 9738 12260
rect 10502 12248 10508 12260
rect 10560 12248 10566 12300
rect 11808 12260 12002 12288
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2406 12220 2412 12232
rect 2179 12192 2412 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2406 12180 2412 12192
rect 2464 12180 2470 12232
rect 4615 12223 4673 12229
rect 4615 12189 4627 12223
rect 4661 12220 4673 12223
rect 5626 12220 5632 12232
rect 4661 12192 5632 12220
rect 4661 12189 4673 12192
rect 4615 12183 4673 12189
rect 5626 12180 5632 12192
rect 5684 12180 5690 12232
rect 5721 12223 5779 12229
rect 5721 12189 5733 12223
rect 5767 12189 5779 12223
rect 5721 12183 5779 12189
rect 5995 12223 6053 12229
rect 5995 12189 6007 12223
rect 6041 12220 6053 12223
rect 7006 12220 7012 12232
rect 6041 12192 7012 12220
rect 6041 12189 6053 12192
rect 5995 12183 6053 12189
rect 1489 12155 1547 12161
rect 1489 12121 1501 12155
rect 1535 12152 1547 12155
rect 1535 12124 1992 12152
rect 1535 12121 1547 12124
rect 1489 12115 1547 12121
rect 842 12044 848 12096
rect 900 12084 906 12096
rect 1964 12093 1992 12124
rect 4706 12112 4712 12164
rect 4764 12152 4770 12164
rect 5736 12152 5764 12183
rect 7006 12180 7012 12192
rect 7064 12180 7070 12232
rect 7374 12220 7380 12232
rect 7335 12192 7380 12220
rect 7374 12180 7380 12192
rect 7432 12180 7438 12232
rect 9214 12180 9220 12232
rect 9272 12180 9278 12232
rect 10747 12223 10805 12229
rect 10747 12220 10759 12223
rect 10152 12192 10759 12220
rect 4764 12124 5764 12152
rect 4764 12112 4770 12124
rect 1581 12087 1639 12093
rect 1581 12084 1593 12087
rect 900 12056 1593 12084
rect 900 12044 906 12056
rect 1581 12053 1593 12056
rect 1627 12053 1639 12087
rect 1581 12047 1639 12053
rect 1949 12087 2007 12093
rect 1949 12053 1961 12087
rect 1995 12053 2007 12087
rect 1949 12047 2007 12053
rect 5353 12087 5411 12093
rect 5353 12053 5365 12087
rect 5399 12084 5411 12087
rect 5626 12084 5632 12096
rect 5399 12056 5632 12084
rect 5399 12053 5411 12056
rect 5353 12047 5411 12053
rect 5626 12044 5632 12056
rect 5684 12044 5690 12096
rect 6733 12087 6791 12093
rect 6733 12053 6745 12087
rect 6779 12084 6791 12087
rect 7190 12084 7196 12096
rect 6779 12056 7196 12084
rect 6779 12053 6791 12056
rect 6733 12047 6791 12053
rect 7190 12044 7196 12056
rect 7248 12044 7254 12096
rect 8110 12044 8116 12096
rect 8168 12044 8174 12096
rect 9232 12084 9260 12180
rect 10152 12164 10180 12192
rect 10747 12189 10759 12192
rect 10793 12220 10805 12223
rect 11808 12220 11836 12260
rect 10793 12192 11836 12220
rect 11885 12223 11943 12229
rect 10793 12189 10805 12192
rect 10747 12183 10805 12189
rect 11885 12189 11897 12223
rect 11931 12189 11943 12223
rect 11974 12220 12002 12260
rect 12066 12248 12072 12300
rect 12124 12288 12130 12300
rect 12161 12291 12219 12297
rect 12161 12288 12173 12291
rect 12124 12260 12173 12288
rect 12124 12248 12130 12260
rect 12161 12257 12173 12260
rect 12207 12257 12219 12291
rect 12161 12251 12219 12257
rect 12403 12223 12461 12229
rect 12403 12220 12415 12223
rect 11974 12192 12415 12220
rect 11885 12183 11943 12189
rect 12403 12189 12415 12192
rect 12449 12189 12461 12223
rect 12403 12183 12461 12189
rect 10134 12112 10140 12164
rect 10192 12112 10198 12164
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 11900 12152 11928 12183
rect 13722 12180 13728 12232
rect 13780 12180 13786 12232
rect 11664 12124 11928 12152
rect 11664 12112 11670 12124
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 12158 12152 12164 12164
rect 12032 12124 12164 12152
rect 12032 12112 12038 12124
rect 12158 12112 12164 12124
rect 12216 12112 12222 12164
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 9232 12056 12081 12084
rect 12069 12053 12081 12056
rect 12115 12053 12127 12087
rect 12069 12047 12127 12053
rect 13446 12044 13452 12096
rect 13504 12084 13510 12096
rect 13630 12084 13636 12096
rect 13504 12056 13636 12084
rect 13504 12044 13510 12056
rect 13630 12044 13636 12056
rect 13688 12084 13694 12096
rect 13817 12087 13875 12093
rect 13817 12084 13829 12087
rect 13688 12056 13829 12084
rect 13688 12044 13694 12056
rect 13817 12053 13829 12056
rect 13863 12053 13875 12087
rect 13817 12047 13875 12053
rect 1104 11994 14696 12016
rect 1104 11942 4308 11994
rect 4360 11942 4372 11994
rect 4424 11942 4436 11994
rect 4488 11942 4500 11994
rect 4552 11942 4564 11994
rect 4616 11942 7666 11994
rect 7718 11942 7730 11994
rect 7782 11942 7794 11994
rect 7846 11942 7858 11994
rect 7910 11942 7922 11994
rect 7974 11942 11024 11994
rect 11076 11942 11088 11994
rect 11140 11942 11152 11994
rect 11204 11942 11216 11994
rect 11268 11942 11280 11994
rect 11332 11942 14382 11994
rect 14434 11942 14446 11994
rect 14498 11942 14510 11994
rect 14562 11942 14574 11994
rect 14626 11942 14638 11994
rect 14690 11942 14696 11994
rect 1104 11920 14696 11942
rect 5810 11840 5816 11892
rect 5868 11880 5874 11892
rect 10134 11880 10140 11892
rect 5868 11852 10140 11880
rect 5868 11840 5874 11852
rect 10134 11840 10140 11852
rect 10192 11840 10198 11892
rect 12342 11880 12348 11892
rect 10520 11852 12348 11880
rect 5151 11777 5209 11783
rect 1486 11704 1492 11756
rect 1544 11704 1550 11756
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4893 11747 4951 11753
rect 4893 11744 4905 11747
rect 4764 11716 4905 11744
rect 4764 11704 4770 11716
rect 4893 11713 4905 11716
rect 4939 11713 4951 11747
rect 5151 11743 5163 11777
rect 5197 11774 5209 11777
rect 5197 11744 5212 11774
rect 5902 11772 5908 11824
rect 5960 11812 5966 11824
rect 7742 11812 7748 11824
rect 5960 11784 7748 11812
rect 5960 11772 5966 11784
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 8018 11812 8024 11824
rect 7944 11784 8024 11812
rect 7944 11783 7972 11784
rect 7911 11777 7972 11783
rect 5534 11744 5540 11756
rect 5197 11743 5540 11744
rect 5151 11737 5540 11743
rect 5184 11716 5540 11737
rect 4893 11707 4951 11713
rect 5534 11704 5540 11716
rect 5592 11704 5598 11756
rect 6914 11704 6920 11756
rect 6972 11744 6978 11756
rect 7282 11744 7288 11756
rect 6972 11716 7288 11744
rect 6972 11704 6978 11716
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 7911 11743 7923 11777
rect 7957 11746 7972 11777
rect 8018 11772 8024 11784
rect 8076 11772 8082 11824
rect 8202 11772 8208 11824
rect 8260 11812 8266 11824
rect 8260 11784 8340 11812
rect 8260 11772 8266 11784
rect 7957 11743 7969 11746
rect 7911 11737 7969 11743
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7653 11679 7711 11685
rect 7653 11676 7665 11679
rect 7156 11648 7665 11676
rect 7156 11636 7162 11648
rect 7653 11645 7665 11648
rect 7699 11645 7711 11679
rect 8312 11676 8340 11784
rect 10520 11753 10548 11852
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 13538 11840 13544 11892
rect 13596 11880 13602 11892
rect 13633 11883 13691 11889
rect 13633 11880 13645 11883
rect 13596 11852 13645 11880
rect 13596 11840 13602 11852
rect 13633 11849 13645 11852
rect 13679 11849 13691 11883
rect 13633 11843 13691 11849
rect 12066 11812 12072 11824
rect 11716 11784 12072 11812
rect 10505 11747 10563 11753
rect 10505 11713 10517 11747
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 11716 11753 11744 11784
rect 12066 11772 12072 11784
rect 12124 11772 12130 11824
rect 12544 11784 12906 11812
rect 11701 11747 11759 11753
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11790 11704 11796 11756
rect 11848 11744 11854 11756
rect 12544 11744 12572 11784
rect 12878 11783 12906 11784
rect 12878 11777 12937 11783
rect 12878 11746 12891 11777
rect 11848 11716 12572 11744
rect 12879 11743 12891 11746
rect 12925 11743 12937 11777
rect 12879 11737 12937 11743
rect 11848 11704 11854 11716
rect 13998 11704 14004 11756
rect 14056 11704 14062 11756
rect 11977 11679 12035 11685
rect 11977 11676 11989 11679
rect 8312 11648 11989 11676
rect 7653 11639 7711 11645
rect 11977 11645 11989 11648
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12621 11679 12679 11685
rect 12621 11645 12633 11679
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 842 11500 848 11552
rect 900 11540 906 11552
rect 1581 11543 1639 11549
rect 1581 11540 1593 11543
rect 900 11512 1593 11540
rect 900 11500 906 11512
rect 1581 11509 1593 11512
rect 1627 11509 1639 11543
rect 1581 11503 1639 11509
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 7282 11540 7288 11552
rect 5960 11512 7288 11540
rect 5960 11500 5966 11512
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 7668 11540 7696 11639
rect 11882 11608 11888 11620
rect 8312 11580 11888 11608
rect 8312 11540 8340 11580
rect 11882 11568 11888 11580
rect 11940 11608 11946 11620
rect 12342 11608 12348 11620
rect 11940 11580 12348 11608
rect 11940 11568 11946 11580
rect 12342 11568 12348 11580
rect 12400 11608 12406 11620
rect 12636 11608 12664 11639
rect 12400 11580 12664 11608
rect 13280 11580 14228 11608
rect 12400 11568 12406 11580
rect 7668 11512 8340 11540
rect 8662 11500 8668 11552
rect 8720 11500 8726 11552
rect 11422 11500 11428 11552
rect 11480 11540 11486 11552
rect 13280 11540 13308 11580
rect 14200 11549 14228 11580
rect 11480 11512 13308 11540
rect 14185 11543 14243 11549
rect 11480 11500 11486 11512
rect 14185 11509 14197 11543
rect 14231 11509 14243 11543
rect 14185 11503 14243 11509
rect 1104 11450 14536 11472
rect 1104 11398 2629 11450
rect 2681 11398 2693 11450
rect 2745 11398 2757 11450
rect 2809 11398 2821 11450
rect 2873 11398 2885 11450
rect 2937 11398 5987 11450
rect 6039 11398 6051 11450
rect 6103 11398 6115 11450
rect 6167 11398 6179 11450
rect 6231 11398 6243 11450
rect 6295 11398 9345 11450
rect 9397 11398 9409 11450
rect 9461 11398 9473 11450
rect 9525 11398 9537 11450
rect 9589 11398 9601 11450
rect 9653 11398 12703 11450
rect 12755 11398 12767 11450
rect 12819 11398 12831 11450
rect 12883 11398 12895 11450
rect 12947 11398 12959 11450
rect 13011 11398 14536 11450
rect 1104 11376 14536 11398
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 7837 11339 7895 11345
rect 7837 11336 7849 11339
rect 6696 11308 7849 11336
rect 6696 11296 6702 11308
rect 7837 11305 7849 11308
rect 7883 11305 7895 11339
rect 7837 11299 7895 11305
rect 10502 11296 10508 11348
rect 10560 11336 10566 11348
rect 11514 11336 11520 11348
rect 10560 11308 11520 11336
rect 10560 11296 10566 11308
rect 11514 11296 11520 11308
rect 11572 11336 11578 11348
rect 13170 11336 13176 11348
rect 11572 11308 13176 11336
rect 11572 11296 11578 11308
rect 6012 11240 6776 11268
rect 5718 11160 5724 11212
rect 5776 11160 5782 11212
rect 5736 11132 5764 11160
rect 6012 11141 6040 11240
rect 6086 11160 6092 11212
rect 6144 11200 6150 11212
rect 6641 11203 6699 11209
rect 6641 11200 6653 11203
rect 6144 11172 6653 11200
rect 6144 11160 6150 11172
rect 6641 11169 6653 11172
rect 6687 11169 6699 11203
rect 6748 11200 6776 11240
rect 7742 11228 7748 11280
rect 7800 11268 7806 11280
rect 8478 11268 8484 11280
rect 7800 11240 8484 11268
rect 7800 11228 7806 11240
rect 8478 11228 8484 11240
rect 8536 11228 8542 11280
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 11149 11271 11207 11277
rect 11149 11268 11161 11271
rect 10744 11240 11161 11268
rect 10744 11228 10750 11240
rect 11149 11237 11161 11240
rect 11195 11237 11207 11271
rect 11149 11231 11207 11237
rect 8386 11200 8392 11212
rect 6748 11172 8392 11200
rect 6641 11163 6699 11169
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 12452 11209 12480 11308
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 12345 11203 12403 11209
rect 12345 11200 12357 11203
rect 9692 11172 12357 11200
rect 5997 11135 6055 11141
rect 5997 11132 6009 11135
rect 5736 11104 6009 11132
rect 5997 11101 6009 11104
rect 6043 11101 6055 11135
rect 5997 11095 6055 11101
rect 6181 11135 6239 11141
rect 6181 11101 6193 11135
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 5810 11024 5816 11076
rect 5868 11064 5874 11076
rect 6196 11064 6224 11095
rect 6914 11092 6920 11144
rect 6972 11092 6978 11144
rect 7098 11141 7104 11144
rect 7055 11135 7104 11141
rect 7055 11101 7067 11135
rect 7101 11101 7104 11135
rect 7055 11095 7104 11101
rect 7098 11092 7104 11095
rect 7156 11092 7162 11144
rect 7190 11092 7196 11144
rect 7248 11092 7254 11144
rect 8846 11092 8852 11144
rect 8904 11132 8910 11144
rect 9030 11132 9036 11144
rect 8904 11104 9036 11132
rect 8904 11092 8910 11104
rect 9030 11092 9036 11104
rect 9088 11092 9094 11144
rect 5868 11036 6224 11064
rect 7760 11036 7972 11064
rect 5868 11024 5874 11036
rect 2130 10956 2136 11008
rect 2188 10996 2194 11008
rect 7760 10996 7788 11036
rect 2188 10968 7788 10996
rect 7944 10996 7972 11036
rect 9692 10996 9720 11172
rect 12345 11169 12357 11172
rect 12391 11169 12403 11203
rect 12345 11163 12403 11169
rect 12437 11203 12495 11209
rect 12437 11169 12449 11203
rect 12483 11169 12495 11203
rect 12437 11163 12495 11169
rect 10502 11092 10508 11144
rect 10560 11092 10566 11144
rect 10689 11135 10747 11141
rect 10689 11101 10701 11135
rect 10735 11132 10747 11135
rect 10870 11132 10876 11144
rect 10735 11104 10876 11132
rect 10735 11101 10747 11104
rect 10689 11095 10747 11101
rect 10870 11092 10876 11104
rect 10928 11092 10934 11144
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 11606 11141 11612 11144
rect 11563 11135 11612 11141
rect 11563 11101 11575 11135
rect 11609 11101 11612 11135
rect 11563 11095 11612 11101
rect 11578 11094 11612 11095
rect 11606 11092 11612 11094
rect 11664 11092 11670 11144
rect 11698 11092 11704 11144
rect 11756 11092 11762 11144
rect 12710 11111 12716 11144
rect 12695 11105 12716 11111
rect 12695 11071 12707 11105
rect 12768 11092 12774 11144
rect 12741 11074 12756 11092
rect 12741 11071 12753 11074
rect 12695 11065 12753 11071
rect 7944 10968 9720 10996
rect 2188 10956 2194 10968
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13449 10999 13507 11005
rect 13449 10996 13461 10999
rect 12952 10968 13461 10996
rect 12952 10956 12958 10968
rect 13449 10965 13461 10968
rect 13495 10965 13507 10999
rect 13449 10959 13507 10965
rect 1104 10906 14696 10928
rect 1104 10854 4308 10906
rect 4360 10854 4372 10906
rect 4424 10854 4436 10906
rect 4488 10854 4500 10906
rect 4552 10854 4564 10906
rect 4616 10854 7666 10906
rect 7718 10854 7730 10906
rect 7782 10854 7794 10906
rect 7846 10854 7858 10906
rect 7910 10854 7922 10906
rect 7974 10854 11024 10906
rect 11076 10854 11088 10906
rect 11140 10854 11152 10906
rect 11204 10854 11216 10906
rect 11268 10854 11280 10906
rect 11332 10854 14382 10906
rect 14434 10854 14446 10906
rect 14498 10854 14510 10906
rect 14562 10854 14574 10906
rect 14626 10854 14638 10906
rect 14690 10854 14696 10906
rect 1104 10832 14696 10854
rect 1486 10752 1492 10804
rect 1544 10792 1550 10804
rect 1949 10795 2007 10801
rect 1949 10792 1961 10795
rect 1544 10764 1961 10792
rect 1544 10752 1550 10764
rect 1949 10761 1961 10764
rect 1995 10761 2007 10795
rect 1949 10755 2007 10761
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7285 10795 7343 10801
rect 7285 10792 7297 10795
rect 6972 10764 7297 10792
rect 6972 10752 6978 10764
rect 7285 10761 7297 10764
rect 7331 10761 7343 10795
rect 7285 10755 7343 10761
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 8113 10795 8171 10801
rect 8113 10792 8125 10795
rect 7616 10764 8125 10792
rect 7616 10752 7622 10764
rect 8113 10761 8125 10764
rect 8159 10761 8171 10795
rect 8113 10755 8171 10761
rect 8202 10752 8208 10804
rect 8260 10792 8266 10804
rect 10318 10792 10324 10804
rect 8260 10764 10324 10792
rect 8260 10752 8266 10764
rect 10318 10752 10324 10764
rect 10376 10752 10382 10804
rect 10594 10752 10600 10804
rect 10652 10752 10658 10804
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 11057 10795 11115 10801
rect 11057 10792 11069 10795
rect 10744 10764 11069 10792
rect 10744 10752 10750 10764
rect 11057 10761 11069 10764
rect 11103 10761 11115 10795
rect 11057 10755 11115 10761
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11480 10764 11713 10792
rect 11480 10752 11486 10764
rect 11701 10761 11713 10764
rect 11747 10792 11759 10795
rect 11882 10792 11888 10804
rect 11747 10764 11888 10792
rect 11747 10761 11759 10764
rect 11701 10755 11759 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 11977 10795 12035 10801
rect 11977 10761 11989 10795
rect 12023 10761 12035 10795
rect 11977 10755 12035 10761
rect 5644 10696 6684 10724
rect 5644 10668 5672 10696
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10656 1547 10659
rect 2038 10656 2044 10668
rect 1535 10628 2044 10656
rect 1535 10625 1547 10628
rect 1489 10619 1547 10625
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2130 10616 2136 10668
rect 2188 10616 2194 10668
rect 5626 10616 5632 10668
rect 5684 10616 5690 10668
rect 6362 10616 6368 10668
rect 6420 10616 6426 10668
rect 6656 10665 6684 10696
rect 8386 10684 8392 10736
rect 8444 10684 8450 10736
rect 8481 10727 8539 10733
rect 8481 10693 8493 10727
rect 8527 10724 8539 10727
rect 8662 10724 8668 10736
rect 8527 10696 8668 10724
rect 8527 10693 8539 10696
rect 8481 10687 8539 10693
rect 8662 10684 8668 10696
rect 8720 10684 8726 10736
rect 9217 10727 9275 10733
rect 9217 10724 9229 10727
rect 8772 10696 9229 10724
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10625 6699 10659
rect 6641 10619 6699 10625
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10625 6883 10659
rect 6825 10619 6883 10625
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6840 10588 6868 10619
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 7156 10628 7205 10656
rect 7156 10616 7162 10628
rect 7193 10625 7205 10628
rect 7239 10625 7251 10659
rect 8036 10656 8248 10660
rect 8772 10656 8800 10696
rect 9217 10693 9229 10696
rect 9263 10724 9275 10727
rect 9263 10696 9812 10724
rect 9263 10693 9275 10696
rect 9217 10687 9275 10693
rect 7193 10619 7251 10625
rect 7668 10632 8800 10656
rect 7668 10628 8064 10632
rect 8220 10628 8800 10632
rect 8849 10659 8907 10665
rect 6604 10560 6868 10588
rect 6604 10548 6610 10560
rect 7668 10464 7696 10628
rect 8849 10625 8861 10659
rect 8895 10656 8907 10659
rect 9674 10656 9680 10668
rect 8895 10628 9680 10656
rect 8895 10625 8907 10628
rect 8849 10619 8907 10625
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 8128 10464 8156 10574
rect 842 10412 848 10464
rect 900 10452 906 10464
rect 1581 10455 1639 10461
rect 1581 10452 1593 10455
rect 900 10424 1593 10452
rect 900 10412 906 10424
rect 1581 10421 1593 10424
rect 1627 10421 1639 10455
rect 1581 10415 1639 10421
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 5776 10424 6469 10452
rect 5776 10412 5782 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 6730 10412 6736 10464
rect 6788 10412 6794 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7650 10452 7656 10464
rect 6972 10424 7656 10452
rect 6972 10412 6978 10424
rect 7650 10412 7656 10424
rect 7708 10412 7714 10464
rect 8110 10412 8116 10464
rect 8168 10412 8174 10464
rect 9398 10412 9404 10464
rect 9456 10412 9462 10464
rect 9784 10452 9812 10696
rect 10336 10695 10364 10752
rect 10612 10724 10640 10752
rect 11992 10724 12020 10755
rect 12250 10752 12256 10804
rect 12308 10752 12314 10804
rect 12342 10752 12348 10804
rect 12400 10792 12406 10804
rect 13078 10792 13084 10804
rect 12400 10764 13084 10792
rect 12400 10752 12406 10764
rect 13078 10752 13084 10764
rect 13136 10752 13142 10804
rect 14185 10795 14243 10801
rect 14185 10761 14197 10795
rect 14231 10792 14243 10795
rect 14274 10792 14280 10804
rect 14231 10764 14280 10792
rect 14231 10761 14243 10764
rect 14185 10755 14243 10761
rect 14274 10752 14280 10764
rect 14332 10752 14338 10804
rect 10612 10696 12020 10724
rect 10303 10689 10364 10695
rect 10303 10655 10315 10689
rect 10349 10658 10364 10689
rect 11517 10659 11575 10665
rect 10349 10655 10361 10658
rect 10303 10649 10361 10655
rect 11517 10625 11529 10659
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 9858 10548 9864 10600
rect 9916 10588 9922 10600
rect 10045 10591 10103 10597
rect 10045 10588 10057 10591
rect 9916 10560 10057 10588
rect 9916 10548 9922 10560
rect 10045 10557 10057 10560
rect 10091 10557 10103 10591
rect 10045 10551 10103 10557
rect 11054 10520 11060 10532
rect 10704 10492 11060 10520
rect 10704 10452 10732 10492
rect 11054 10480 11060 10492
rect 11112 10480 11118 10532
rect 11532 10520 11560 10619
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 11882 10616 11888 10668
rect 11940 10616 11946 10668
rect 12066 10616 12072 10668
rect 12124 10616 12130 10668
rect 13262 10616 13268 10668
rect 13320 10616 13326 10668
rect 13354 10616 13360 10668
rect 13412 10665 13418 10668
rect 13412 10659 13440 10665
rect 13428 10625 13440 10659
rect 13412 10619 13440 10625
rect 13412 10616 13418 10619
rect 11900 10588 11928 10616
rect 12345 10591 12403 10597
rect 12345 10588 12357 10591
rect 11900 10560 12357 10588
rect 12345 10557 12357 10560
rect 12391 10557 12403 10591
rect 12345 10551 12403 10557
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12492 10560 12541 10588
rect 12492 10548 12498 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 12894 10548 12900 10600
rect 12952 10588 12958 10600
rect 12989 10591 13047 10597
rect 12989 10588 13001 10591
rect 12952 10560 13001 10588
rect 12952 10548 12958 10560
rect 12989 10557 13001 10560
rect 13035 10557 13047 10591
rect 12989 10551 13047 10557
rect 13538 10548 13544 10600
rect 13596 10548 13602 10600
rect 11532 10492 13124 10520
rect 9784 10424 10732 10452
rect 10778 10412 10784 10464
rect 10836 10452 10842 10464
rect 12526 10452 12532 10464
rect 10836 10424 12532 10452
rect 10836 10412 10842 10424
rect 12526 10412 12532 10424
rect 12584 10412 12590 10464
rect 13096 10452 13124 10492
rect 13998 10452 14004 10464
rect 13096 10424 14004 10452
rect 13998 10412 14004 10424
rect 14056 10412 14062 10464
rect 1104 10362 14536 10384
rect 1104 10310 2629 10362
rect 2681 10310 2693 10362
rect 2745 10310 2757 10362
rect 2809 10310 2821 10362
rect 2873 10310 2885 10362
rect 2937 10310 5987 10362
rect 6039 10310 6051 10362
rect 6103 10310 6115 10362
rect 6167 10310 6179 10362
rect 6231 10310 6243 10362
rect 6295 10310 9345 10362
rect 9397 10310 9409 10362
rect 9461 10310 9473 10362
rect 9525 10310 9537 10362
rect 9589 10310 9601 10362
rect 9653 10310 12703 10362
rect 12755 10310 12767 10362
rect 12819 10310 12831 10362
rect 12883 10310 12895 10362
rect 12947 10310 12959 10362
rect 13011 10310 14536 10362
rect 1104 10288 14536 10310
rect 2958 10208 2964 10260
rect 3016 10208 3022 10260
rect 5718 10208 5724 10260
rect 5776 10208 5782 10260
rect 6546 10208 6552 10260
rect 6604 10208 6610 10260
rect 6730 10208 6736 10260
rect 6788 10208 6794 10260
rect 10502 10208 10508 10260
rect 10560 10248 10566 10260
rect 10781 10251 10839 10257
rect 10781 10248 10793 10251
rect 10560 10220 10793 10248
rect 10560 10208 10566 10220
rect 10781 10217 10793 10220
rect 10827 10217 10839 10251
rect 10781 10211 10839 10217
rect 11606 10208 11612 10260
rect 11664 10248 11670 10260
rect 12713 10251 12771 10257
rect 12713 10248 12725 10251
rect 11664 10220 12725 10248
rect 11664 10208 11670 10220
rect 12713 10217 12725 10220
rect 12759 10217 12771 10251
rect 12713 10211 12771 10217
rect 6365 10183 6423 10189
rect 6365 10149 6377 10183
rect 6411 10180 6423 10183
rect 6564 10180 6592 10208
rect 6411 10152 6592 10180
rect 6411 10149 6423 10152
rect 6365 10143 6423 10149
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6748 10112 6776 10208
rect 7098 10180 7104 10192
rect 7024 10152 7104 10180
rect 5951 10084 6776 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6822 10072 6828 10124
rect 6880 10072 6886 10124
rect 1394 10004 1400 10056
rect 1452 10004 1458 10056
rect 1671 10047 1729 10053
rect 1671 10013 1683 10047
rect 1717 10044 1729 10047
rect 1717 10016 1900 10044
rect 1717 10013 1729 10016
rect 1671 10007 1729 10013
rect 1872 9988 1900 10016
rect 2774 10004 2780 10056
rect 2832 10004 2838 10056
rect 5626 10004 5632 10056
rect 5684 10004 5690 10056
rect 6273 10047 6331 10053
rect 6273 10013 6285 10047
rect 6319 10044 6331 10047
rect 6319 10016 6500 10044
rect 6319 10013 6331 10016
rect 6273 10007 6331 10013
rect 1854 9936 1860 9988
rect 1912 9936 1918 9988
rect 6362 9936 6368 9988
rect 6420 9936 6426 9988
rect 2409 9911 2467 9917
rect 2409 9877 2421 9911
rect 2455 9908 2467 9911
rect 2498 9908 2504 9920
rect 2455 9880 2504 9908
rect 2455 9877 2467 9880
rect 2409 9871 2467 9877
rect 2498 9868 2504 9880
rect 2556 9868 2562 9920
rect 4706 9868 4712 9920
rect 4764 9908 4770 9920
rect 5905 9911 5963 9917
rect 5905 9908 5917 9911
rect 4764 9880 5917 9908
rect 4764 9868 4770 9880
rect 5905 9877 5917 9880
rect 5951 9877 5963 9911
rect 5905 9871 5963 9877
rect 6089 9911 6147 9917
rect 6089 9877 6101 9911
rect 6135 9908 6147 9911
rect 6380 9908 6408 9936
rect 6135 9880 6408 9908
rect 6472 9908 6500 10016
rect 6546 10004 6552 10056
rect 6604 10004 6610 10056
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 7024 10044 7052 10152
rect 7098 10140 7104 10152
rect 7156 10140 7162 10192
rect 7208 10152 7420 10180
rect 7208 10124 7236 10152
rect 7190 10072 7196 10124
rect 7248 10072 7254 10124
rect 7282 10072 7288 10124
rect 7340 10072 7346 10124
rect 7392 10112 7420 10152
rect 9582 10140 9588 10192
rect 9640 10140 9646 10192
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7392 10084 7849 10112
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 8662 10072 8668 10124
rect 8720 10112 8726 10124
rect 9125 10115 9183 10121
rect 9125 10112 9137 10115
rect 8720 10084 9137 10112
rect 8720 10072 8726 10084
rect 9125 10081 9137 10084
rect 9171 10112 9183 10115
rect 9214 10112 9220 10124
rect 9171 10084 9220 10112
rect 9171 10081 9183 10084
rect 9125 10075 9183 10081
rect 9214 10072 9220 10084
rect 9272 10072 9278 10124
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 9876 10112 10042 10120
rect 9548 10092 10042 10112
rect 9548 10084 9904 10092
rect 9548 10072 9554 10084
rect 6687 10016 7052 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 7558 10004 7564 10056
rect 7616 10004 7622 10056
rect 7650 10004 7656 10056
rect 7708 10053 7714 10056
rect 7708 10047 7736 10053
rect 7724 10013 7736 10047
rect 7708 10007 7736 10013
rect 7708 10004 7714 10007
rect 8846 10004 8852 10056
rect 8904 10044 8910 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8904 10016 8953 10044
rect 8904 10004 8910 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 9858 10004 9864 10056
rect 9916 10004 9922 10056
rect 10014 10053 10042 10092
rect 10778 10072 10784 10124
rect 10836 10072 10842 10124
rect 11517 10115 11575 10121
rect 11517 10112 11529 10115
rect 10980 10084 11529 10112
rect 9999 10047 10057 10053
rect 9999 10013 10011 10047
rect 10045 10013 10057 10047
rect 9999 10007 10057 10013
rect 10134 10004 10140 10056
rect 10192 10004 10198 10056
rect 10796 10020 10824 10072
rect 10873 10047 10931 10053
rect 10873 10020 10885 10047
rect 10796 10013 10885 10020
rect 10919 10013 10931 10047
rect 10796 10007 10931 10013
rect 10796 9992 10916 10007
rect 8481 9911 8539 9917
rect 8481 9908 8493 9911
rect 6472 9880 8493 9908
rect 6135 9877 6147 9880
rect 6089 9871 6147 9877
rect 8481 9877 8493 9880
rect 8527 9877 8539 9911
rect 8481 9871 8539 9877
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 9858 9908 9864 9920
rect 9640 9880 9864 9908
rect 9640 9868 9646 9880
rect 9858 9868 9864 9880
rect 9916 9908 9922 9920
rect 10980 9908 11008 10084
rect 11517 10081 11529 10084
rect 11563 10081 11575 10115
rect 11517 10075 11575 10081
rect 11606 10072 11612 10124
rect 11664 10112 11670 10124
rect 11808 10112 11928 10120
rect 11664 10092 11928 10112
rect 11664 10084 11836 10092
rect 11664 10072 11670 10084
rect 11054 10004 11060 10056
rect 11112 10004 11118 10056
rect 11790 10004 11796 10056
rect 11848 10004 11854 10056
rect 11900 10053 11928 10092
rect 12805 10115 12863 10121
rect 12805 10081 12817 10115
rect 12851 10112 12863 10115
rect 14090 10112 14096 10124
rect 12851 10084 14096 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 14090 10072 14096 10084
rect 14148 10072 14154 10124
rect 11900 10047 11968 10053
rect 11900 10016 11922 10047
rect 11910 10013 11922 10016
rect 11956 10013 11968 10047
rect 11910 10007 11968 10013
rect 12066 10004 12072 10056
rect 12124 10004 12130 10056
rect 13081 10047 13139 10053
rect 13081 10013 13093 10047
rect 13127 10013 13139 10047
rect 13081 10007 13139 10013
rect 9916 9880 11008 9908
rect 11072 9908 11100 10004
rect 11606 9908 11612 9920
rect 11072 9880 11612 9908
rect 9916 9868 9922 9880
rect 11606 9868 11612 9880
rect 11664 9868 11670 9920
rect 11790 9868 11796 9920
rect 11848 9908 11854 9920
rect 12158 9908 12164 9920
rect 11848 9880 12164 9908
rect 11848 9868 11854 9880
rect 12158 9868 12164 9880
rect 12216 9868 12222 9920
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 13096 9908 13124 10007
rect 12400 9880 13124 9908
rect 12400 9868 12406 9880
rect 1104 9818 14696 9840
rect 1104 9766 4308 9818
rect 4360 9766 4372 9818
rect 4424 9766 4436 9818
rect 4488 9766 4500 9818
rect 4552 9766 4564 9818
rect 4616 9766 7666 9818
rect 7718 9766 7730 9818
rect 7782 9766 7794 9818
rect 7846 9766 7858 9818
rect 7910 9766 7922 9818
rect 7974 9766 11024 9818
rect 11076 9766 11088 9818
rect 11140 9766 11152 9818
rect 11204 9766 11216 9818
rect 11268 9766 11280 9818
rect 11332 9766 14382 9818
rect 14434 9766 14446 9818
rect 14498 9766 14510 9818
rect 14562 9766 14574 9818
rect 14626 9766 14638 9818
rect 14690 9766 14696 9818
rect 1104 9744 14696 9766
rect 6822 9664 6828 9716
rect 6880 9704 6886 9716
rect 6880 9676 8156 9704
rect 6880 9664 6886 9676
rect 1762 9636 1768 9648
rect 1688 9608 1768 9636
rect 1688 9607 1716 9608
rect 1655 9601 1716 9607
rect 1655 9567 1667 9601
rect 1701 9570 1716 9601
rect 1762 9596 1768 9608
rect 1820 9596 1826 9648
rect 8128 9636 8156 9676
rect 8202 9664 8208 9716
rect 8260 9704 8266 9716
rect 8570 9704 8576 9716
rect 8260 9676 8576 9704
rect 8260 9664 8266 9676
rect 8570 9664 8576 9676
rect 8628 9664 8634 9716
rect 9582 9704 9588 9716
rect 8772 9676 9588 9704
rect 8772 9636 8800 9676
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 9674 9664 9680 9716
rect 9732 9704 9738 9716
rect 12434 9704 12440 9716
rect 9732 9676 12440 9704
rect 9732 9664 9738 9676
rect 12434 9664 12440 9676
rect 12492 9704 12498 9716
rect 13814 9704 13820 9716
rect 12492 9676 13820 9704
rect 12492 9664 12498 9676
rect 13814 9664 13820 9676
rect 13872 9664 13878 9716
rect 8128 9608 8800 9636
rect 11606 9596 11612 9648
rect 11664 9636 11670 9648
rect 11664 9608 12204 9636
rect 11664 9596 11670 9608
rect 1701 9567 1713 9570
rect 1655 9561 1713 9567
rect 8294 9528 8300 9580
rect 8352 9568 8358 9580
rect 8570 9568 8576 9580
rect 8352 9540 8576 9568
rect 8352 9528 8358 9540
rect 8570 9528 8576 9540
rect 8628 9568 8634 9580
rect 9401 9571 9459 9577
rect 9401 9568 9413 9571
rect 8628 9540 9413 9568
rect 8628 9528 8634 9540
rect 9401 9537 9413 9540
rect 9447 9537 9459 9571
rect 9401 9531 9459 9537
rect 10134 9528 10140 9580
rect 10192 9528 10198 9580
rect 10226 9528 10232 9580
rect 10284 9577 10290 9580
rect 10284 9571 10312 9577
rect 10300 9537 10312 9571
rect 10284 9531 10312 9537
rect 10284 9528 10290 9531
rect 10410 9528 10416 9580
rect 10468 9528 10474 9580
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9537 12127 9571
rect 12069 9531 12127 9537
rect 1394 9460 1400 9512
rect 1452 9460 1458 9512
rect 9214 9460 9220 9512
rect 9272 9460 9278 9512
rect 9766 9500 9772 9512
rect 9646 9472 9772 9500
rect 9646 9432 9674 9472
rect 9766 9460 9772 9472
rect 9824 9500 9830 9512
rect 9824 9472 11376 9500
rect 9824 9460 9830 9472
rect 11348 9444 11376 9472
rect 7392 9404 9674 9432
rect 7392 9376 7420 9404
rect 9858 9392 9864 9444
rect 9916 9392 9922 9444
rect 10870 9392 10876 9444
rect 10928 9432 10934 9444
rect 11057 9435 11115 9441
rect 11057 9432 11069 9435
rect 10928 9404 11069 9432
rect 10928 9392 10934 9404
rect 11057 9401 11069 9404
rect 11103 9401 11115 9435
rect 11057 9395 11115 9401
rect 11330 9392 11336 9444
rect 11388 9392 11394 9444
rect 12084 9432 12112 9531
rect 12176 9512 12204 9608
rect 14182 9596 14188 9648
rect 14240 9596 14246 9648
rect 12342 9528 12348 9580
rect 12400 9528 12406 9580
rect 13446 9577 13452 9580
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 13403 9571 13452 9577
rect 13403 9537 13415 9571
rect 13449 9537 13452 9571
rect 13403 9531 13452 9537
rect 12158 9460 12164 9512
rect 12216 9500 12222 9512
rect 12529 9503 12587 9509
rect 12529 9500 12541 9503
rect 12216 9472 12541 9500
rect 12216 9460 12222 9472
rect 12529 9469 12541 9472
rect 12575 9469 12587 9503
rect 12529 9463 12587 9469
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 13280 9500 13308 9531
rect 13446 9528 13452 9531
rect 13504 9528 13510 9580
rect 12676 9472 13308 9500
rect 13541 9503 13599 9509
rect 12676 9460 12682 9472
rect 13541 9469 13553 9503
rect 13587 9500 13599 9503
rect 13722 9500 13728 9512
rect 13587 9472 13728 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 13722 9460 13728 9472
rect 13780 9460 13786 9512
rect 12989 9435 13047 9441
rect 12084 9404 12940 9432
rect 2406 9324 2412 9376
rect 2464 9324 2470 9376
rect 7374 9324 7380 9376
rect 7432 9324 7438 9376
rect 9766 9324 9772 9376
rect 9824 9364 9830 9376
rect 12161 9367 12219 9373
rect 12161 9364 12173 9367
rect 9824 9336 12173 9364
rect 9824 9324 9830 9336
rect 12161 9333 12173 9336
rect 12207 9364 12219 9367
rect 12618 9364 12624 9376
rect 12207 9336 12624 9364
rect 12207 9333 12219 9336
rect 12161 9327 12219 9333
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 12912 9364 12940 9404
rect 12989 9401 13001 9435
rect 13035 9432 13047 9435
rect 13078 9432 13084 9444
rect 13035 9404 13084 9432
rect 13035 9401 13047 9404
rect 12989 9395 13047 9401
rect 13078 9392 13084 9404
rect 13136 9392 13142 9444
rect 13998 9364 14004 9376
rect 12912 9336 14004 9364
rect 13998 9324 14004 9336
rect 14056 9324 14062 9376
rect 1104 9274 14536 9296
rect 1104 9222 2629 9274
rect 2681 9222 2693 9274
rect 2745 9222 2757 9274
rect 2809 9222 2821 9274
rect 2873 9222 2885 9274
rect 2937 9222 5987 9274
rect 6039 9222 6051 9274
rect 6103 9222 6115 9274
rect 6167 9222 6179 9274
rect 6231 9222 6243 9274
rect 6295 9222 9345 9274
rect 9397 9222 9409 9274
rect 9461 9222 9473 9274
rect 9525 9222 9537 9274
rect 9589 9222 9601 9274
rect 9653 9222 12703 9274
rect 12755 9222 12767 9274
rect 12819 9222 12831 9274
rect 12883 9222 12895 9274
rect 12947 9222 12959 9274
rect 13011 9222 14536 9274
rect 1104 9200 14536 9222
rect 1762 9120 1768 9172
rect 1820 9160 1826 9172
rect 11333 9163 11391 9169
rect 1820 9132 11284 9160
rect 1820 9120 1826 9132
rect 2406 9052 2412 9104
rect 2464 9052 2470 9104
rect 8481 9095 8539 9101
rect 8481 9061 8493 9095
rect 8527 9092 8539 9095
rect 8527 9064 10297 9092
rect 8527 9061 8539 9064
rect 8481 9055 8539 9061
rect 2038 8916 2044 8968
rect 2096 8956 2102 8968
rect 2225 8959 2283 8965
rect 2096 8928 2176 8956
rect 2096 8916 2102 8928
rect 1489 8891 1547 8897
rect 1489 8857 1501 8891
rect 1535 8888 1547 8891
rect 2148 8888 2176 8928
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 2424 8956 2452 9052
rect 9677 9027 9735 9033
rect 9677 8993 9689 9027
rect 9723 9024 9735 9027
rect 9766 9024 9772 9036
rect 9723 8996 9772 9024
rect 9723 8993 9735 8996
rect 9677 8987 9735 8993
rect 9766 8984 9772 8996
rect 9824 8984 9830 9036
rect 9858 8984 9864 9036
rect 9916 9024 9922 9036
rect 10137 9027 10195 9033
rect 10137 9024 10149 9027
rect 9916 8996 10149 9024
rect 9916 8984 9922 8996
rect 10137 8993 10149 8996
rect 10183 8993 10195 9027
rect 10269 9024 10297 9064
rect 10686 9024 10692 9036
rect 10269 8996 10692 9024
rect 10137 8987 10195 8993
rect 10686 8984 10692 8996
rect 10744 8984 10750 9036
rect 2271 8928 2452 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 2498 8916 2504 8968
rect 2556 8916 2562 8968
rect 2590 8916 2596 8968
rect 2648 8916 2654 8968
rect 4798 8916 4804 8968
rect 4856 8956 4862 8968
rect 7374 8956 7380 8968
rect 4856 8928 7380 8956
rect 4856 8916 4862 8928
rect 7374 8916 7380 8928
rect 7432 8956 7438 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 7432 8928 7481 8956
rect 7432 8916 7438 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7727 8959 7785 8965
rect 7727 8956 7739 8959
rect 7469 8919 7527 8925
rect 7668 8928 7739 8956
rect 2685 8891 2743 8897
rect 2685 8888 2697 8891
rect 1535 8860 2084 8888
rect 2148 8860 2697 8888
rect 1535 8857 1547 8860
rect 1489 8851 1547 8857
rect 842 8780 848 8832
rect 900 8820 906 8832
rect 2056 8829 2084 8860
rect 2685 8857 2697 8860
rect 2731 8857 2743 8891
rect 2685 8851 2743 8857
rect 1581 8823 1639 8829
rect 1581 8820 1593 8823
rect 900 8792 1593 8820
rect 900 8780 906 8792
rect 1581 8789 1593 8792
rect 1627 8789 1639 8823
rect 1581 8783 1639 8789
rect 2041 8823 2099 8829
rect 2041 8789 2053 8823
rect 2087 8789 2099 8823
rect 2041 8783 2099 8789
rect 2314 8780 2320 8832
rect 2372 8780 2378 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 7282 8820 7288 8832
rect 5592 8792 7288 8820
rect 5592 8780 5598 8792
rect 7282 8780 7288 8792
rect 7340 8820 7346 8832
rect 7668 8820 7696 8928
rect 7727 8925 7739 8928
rect 7773 8925 7785 8959
rect 7727 8919 7785 8925
rect 8478 8916 8484 8968
rect 8536 8956 8542 8968
rect 9493 8959 9551 8965
rect 9493 8956 9505 8959
rect 8536 8928 9505 8956
rect 8536 8916 8542 8928
rect 9493 8925 9505 8928
rect 9539 8925 9551 8959
rect 9493 8919 9551 8925
rect 10410 8916 10416 8968
rect 10468 8916 10474 8968
rect 10502 8916 10508 8968
rect 10560 8965 10566 8968
rect 10560 8959 10588 8965
rect 10576 8925 10588 8959
rect 11256 8956 11284 9132
rect 11333 9129 11345 9163
rect 11379 9160 11391 9163
rect 11514 9160 11520 9172
rect 11379 9132 11520 9160
rect 11379 9129 11391 9132
rect 11333 9123 11391 9129
rect 11514 9120 11520 9132
rect 11572 9120 11578 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12437 9163 12495 9169
rect 12437 9160 12449 9163
rect 11756 9132 12449 9160
rect 11756 9120 11762 9132
rect 12437 9129 12449 9132
rect 12483 9129 12495 9163
rect 12437 9123 12495 9129
rect 13814 9120 13820 9172
rect 13872 9160 13878 9172
rect 13909 9163 13967 9169
rect 13909 9160 13921 9163
rect 13872 9132 13921 9160
rect 13872 9120 13878 9132
rect 13909 9129 13921 9132
rect 13955 9129 13967 9163
rect 13909 9123 13967 9129
rect 12618 9052 12624 9104
rect 12676 9092 12682 9104
rect 12676 9064 13952 9092
rect 12676 9052 12682 9064
rect 13924 9036 13952 9064
rect 11330 8984 11336 9036
rect 11388 9024 11394 9036
rect 11425 9027 11483 9033
rect 11425 9024 11437 9027
rect 11388 8996 11437 9024
rect 11388 8984 11394 8996
rect 11425 8993 11437 8996
rect 11471 8993 11483 9027
rect 11425 8987 11483 8993
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 13081 9027 13139 9033
rect 13081 9024 13093 9027
rect 12584 8996 13093 9024
rect 12584 8984 12590 8996
rect 13081 8993 13093 8996
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 13906 8984 13912 9036
rect 13964 8984 13970 9036
rect 11667 8959 11725 8965
rect 11667 8956 11679 8959
rect 11256 8928 11679 8956
rect 10560 8919 10588 8925
rect 11667 8925 11679 8928
rect 11713 8956 11725 8959
rect 12618 8956 12624 8968
rect 11713 8928 12624 8956
rect 11713 8925 11725 8928
rect 11667 8919 11725 8925
rect 10560 8916 10566 8919
rect 12618 8916 12624 8928
rect 12676 8916 12682 8968
rect 12805 8959 12863 8965
rect 12805 8925 12817 8959
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 13725 8959 13783 8965
rect 13725 8925 13737 8959
rect 13771 8956 13783 8959
rect 14826 8956 14832 8968
rect 13771 8928 14832 8956
rect 13771 8925 13783 8928
rect 13725 8919 13783 8925
rect 12820 8888 12848 8919
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 14182 8888 14188 8900
rect 12820 8860 14188 8888
rect 14182 8848 14188 8860
rect 14240 8848 14246 8900
rect 7340 8792 7696 8820
rect 7340 8780 7346 8792
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 10502 8820 10508 8832
rect 8444 8792 10508 8820
rect 8444 8780 8450 8792
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10686 8780 10692 8832
rect 10744 8820 10750 8832
rect 12066 8820 12072 8832
rect 10744 8792 12072 8820
rect 10744 8780 10750 8792
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12526 8780 12532 8832
rect 12584 8820 12590 8832
rect 13170 8820 13176 8832
rect 12584 8792 13176 8820
rect 12584 8780 12590 8792
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 1104 8730 14696 8752
rect 1104 8678 4308 8730
rect 4360 8678 4372 8730
rect 4424 8678 4436 8730
rect 4488 8678 4500 8730
rect 4552 8678 4564 8730
rect 4616 8678 7666 8730
rect 7718 8678 7730 8730
rect 7782 8678 7794 8730
rect 7846 8678 7858 8730
rect 7910 8678 7922 8730
rect 7974 8678 11024 8730
rect 11076 8678 11088 8730
rect 11140 8678 11152 8730
rect 11204 8678 11216 8730
rect 11268 8678 11280 8730
rect 11332 8678 14382 8730
rect 14434 8678 14446 8730
rect 14498 8678 14510 8730
rect 14562 8678 14574 8730
rect 14626 8678 14638 8730
rect 14690 8678 14696 8730
rect 1104 8656 14696 8678
rect 2314 8576 2320 8628
rect 2372 8576 2378 8628
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 6641 8619 6699 8625
rect 6641 8616 6653 8619
rect 2648 8588 6653 8616
rect 2648 8576 2654 8588
rect 6641 8585 6653 8588
rect 6687 8585 6699 8619
rect 6641 8579 6699 8585
rect 8846 8576 8852 8628
rect 8904 8576 8910 8628
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 10735 8619 10793 8625
rect 10735 8616 10747 8619
rect 10376 8588 10747 8616
rect 10376 8576 10382 8588
rect 10735 8585 10747 8588
rect 10781 8616 10793 8619
rect 11790 8616 11796 8628
rect 10781 8588 11796 8616
rect 10781 8585 10793 8588
rect 10735 8579 10793 8585
rect 11790 8576 11796 8588
rect 11848 8576 11854 8628
rect 12406 8588 13308 8616
rect 1489 8551 1547 8557
rect 1489 8517 1501 8551
rect 1535 8548 1547 8551
rect 2332 8548 2360 8576
rect 5902 8548 5908 8560
rect 1535 8520 2360 8548
rect 5184 8520 5908 8548
rect 1535 8517 1547 8520
rect 5184 8519 5212 8520
rect 1489 8511 1547 8517
rect 5151 8513 5212 8519
rect 4798 8440 4804 8492
rect 4856 8480 4862 8492
rect 4893 8483 4951 8489
rect 4893 8480 4905 8483
rect 4856 8452 4905 8480
rect 4856 8440 4862 8452
rect 4893 8449 4905 8452
rect 4939 8449 4951 8483
rect 5151 8479 5163 8513
rect 5197 8482 5212 8513
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 8864 8548 8892 8576
rect 11698 8548 11704 8560
rect 6380 8520 7052 8548
rect 8864 8520 9996 8548
rect 6380 8489 6408 8520
rect 6365 8483 6423 8489
rect 5197 8479 5209 8482
rect 6365 8480 6377 8483
rect 5151 8473 5209 8479
rect 4893 8443 4951 8449
rect 5920 8452 6377 8480
rect 1670 8304 1676 8356
rect 1728 8304 1734 8356
rect 5920 8353 5948 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 6730 8440 6736 8492
rect 6788 8440 6794 8492
rect 7024 8489 7052 8520
rect 7009 8483 7067 8489
rect 7009 8449 7021 8483
rect 7055 8449 7067 8483
rect 7009 8443 7067 8449
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 9861 8483 9919 8489
rect 9861 8449 9873 8483
rect 9907 8449 9919 8483
rect 9861 8443 9919 8449
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 7101 8415 7159 8421
rect 7101 8412 7113 8415
rect 6687 8384 7113 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 7101 8381 7113 8384
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 8294 8372 8300 8424
rect 8352 8412 8358 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8352 8384 8585 8412
rect 8352 8372 8358 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 5905 8347 5963 8353
rect 5905 8313 5917 8347
rect 5951 8313 5963 8347
rect 5905 8307 5963 8313
rect 6457 8347 6515 8353
rect 6457 8313 6469 8347
rect 6503 8344 6515 8347
rect 6825 8347 6883 8353
rect 6825 8344 6837 8347
rect 6503 8316 6837 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 6825 8313 6837 8316
rect 6871 8313 6883 8347
rect 6825 8307 6883 8313
rect 8202 8304 8208 8356
rect 8260 8344 8266 8356
rect 8481 8347 8539 8353
rect 8481 8344 8493 8347
rect 8260 8316 8493 8344
rect 8260 8304 8266 8316
rect 8481 8313 8493 8316
rect 8527 8313 8539 8347
rect 9876 8344 9904 8443
rect 9968 8412 9996 8520
rect 10244 8520 11704 8548
rect 10244 8489 10272 8520
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 10229 8483 10287 8489
rect 10229 8449 10241 8483
rect 10275 8449 10287 8483
rect 10229 8443 10287 8449
rect 10505 8483 10563 8489
rect 10505 8449 10517 8483
rect 10551 8480 10563 8483
rect 11422 8480 11428 8492
rect 10551 8452 11428 8480
rect 10551 8449 10563 8452
rect 10505 8443 10563 8449
rect 11422 8440 11428 8452
rect 11480 8440 11486 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8480 11851 8483
rect 12158 8480 12164 8492
rect 11839 8452 12164 8480
rect 11839 8449 11851 8452
rect 11793 8443 11851 8449
rect 12158 8440 12164 8452
rect 12216 8440 12222 8492
rect 10413 8415 10471 8421
rect 10413 8412 10425 8415
rect 9968 8384 10425 8412
rect 10413 8381 10425 8384
rect 10459 8412 10471 8415
rect 10870 8412 10876 8424
rect 10459 8384 10876 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 11296 8384 11529 8412
rect 11296 8372 11302 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 11146 8344 11152 8356
rect 9876 8316 11152 8344
rect 8481 8307 8539 8313
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 12406 8344 12434 8588
rect 12618 8508 12624 8560
rect 12676 8508 12682 8560
rect 13280 8548 13308 8588
rect 13538 8576 13544 8628
rect 13596 8576 13602 8628
rect 14093 8619 14151 8625
rect 14093 8585 14105 8619
rect 14139 8585 14151 8619
rect 14093 8579 14151 8585
rect 14108 8548 14136 8579
rect 13280 8520 14136 8548
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12636 8480 12664 8508
rect 12771 8483 12829 8489
rect 12771 8480 12783 8483
rect 12636 8452 12783 8480
rect 12771 8449 12783 8452
rect 12817 8449 12829 8483
rect 12771 8443 12829 8449
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14001 8483 14059 8489
rect 14001 8480 14013 8483
rect 13688 8452 14013 8480
rect 13688 8440 13694 8452
rect 14001 8449 14013 8452
rect 14047 8449 14059 8483
rect 14001 8443 14059 8449
rect 11256 8316 12434 8344
rect 8110 8236 8116 8288
rect 8168 8276 8174 8288
rect 8386 8276 8392 8288
rect 8168 8248 8392 8276
rect 8168 8236 8174 8248
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 9950 8236 9956 8288
rect 10008 8236 10014 8288
rect 10594 8236 10600 8288
rect 10652 8276 10658 8288
rect 11256 8276 11284 8316
rect 10652 8248 11284 8276
rect 10652 8236 10658 8248
rect 1104 8186 14536 8208
rect 1104 8134 2629 8186
rect 2681 8134 2693 8186
rect 2745 8134 2757 8186
rect 2809 8134 2821 8186
rect 2873 8134 2885 8186
rect 2937 8134 5987 8186
rect 6039 8134 6051 8186
rect 6103 8134 6115 8186
rect 6167 8134 6179 8186
rect 6231 8134 6243 8186
rect 6295 8134 9345 8186
rect 9397 8134 9409 8186
rect 9461 8134 9473 8186
rect 9525 8134 9537 8186
rect 9589 8134 9601 8186
rect 9653 8134 12703 8186
rect 12755 8134 12767 8186
rect 12819 8134 12831 8186
rect 12883 8134 12895 8186
rect 12947 8134 12959 8186
rect 13011 8134 14536 8186
rect 1104 8112 14536 8134
rect 6365 8075 6423 8081
rect 6365 8041 6377 8075
rect 6411 8072 6423 8075
rect 6730 8072 6736 8084
rect 6411 8044 6736 8072
rect 6411 8041 6423 8044
rect 6365 8035 6423 8041
rect 6730 8032 6736 8044
rect 6788 8032 6794 8084
rect 7190 8032 7196 8084
rect 7248 8032 7254 8084
rect 7926 8032 7932 8084
rect 7984 8072 7990 8084
rect 8938 8072 8944 8084
rect 7984 8044 8944 8072
rect 7984 8032 7990 8044
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9180 8044 11376 8072
rect 9180 8032 9186 8044
rect 6641 8007 6699 8013
rect 6641 7973 6653 8007
rect 6687 8004 6699 8007
rect 7208 8004 7236 8032
rect 6687 7976 7236 8004
rect 6687 7973 6699 7976
rect 6641 7967 6699 7973
rect 9582 7964 9588 8016
rect 9640 8004 9646 8016
rect 10134 8004 10140 8016
rect 9640 7976 10140 8004
rect 9640 7964 9646 7976
rect 10134 7964 10140 7976
rect 10192 7964 10198 8016
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 6972 7908 7328 7936
rect 6972 7896 6978 7908
rect 7300 7880 7328 7908
rect 7558 7896 7564 7948
rect 7616 7896 7622 7948
rect 7834 7896 7840 7948
rect 7892 7896 7898 7948
rect 8018 7945 8024 7948
rect 7975 7939 8024 7945
rect 7975 7905 7987 7939
rect 8021 7905 8024 7939
rect 7975 7899 8024 7905
rect 8018 7896 8024 7899
rect 8076 7896 8082 7948
rect 8110 7896 8116 7948
rect 8168 7896 8174 7948
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 9674 7936 9680 7948
rect 9364 7908 9680 7936
rect 9364 7896 9370 7908
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10008 7908 10241 7936
rect 10008 7896 10014 7908
rect 10229 7905 10241 7908
rect 10275 7905 10287 7939
rect 10229 7899 10287 7905
rect 10502 7896 10508 7948
rect 10560 7896 10566 7948
rect 10594 7896 10600 7948
rect 10652 7945 10658 7948
rect 10652 7939 10680 7945
rect 10668 7905 10680 7939
rect 10652 7899 10680 7905
rect 10652 7896 10658 7899
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 1671 7871 1729 7877
rect 1671 7837 1683 7871
rect 1717 7868 1729 7871
rect 5534 7868 5540 7880
rect 1717 7840 5540 7868
rect 1717 7837 1729 7840
rect 1671 7831 1729 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 6549 7871 6607 7877
rect 6549 7837 6561 7871
rect 6595 7868 6607 7871
rect 6595 7840 6776 7868
rect 6595 7837 6607 7840
rect 6549 7831 6607 7837
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 6748 7732 6776 7840
rect 6822 7828 6828 7880
rect 6880 7828 6886 7880
rect 7098 7828 7104 7880
rect 7156 7828 7162 7880
rect 7282 7828 7288 7880
rect 7340 7828 7346 7880
rect 9490 7828 9496 7880
rect 9548 7868 9554 7880
rect 9585 7871 9643 7877
rect 9585 7868 9597 7871
rect 9548 7840 9597 7868
rect 9548 7828 9554 7840
rect 9585 7837 9597 7840
rect 9631 7837 9643 7871
rect 9585 7831 9643 7837
rect 8757 7735 8815 7741
rect 8757 7732 8769 7735
rect 6748 7704 8769 7732
rect 8757 7701 8769 7704
rect 8803 7701 8815 7735
rect 9692 7732 9720 7896
rect 9766 7828 9772 7880
rect 9824 7828 9830 7880
rect 10778 7828 10784 7880
rect 10836 7828 10842 7880
rect 11348 7800 11376 8044
rect 11974 8032 11980 8084
rect 12032 8032 12038 8084
rect 13633 8075 13691 8081
rect 13633 8041 13645 8075
rect 13679 8072 13691 8075
rect 13722 8072 13728 8084
rect 13679 8044 13728 8072
rect 13679 8041 13691 8044
rect 13633 8035 13691 8041
rect 13722 8032 13728 8044
rect 13780 8032 13786 8084
rect 11701 7939 11759 7945
rect 11701 7905 11713 7939
rect 11747 7936 11759 7939
rect 11992 7936 12020 8032
rect 11747 7908 12020 7936
rect 11747 7905 11759 7908
rect 11701 7899 11759 7905
rect 12526 7896 12532 7948
rect 12584 7936 12590 7948
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12584 7908 12633 7936
rect 12584 7896 12590 7908
rect 12621 7905 12633 7908
rect 12667 7905 12679 7939
rect 12621 7899 12679 7905
rect 11425 7871 11483 7877
rect 11425 7837 11437 7871
rect 11471 7868 11483 7871
rect 11514 7868 11520 7880
rect 11471 7840 11520 7868
rect 11471 7837 11483 7840
rect 11425 7831 11483 7837
rect 11514 7828 11520 7840
rect 11572 7828 11578 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 11977 7871 12035 7877
rect 11977 7868 11989 7871
rect 11940 7840 11989 7868
rect 11940 7828 11946 7840
rect 11977 7837 11989 7840
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 12895 7871 12953 7877
rect 12895 7837 12907 7871
rect 12941 7868 12953 7871
rect 13262 7868 13268 7880
rect 12941 7840 13268 7868
rect 12941 7837 12953 7840
rect 12895 7831 12953 7837
rect 13262 7828 13268 7840
rect 13320 7828 13326 7880
rect 13630 7800 13636 7812
rect 11348 7772 13636 7800
rect 13630 7760 13636 7772
rect 13688 7760 13694 7812
rect 10502 7732 10508 7744
rect 9692 7704 10508 7732
rect 8757 7695 8815 7701
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 10778 7692 10784 7744
rect 10836 7732 10842 7744
rect 13170 7732 13176 7744
rect 10836 7704 13176 7732
rect 10836 7692 10842 7704
rect 13170 7692 13176 7704
rect 13228 7732 13234 7744
rect 13722 7732 13728 7744
rect 13228 7704 13728 7732
rect 13228 7692 13234 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 1104 7642 14696 7664
rect 1104 7590 4308 7642
rect 4360 7590 4372 7642
rect 4424 7590 4436 7642
rect 4488 7590 4500 7642
rect 4552 7590 4564 7642
rect 4616 7590 7666 7642
rect 7718 7590 7730 7642
rect 7782 7590 7794 7642
rect 7846 7590 7858 7642
rect 7910 7590 7922 7642
rect 7974 7590 11024 7642
rect 11076 7590 11088 7642
rect 11140 7590 11152 7642
rect 11204 7590 11216 7642
rect 11268 7590 11280 7642
rect 11332 7590 14382 7642
rect 14434 7590 14446 7642
rect 14498 7590 14510 7642
rect 14562 7590 14574 7642
rect 14626 7590 14638 7642
rect 14690 7590 14696 7642
rect 1104 7568 14696 7590
rect 1949 7531 2007 7537
rect 1949 7497 1961 7531
rect 1995 7497 2007 7531
rect 1949 7491 2007 7497
rect 1489 7463 1547 7469
rect 1489 7429 1501 7463
rect 1535 7460 1547 7463
rect 1964 7460 1992 7491
rect 2406 7488 2412 7540
rect 2464 7488 2470 7540
rect 6822 7488 6828 7540
rect 6880 7528 6886 7540
rect 9033 7531 9091 7537
rect 9033 7528 9045 7531
rect 6880 7500 9045 7528
rect 6880 7488 6886 7500
rect 9033 7497 9045 7500
rect 9079 7497 9091 7531
rect 9033 7491 9091 7497
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 11974 7528 11980 7540
rect 9180 7500 11980 7528
rect 9180 7488 9186 7500
rect 11974 7488 11980 7500
rect 12032 7528 12038 7540
rect 12526 7528 12532 7540
rect 12032 7500 12532 7528
rect 12032 7488 12038 7500
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 12989 7531 13047 7537
rect 12989 7497 13001 7531
rect 13035 7528 13047 7531
rect 13078 7528 13084 7540
rect 13035 7500 13084 7528
rect 13035 7497 13047 7500
rect 12989 7491 13047 7497
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 14274 7528 14280 7540
rect 13228 7500 14280 7528
rect 13228 7488 13234 7500
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 1535 7432 1992 7460
rect 1535 7429 1547 7432
rect 1489 7423 1547 7429
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2424 7392 2452 7488
rect 8938 7420 8944 7472
rect 8996 7460 9002 7472
rect 11701 7463 11759 7469
rect 8996 7432 9536 7460
rect 8996 7420 9002 7432
rect 2179 7364 2452 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 7190 7352 7196 7404
rect 7248 7352 7254 7404
rect 7377 7395 7435 7401
rect 7377 7361 7389 7395
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 842 7148 848 7200
rect 900 7188 906 7200
rect 1581 7191 1639 7197
rect 1581 7188 1593 7191
rect 900 7160 1593 7188
rect 900 7148 906 7160
rect 1581 7157 1593 7160
rect 1627 7157 1639 7191
rect 7392 7188 7420 7355
rect 8202 7352 8208 7404
rect 8260 7401 8266 7404
rect 8260 7395 8309 7401
rect 8260 7361 8263 7395
rect 8297 7361 8309 7395
rect 8260 7355 8309 7361
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9306 7392 9312 7404
rect 9263 7364 9312 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 8260 7352 8266 7355
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9508 7401 9536 7432
rect 11701 7429 11713 7463
rect 11747 7460 11759 7463
rect 14826 7460 14832 7472
rect 11747 7432 14832 7460
rect 11747 7429 11759 7432
rect 11701 7423 11759 7429
rect 14826 7420 14832 7432
rect 14884 7420 14890 7472
rect 9493 7395 9551 7401
rect 9493 7361 9505 7395
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 9582 7364 9812 7392
rect 7558 7284 7564 7336
rect 7616 7324 7622 7336
rect 7837 7327 7895 7333
rect 7837 7324 7849 7327
rect 7616 7296 7849 7324
rect 7616 7284 7622 7296
rect 7837 7293 7849 7296
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 7926 7284 7932 7336
rect 7984 7324 7990 7336
rect 8113 7327 8171 7333
rect 8113 7324 8125 7327
rect 7984 7296 8125 7324
rect 7984 7284 7990 7296
rect 8113 7293 8125 7296
rect 8159 7293 8171 7327
rect 8113 7287 8171 7293
rect 8386 7284 8392 7336
rect 8444 7284 8450 7336
rect 9582 7324 9610 7364
rect 9784 7358 9812 7364
rect 9048 7296 9610 7324
rect 9048 7188 9076 7296
rect 9674 7284 9680 7336
rect 9732 7284 9738 7336
rect 9784 7330 9904 7358
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 10502 7352 10508 7404
rect 10560 7401 10566 7404
rect 10560 7395 10588 7401
rect 10576 7361 10588 7395
rect 10560 7355 10588 7361
rect 10560 7352 10566 7355
rect 11422 7352 11428 7404
rect 11480 7392 11486 7404
rect 12219 7395 12277 7401
rect 12219 7392 12231 7395
rect 11480 7364 12231 7392
rect 11480 7352 11486 7364
rect 12219 7361 12231 7364
rect 12265 7361 12277 7395
rect 12219 7355 12277 7361
rect 13630 7352 13636 7404
rect 13688 7352 13694 7404
rect 9876 7324 9904 7330
rect 10428 7324 10456 7352
rect 9876 7296 10456 7324
rect 10686 7284 10692 7336
rect 10744 7284 10750 7336
rect 11974 7284 11980 7336
rect 12032 7284 12038 7336
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 9582 7216 9588 7268
rect 9640 7256 9646 7268
rect 9766 7256 9772 7268
rect 9640 7228 9772 7256
rect 9640 7216 9646 7228
rect 9766 7216 9772 7228
rect 9824 7216 9830 7268
rect 9950 7216 9956 7268
rect 10008 7256 10014 7268
rect 10134 7256 10140 7268
rect 10008 7228 10140 7256
rect 10008 7216 10014 7228
rect 10134 7216 10140 7228
rect 10192 7216 10198 7268
rect 7392 7160 9076 7188
rect 9401 7191 9459 7197
rect 1581 7151 1639 7157
rect 9401 7157 9413 7191
rect 9447 7188 9459 7191
rect 9674 7188 9680 7200
rect 9447 7160 9680 7188
rect 9447 7157 9459 7160
rect 9401 7151 9459 7157
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 10042 7148 10048 7200
rect 10100 7188 10106 7200
rect 10594 7188 10600 7200
rect 10100 7160 10600 7188
rect 10100 7148 10106 7160
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 11606 7188 11612 7200
rect 11379 7160 11612 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 11793 7191 11851 7197
rect 11793 7157 11805 7191
rect 11839 7188 11851 7191
rect 11882 7188 11888 7200
rect 11839 7160 11888 7188
rect 11839 7157 11851 7160
rect 11793 7151 11851 7157
rect 11882 7148 11888 7160
rect 11940 7148 11946 7200
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 13372 7188 13400 7287
rect 12308 7160 13400 7188
rect 12308 7148 12314 7160
rect 1104 7098 14536 7120
rect 1104 7046 2629 7098
rect 2681 7046 2693 7098
rect 2745 7046 2757 7098
rect 2809 7046 2821 7098
rect 2873 7046 2885 7098
rect 2937 7046 5987 7098
rect 6039 7046 6051 7098
rect 6103 7046 6115 7098
rect 6167 7046 6179 7098
rect 6231 7046 6243 7098
rect 6295 7046 9345 7098
rect 9397 7046 9409 7098
rect 9461 7046 9473 7098
rect 9525 7046 9537 7098
rect 9589 7046 9601 7098
rect 9653 7046 12703 7098
rect 12755 7046 12767 7098
rect 12819 7046 12831 7098
rect 12883 7046 12895 7098
rect 12947 7046 12959 7098
rect 13011 7046 14536 7098
rect 1104 7024 14536 7046
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 7837 6987 7895 6993
rect 7837 6984 7849 6987
rect 7616 6956 7849 6984
rect 7616 6944 7622 6956
rect 7837 6953 7849 6956
rect 7883 6953 7895 6987
rect 7837 6947 7895 6953
rect 7926 6944 7932 6996
rect 7984 6984 7990 6996
rect 8294 6984 8300 6996
rect 7984 6956 8300 6984
rect 7984 6944 7990 6956
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 9858 6984 9864 6996
rect 9692 6956 9864 6984
rect 8662 6808 8668 6860
rect 8720 6808 8726 6860
rect 8846 6808 8852 6860
rect 8904 6848 8910 6860
rect 8941 6851 8999 6857
rect 8941 6848 8953 6851
rect 8904 6820 8953 6848
rect 8904 6808 8910 6820
rect 8941 6817 8953 6820
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 9582 6808 9588 6860
rect 9640 6808 9646 6860
rect 9692 6848 9720 6956
rect 9858 6944 9864 6956
rect 9916 6984 9922 6996
rect 9916 6956 11836 6984
rect 9916 6944 9922 6956
rect 11808 6928 11836 6956
rect 11790 6876 11796 6928
rect 11848 6876 11854 6928
rect 11977 6919 12035 6925
rect 11977 6885 11989 6919
rect 12023 6885 12035 6919
rect 11977 6879 12035 6885
rect 9861 6851 9919 6857
rect 9861 6848 9873 6851
rect 9692 6820 9873 6848
rect 9861 6817 9873 6820
rect 9907 6817 9919 6851
rect 9861 6811 9919 6817
rect 10147 6851 10205 6857
rect 10147 6817 10159 6851
rect 10193 6848 10205 6851
rect 10502 6848 10508 6860
rect 10193 6820 10508 6848
rect 10193 6817 10205 6820
rect 10147 6811 10205 6817
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 11992 6848 12020 6879
rect 11992 6820 12374 6848
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 7099 6783 7157 6789
rect 7099 6749 7111 6783
rect 7145 6780 7157 6783
rect 8680 6780 8708 6808
rect 9125 6783 9183 6789
rect 9125 6780 9137 6783
rect 7145 6752 8248 6780
rect 8680 6752 9137 6780
rect 7145 6749 7157 6752
rect 7099 6743 7157 6749
rect 1486 6672 1492 6724
rect 1544 6672 1550 6724
rect 842 6604 848 6656
rect 900 6644 906 6656
rect 1581 6647 1639 6653
rect 1581 6644 1593 6647
rect 900 6616 1593 6644
rect 900 6604 906 6616
rect 1581 6613 1593 6616
rect 1627 6613 1639 6647
rect 6840 6644 6868 6743
rect 8220 6724 8248 6752
rect 9125 6749 9137 6752
rect 9171 6749 9183 6783
rect 9125 6743 9183 6749
rect 9950 6740 9956 6792
rect 10008 6789 10014 6792
rect 10008 6783 10036 6789
rect 10024 6749 10036 6783
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10008 6743 10036 6749
rect 10704 6752 10977 6780
rect 10008 6740 10014 6743
rect 8202 6672 8208 6724
rect 8260 6672 8266 6724
rect 7374 6644 7380 6656
rect 6840 6616 7380 6644
rect 1581 6607 1639 6613
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 10704 6644 10732 6752
rect 10965 6749 10977 6752
rect 11011 6749 11023 6783
rect 11238 6780 11244 6792
rect 11199 6752 11244 6780
rect 10965 6743 11023 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 11348 6752 13277 6780
rect 10870 6672 10876 6724
rect 10928 6712 10934 6724
rect 11348 6712 11376 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 10928 6684 11376 6712
rect 10928 6672 10934 6684
rect 11790 6672 11796 6724
rect 11848 6712 11854 6724
rect 12805 6715 12863 6721
rect 12805 6712 12817 6715
rect 11848 6684 12817 6712
rect 11848 6672 11854 6684
rect 12805 6681 12817 6684
rect 12851 6681 12863 6715
rect 12805 6675 12863 6681
rect 12897 6715 12955 6721
rect 12897 6681 12909 6715
rect 12943 6712 12955 6715
rect 13354 6712 13360 6724
rect 12943 6684 13360 6712
rect 12943 6681 12955 6684
rect 12897 6675 12955 6681
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 13446 6672 13452 6724
rect 13504 6712 13510 6724
rect 13633 6715 13691 6721
rect 13633 6712 13645 6715
rect 13504 6684 13645 6712
rect 13504 6672 13510 6684
rect 13633 6681 13645 6684
rect 13679 6681 13691 6715
rect 13633 6675 13691 6681
rect 9088 6616 10732 6644
rect 9088 6604 9094 6616
rect 10778 6604 10784 6656
rect 10836 6604 10842 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 12529 6647 12587 6653
rect 12529 6644 12541 6647
rect 11020 6616 12541 6644
rect 11020 6604 11026 6616
rect 12529 6613 12541 6616
rect 12575 6613 12587 6647
rect 12529 6607 12587 6613
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 13464 6644 13492 6672
rect 12676 6616 13492 6644
rect 13817 6647 13875 6653
rect 12676 6604 12682 6616
rect 13817 6613 13829 6647
rect 13863 6644 13875 6647
rect 15010 6644 15016 6656
rect 13863 6616 15016 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 1104 6554 14696 6576
rect 1104 6502 4308 6554
rect 4360 6502 4372 6554
rect 4424 6502 4436 6554
rect 4488 6502 4500 6554
rect 4552 6502 4564 6554
rect 4616 6502 7666 6554
rect 7718 6502 7730 6554
rect 7782 6502 7794 6554
rect 7846 6502 7858 6554
rect 7910 6502 7922 6554
rect 7974 6502 11024 6554
rect 11076 6502 11088 6554
rect 11140 6502 11152 6554
rect 11204 6502 11216 6554
rect 11268 6502 11280 6554
rect 11332 6502 14382 6554
rect 14434 6502 14446 6554
rect 14498 6502 14510 6554
rect 14562 6502 14574 6554
rect 14626 6502 14638 6554
rect 14690 6502 14696 6554
rect 1104 6480 14696 6502
rect 8941 6443 8999 6449
rect 8941 6409 8953 6443
rect 8987 6440 8999 6443
rect 9766 6440 9772 6452
rect 8987 6412 9772 6440
rect 8987 6409 8999 6412
rect 8941 6403 8999 6409
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 11882 6440 11888 6452
rect 10008 6412 11888 6440
rect 10008 6400 10014 6412
rect 11882 6400 11888 6412
rect 11940 6440 11946 6452
rect 14093 6443 14151 6449
rect 11940 6412 13124 6440
rect 11940 6400 11946 6412
rect 6454 6372 6460 6384
rect 1686 6344 6460 6372
rect 1686 6343 1714 6344
rect 1655 6337 1714 6343
rect 1655 6303 1667 6337
rect 1701 6306 1714 6337
rect 6454 6332 6460 6344
rect 6512 6372 6518 6384
rect 13096 6381 13124 6412
rect 14093 6409 14105 6443
rect 14139 6440 14151 6443
rect 15102 6440 15108 6452
rect 14139 6412 15108 6440
rect 14139 6409 14151 6412
rect 14093 6403 14151 6409
rect 15102 6400 15108 6412
rect 15160 6400 15166 6452
rect 12805 6375 12863 6381
rect 12805 6372 12817 6375
rect 6512 6344 8064 6372
rect 6512 6332 6518 6344
rect 1701 6303 1713 6306
rect 1655 6297 1713 6303
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7432 6276 7941 6304
rect 7432 6264 7438 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 8036 6304 8064 6344
rect 12802 6341 12817 6372
rect 12851 6341 12863 6375
rect 12802 6335 12863 6341
rect 13081 6375 13139 6381
rect 13081 6341 13093 6375
rect 13127 6341 13139 6375
rect 13081 6335 13139 6341
rect 8171 6307 8229 6313
rect 8171 6304 8183 6307
rect 8036 6276 8183 6304
rect 7929 6267 7987 6273
rect 8171 6273 8183 6276
rect 8217 6273 8229 6307
rect 8171 6267 8229 6273
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 8628 6276 9505 6304
rect 8628 6264 8634 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9674 6264 9680 6316
rect 9732 6264 9738 6316
rect 10318 6264 10324 6316
rect 10376 6313 10382 6316
rect 10376 6307 10404 6313
rect 10392 6273 10404 6307
rect 10376 6267 10404 6273
rect 10376 6264 10382 6267
rect 10502 6264 10508 6316
rect 10560 6264 10566 6316
rect 11701 6307 11759 6313
rect 11701 6273 11713 6307
rect 11747 6304 11759 6307
rect 12066 6304 12072 6316
rect 11747 6276 12072 6304
rect 11747 6273 11759 6276
rect 11701 6267 11759 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 12802 6304 12830 6335
rect 13446 6332 13452 6384
rect 13504 6372 13510 6384
rect 13541 6375 13599 6381
rect 13541 6372 13553 6375
rect 13504 6344 13553 6372
rect 13504 6332 13510 6344
rect 13541 6341 13553 6344
rect 13587 6341 13599 6375
rect 13541 6335 13599 6341
rect 13630 6332 13636 6384
rect 13688 6372 13694 6384
rect 13909 6375 13967 6381
rect 13909 6372 13921 6375
rect 13688 6344 13921 6372
rect 13688 6332 13694 6344
rect 13909 6341 13921 6344
rect 13955 6341 13967 6375
rect 13909 6335 13967 6341
rect 12544 6276 12830 6304
rect 1394 6196 1400 6248
rect 1452 6196 1458 6248
rect 9214 6196 9220 6248
rect 9272 6236 9278 6248
rect 9309 6239 9367 6245
rect 9309 6236 9321 6239
rect 9272 6208 9321 6236
rect 9272 6196 9278 6208
rect 9309 6205 9321 6208
rect 9355 6205 9367 6239
rect 9692 6236 9720 6264
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 9692 6208 10241 6236
rect 9309 6199 9367 6205
rect 10229 6205 10241 6208
rect 10275 6236 10287 6239
rect 10870 6236 10876 6248
rect 10275 6208 10876 6236
rect 10275 6205 10287 6208
rect 10229 6199 10287 6205
rect 1412 6100 1440 6196
rect 2314 6100 2320 6112
rect 1412 6072 2320 6100
rect 2314 6060 2320 6072
rect 2372 6060 2378 6112
rect 2406 6060 2412 6112
rect 2464 6060 2470 6112
rect 9324 6100 9352 6199
rect 10870 6196 10876 6208
rect 10928 6196 10934 6248
rect 11977 6239 12035 6245
rect 11977 6236 11989 6239
rect 10980 6208 11989 6236
rect 10980 6180 11008 6208
rect 11977 6205 11989 6208
rect 12023 6236 12035 6239
rect 12544 6236 12572 6276
rect 13170 6264 13176 6316
rect 13228 6264 13234 6316
rect 13722 6264 13728 6316
rect 13780 6264 13786 6316
rect 12023 6208 12572 6236
rect 13740 6222 13768 6264
rect 12023 6205 12035 6208
rect 11977 6199 12035 6205
rect 9950 6128 9956 6180
rect 10008 6128 10014 6180
rect 10962 6128 10968 6180
rect 11020 6128 11026 6180
rect 11072 6140 12664 6168
rect 11072 6100 11100 6140
rect 12636 6112 12664 6140
rect 9324 6072 11100 6100
rect 11146 6060 11152 6112
rect 11204 6060 11210 6112
rect 12618 6060 12624 6112
rect 12676 6060 12682 6112
rect 1104 6010 14536 6032
rect 1104 5958 2629 6010
rect 2681 5958 2693 6010
rect 2745 5958 2757 6010
rect 2809 5958 2821 6010
rect 2873 5958 2885 6010
rect 2937 5958 5987 6010
rect 6039 5958 6051 6010
rect 6103 5958 6115 6010
rect 6167 5958 6179 6010
rect 6231 5958 6243 6010
rect 6295 5958 9345 6010
rect 9397 5958 9409 6010
rect 9461 5958 9473 6010
rect 9525 5958 9537 6010
rect 9589 5958 9601 6010
rect 9653 5958 12703 6010
rect 12755 5958 12767 6010
rect 12819 5958 12831 6010
rect 12883 5958 12895 6010
rect 12947 5958 12959 6010
rect 13011 5958 14536 6010
rect 1104 5936 14536 5958
rect 1486 5856 1492 5908
rect 1544 5896 1550 5908
rect 2317 5899 2375 5905
rect 2317 5896 2329 5899
rect 1544 5868 2329 5896
rect 1544 5856 1550 5868
rect 2317 5865 2329 5868
rect 2363 5865 2375 5899
rect 2317 5859 2375 5865
rect 2406 5856 2412 5908
rect 2464 5856 2470 5908
rect 7374 5856 7380 5908
rect 7432 5856 7438 5908
rect 8297 5899 8355 5905
rect 8297 5865 8309 5899
rect 8343 5896 8355 5899
rect 8386 5896 8392 5908
rect 8343 5868 8392 5896
rect 8343 5865 8355 5868
rect 8297 5859 8355 5865
rect 8386 5856 8392 5868
rect 8444 5856 8450 5908
rect 8570 5856 8576 5908
rect 8628 5896 8634 5908
rect 12894 5896 12900 5908
rect 8628 5868 12900 5896
rect 8628 5856 8634 5868
rect 12894 5856 12900 5868
rect 12952 5896 12958 5908
rect 12952 5868 13216 5896
rect 12952 5856 12958 5868
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2424 5692 2452 5856
rect 7392 5828 7420 5856
rect 7300 5800 7420 5828
rect 7300 5769 7328 5800
rect 8662 5788 8668 5840
rect 8720 5828 8726 5840
rect 10962 5828 10968 5840
rect 8720 5800 10968 5828
rect 8720 5788 8726 5800
rect 10962 5788 10968 5800
rect 11020 5788 11026 5840
rect 13188 5828 13216 5868
rect 13630 5856 13636 5908
rect 13688 5856 13694 5908
rect 13648 5828 13676 5856
rect 13188 5800 13676 5828
rect 7285 5763 7343 5769
rect 7285 5729 7297 5763
rect 7331 5729 7343 5763
rect 10597 5763 10655 5769
rect 7285 5723 7343 5729
rect 8220 5732 8984 5760
rect 2501 5695 2559 5701
rect 2501 5692 2513 5695
rect 2424 5664 2513 5692
rect 2225 5655 2283 5661
rect 2501 5661 2513 5664
rect 2547 5661 2559 5695
rect 2501 5655 2559 5661
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5624 1547 5627
rect 2240 5624 2268 5655
rect 2590 5652 2596 5704
rect 2648 5692 2654 5704
rect 7300 5692 7328 5723
rect 2648 5664 7328 5692
rect 7559 5695 7617 5701
rect 2648 5652 2654 5664
rect 7559 5661 7571 5695
rect 7605 5692 7617 5695
rect 8220 5692 8248 5732
rect 8956 5704 8984 5732
rect 10597 5729 10609 5763
rect 10643 5760 10655 5763
rect 10686 5760 10692 5772
rect 10643 5732 10692 5760
rect 10643 5729 10655 5732
rect 10597 5723 10655 5729
rect 10686 5720 10692 5732
rect 10744 5720 10750 5772
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11146 5760 11152 5772
rect 10827 5732 11152 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5760 11299 5763
rect 11330 5760 11336 5772
rect 11287 5732 11336 5760
rect 11287 5729 11299 5732
rect 11241 5723 11299 5729
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 11514 5720 11520 5772
rect 11572 5720 11578 5772
rect 11606 5720 11612 5772
rect 11664 5769 11670 5772
rect 11664 5763 11692 5769
rect 11680 5729 11692 5763
rect 11664 5723 11692 5729
rect 11664 5720 11670 5723
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12492 5732 12541 5760
rect 12492 5720 12498 5732
rect 12529 5729 12541 5732
rect 12575 5729 12587 5763
rect 12529 5723 12587 5729
rect 7605 5664 8248 5692
rect 7605 5661 7617 5664
rect 7559 5655 7617 5661
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8938 5652 8944 5704
rect 8996 5652 9002 5704
rect 11790 5652 11796 5704
rect 11848 5652 11854 5704
rect 8312 5624 8340 5652
rect 1535 5596 2084 5624
rect 2240 5596 8340 5624
rect 1535 5593 1547 5596
rect 1489 5587 1547 5593
rect 1578 5516 1584 5568
rect 1636 5516 1642 5568
rect 2056 5565 2084 5596
rect 12434 5584 12440 5636
rect 12492 5584 12498 5636
rect 2041 5559 2099 5565
rect 2041 5525 2053 5559
rect 2087 5525 2099 5559
rect 12544 5556 12572 5723
rect 12802 5701 12808 5704
rect 12771 5695 12808 5701
rect 12771 5661 12783 5695
rect 12771 5655 12808 5661
rect 12802 5652 12808 5655
rect 12860 5652 12866 5704
rect 13722 5652 13728 5704
rect 13780 5652 13786 5704
rect 12710 5556 12716 5568
rect 12544 5528 12716 5556
rect 2041 5519 2099 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 13740 5556 13768 5652
rect 13587 5528 13768 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 1104 5466 14696 5488
rect 1104 5414 4308 5466
rect 4360 5414 4372 5466
rect 4424 5414 4436 5466
rect 4488 5414 4500 5466
rect 4552 5414 4564 5466
rect 4616 5414 7666 5466
rect 7718 5414 7730 5466
rect 7782 5414 7794 5466
rect 7846 5414 7858 5466
rect 7910 5414 7922 5466
rect 7974 5414 11024 5466
rect 11076 5414 11088 5466
rect 11140 5414 11152 5466
rect 11204 5414 11216 5466
rect 11268 5414 11280 5466
rect 11332 5414 14382 5466
rect 14434 5414 14446 5466
rect 14498 5414 14510 5466
rect 14562 5414 14574 5466
rect 14626 5414 14638 5466
rect 14690 5414 14696 5466
rect 1104 5392 14696 5414
rect 8754 5312 8760 5364
rect 8812 5352 8818 5364
rect 10321 5355 10379 5361
rect 8812 5324 10272 5352
rect 8812 5312 8818 5324
rect 1489 5287 1547 5293
rect 1489 5253 1501 5287
rect 1535 5284 1547 5287
rect 2041 5287 2099 5293
rect 2041 5284 2053 5287
rect 1535 5256 2053 5284
rect 1535 5253 1547 5256
rect 1489 5247 1547 5253
rect 2041 5253 2053 5256
rect 2087 5253 2099 5287
rect 2041 5247 2099 5253
rect 9567 5249 9625 5255
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 4706 5216 4712 5228
rect 1995 5188 4712 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 4706 5176 4712 5188
rect 4764 5176 4770 5228
rect 7006 5176 7012 5228
rect 7064 5216 7070 5228
rect 9567 5216 9579 5249
rect 7064 5215 9579 5216
rect 9613 5246 9625 5249
rect 9613 5215 9628 5246
rect 7064 5188 9628 5215
rect 10244 5216 10272 5324
rect 10321 5321 10333 5355
rect 10367 5352 10379 5355
rect 10502 5352 10508 5364
rect 10367 5324 10508 5352
rect 10367 5321 10379 5324
rect 10321 5315 10379 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 11790 5312 11796 5364
rect 11848 5352 11854 5364
rect 12529 5355 12587 5361
rect 12529 5352 12541 5355
rect 11848 5324 12541 5352
rect 11848 5312 11854 5324
rect 12529 5321 12541 5324
rect 12575 5321 12587 5355
rect 12529 5315 12587 5321
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 13909 5355 13967 5361
rect 13909 5352 13921 5355
rect 13228 5324 13921 5352
rect 13228 5312 13234 5324
rect 13909 5321 13921 5324
rect 13955 5321 13967 5355
rect 13909 5315 13967 5321
rect 11759 5229 11817 5235
rect 11759 5216 11771 5229
rect 10244 5195 11771 5216
rect 11805 5226 11817 5229
rect 11805 5195 11818 5226
rect 13139 5219 13197 5225
rect 13139 5216 13151 5219
rect 10244 5188 11818 5195
rect 12406 5188 13151 5216
rect 7064 5176 7070 5188
rect 7374 5108 7380 5160
rect 7432 5148 7438 5160
rect 8202 5148 8208 5160
rect 7432 5120 8208 5148
rect 7432 5108 7438 5120
rect 8202 5108 8208 5120
rect 8260 5148 8266 5160
rect 9309 5151 9367 5157
rect 9309 5148 9321 5151
rect 8260 5120 9321 5148
rect 8260 5108 8266 5120
rect 9309 5117 9321 5120
rect 9355 5117 9367 5151
rect 9309 5111 9367 5117
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 11517 5151 11575 5157
rect 11517 5148 11529 5151
rect 10284 5120 11529 5148
rect 10284 5108 10290 5120
rect 11517 5117 11529 5120
rect 11563 5117 11575 5151
rect 11517 5111 11575 5117
rect 8938 5040 8944 5092
rect 8996 5040 9002 5092
rect 842 4972 848 5024
rect 900 5012 906 5024
rect 1581 5015 1639 5021
rect 1581 5012 1593 5015
rect 900 4984 1593 5012
rect 900 4972 906 4984
rect 1581 4981 1593 4984
rect 1627 4981 1639 5015
rect 8956 5012 8984 5040
rect 12406 5012 12434 5188
rect 13139 5185 13151 5188
rect 13185 5185 13197 5219
rect 13139 5179 13197 5185
rect 12710 5108 12716 5160
rect 12768 5148 12774 5160
rect 12897 5151 12955 5157
rect 12897 5148 12909 5151
rect 12768 5120 12909 5148
rect 12768 5108 12774 5120
rect 12897 5117 12909 5120
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 8956 4984 12434 5012
rect 1581 4975 1639 4981
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12894 5012 12900 5024
rect 12584 4984 12900 5012
rect 12584 4972 12590 4984
rect 12894 4972 12900 4984
rect 12952 4972 12958 5024
rect 1104 4922 14536 4944
rect 1104 4870 2629 4922
rect 2681 4870 2693 4922
rect 2745 4870 2757 4922
rect 2809 4870 2821 4922
rect 2873 4870 2885 4922
rect 2937 4870 5987 4922
rect 6039 4870 6051 4922
rect 6103 4870 6115 4922
rect 6167 4870 6179 4922
rect 6231 4870 6243 4922
rect 6295 4870 9345 4922
rect 9397 4870 9409 4922
rect 9461 4870 9473 4922
rect 9525 4870 9537 4922
rect 9589 4870 9601 4922
rect 9653 4870 12703 4922
rect 12755 4870 12767 4922
rect 12819 4870 12831 4922
rect 12883 4870 12895 4922
rect 12947 4870 12959 4922
rect 13011 4870 14536 4922
rect 1104 4848 14536 4870
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5040 4780 9628 4808
rect 5040 4768 5046 4780
rect 9600 4740 9628 4780
rect 9950 4768 9956 4820
rect 10008 4768 10014 4820
rect 11238 4808 11244 4820
rect 10060 4780 11244 4808
rect 10060 4740 10088 4780
rect 11238 4768 11244 4780
rect 11296 4768 11302 4820
rect 11333 4811 11391 4817
rect 11333 4777 11345 4811
rect 11379 4808 11391 4811
rect 11422 4808 11428 4820
rect 11379 4780 11428 4808
rect 11379 4777 11391 4780
rect 11333 4771 11391 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 12437 4811 12495 4817
rect 12437 4777 12449 4811
rect 12483 4808 12495 4811
rect 12526 4808 12532 4820
rect 12483 4780 12532 4808
rect 12483 4777 12495 4780
rect 12437 4771 12495 4777
rect 12526 4768 12532 4780
rect 12584 4768 12590 4820
rect 13354 4768 13360 4820
rect 13412 4808 13418 4820
rect 13633 4811 13691 4817
rect 13633 4808 13645 4811
rect 13412 4780 13645 4808
rect 13412 4768 13418 4780
rect 13633 4777 13645 4780
rect 13679 4777 13691 4811
rect 13633 4771 13691 4777
rect 9600 4712 10088 4740
rect 8202 4632 8208 4684
rect 8260 4672 8266 4684
rect 8941 4675 8999 4681
rect 8941 4672 8953 4675
rect 8260 4644 8953 4672
rect 8260 4632 8266 4644
rect 8864 4536 8892 4644
rect 8941 4641 8953 4644
rect 8987 4641 8999 4675
rect 10226 4672 10232 4684
rect 8941 4635 8999 4641
rect 9646 4644 10232 4672
rect 9214 4604 9220 4616
rect 9175 4576 9220 4604
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 9646 4604 9674 4644
rect 10226 4632 10232 4644
rect 10284 4672 10290 4684
rect 10321 4675 10379 4681
rect 10321 4672 10333 4675
rect 10284 4644 10333 4672
rect 10284 4632 10290 4644
rect 10321 4641 10333 4644
rect 10367 4641 10379 4675
rect 10321 4635 10379 4641
rect 11330 4632 11336 4684
rect 11388 4672 11394 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 11388 4644 12173 4672
rect 11388 4632 11394 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 10594 4613 10600 4616
rect 9324 4576 9674 4604
rect 10563 4607 10600 4613
rect 9324 4536 9352 4576
rect 10563 4573 10575 4607
rect 10563 4567 10600 4573
rect 10594 4564 10600 4567
rect 10652 4564 10658 4616
rect 11974 4564 11980 4616
rect 12032 4564 12038 4616
rect 12618 4604 12624 4616
rect 12452 4576 12624 4604
rect 8864 4508 9352 4536
rect 12342 4496 12348 4548
rect 12400 4496 12406 4548
rect 9030 4428 9036 4480
rect 9088 4468 9094 4480
rect 12452 4468 12480 4576
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 13262 4604 13268 4616
rect 12910 4583 13268 4604
rect 12879 4577 13268 4583
rect 12879 4574 12891 4577
rect 12526 4496 12532 4548
rect 12584 4536 12590 4548
rect 12802 4546 12891 4574
rect 12802 4536 12830 4546
rect 12879 4543 12891 4546
rect 12925 4576 13268 4577
rect 12925 4546 12938 4576
rect 13262 4564 13268 4576
rect 13320 4564 13326 4616
rect 12925 4543 12937 4546
rect 12879 4537 12937 4543
rect 12584 4508 12830 4536
rect 12584 4496 12590 4508
rect 9088 4440 12480 4468
rect 9088 4428 9094 4440
rect 1104 4378 14696 4400
rect 1104 4326 4308 4378
rect 4360 4326 4372 4378
rect 4424 4326 4436 4378
rect 4488 4326 4500 4378
rect 4552 4326 4564 4378
rect 4616 4326 7666 4378
rect 7718 4326 7730 4378
rect 7782 4326 7794 4378
rect 7846 4326 7858 4378
rect 7910 4326 7922 4378
rect 7974 4326 11024 4378
rect 11076 4326 11088 4378
rect 11140 4326 11152 4378
rect 11204 4326 11216 4378
rect 11268 4326 11280 4378
rect 11332 4326 14382 4378
rect 14434 4326 14446 4378
rect 14498 4326 14510 4378
rect 14562 4326 14574 4378
rect 14626 4326 14638 4378
rect 14690 4326 14696 4378
rect 1104 4304 14696 4326
rect 9214 4224 9220 4276
rect 9272 4264 9278 4276
rect 12526 4264 12532 4276
rect 9272 4236 12532 4264
rect 9272 4224 9278 4236
rect 12526 4224 12532 4236
rect 12584 4224 12590 4276
rect 10318 4156 10324 4208
rect 10376 4156 10382 4208
rect 12342 4156 12348 4208
rect 12400 4156 12406 4208
rect 13081 4199 13139 4205
rect 13081 4165 13093 4199
rect 13127 4196 13139 4199
rect 13906 4196 13912 4208
rect 13127 4168 13912 4196
rect 13127 4165 13139 4168
rect 13081 4159 13139 4165
rect 13906 4156 13912 4168
rect 13964 4156 13970 4208
rect 14001 4199 14059 4205
rect 14001 4165 14013 4199
rect 14047 4196 14059 4199
rect 15286 4196 15292 4208
rect 14047 4168 15292 4196
rect 14047 4165 14059 4168
rect 14001 4159 14059 4165
rect 15286 4156 15292 4168
rect 15344 4156 15350 4208
rect 750 4088 756 4140
rect 808 4128 814 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 808 4100 1409 4128
rect 808 4088 814 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 10336 4060 10364 4156
rect 10505 4131 10563 4137
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 11698 4128 11704 4140
rect 10551 4100 11704 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 13446 4088 13452 4140
rect 13504 4088 13510 4140
rect 13630 4088 13636 4140
rect 13688 4088 13694 4140
rect 15378 4088 15384 4140
rect 15436 4088 15442 4140
rect 10781 4063 10839 4069
rect 10781 4060 10793 4063
rect 10336 4032 10793 4060
rect 10781 4029 10793 4032
rect 10827 4029 10839 4063
rect 10781 4023 10839 4029
rect 12529 4063 12587 4069
rect 12529 4029 12541 4063
rect 12575 4060 12587 4063
rect 13464 4060 13492 4088
rect 12575 4032 13492 4060
rect 13817 4063 13875 4069
rect 12575 4029 12587 4032
rect 12529 4023 12587 4029
rect 13817 4029 13829 4063
rect 13863 4060 13875 4063
rect 15396 4060 15424 4088
rect 13863 4032 15424 4060
rect 13863 4029 13875 4032
rect 13817 4023 13875 4029
rect 5074 3952 5080 4004
rect 5132 3992 5138 4004
rect 5132 3964 13216 3992
rect 5132 3952 5138 3964
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 3418 3924 3424 3936
rect 1627 3896 3424 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 13188 3933 13216 3964
rect 13173 3927 13231 3933
rect 13173 3893 13185 3927
rect 13219 3893 13231 3927
rect 13173 3887 13231 3893
rect 13814 3884 13820 3936
rect 13872 3924 13878 3936
rect 14093 3927 14151 3933
rect 14093 3924 14105 3927
rect 13872 3896 14105 3924
rect 13872 3884 13878 3896
rect 14093 3893 14105 3896
rect 14139 3893 14151 3927
rect 14093 3887 14151 3893
rect 1104 3834 14536 3856
rect 1104 3782 2629 3834
rect 2681 3782 2693 3834
rect 2745 3782 2757 3834
rect 2809 3782 2821 3834
rect 2873 3782 2885 3834
rect 2937 3782 5987 3834
rect 6039 3782 6051 3834
rect 6103 3782 6115 3834
rect 6167 3782 6179 3834
rect 6231 3782 6243 3834
rect 6295 3782 9345 3834
rect 9397 3782 9409 3834
rect 9461 3782 9473 3834
rect 9525 3782 9537 3834
rect 9589 3782 9601 3834
rect 9653 3782 12703 3834
rect 12755 3782 12767 3834
rect 12819 3782 12831 3834
rect 12883 3782 12895 3834
rect 12947 3782 12959 3834
rect 13011 3782 14536 3834
rect 1104 3760 14536 3782
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 13817 3723 13875 3729
rect 13817 3720 13829 3723
rect 8536 3692 13829 3720
rect 8536 3680 8542 3692
rect 13817 3689 13829 3692
rect 13863 3689 13875 3723
rect 13817 3683 13875 3689
rect 13722 3476 13728 3528
rect 13780 3476 13786 3528
rect 1104 3290 14696 3312
rect 1104 3238 4308 3290
rect 4360 3238 4372 3290
rect 4424 3238 4436 3290
rect 4488 3238 4500 3290
rect 4552 3238 4564 3290
rect 4616 3238 7666 3290
rect 7718 3238 7730 3290
rect 7782 3238 7794 3290
rect 7846 3238 7858 3290
rect 7910 3238 7922 3290
rect 7974 3238 11024 3290
rect 11076 3238 11088 3290
rect 11140 3238 11152 3290
rect 11204 3238 11216 3290
rect 11268 3238 11280 3290
rect 11332 3238 14382 3290
rect 14434 3238 14446 3290
rect 14498 3238 14510 3290
rect 14562 3238 14574 3290
rect 14626 3238 14638 3290
rect 14690 3238 14696 3290
rect 1104 3216 14696 3238
rect 13078 2796 13084 2848
rect 13136 2836 13142 2848
rect 13354 2836 13360 2848
rect 13136 2808 13360 2836
rect 13136 2796 13142 2808
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 1104 2746 14536 2768
rect 1104 2694 2629 2746
rect 2681 2694 2693 2746
rect 2745 2694 2757 2746
rect 2809 2694 2821 2746
rect 2873 2694 2885 2746
rect 2937 2694 5987 2746
rect 6039 2694 6051 2746
rect 6103 2694 6115 2746
rect 6167 2694 6179 2746
rect 6231 2694 6243 2746
rect 6295 2694 9345 2746
rect 9397 2694 9409 2746
rect 9461 2694 9473 2746
rect 9525 2694 9537 2746
rect 9589 2694 9601 2746
rect 9653 2694 12703 2746
rect 12755 2694 12767 2746
rect 12819 2694 12831 2746
rect 12883 2694 12895 2746
rect 12947 2694 12959 2746
rect 13011 2694 14536 2746
rect 1104 2672 14536 2694
rect 1104 2202 14696 2224
rect 1104 2150 4308 2202
rect 4360 2150 4372 2202
rect 4424 2150 4436 2202
rect 4488 2150 4500 2202
rect 4552 2150 4564 2202
rect 4616 2150 7666 2202
rect 7718 2150 7730 2202
rect 7782 2150 7794 2202
rect 7846 2150 7858 2202
rect 7910 2150 7922 2202
rect 7974 2150 11024 2202
rect 11076 2150 11088 2202
rect 11140 2150 11152 2202
rect 11204 2150 11216 2202
rect 11268 2150 11280 2202
rect 11332 2150 14382 2202
rect 14434 2150 14446 2202
rect 14498 2150 14510 2202
rect 14562 2150 14574 2202
rect 14626 2150 14638 2202
rect 14690 2150 14696 2202
rect 1104 2128 14696 2150
rect 6549 2091 6607 2097
rect 6549 2057 6561 2091
rect 6595 2088 6607 2091
rect 6638 2088 6644 2100
rect 6595 2060 6644 2088
rect 6595 2057 6607 2060
rect 6549 2051 6607 2057
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 7190 2048 7196 2100
rect 7248 2048 7254 2100
rect 7466 2048 7472 2100
rect 7524 2088 7530 2100
rect 7929 2091 7987 2097
rect 7929 2088 7941 2091
rect 7524 2060 7941 2088
rect 7524 2048 7530 2060
rect 7929 2057 7941 2060
rect 7975 2057 7987 2091
rect 7929 2051 7987 2057
rect 8662 2048 8668 2100
rect 8720 2048 8726 2100
rect 9398 2048 9404 2100
rect 9456 2048 9462 2100
rect 10134 2048 10140 2100
rect 10192 2048 10198 2100
rect 10870 2048 10876 2100
rect 10928 2048 10934 2100
rect 13446 2048 13452 2100
rect 13504 2048 13510 2100
rect 14001 2091 14059 2097
rect 14001 2057 14013 2091
rect 14047 2057 14059 2091
rect 14001 2051 14059 2057
rect 2869 2023 2927 2029
rect 2869 1989 2881 2023
rect 2915 2020 2927 2023
rect 9030 2020 9036 2032
rect 2915 1992 9036 2020
rect 2915 1989 2927 1992
rect 2869 1983 2927 1989
rect 9030 1980 9036 1992
rect 9088 1980 9094 2032
rect 13357 2023 13415 2029
rect 13357 1989 13369 2023
rect 13403 2020 13415 2023
rect 14016 2020 14044 2051
rect 13403 1992 14044 2020
rect 13403 1989 13415 1992
rect 13357 1983 13415 1989
rect 2038 1912 2044 1964
rect 2096 1912 2102 1964
rect 6454 1912 6460 1964
rect 6512 1912 6518 1964
rect 7098 1912 7104 1964
rect 7156 1912 7162 1964
rect 7834 1912 7840 1964
rect 7892 1912 7898 1964
rect 8570 1912 8576 1964
rect 8628 1912 8634 1964
rect 9214 1912 9220 1964
rect 9272 1952 9278 1964
rect 9309 1955 9367 1961
rect 9309 1952 9321 1955
rect 9272 1924 9321 1952
rect 9272 1912 9278 1924
rect 9309 1921 9321 1924
rect 9355 1921 9367 1955
rect 9309 1915 9367 1921
rect 10042 1912 10048 1964
rect 10100 1912 10106 1964
rect 10778 1912 10784 1964
rect 10836 1912 10842 1964
rect 11606 1912 11612 1964
rect 11664 1912 11670 1964
rect 12250 1912 12256 1964
rect 12308 1912 12314 1964
rect 12897 1955 12955 1961
rect 12897 1921 12909 1955
rect 12943 1952 12955 1955
rect 13078 1952 13084 1964
rect 12943 1924 13084 1952
rect 12943 1921 12955 1924
rect 12897 1915 12955 1921
rect 13078 1912 13084 1924
rect 13136 1912 13142 1964
rect 13722 1912 13728 1964
rect 13780 1912 13786 1964
rect 14182 1912 14188 1964
rect 14240 1912 14246 1964
rect 11793 1887 11851 1893
rect 11793 1853 11805 1887
rect 11839 1884 11851 1887
rect 13909 1887 13967 1893
rect 11839 1856 13676 1884
rect 11839 1853 11851 1856
rect 11793 1847 11851 1853
rect 4154 1776 4160 1828
rect 4212 1816 4218 1828
rect 13648 1816 13676 1856
rect 13909 1853 13921 1887
rect 13955 1884 13967 1887
rect 14734 1884 14740 1896
rect 13955 1856 14740 1884
rect 13955 1853 13967 1856
rect 13909 1847 13967 1853
rect 14734 1844 14740 1856
rect 14792 1844 14798 1896
rect 15562 1844 15568 1896
rect 15620 1844 15626 1896
rect 15580 1816 15608 1844
rect 4212 1788 12388 1816
rect 13648 1788 15608 1816
rect 4212 1776 4218 1788
rect 12360 1757 12388 1788
rect 12345 1751 12403 1757
rect 12345 1717 12357 1751
rect 12391 1717 12403 1751
rect 12345 1711 12403 1717
rect 12989 1751 13047 1757
rect 12989 1717 13001 1751
rect 13035 1748 13047 1751
rect 14826 1748 14832 1760
rect 13035 1720 14832 1748
rect 13035 1717 13047 1720
rect 12989 1711 13047 1717
rect 14826 1708 14832 1720
rect 14884 1708 14890 1760
rect 1104 1658 14536 1680
rect 1104 1606 2629 1658
rect 2681 1606 2693 1658
rect 2745 1606 2757 1658
rect 2809 1606 2821 1658
rect 2873 1606 2885 1658
rect 2937 1606 5987 1658
rect 6039 1606 6051 1658
rect 6103 1606 6115 1658
rect 6167 1606 6179 1658
rect 6231 1606 6243 1658
rect 6295 1606 9345 1658
rect 9397 1606 9409 1658
rect 9461 1606 9473 1658
rect 9525 1606 9537 1658
rect 9589 1606 9601 1658
rect 9653 1606 12703 1658
rect 12755 1606 12767 1658
rect 12819 1606 12831 1658
rect 12883 1606 12895 1658
rect 12947 1606 12959 1658
rect 13011 1606 14536 1658
rect 1104 1584 14536 1606
rect 5997 1547 6055 1553
rect 5997 1513 6009 1547
rect 6043 1544 6055 1547
rect 6454 1544 6460 1556
rect 6043 1516 6460 1544
rect 6043 1513 6055 1516
rect 5997 1507 6055 1513
rect 6454 1504 6460 1516
rect 6512 1504 6518 1556
rect 7098 1504 7104 1556
rect 7156 1544 7162 1556
rect 7285 1547 7343 1553
rect 7285 1544 7297 1547
rect 7156 1516 7297 1544
rect 7156 1504 7162 1516
rect 7285 1513 7297 1516
rect 7331 1513 7343 1547
rect 7285 1507 7343 1513
rect 7834 1504 7840 1556
rect 7892 1544 7898 1556
rect 7929 1547 7987 1553
rect 7929 1544 7941 1547
rect 7892 1516 7941 1544
rect 7892 1504 7898 1516
rect 7929 1513 7941 1516
rect 7975 1513 7987 1547
rect 7929 1507 7987 1513
rect 8570 1504 8576 1556
rect 8628 1544 8634 1556
rect 8941 1547 8999 1553
rect 8941 1544 8953 1547
rect 8628 1516 8953 1544
rect 8628 1504 8634 1516
rect 8941 1513 8953 1516
rect 8987 1513 8999 1547
rect 8941 1507 8999 1513
rect 9214 1504 9220 1556
rect 9272 1544 9278 1556
rect 9401 1547 9459 1553
rect 9401 1544 9413 1547
rect 9272 1516 9413 1544
rect 9272 1504 9278 1516
rect 9401 1513 9413 1516
rect 9447 1513 9459 1547
rect 9401 1507 9459 1513
rect 10042 1504 10048 1556
rect 10100 1544 10106 1556
rect 10137 1547 10195 1553
rect 10137 1544 10149 1547
rect 10100 1516 10149 1544
rect 10100 1504 10106 1516
rect 10137 1513 10149 1516
rect 10183 1513 10195 1547
rect 10137 1507 10195 1513
rect 10778 1504 10784 1556
rect 10836 1544 10842 1556
rect 10873 1547 10931 1553
rect 10873 1544 10885 1547
rect 10836 1516 10885 1544
rect 10836 1504 10842 1516
rect 10873 1513 10885 1516
rect 10919 1513 10931 1547
rect 10873 1507 10931 1513
rect 11606 1504 11612 1556
rect 11664 1504 11670 1556
rect 12250 1504 12256 1556
rect 12308 1544 12314 1556
rect 12345 1547 12403 1553
rect 12345 1544 12357 1547
rect 12308 1516 12357 1544
rect 12308 1504 12314 1516
rect 12345 1513 12357 1516
rect 12391 1513 12403 1547
rect 12345 1507 12403 1513
rect 13078 1504 13084 1556
rect 13136 1504 13142 1556
rect 13357 1547 13415 1553
rect 13357 1513 13369 1547
rect 13403 1544 13415 1547
rect 13722 1544 13728 1556
rect 13403 1516 13728 1544
rect 13403 1513 13415 1516
rect 13357 1507 13415 1513
rect 13722 1504 13728 1516
rect 13780 1504 13786 1556
rect 9122 1476 9128 1488
rect 3436 1448 9128 1476
rect 3436 1417 3464 1448
rect 9122 1436 9128 1448
rect 9180 1436 9186 1488
rect 3421 1411 3479 1417
rect 3421 1377 3433 1411
rect 3467 1377 3479 1411
rect 3421 1371 3479 1377
rect 13188 1380 13676 1408
rect 1210 1300 1216 1352
rect 1268 1340 1274 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 1268 1312 1409 1340
rect 1268 1300 1274 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 2225 1343 2283 1349
rect 2225 1309 2237 1343
rect 2271 1340 2283 1343
rect 2498 1340 2504 1352
rect 2271 1312 2504 1340
rect 2271 1309 2283 1312
rect 2225 1303 2283 1309
rect 2498 1300 2504 1312
rect 2556 1300 2562 1352
rect 2682 1300 2688 1352
rect 2740 1300 2746 1352
rect 2792 1312 3556 1340
rect 2314 1232 2320 1284
rect 2372 1272 2378 1284
rect 2792 1272 2820 1312
rect 2372 1244 2820 1272
rect 3528 1272 3556 1312
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 4614 1300 4620 1352
rect 4672 1300 4678 1352
rect 5166 1300 5172 1352
rect 5224 1340 5230 1352
rect 5261 1343 5319 1349
rect 5261 1340 5273 1343
rect 5224 1312 5273 1340
rect 5224 1300 5230 1312
rect 5261 1309 5273 1312
rect 5307 1309 5319 1343
rect 5261 1303 5319 1309
rect 6178 1300 6184 1352
rect 6236 1300 6242 1352
rect 6365 1343 6423 1349
rect 6365 1309 6377 1343
rect 6411 1309 6423 1343
rect 6365 1303 6423 1309
rect 4065 1275 4123 1281
rect 4065 1272 4077 1275
rect 3528 1244 4077 1272
rect 2372 1232 2378 1244
rect 4065 1241 4077 1244
rect 4111 1241 4123 1275
rect 4065 1235 4123 1241
rect 4154 1232 4160 1284
rect 4212 1272 4218 1284
rect 4433 1275 4491 1281
rect 4433 1272 4445 1275
rect 4212 1244 4445 1272
rect 4212 1232 4218 1244
rect 4433 1241 4445 1244
rect 4479 1241 4491 1275
rect 4433 1235 4491 1241
rect 5074 1232 5080 1284
rect 5132 1232 5138 1284
rect 5626 1232 5632 1284
rect 5684 1272 5690 1284
rect 6380 1272 6408 1303
rect 6638 1300 6644 1352
rect 6696 1300 6702 1352
rect 7098 1300 7104 1352
rect 7156 1340 7162 1352
rect 7469 1343 7527 1349
rect 7469 1340 7481 1343
rect 7156 1312 7481 1340
rect 7156 1300 7162 1312
rect 7469 1309 7481 1312
rect 7515 1309 7527 1343
rect 7469 1303 7527 1309
rect 8110 1300 8116 1352
rect 8168 1300 8174 1352
rect 8570 1300 8576 1352
rect 8628 1340 8634 1352
rect 9125 1343 9183 1349
rect 9125 1340 9137 1343
rect 8628 1312 9137 1340
rect 8628 1300 8634 1312
rect 9125 1309 9137 1312
rect 9171 1309 9183 1343
rect 9125 1303 9183 1309
rect 9306 1300 9312 1352
rect 9364 1340 9370 1352
rect 9585 1343 9643 1349
rect 9585 1340 9597 1343
rect 9364 1312 9597 1340
rect 9364 1300 9370 1312
rect 9585 1309 9597 1312
rect 9631 1309 9643 1343
rect 9585 1303 9643 1309
rect 10042 1300 10048 1352
rect 10100 1340 10106 1352
rect 10321 1343 10379 1349
rect 10321 1340 10333 1343
rect 10100 1312 10333 1340
rect 10100 1300 10106 1312
rect 10321 1309 10333 1312
rect 10367 1309 10379 1343
rect 10321 1303 10379 1309
rect 10778 1300 10784 1352
rect 10836 1340 10842 1352
rect 11057 1343 11115 1349
rect 11057 1340 11069 1343
rect 10836 1312 11069 1340
rect 10836 1300 10842 1312
rect 11057 1309 11069 1312
rect 11103 1309 11115 1343
rect 11057 1303 11115 1309
rect 11514 1300 11520 1352
rect 11572 1340 11578 1352
rect 11793 1343 11851 1349
rect 11793 1340 11805 1343
rect 11572 1312 11805 1340
rect 11572 1300 11578 1312
rect 11793 1309 11805 1312
rect 11839 1309 11851 1343
rect 11793 1303 11851 1309
rect 12250 1300 12256 1352
rect 12308 1340 12314 1352
rect 12529 1343 12587 1349
rect 12529 1340 12541 1343
rect 12308 1312 12541 1340
rect 12308 1300 12314 1312
rect 12529 1309 12541 1312
rect 12575 1309 12587 1343
rect 12529 1303 12587 1309
rect 12989 1343 13047 1349
rect 12989 1309 13001 1343
rect 13035 1340 13047 1343
rect 13188 1340 13216 1380
rect 13035 1312 13216 1340
rect 13035 1309 13047 1312
rect 12989 1303 13047 1309
rect 13262 1300 13268 1352
rect 13320 1300 13326 1352
rect 13538 1300 13544 1352
rect 13596 1300 13602 1352
rect 13648 1340 13676 1380
rect 15194 1340 15200 1352
rect 13648 1312 15200 1340
rect 15194 1300 15200 1312
rect 15252 1300 15258 1352
rect 13725 1275 13783 1281
rect 13725 1272 13737 1275
rect 5684 1244 6408 1272
rect 12820 1244 13737 1272
rect 5684 1232 5690 1244
rect 12820 1213 12848 1244
rect 13725 1241 13737 1244
rect 13771 1241 13783 1275
rect 13725 1235 13783 1241
rect 12805 1207 12863 1213
rect 12805 1173 12817 1207
rect 12851 1173 12863 1207
rect 12805 1167 12863 1173
rect 13814 1164 13820 1216
rect 13872 1164 13878 1216
rect 1104 1114 14696 1136
rect 1104 1062 4308 1114
rect 4360 1062 4372 1114
rect 4424 1062 4436 1114
rect 4488 1062 4500 1114
rect 4552 1062 4564 1114
rect 4616 1062 7666 1114
rect 7718 1062 7730 1114
rect 7782 1062 7794 1114
rect 7846 1062 7858 1114
rect 7910 1062 7922 1114
rect 7974 1062 11024 1114
rect 11076 1062 11088 1114
rect 11140 1062 11152 1114
rect 11204 1062 11216 1114
rect 11268 1062 11280 1114
rect 11332 1062 14382 1114
rect 14434 1062 14446 1114
rect 14498 1062 14510 1114
rect 14562 1062 14574 1114
rect 14626 1062 14638 1114
rect 14690 1062 14696 1114
rect 1104 1040 14696 1062
<< via1 >>
rect 4308 43494 4360 43546
rect 4372 43494 4424 43546
rect 4436 43494 4488 43546
rect 4500 43494 4552 43546
rect 4564 43494 4616 43546
rect 7666 43494 7718 43546
rect 7730 43494 7782 43546
rect 7794 43494 7846 43546
rect 7858 43494 7910 43546
rect 7922 43494 7974 43546
rect 11024 43494 11076 43546
rect 11088 43494 11140 43546
rect 11152 43494 11204 43546
rect 11216 43494 11268 43546
rect 11280 43494 11332 43546
rect 14382 43494 14434 43546
rect 14446 43494 14498 43546
rect 14510 43494 14562 43546
rect 14574 43494 14626 43546
rect 14638 43494 14690 43546
rect 480 43392 532 43444
rect 3424 43392 3476 43444
rect 4160 43392 4212 43444
rect 4896 43392 4948 43444
rect 5632 43392 5684 43444
rect 6368 43392 6420 43444
rect 7104 43392 7156 43444
rect 8024 43392 8076 43444
rect 8576 43392 8628 43444
rect 9312 43392 9364 43444
rect 10048 43392 10100 43444
rect 10784 43392 10836 43444
rect 11520 43392 11572 43444
rect 12256 43392 12308 43444
rect 12992 43392 13044 43444
rect 15200 43392 15252 43444
rect 1768 43256 1820 43308
rect 2044 43299 2096 43308
rect 2044 43265 2053 43299
rect 2053 43265 2087 43299
rect 2087 43265 2096 43299
rect 2044 43256 2096 43265
rect 3056 43256 3108 43308
rect 3148 43299 3200 43308
rect 3148 43265 3157 43299
rect 3157 43265 3191 43299
rect 3191 43265 3200 43299
rect 3148 43256 3200 43265
rect 3792 43299 3844 43308
rect 3792 43265 3801 43299
rect 3801 43265 3835 43299
rect 3835 43265 3844 43299
rect 3792 43256 3844 43265
rect 4344 43299 4396 43308
rect 4344 43265 4353 43299
rect 4353 43265 4387 43299
rect 4387 43265 4396 43299
rect 4344 43256 4396 43265
rect 4988 43299 5040 43308
rect 4988 43265 4997 43299
rect 4997 43265 5031 43299
rect 5031 43265 5040 43299
rect 4988 43256 5040 43265
rect 5724 43299 5776 43308
rect 5724 43265 5733 43299
rect 5733 43265 5767 43299
rect 5767 43265 5776 43299
rect 5724 43256 5776 43265
rect 6460 43299 6512 43308
rect 6460 43265 6469 43299
rect 6469 43265 6503 43299
rect 6503 43265 6512 43299
rect 6460 43256 6512 43265
rect 7196 43299 7248 43308
rect 7196 43265 7205 43299
rect 7205 43265 7239 43299
rect 7239 43265 7248 43299
rect 7196 43256 7248 43265
rect 7932 43299 7984 43308
rect 7932 43265 7941 43299
rect 7941 43265 7975 43299
rect 7975 43265 7984 43299
rect 7932 43256 7984 43265
rect 8944 43299 8996 43308
rect 8944 43265 8953 43299
rect 8953 43265 8987 43299
rect 8987 43265 8996 43299
rect 8944 43256 8996 43265
rect 9220 43256 9272 43308
rect 10140 43299 10192 43308
rect 10140 43265 10149 43299
rect 10149 43265 10183 43299
rect 10183 43265 10192 43299
rect 10140 43256 10192 43265
rect 10968 43299 11020 43308
rect 10968 43265 10977 43299
rect 10977 43265 11011 43299
rect 11011 43265 11020 43299
rect 10968 43256 11020 43265
rect 11612 43299 11664 43308
rect 11612 43265 11621 43299
rect 11621 43265 11655 43299
rect 11655 43265 11664 43299
rect 11612 43256 11664 43265
rect 12440 43299 12492 43308
rect 12440 43265 12449 43299
rect 12449 43265 12483 43299
rect 12483 43265 12492 43299
rect 12440 43256 12492 43265
rect 13084 43299 13136 43308
rect 13084 43265 13093 43299
rect 13093 43265 13127 43299
rect 13127 43265 13136 43299
rect 13084 43256 13136 43265
rect 13544 43299 13596 43308
rect 13544 43265 13553 43299
rect 13553 43265 13587 43299
rect 13587 43265 13596 43299
rect 13544 43256 13596 43265
rect 1952 43120 2004 43172
rect 1400 43052 1452 43104
rect 2780 43095 2832 43104
rect 2780 43061 2789 43095
rect 2789 43061 2823 43095
rect 2823 43061 2832 43095
rect 2780 43052 2832 43061
rect 2629 42950 2681 43002
rect 2693 42950 2745 43002
rect 2757 42950 2809 43002
rect 2821 42950 2873 43002
rect 2885 42950 2937 43002
rect 5987 42950 6039 43002
rect 6051 42950 6103 43002
rect 6115 42950 6167 43002
rect 6179 42950 6231 43002
rect 6243 42950 6295 43002
rect 9345 42950 9397 43002
rect 9409 42950 9461 43002
rect 9473 42950 9525 43002
rect 9537 42950 9589 43002
rect 9601 42950 9653 43002
rect 12703 42950 12755 43002
rect 12767 42950 12819 43002
rect 12831 42950 12883 43002
rect 12895 42950 12947 43002
rect 12959 42950 13011 43002
rect 3148 42848 3200 42900
rect 3792 42848 3844 42900
rect 4344 42848 4396 42900
rect 4988 42848 5040 42900
rect 6460 42848 6512 42900
rect 7196 42848 7248 42900
rect 7932 42848 7984 42900
rect 8944 42848 8996 42900
rect 9220 42891 9272 42900
rect 9220 42857 9229 42891
rect 9229 42857 9263 42891
rect 9263 42857 9272 42891
rect 9220 42848 9272 42857
rect 10140 42848 10192 42900
rect 10968 42848 11020 42900
rect 11612 42848 11664 42900
rect 12440 42848 12492 42900
rect 13084 42848 13136 42900
rect 14280 42712 14332 42764
rect 3424 42687 3476 42696
rect 3424 42653 3433 42687
rect 3433 42653 3467 42687
rect 3467 42653 3476 42687
rect 3424 42644 3476 42653
rect 4068 42644 4120 42696
rect 4988 42687 5040 42696
rect 4988 42653 4997 42687
rect 4997 42653 5031 42687
rect 5031 42653 5040 42687
rect 4988 42644 5040 42653
rect 6460 42687 6512 42696
rect 6460 42653 6469 42687
rect 6469 42653 6503 42687
rect 6503 42653 6512 42687
rect 6460 42644 6512 42653
rect 7196 42687 7248 42696
rect 7196 42653 7205 42687
rect 7205 42653 7239 42687
rect 7239 42653 7248 42687
rect 7196 42644 7248 42653
rect 7932 42687 7984 42696
rect 7932 42653 7941 42687
rect 7941 42653 7975 42687
rect 7975 42653 7984 42687
rect 7932 42644 7984 42653
rect 8668 42687 8720 42696
rect 8668 42653 8677 42687
rect 8677 42653 8711 42687
rect 8711 42653 8720 42687
rect 8668 42644 8720 42653
rect 1400 42619 1452 42628
rect 1400 42585 1409 42619
rect 1409 42585 1443 42619
rect 1443 42585 1452 42619
rect 1400 42576 1452 42585
rect 3608 42576 3660 42628
rect 10048 42687 10100 42696
rect 10048 42653 10057 42687
rect 10057 42653 10091 42687
rect 10091 42653 10100 42687
rect 10048 42644 10100 42653
rect 10324 42551 10376 42560
rect 10324 42517 10333 42551
rect 10333 42517 10367 42551
rect 10367 42517 10376 42551
rect 10324 42508 10376 42517
rect 12348 42687 12400 42696
rect 12348 42653 12357 42687
rect 12357 42653 12391 42687
rect 12391 42653 12400 42687
rect 12348 42644 12400 42653
rect 13820 42687 13872 42696
rect 13820 42653 13829 42687
rect 13829 42653 13863 42687
rect 13863 42653 13872 42687
rect 13820 42644 13872 42653
rect 13176 42619 13228 42628
rect 13176 42585 13185 42619
rect 13185 42585 13219 42619
rect 13219 42585 13228 42619
rect 13176 42576 13228 42585
rect 15568 42508 15620 42560
rect 4308 42406 4360 42458
rect 4372 42406 4424 42458
rect 4436 42406 4488 42458
rect 4500 42406 4552 42458
rect 4564 42406 4616 42458
rect 7666 42406 7718 42458
rect 7730 42406 7782 42458
rect 7794 42406 7846 42458
rect 7858 42406 7910 42458
rect 7922 42406 7974 42458
rect 11024 42406 11076 42458
rect 11088 42406 11140 42458
rect 11152 42406 11204 42458
rect 11216 42406 11268 42458
rect 11280 42406 11332 42458
rect 14382 42406 14434 42458
rect 14446 42406 14498 42458
rect 14510 42406 14562 42458
rect 14574 42406 14626 42458
rect 14638 42406 14690 42458
rect 2044 42304 2096 42356
rect 4068 42347 4120 42356
rect 4068 42313 4077 42347
rect 4077 42313 4111 42347
rect 4111 42313 4120 42347
rect 4068 42304 4120 42313
rect 4988 42304 5040 42356
rect 5632 42304 5684 42356
rect 12348 42304 12400 42356
rect 13544 42304 13596 42356
rect 13728 42304 13780 42356
rect 3976 42236 4028 42288
rect 10324 42236 10376 42288
rect 2136 42211 2188 42220
rect 2136 42177 2145 42211
rect 2145 42177 2179 42211
rect 2179 42177 2188 42211
rect 2136 42168 2188 42177
rect 4252 42211 4304 42220
rect 4252 42177 4261 42211
rect 4261 42177 4295 42211
rect 4295 42177 4304 42211
rect 4252 42168 4304 42177
rect 4896 42211 4948 42220
rect 4896 42177 4905 42211
rect 4905 42177 4939 42211
rect 4939 42177 4948 42211
rect 4896 42168 4948 42177
rect 13728 42211 13780 42220
rect 13728 42177 13737 42211
rect 13737 42177 13771 42211
rect 13771 42177 13780 42211
rect 13728 42168 13780 42177
rect 15476 42032 15528 42084
rect 2629 41862 2681 41914
rect 2693 41862 2745 41914
rect 2757 41862 2809 41914
rect 2821 41862 2873 41914
rect 2885 41862 2937 41914
rect 5987 41862 6039 41914
rect 6051 41862 6103 41914
rect 6115 41862 6167 41914
rect 6179 41862 6231 41914
rect 6243 41862 6295 41914
rect 9345 41862 9397 41914
rect 9409 41862 9461 41914
rect 9473 41862 9525 41914
rect 9537 41862 9589 41914
rect 9601 41862 9653 41914
rect 12703 41862 12755 41914
rect 12767 41862 12819 41914
rect 12831 41862 12883 41914
rect 12895 41862 12947 41914
rect 12959 41862 13011 41914
rect 13176 41760 13228 41812
rect 13728 41760 13780 41812
rect 14740 41556 14792 41608
rect 14004 41488 14056 41540
rect 4308 41318 4360 41370
rect 4372 41318 4424 41370
rect 4436 41318 4488 41370
rect 4500 41318 4552 41370
rect 4564 41318 4616 41370
rect 7666 41318 7718 41370
rect 7730 41318 7782 41370
rect 7794 41318 7846 41370
rect 7858 41318 7910 41370
rect 7922 41318 7974 41370
rect 11024 41318 11076 41370
rect 11088 41318 11140 41370
rect 11152 41318 11204 41370
rect 11216 41318 11268 41370
rect 11280 41318 11332 41370
rect 14382 41318 14434 41370
rect 14446 41318 14498 41370
rect 14510 41318 14562 41370
rect 14574 41318 14626 41370
rect 14638 41318 14690 41370
rect 756 41080 808 41132
rect 6368 40876 6420 40928
rect 2629 40774 2681 40826
rect 2693 40774 2745 40826
rect 2757 40774 2809 40826
rect 2821 40774 2873 40826
rect 2885 40774 2937 40826
rect 5987 40774 6039 40826
rect 6051 40774 6103 40826
rect 6115 40774 6167 40826
rect 6179 40774 6231 40826
rect 6243 40774 6295 40826
rect 9345 40774 9397 40826
rect 9409 40774 9461 40826
rect 9473 40774 9525 40826
rect 9537 40774 9589 40826
rect 9601 40774 9653 40826
rect 12703 40774 12755 40826
rect 12767 40774 12819 40826
rect 12831 40774 12883 40826
rect 12895 40774 12947 40826
rect 12959 40774 13011 40826
rect 4308 40230 4360 40282
rect 4372 40230 4424 40282
rect 4436 40230 4488 40282
rect 4500 40230 4552 40282
rect 4564 40230 4616 40282
rect 7666 40230 7718 40282
rect 7730 40230 7782 40282
rect 7794 40230 7846 40282
rect 7858 40230 7910 40282
rect 7922 40230 7974 40282
rect 11024 40230 11076 40282
rect 11088 40230 11140 40282
rect 11152 40230 11204 40282
rect 11216 40230 11268 40282
rect 11280 40230 11332 40282
rect 14382 40230 14434 40282
rect 14446 40230 14498 40282
rect 14510 40230 14562 40282
rect 14574 40230 14626 40282
rect 14638 40230 14690 40282
rect 1492 40103 1544 40112
rect 1492 40069 1501 40103
rect 1501 40069 1535 40103
rect 1535 40069 1544 40103
rect 1492 40060 1544 40069
rect 7472 39992 7524 40044
rect 13820 40035 13872 40044
rect 13820 40001 13829 40035
rect 13829 40001 13863 40035
rect 13863 40001 13872 40035
rect 13820 39992 13872 40001
rect 4712 39856 4764 39908
rect 13268 39831 13320 39840
rect 13268 39797 13277 39831
rect 13277 39797 13311 39831
rect 13311 39797 13320 39831
rect 13268 39788 13320 39797
rect 14096 39831 14148 39840
rect 14096 39797 14105 39831
rect 14105 39797 14139 39831
rect 14139 39797 14148 39831
rect 14096 39788 14148 39797
rect 2629 39686 2681 39738
rect 2693 39686 2745 39738
rect 2757 39686 2809 39738
rect 2821 39686 2873 39738
rect 2885 39686 2937 39738
rect 5987 39686 6039 39738
rect 6051 39686 6103 39738
rect 6115 39686 6167 39738
rect 6179 39686 6231 39738
rect 6243 39686 6295 39738
rect 9345 39686 9397 39738
rect 9409 39686 9461 39738
rect 9473 39686 9525 39738
rect 9537 39686 9589 39738
rect 9601 39686 9653 39738
rect 12703 39686 12755 39738
rect 12767 39686 12819 39738
rect 12831 39686 12883 39738
rect 12895 39686 12947 39738
rect 12959 39686 13011 39738
rect 6368 39584 6420 39636
rect 6736 39584 6788 39636
rect 4712 39380 4764 39432
rect 13820 39584 13872 39636
rect 12900 39423 12952 39432
rect 12900 39389 12909 39423
rect 12909 39389 12943 39423
rect 12943 39389 12952 39423
rect 12900 39380 12952 39389
rect 756 39312 808 39364
rect 7472 39312 7524 39364
rect 14832 39312 14884 39364
rect 14280 39244 14332 39296
rect 4308 39142 4360 39194
rect 4372 39142 4424 39194
rect 4436 39142 4488 39194
rect 4500 39142 4552 39194
rect 4564 39142 4616 39194
rect 7666 39142 7718 39194
rect 7730 39142 7782 39194
rect 7794 39142 7846 39194
rect 7858 39142 7910 39194
rect 7922 39142 7974 39194
rect 11024 39142 11076 39194
rect 11088 39142 11140 39194
rect 11152 39142 11204 39194
rect 11216 39142 11268 39194
rect 11280 39142 11332 39194
rect 14382 39142 14434 39194
rect 14446 39142 14498 39194
rect 14510 39142 14562 39194
rect 14574 39142 14626 39194
rect 14638 39142 14690 39194
rect 12900 39040 12952 39092
rect 13268 39040 13320 39092
rect 12256 38836 12308 38888
rect 12440 38768 12492 38820
rect 13636 38947 13688 38956
rect 13636 38913 13645 38947
rect 13645 38913 13679 38947
rect 13679 38913 13688 38947
rect 13636 38904 13688 38913
rect 13084 38700 13136 38752
rect 13360 38743 13412 38752
rect 13360 38709 13369 38743
rect 13369 38709 13403 38743
rect 13403 38709 13412 38743
rect 13360 38700 13412 38709
rect 13912 38743 13964 38752
rect 13912 38709 13921 38743
rect 13921 38709 13955 38743
rect 13955 38709 13964 38743
rect 13912 38700 13964 38709
rect 2629 38598 2681 38650
rect 2693 38598 2745 38650
rect 2757 38598 2809 38650
rect 2821 38598 2873 38650
rect 2885 38598 2937 38650
rect 5987 38598 6039 38650
rect 6051 38598 6103 38650
rect 6115 38598 6167 38650
rect 6179 38598 6231 38650
rect 6243 38598 6295 38650
rect 9345 38598 9397 38650
rect 9409 38598 9461 38650
rect 9473 38598 9525 38650
rect 9537 38598 9589 38650
rect 9601 38598 9653 38650
rect 12703 38598 12755 38650
rect 12767 38598 12819 38650
rect 12831 38598 12883 38650
rect 12895 38598 12947 38650
rect 12959 38598 13011 38650
rect 13636 38496 13688 38548
rect 12164 38428 12216 38480
rect 13452 38428 13504 38480
rect 756 38292 808 38344
rect 11796 38292 11848 38344
rect 12624 38292 12676 38344
rect 11888 38224 11940 38276
rect 13360 38267 13412 38276
rect 13360 38233 13369 38267
rect 13369 38233 13403 38267
rect 13403 38233 13412 38267
rect 13360 38224 13412 38233
rect 14832 38224 14884 38276
rect 12624 38199 12676 38208
rect 12624 38165 12633 38199
rect 12633 38165 12667 38199
rect 12667 38165 12676 38199
rect 12624 38156 12676 38165
rect 14280 38156 14332 38208
rect 4308 38054 4360 38106
rect 4372 38054 4424 38106
rect 4436 38054 4488 38106
rect 4500 38054 4552 38106
rect 4564 38054 4616 38106
rect 7666 38054 7718 38106
rect 7730 38054 7782 38106
rect 7794 38054 7846 38106
rect 7858 38054 7910 38106
rect 7922 38054 7974 38106
rect 11024 38054 11076 38106
rect 11088 38054 11140 38106
rect 11152 38054 11204 38106
rect 11216 38054 11268 38106
rect 11280 38054 11332 38106
rect 14382 38054 14434 38106
rect 14446 38054 14498 38106
rect 14510 38054 14562 38106
rect 14574 38054 14626 38106
rect 14638 38054 14690 38106
rect 11888 37995 11940 38004
rect 11888 37961 11897 37995
rect 11897 37961 11931 37995
rect 11931 37961 11940 37995
rect 11888 37952 11940 37961
rect 12348 37952 12400 38004
rect 12624 37952 12676 38004
rect 13360 37952 13412 38004
rect 13452 37952 13504 38004
rect 756 37816 808 37868
rect 10324 37816 10376 37868
rect 10416 37748 10468 37800
rect 12624 37859 12676 37868
rect 12624 37825 12633 37859
rect 12633 37825 12667 37859
rect 12667 37825 12676 37859
rect 12624 37816 12676 37825
rect 13084 37884 13136 37936
rect 14372 37748 14424 37800
rect 14188 37680 14240 37732
rect 13728 37612 13780 37664
rect 2629 37510 2681 37562
rect 2693 37510 2745 37562
rect 2757 37510 2809 37562
rect 2821 37510 2873 37562
rect 2885 37510 2937 37562
rect 5987 37510 6039 37562
rect 6051 37510 6103 37562
rect 6115 37510 6167 37562
rect 6179 37510 6231 37562
rect 6243 37510 6295 37562
rect 9345 37510 9397 37562
rect 9409 37510 9461 37562
rect 9473 37510 9525 37562
rect 9537 37510 9589 37562
rect 9601 37510 9653 37562
rect 12703 37510 12755 37562
rect 12767 37510 12819 37562
rect 12831 37510 12883 37562
rect 12895 37510 12947 37562
rect 12959 37510 13011 37562
rect 10324 37451 10376 37460
rect 10324 37417 10333 37451
rect 10333 37417 10367 37451
rect 10367 37417 10376 37451
rect 10324 37408 10376 37417
rect 10508 37408 10560 37460
rect 12624 37408 12676 37460
rect 12256 37383 12308 37392
rect 12256 37349 12265 37383
rect 12265 37349 12299 37383
rect 12299 37349 12308 37383
rect 12256 37340 12308 37349
rect 12348 37272 12400 37324
rect 8300 37204 8352 37256
rect 11888 37247 11940 37256
rect 11888 37213 11897 37247
rect 11897 37213 11931 37247
rect 11931 37213 11940 37247
rect 11888 37204 11940 37213
rect 12624 37204 12676 37256
rect 12716 37247 12768 37256
rect 12716 37213 12725 37247
rect 12725 37213 12759 37247
rect 12759 37213 12768 37247
rect 12716 37204 12768 37213
rect 1584 37136 1636 37188
rect 13360 37179 13412 37188
rect 13360 37145 13369 37179
rect 13369 37145 13403 37179
rect 13403 37145 13412 37179
rect 13360 37136 13412 37145
rect 13544 37179 13596 37188
rect 13544 37145 13553 37179
rect 13553 37145 13587 37179
rect 13587 37145 13596 37179
rect 13544 37136 13596 37145
rect 11704 37111 11756 37120
rect 11704 37077 11713 37111
rect 11713 37077 11747 37111
rect 11747 37077 11756 37111
rect 11704 37068 11756 37077
rect 11980 37111 12032 37120
rect 11980 37077 11989 37111
rect 11989 37077 12023 37111
rect 12023 37077 12032 37111
rect 11980 37068 12032 37077
rect 12072 37068 12124 37120
rect 13636 37111 13688 37120
rect 13636 37077 13645 37111
rect 13645 37077 13679 37111
rect 13679 37077 13688 37111
rect 13636 37068 13688 37077
rect 4308 36966 4360 37018
rect 4372 36966 4424 37018
rect 4436 36966 4488 37018
rect 4500 36966 4552 37018
rect 4564 36966 4616 37018
rect 7666 36966 7718 37018
rect 7730 36966 7782 37018
rect 7794 36966 7846 37018
rect 7858 36966 7910 37018
rect 7922 36966 7974 37018
rect 11024 36966 11076 37018
rect 11088 36966 11140 37018
rect 11152 36966 11204 37018
rect 11216 36966 11268 37018
rect 11280 36966 11332 37018
rect 14382 36966 14434 37018
rect 14446 36966 14498 37018
rect 14510 36966 14562 37018
rect 14574 36966 14626 37018
rect 14638 36966 14690 37018
rect 8300 36864 8352 36916
rect 13544 36864 13596 36916
rect 10600 36796 10652 36848
rect 756 36728 808 36780
rect 1952 36771 2004 36780
rect 1952 36737 1961 36771
rect 1961 36737 1995 36771
rect 1995 36737 2004 36771
rect 1952 36728 2004 36737
rect 9772 36728 9824 36780
rect 11980 36728 12032 36780
rect 12440 36771 12492 36780
rect 12440 36737 12449 36771
rect 12449 36737 12483 36771
rect 12483 36737 12492 36771
rect 12440 36728 12492 36737
rect 12532 36728 12584 36780
rect 10232 36660 10284 36712
rect 15016 36728 15068 36780
rect 1768 36635 1820 36644
rect 1768 36601 1777 36635
rect 1777 36601 1811 36635
rect 1811 36601 1820 36635
rect 1768 36592 1820 36601
rect 12808 36592 12860 36644
rect 12164 36524 12216 36576
rect 14188 36592 14240 36644
rect 13544 36524 13596 36576
rect 2629 36422 2681 36474
rect 2693 36422 2745 36474
rect 2757 36422 2809 36474
rect 2821 36422 2873 36474
rect 2885 36422 2937 36474
rect 5987 36422 6039 36474
rect 6051 36422 6103 36474
rect 6115 36422 6167 36474
rect 6179 36422 6231 36474
rect 6243 36422 6295 36474
rect 9345 36422 9397 36474
rect 9409 36422 9461 36474
rect 9473 36422 9525 36474
rect 9537 36422 9589 36474
rect 9601 36422 9653 36474
rect 12703 36422 12755 36474
rect 12767 36422 12819 36474
rect 12831 36422 12883 36474
rect 12895 36422 12947 36474
rect 12959 36422 13011 36474
rect 1952 36363 2004 36372
rect 1952 36329 1961 36363
rect 1961 36329 1995 36363
rect 1995 36329 2004 36363
rect 1952 36320 2004 36329
rect 3700 36320 3752 36372
rect 10508 36320 10560 36372
rect 12440 36320 12492 36372
rect 10508 36184 10560 36236
rect 7380 36116 7432 36168
rect 10876 36116 10928 36168
rect 1492 36091 1544 36100
rect 1492 36057 1501 36091
rect 1501 36057 1535 36091
rect 1535 36057 1544 36091
rect 1492 36048 1544 36057
rect 12256 36091 12308 36100
rect 12256 36057 12265 36091
rect 12265 36057 12299 36091
rect 12299 36057 12308 36091
rect 12256 36048 12308 36057
rect 12624 36091 12676 36100
rect 12624 36057 12633 36091
rect 12633 36057 12667 36091
rect 12667 36057 12676 36091
rect 12624 36048 12676 36057
rect 13176 36091 13228 36100
rect 13176 36057 13185 36091
rect 13185 36057 13219 36091
rect 13219 36057 13228 36091
rect 13176 36048 13228 36057
rect 13360 36091 13412 36100
rect 13360 36057 13369 36091
rect 13369 36057 13403 36091
rect 13403 36057 13412 36091
rect 13360 36048 13412 36057
rect 13728 36091 13780 36100
rect 13728 36057 13737 36091
rect 13737 36057 13771 36091
rect 13771 36057 13780 36091
rect 13728 36048 13780 36057
rect 11796 35980 11848 36032
rect 11888 35980 11940 36032
rect 4308 35878 4360 35930
rect 4372 35878 4424 35930
rect 4436 35878 4488 35930
rect 4500 35878 4552 35930
rect 4564 35878 4616 35930
rect 7666 35878 7718 35930
rect 7730 35878 7782 35930
rect 7794 35878 7846 35930
rect 7858 35878 7910 35930
rect 7922 35878 7974 35930
rect 11024 35878 11076 35930
rect 11088 35878 11140 35930
rect 11152 35878 11204 35930
rect 11216 35878 11268 35930
rect 11280 35878 11332 35930
rect 14382 35878 14434 35930
rect 14446 35878 14498 35930
rect 14510 35878 14562 35930
rect 14574 35878 14626 35930
rect 14638 35878 14690 35930
rect 10232 35819 10284 35828
rect 10232 35785 10241 35819
rect 10241 35785 10275 35819
rect 10275 35785 10284 35819
rect 10232 35776 10284 35785
rect 10600 35819 10652 35828
rect 10600 35785 10609 35819
rect 10609 35785 10643 35819
rect 10643 35785 10652 35819
rect 10600 35776 10652 35785
rect 10876 35819 10928 35828
rect 10876 35785 10885 35819
rect 10885 35785 10919 35819
rect 10919 35785 10928 35819
rect 10876 35776 10928 35785
rect 11244 35776 11296 35828
rect 11428 35776 11480 35828
rect 12164 35776 12216 35828
rect 8944 35640 8996 35692
rect 10416 35683 10468 35692
rect 10416 35649 10425 35683
rect 10425 35649 10459 35683
rect 10459 35649 10468 35683
rect 10416 35640 10468 35649
rect 11704 35708 11756 35760
rect 11428 35640 11480 35692
rect 11796 35683 11848 35692
rect 11796 35649 11805 35683
rect 11805 35649 11839 35683
rect 11839 35649 11848 35683
rect 11796 35640 11848 35649
rect 12072 35683 12124 35692
rect 12072 35649 12081 35683
rect 12081 35649 12115 35683
rect 12115 35649 12124 35683
rect 12072 35640 12124 35649
rect 12348 35708 12400 35760
rect 10968 35572 11020 35624
rect 12440 35640 12492 35692
rect 12532 35640 12584 35692
rect 13820 35640 13872 35692
rect 14096 35683 14148 35692
rect 14096 35649 14105 35683
rect 14105 35649 14139 35683
rect 14139 35649 14148 35683
rect 14096 35640 14148 35649
rect 12256 35572 12308 35624
rect 11520 35504 11572 35556
rect 14004 35504 14056 35556
rect 10876 35436 10928 35488
rect 13268 35436 13320 35488
rect 13452 35479 13504 35488
rect 13452 35445 13461 35479
rect 13461 35445 13495 35479
rect 13495 35445 13504 35479
rect 13452 35436 13504 35445
rect 2629 35334 2681 35386
rect 2693 35334 2745 35386
rect 2757 35334 2809 35386
rect 2821 35334 2873 35386
rect 2885 35334 2937 35386
rect 5987 35334 6039 35386
rect 6051 35334 6103 35386
rect 6115 35334 6167 35386
rect 6179 35334 6231 35386
rect 6243 35334 6295 35386
rect 9345 35334 9397 35386
rect 9409 35334 9461 35386
rect 9473 35334 9525 35386
rect 9537 35334 9589 35386
rect 9601 35334 9653 35386
rect 12703 35334 12755 35386
rect 12767 35334 12819 35386
rect 12831 35334 12883 35386
rect 12895 35334 12947 35386
rect 12959 35334 13011 35386
rect 5540 35275 5592 35284
rect 5540 35241 5549 35275
rect 5549 35241 5583 35275
rect 5583 35241 5592 35275
rect 5540 35232 5592 35241
rect 8944 35275 8996 35284
rect 8944 35241 8953 35275
rect 8953 35241 8987 35275
rect 8987 35241 8996 35275
rect 8944 35232 8996 35241
rect 10416 35232 10468 35284
rect 10968 35232 11020 35284
rect 13360 35232 13412 35284
rect 9864 35164 9916 35216
rect 11244 35164 11296 35216
rect 756 35028 808 35080
rect 5724 35071 5776 35080
rect 5724 35037 5733 35071
rect 5733 35037 5767 35071
rect 5767 35037 5776 35071
rect 5724 35028 5776 35037
rect 8116 35028 8168 35080
rect 9680 35071 9732 35080
rect 9680 35037 9689 35071
rect 9689 35037 9723 35071
rect 9723 35037 9732 35071
rect 9680 35028 9732 35037
rect 10600 35028 10652 35080
rect 10416 34960 10468 35012
rect 11520 35071 11572 35080
rect 11520 35037 11529 35071
rect 11529 35037 11563 35071
rect 11563 35037 11572 35071
rect 11520 35028 11572 35037
rect 13084 35071 13136 35080
rect 13084 35037 13093 35071
rect 13093 35037 13127 35071
rect 13127 35037 13136 35071
rect 13084 35028 13136 35037
rect 6460 34892 6512 34944
rect 13176 34960 13228 35012
rect 11888 34892 11940 34944
rect 12440 34892 12492 34944
rect 12624 34892 12676 34944
rect 13636 34935 13688 34944
rect 13636 34901 13645 34935
rect 13645 34901 13679 34935
rect 13679 34901 13688 34935
rect 13636 34892 13688 34901
rect 4308 34790 4360 34842
rect 4372 34790 4424 34842
rect 4436 34790 4488 34842
rect 4500 34790 4552 34842
rect 4564 34790 4616 34842
rect 7666 34790 7718 34842
rect 7730 34790 7782 34842
rect 7794 34790 7846 34842
rect 7858 34790 7910 34842
rect 7922 34790 7974 34842
rect 11024 34790 11076 34842
rect 11088 34790 11140 34842
rect 11152 34790 11204 34842
rect 11216 34790 11268 34842
rect 11280 34790 11332 34842
rect 14382 34790 14434 34842
rect 14446 34790 14498 34842
rect 14510 34790 14562 34842
rect 14574 34790 14626 34842
rect 14638 34790 14690 34842
rect 5724 34688 5776 34740
rect 10600 34731 10652 34740
rect 10600 34697 10609 34731
rect 10609 34697 10643 34731
rect 10643 34697 10652 34731
rect 10600 34688 10652 34697
rect 12992 34688 13044 34740
rect 13820 34688 13872 34740
rect 5356 34620 5408 34672
rect 9772 34620 9824 34672
rect 11244 34620 11296 34672
rect 1400 34595 1452 34604
rect 1400 34561 1409 34595
rect 1409 34561 1443 34595
rect 1443 34561 1452 34595
rect 1400 34552 1452 34561
rect 5724 34595 5776 34604
rect 5724 34561 5733 34595
rect 5733 34561 5767 34595
rect 5767 34561 5776 34595
rect 5724 34552 5776 34561
rect 8208 34552 8260 34604
rect 10968 34595 11020 34604
rect 10968 34561 10977 34595
rect 10977 34561 11011 34595
rect 11011 34561 11020 34595
rect 10968 34552 11020 34561
rect 11336 34595 11388 34604
rect 11336 34561 11345 34595
rect 11345 34561 11379 34595
rect 11379 34561 11388 34595
rect 11336 34552 11388 34561
rect 11428 34552 11480 34604
rect 13820 34595 13872 34604
rect 13820 34561 13829 34595
rect 13829 34561 13863 34595
rect 13863 34561 13872 34595
rect 13820 34552 13872 34561
rect 14924 34552 14976 34604
rect 11520 34484 11572 34536
rect 13544 34484 13596 34536
rect 9772 34348 9824 34400
rect 13360 34391 13412 34400
rect 13360 34357 13369 34391
rect 13369 34357 13403 34391
rect 13403 34357 13412 34391
rect 13360 34348 13412 34357
rect 2629 34246 2681 34298
rect 2693 34246 2745 34298
rect 2757 34246 2809 34298
rect 2821 34246 2873 34298
rect 2885 34246 2937 34298
rect 5987 34246 6039 34298
rect 6051 34246 6103 34298
rect 6115 34246 6167 34298
rect 6179 34246 6231 34298
rect 6243 34246 6295 34298
rect 9345 34246 9397 34298
rect 9409 34246 9461 34298
rect 9473 34246 9525 34298
rect 9537 34246 9589 34298
rect 9601 34246 9653 34298
rect 12703 34246 12755 34298
rect 12767 34246 12819 34298
rect 12831 34246 12883 34298
rect 12895 34246 12947 34298
rect 12959 34246 13011 34298
rect 4988 34144 5040 34196
rect 9864 34144 9916 34196
rect 10416 34187 10468 34196
rect 10416 34153 10425 34187
rect 10425 34153 10459 34187
rect 10459 34153 10468 34187
rect 10416 34144 10468 34153
rect 10968 34187 11020 34196
rect 10968 34153 10977 34187
rect 10977 34153 11011 34187
rect 11011 34153 11020 34187
rect 10968 34144 11020 34153
rect 11244 34187 11296 34196
rect 11244 34153 11253 34187
rect 11253 34153 11287 34187
rect 11287 34153 11296 34187
rect 11244 34144 11296 34153
rect 12348 34144 12400 34196
rect 12532 34076 12584 34128
rect 9956 34008 10008 34060
rect 9864 33940 9916 33992
rect 10140 33940 10192 33992
rect 10876 33979 10928 33992
rect 10876 33945 10885 33979
rect 10885 33945 10919 33979
rect 10919 33945 10928 33979
rect 12624 34008 12676 34060
rect 13912 34008 13964 34060
rect 10876 33940 10928 33945
rect 9864 33847 9916 33856
rect 9864 33813 9873 33847
rect 9873 33813 9907 33847
rect 9907 33813 9916 33847
rect 9864 33804 9916 33813
rect 11796 33872 11848 33924
rect 12256 33915 12308 33924
rect 12256 33881 12265 33915
rect 12265 33881 12299 33915
rect 12299 33881 12308 33915
rect 12256 33872 12308 33881
rect 11428 33804 11480 33856
rect 11612 33804 11664 33856
rect 13268 33872 13320 33924
rect 13544 33915 13596 33924
rect 13544 33881 13553 33915
rect 13553 33881 13587 33915
rect 13587 33881 13596 33915
rect 13544 33872 13596 33881
rect 12532 33804 12584 33856
rect 13728 33804 13780 33856
rect 4308 33702 4360 33754
rect 4372 33702 4424 33754
rect 4436 33702 4488 33754
rect 4500 33702 4552 33754
rect 4564 33702 4616 33754
rect 7666 33702 7718 33754
rect 7730 33702 7782 33754
rect 7794 33702 7846 33754
rect 7858 33702 7910 33754
rect 7922 33702 7974 33754
rect 11024 33702 11076 33754
rect 11088 33702 11140 33754
rect 11152 33702 11204 33754
rect 11216 33702 11268 33754
rect 11280 33702 11332 33754
rect 14382 33702 14434 33754
rect 14446 33702 14498 33754
rect 14510 33702 14562 33754
rect 14574 33702 14626 33754
rect 14638 33702 14690 33754
rect 9864 33600 9916 33652
rect 756 33464 808 33516
rect 10692 33464 10744 33516
rect 5540 33396 5592 33448
rect 9680 33396 9732 33448
rect 11612 33532 11664 33584
rect 13176 33600 13228 33652
rect 13728 33600 13780 33652
rect 11336 33507 11388 33516
rect 11336 33473 11345 33507
rect 11345 33473 11379 33507
rect 11379 33473 11388 33507
rect 11336 33464 11388 33473
rect 11428 33464 11480 33516
rect 12164 33464 12216 33516
rect 13176 33507 13228 33516
rect 13176 33473 13185 33507
rect 13185 33473 13219 33507
rect 13219 33473 13228 33507
rect 13176 33464 13228 33473
rect 4988 33260 5040 33312
rect 13728 33507 13780 33516
rect 13728 33473 13737 33507
rect 13737 33473 13771 33507
rect 13771 33473 13780 33507
rect 13728 33464 13780 33473
rect 11520 33439 11572 33448
rect 11520 33405 11529 33439
rect 11529 33405 11563 33439
rect 11563 33405 11572 33439
rect 11520 33396 11572 33405
rect 13636 33396 13688 33448
rect 11980 33260 12032 33312
rect 13544 33328 13596 33380
rect 12532 33303 12584 33312
rect 12532 33269 12541 33303
rect 12541 33269 12575 33303
rect 12575 33269 12584 33303
rect 12532 33260 12584 33269
rect 14188 33328 14240 33380
rect 15016 33260 15068 33312
rect 2629 33158 2681 33210
rect 2693 33158 2745 33210
rect 2757 33158 2809 33210
rect 2821 33158 2873 33210
rect 2885 33158 2937 33210
rect 5987 33158 6039 33210
rect 6051 33158 6103 33210
rect 6115 33158 6167 33210
rect 6179 33158 6231 33210
rect 6243 33158 6295 33210
rect 9345 33158 9397 33210
rect 9409 33158 9461 33210
rect 9473 33158 9525 33210
rect 9537 33158 9589 33210
rect 9601 33158 9653 33210
rect 12703 33158 12755 33210
rect 12767 33158 12819 33210
rect 12831 33158 12883 33210
rect 12895 33158 12947 33210
rect 12959 33158 13011 33210
rect 13544 33056 13596 33108
rect 8760 32988 8812 33040
rect 11152 32988 11204 33040
rect 12440 32988 12492 33040
rect 12900 32988 12952 33040
rect 756 32852 808 32904
rect 9404 32852 9456 32904
rect 10324 32895 10376 32904
rect 10324 32861 10333 32895
rect 10333 32861 10367 32895
rect 10367 32861 10376 32895
rect 10324 32852 10376 32861
rect 11520 32963 11572 32972
rect 11520 32929 11529 32963
rect 11529 32929 11563 32963
rect 11563 32929 11572 32963
rect 11520 32920 11572 32929
rect 13544 32920 13596 32972
rect 6920 32784 6972 32836
rect 10508 32784 10560 32836
rect 1584 32759 1636 32768
rect 1584 32725 1593 32759
rect 1593 32725 1627 32759
rect 1627 32725 1636 32759
rect 1584 32716 1636 32725
rect 1860 32716 1912 32768
rect 10140 32759 10192 32768
rect 10140 32725 10149 32759
rect 10149 32725 10183 32759
rect 10183 32725 10192 32759
rect 10140 32716 10192 32725
rect 10968 32852 11020 32904
rect 10784 32784 10836 32836
rect 11152 32784 11204 32836
rect 11244 32716 11296 32768
rect 12808 32716 12860 32768
rect 13360 32784 13412 32836
rect 14280 32784 14332 32836
rect 4308 32614 4360 32666
rect 4372 32614 4424 32666
rect 4436 32614 4488 32666
rect 4500 32614 4552 32666
rect 4564 32614 4616 32666
rect 7666 32614 7718 32666
rect 7730 32614 7782 32666
rect 7794 32614 7846 32666
rect 7858 32614 7910 32666
rect 7922 32614 7974 32666
rect 11024 32614 11076 32666
rect 11088 32614 11140 32666
rect 11152 32614 11204 32666
rect 11216 32614 11268 32666
rect 11280 32614 11332 32666
rect 14382 32614 14434 32666
rect 14446 32614 14498 32666
rect 14510 32614 14562 32666
rect 14574 32614 14626 32666
rect 14638 32614 14690 32666
rect 10140 32512 10192 32564
rect 13176 32512 13228 32564
rect 13268 32444 13320 32496
rect 8576 32376 8628 32428
rect 9404 32419 9456 32428
rect 9404 32385 9413 32419
rect 9413 32385 9456 32419
rect 9404 32376 9456 32385
rect 10692 32419 10744 32428
rect 10692 32385 10701 32419
rect 10701 32385 10735 32419
rect 10735 32385 10744 32419
rect 10692 32376 10744 32385
rect 7380 32308 7432 32360
rect 9864 32308 9916 32360
rect 11152 32376 11204 32428
rect 12348 32376 12400 32428
rect 11060 32308 11112 32360
rect 11520 32351 11572 32360
rect 11520 32317 11529 32351
rect 11529 32317 11563 32351
rect 11563 32317 11572 32351
rect 11520 32308 11572 32317
rect 15108 32376 15160 32428
rect 13912 32308 13964 32360
rect 4804 32240 4856 32292
rect 11152 32240 11204 32292
rect 10140 32215 10192 32224
rect 10140 32181 10149 32215
rect 10149 32181 10183 32215
rect 10183 32181 10192 32215
rect 10140 32172 10192 32181
rect 12256 32172 12308 32224
rect 12532 32215 12584 32224
rect 12532 32181 12541 32215
rect 12541 32181 12575 32215
rect 12575 32181 12584 32215
rect 12532 32172 12584 32181
rect 13268 32215 13320 32224
rect 13268 32181 13277 32215
rect 13277 32181 13311 32215
rect 13311 32181 13320 32215
rect 13268 32172 13320 32181
rect 15200 32172 15252 32224
rect 2629 32070 2681 32122
rect 2693 32070 2745 32122
rect 2757 32070 2809 32122
rect 2821 32070 2873 32122
rect 2885 32070 2937 32122
rect 5987 32070 6039 32122
rect 6051 32070 6103 32122
rect 6115 32070 6167 32122
rect 6179 32070 6231 32122
rect 6243 32070 6295 32122
rect 9345 32070 9397 32122
rect 9409 32070 9461 32122
rect 9473 32070 9525 32122
rect 9537 32070 9589 32122
rect 9601 32070 9653 32122
rect 12703 32070 12755 32122
rect 12767 32070 12819 32122
rect 12831 32070 12883 32122
rect 12895 32070 12947 32122
rect 12959 32070 13011 32122
rect 10692 31968 10744 32020
rect 10784 32011 10836 32020
rect 10784 31977 10793 32011
rect 10793 31977 10827 32011
rect 10827 31977 10836 32011
rect 10784 31968 10836 31977
rect 11980 31968 12032 32020
rect 12256 31968 12308 32020
rect 15384 31968 15436 32020
rect 7380 31832 7432 31884
rect 11244 31900 11296 31952
rect 11796 31900 11848 31952
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 7196 31764 7248 31816
rect 8208 31764 8260 31816
rect 8852 31764 8904 31816
rect 10140 31807 10192 31816
rect 10140 31773 10149 31807
rect 10149 31773 10183 31807
rect 10183 31773 10192 31807
rect 10140 31764 10192 31773
rect 10508 31764 10560 31816
rect 10784 31764 10836 31816
rect 10876 31696 10928 31748
rect 1768 31628 1820 31680
rect 9220 31628 9272 31680
rect 9680 31628 9732 31680
rect 12072 31832 12124 31884
rect 11336 31807 11388 31816
rect 11336 31773 11345 31807
rect 11345 31773 11379 31807
rect 11379 31773 11388 31807
rect 11336 31764 11388 31773
rect 11704 31807 11756 31816
rect 11704 31773 11713 31807
rect 11713 31773 11747 31807
rect 11747 31773 11756 31807
rect 11704 31764 11756 31773
rect 11796 31696 11848 31748
rect 12256 31764 12308 31816
rect 14004 31832 14056 31884
rect 13636 31764 13688 31816
rect 15292 31764 15344 31816
rect 12992 31628 13044 31680
rect 13544 31628 13596 31680
rect 15568 31696 15620 31748
rect 14280 31628 14332 31680
rect 4308 31526 4360 31578
rect 4372 31526 4424 31578
rect 4436 31526 4488 31578
rect 4500 31526 4552 31578
rect 4564 31526 4616 31578
rect 7666 31526 7718 31578
rect 7730 31526 7782 31578
rect 7794 31526 7846 31578
rect 7858 31526 7910 31578
rect 7922 31526 7974 31578
rect 11024 31526 11076 31578
rect 11088 31526 11140 31578
rect 11152 31526 11204 31578
rect 11216 31526 11268 31578
rect 11280 31526 11332 31578
rect 14382 31526 14434 31578
rect 14446 31526 14498 31578
rect 14510 31526 14562 31578
rect 14574 31526 14626 31578
rect 14638 31526 14690 31578
rect 7012 31424 7064 31476
rect 9864 31467 9916 31476
rect 9864 31433 9873 31467
rect 9873 31433 9907 31467
rect 9907 31433 9916 31467
rect 9864 31424 9916 31433
rect 10784 31424 10836 31476
rect 12716 31424 12768 31476
rect 13360 31424 13412 31476
rect 756 31288 808 31340
rect 6552 31288 6604 31340
rect 8024 31263 8076 31272
rect 8024 31229 8033 31263
rect 8033 31229 8067 31263
rect 8067 31229 8076 31263
rect 8024 31220 8076 31229
rect 8944 31331 8996 31340
rect 8944 31297 8953 31331
rect 8953 31297 8987 31331
rect 8987 31297 8996 31331
rect 8944 31288 8996 31297
rect 9220 31331 9272 31340
rect 9220 31297 9229 31331
rect 9229 31297 9263 31331
rect 9263 31297 9272 31331
rect 9220 31288 9272 31297
rect 10692 31331 10744 31340
rect 10692 31297 10701 31331
rect 10701 31297 10735 31331
rect 10735 31297 10744 31331
rect 10692 31288 10744 31297
rect 12900 31331 12952 31340
rect 12900 31297 12909 31331
rect 12909 31297 12943 31331
rect 12943 31297 12952 31331
rect 12900 31288 12952 31297
rect 14188 31288 14240 31340
rect 3792 31084 3844 31136
rect 9772 31220 9824 31272
rect 10416 31220 10468 31272
rect 11520 31220 11572 31272
rect 11888 31263 11940 31272
rect 11888 31229 11897 31263
rect 11897 31229 11931 31263
rect 11931 31229 11940 31263
rect 11888 31220 11940 31229
rect 12348 31263 12400 31272
rect 12348 31229 12357 31263
rect 12357 31229 12391 31263
rect 12391 31229 12400 31263
rect 12348 31220 12400 31229
rect 12624 31263 12676 31272
rect 12624 31229 12633 31263
rect 12633 31229 12667 31263
rect 12667 31229 12676 31263
rect 12624 31220 12676 31229
rect 8668 31195 8720 31204
rect 8668 31161 8677 31195
rect 8677 31161 8711 31195
rect 8711 31161 8720 31195
rect 8668 31152 8720 31161
rect 11428 31152 11480 31204
rect 9128 31084 9180 31136
rect 9220 31084 9272 31136
rect 11152 31084 11204 31136
rect 11612 31084 11664 31136
rect 12716 31084 12768 31136
rect 13268 31084 13320 31136
rect 13636 31084 13688 31136
rect 14280 31084 14332 31136
rect 15568 31084 15620 31136
rect 2629 30982 2681 31034
rect 2693 30982 2745 31034
rect 2757 30982 2809 31034
rect 2821 30982 2873 31034
rect 2885 30982 2937 31034
rect 5987 30982 6039 31034
rect 6051 30982 6103 31034
rect 6115 30982 6167 31034
rect 6179 30982 6231 31034
rect 6243 30982 6295 31034
rect 9345 30982 9397 31034
rect 9409 30982 9461 31034
rect 9473 30982 9525 31034
rect 9537 30982 9589 31034
rect 9601 30982 9653 31034
rect 12703 30982 12755 31034
rect 12767 30982 12819 31034
rect 12831 30982 12883 31034
rect 12895 30982 12947 31034
rect 12959 30982 13011 31034
rect 7380 30880 7432 30932
rect 8668 30880 8720 30932
rect 9036 30880 9088 30932
rect 9956 30880 10008 30932
rect 10324 30880 10376 30932
rect 11152 30880 11204 30932
rect 12440 30855 12492 30864
rect 12440 30821 12449 30855
rect 12449 30821 12483 30855
rect 12483 30821 12492 30855
rect 12440 30812 12492 30821
rect 13728 30812 13780 30864
rect 8852 30608 8904 30660
rect 9680 30676 9732 30728
rect 10600 30676 10652 30728
rect 11796 30719 11848 30728
rect 11796 30685 11805 30719
rect 11805 30685 11839 30719
rect 11839 30685 11848 30719
rect 11796 30676 11848 30685
rect 11888 30676 11940 30728
rect 12716 30719 12768 30728
rect 12716 30685 12725 30719
rect 12725 30685 12759 30719
rect 12759 30685 12768 30719
rect 12716 30676 12768 30685
rect 12808 30719 12860 30728
rect 12808 30685 12842 30719
rect 12842 30685 12860 30719
rect 12808 30676 12860 30685
rect 12992 30719 13044 30728
rect 12992 30685 13001 30719
rect 13001 30685 13035 30719
rect 13035 30685 13044 30719
rect 12992 30676 13044 30685
rect 7380 30540 7432 30592
rect 9036 30540 9088 30592
rect 9220 30540 9272 30592
rect 9588 30540 9640 30592
rect 12256 30540 12308 30592
rect 14372 30608 14424 30660
rect 15476 30608 15528 30660
rect 4308 30438 4360 30490
rect 4372 30438 4424 30490
rect 4436 30438 4488 30490
rect 4500 30438 4552 30490
rect 4564 30438 4616 30490
rect 7666 30438 7718 30490
rect 7730 30438 7782 30490
rect 7794 30438 7846 30490
rect 7858 30438 7910 30490
rect 7922 30438 7974 30490
rect 11024 30438 11076 30490
rect 11088 30438 11140 30490
rect 11152 30438 11204 30490
rect 11216 30438 11268 30490
rect 11280 30438 11332 30490
rect 14382 30438 14434 30490
rect 14446 30438 14498 30490
rect 14510 30438 14562 30490
rect 14574 30438 14626 30490
rect 14638 30438 14690 30490
rect 8208 30336 8260 30388
rect 10692 30336 10744 30388
rect 12440 30336 12492 30388
rect 12808 30336 12860 30388
rect 11704 30268 11756 30320
rect 13820 30311 13872 30320
rect 13820 30277 13829 30311
rect 13829 30277 13863 30311
rect 13863 30277 13872 30311
rect 13820 30268 13872 30277
rect 756 30200 808 30252
rect 10232 30243 10284 30252
rect 10232 30209 10241 30243
rect 10241 30209 10275 30243
rect 10275 30209 10284 30243
rect 10232 30200 10284 30209
rect 13176 30243 13228 30252
rect 13176 30209 13185 30243
rect 13185 30209 13219 30243
rect 13219 30209 13228 30243
rect 13176 30200 13228 30209
rect 9036 30175 9088 30184
rect 9036 30141 9045 30175
rect 9045 30141 9079 30175
rect 9079 30141 9088 30175
rect 9036 30132 9088 30141
rect 9128 30132 9180 30184
rect 9588 30132 9640 30184
rect 8668 30064 8720 30116
rect 9312 30064 9364 30116
rect 5540 29996 5592 30048
rect 8484 29996 8536 30048
rect 8944 29996 8996 30048
rect 10048 30175 10100 30184
rect 10048 30141 10082 30175
rect 10082 30141 10100 30175
rect 10048 30132 10100 30141
rect 11980 30175 12032 30184
rect 11980 30141 11989 30175
rect 11989 30141 12023 30175
rect 12023 30141 12032 30175
rect 11980 30132 12032 30141
rect 12164 30175 12216 30184
rect 12164 30141 12173 30175
rect 12173 30141 12207 30175
rect 12207 30141 12216 30175
rect 12164 30132 12216 30141
rect 12256 30132 12308 30184
rect 12716 30132 12768 30184
rect 12992 30175 13044 30184
rect 12992 30141 13026 30175
rect 13026 30141 13044 30175
rect 12992 30132 13044 30141
rect 10692 30064 10744 30116
rect 13912 30107 13964 30116
rect 13912 30073 13921 30107
rect 13921 30073 13955 30107
rect 13955 30073 13964 30107
rect 13912 30064 13964 30073
rect 2629 29894 2681 29946
rect 2693 29894 2745 29946
rect 2757 29894 2809 29946
rect 2821 29894 2873 29946
rect 2885 29894 2937 29946
rect 5987 29894 6039 29946
rect 6051 29894 6103 29946
rect 6115 29894 6167 29946
rect 6179 29894 6231 29946
rect 6243 29894 6295 29946
rect 9345 29894 9397 29946
rect 9409 29894 9461 29946
rect 9473 29894 9525 29946
rect 9537 29894 9589 29946
rect 9601 29894 9653 29946
rect 12703 29894 12755 29946
rect 12767 29894 12819 29946
rect 12831 29894 12883 29946
rect 12895 29894 12947 29946
rect 12959 29894 13011 29946
rect 2136 29835 2188 29844
rect 2136 29801 2145 29835
rect 2145 29801 2179 29835
rect 2179 29801 2188 29835
rect 2136 29792 2188 29801
rect 7104 29792 7156 29844
rect 7288 29792 7340 29844
rect 756 29588 808 29640
rect 3792 29588 3844 29640
rect 8116 29656 8168 29708
rect 7288 29588 7340 29640
rect 7472 29588 7524 29640
rect 2044 29452 2096 29504
rect 6828 29452 6880 29504
rect 7472 29452 7524 29504
rect 9680 29588 9732 29640
rect 10508 29588 10560 29640
rect 12072 29792 12124 29844
rect 14924 29792 14976 29844
rect 11796 29656 11848 29708
rect 8944 29520 8996 29572
rect 11428 29520 11480 29572
rect 11704 29520 11756 29572
rect 13176 29520 13228 29572
rect 9680 29452 9732 29504
rect 9772 29452 9824 29504
rect 10692 29452 10744 29504
rect 12072 29452 12124 29504
rect 12256 29495 12308 29504
rect 12256 29461 12265 29495
rect 12265 29461 12299 29495
rect 12299 29461 12308 29495
rect 12256 29452 12308 29461
rect 12348 29452 12400 29504
rect 12532 29452 12584 29504
rect 13544 29452 13596 29504
rect 4308 29350 4360 29402
rect 4372 29350 4424 29402
rect 4436 29350 4488 29402
rect 4500 29350 4552 29402
rect 4564 29350 4616 29402
rect 7666 29350 7718 29402
rect 7730 29350 7782 29402
rect 7794 29350 7846 29402
rect 7858 29350 7910 29402
rect 7922 29350 7974 29402
rect 11024 29350 11076 29402
rect 11088 29350 11140 29402
rect 11152 29350 11204 29402
rect 11216 29350 11268 29402
rect 11280 29350 11332 29402
rect 14382 29350 14434 29402
rect 14446 29350 14498 29402
rect 14510 29350 14562 29402
rect 14574 29350 14626 29402
rect 14638 29350 14690 29402
rect 6828 29248 6880 29300
rect 11888 29248 11940 29300
rect 13360 29248 13412 29300
rect 7104 29155 7156 29164
rect 7104 29121 7113 29155
rect 7113 29121 7147 29155
rect 7147 29121 7156 29155
rect 7104 29112 7156 29121
rect 8392 29112 8444 29164
rect 8668 29112 8720 29164
rect 9772 29112 9824 29164
rect 10232 29180 10284 29232
rect 10508 29180 10560 29232
rect 10784 29180 10836 29232
rect 12624 29180 12676 29232
rect 10140 29155 10192 29164
rect 10140 29121 10147 29155
rect 10147 29121 10181 29155
rect 10181 29121 10192 29155
rect 10140 29112 10192 29121
rect 11060 29112 11112 29164
rect 13636 29112 13688 29164
rect 5540 28908 5592 28960
rect 9680 29044 9732 29096
rect 11612 29044 11664 29096
rect 11796 29087 11848 29096
rect 11796 29053 11805 29087
rect 11805 29053 11839 29087
rect 11839 29053 11848 29087
rect 11796 29044 11848 29053
rect 8116 28951 8168 28960
rect 8116 28917 8125 28951
rect 8125 28917 8159 28951
rect 8159 28917 8168 28951
rect 8116 28908 8168 28917
rect 11336 28976 11388 29028
rect 11704 28976 11756 29028
rect 13820 29019 13872 29028
rect 13820 28985 13829 29019
rect 13829 28985 13863 29019
rect 13863 28985 13872 29019
rect 13820 28976 13872 28985
rect 10140 28908 10192 28960
rect 10876 28951 10928 28960
rect 10876 28917 10885 28951
rect 10885 28917 10919 28951
rect 10919 28917 10928 28951
rect 10876 28908 10928 28917
rect 12256 28908 12308 28960
rect 12716 28908 12768 28960
rect 13084 28908 13136 28960
rect 2629 28806 2681 28858
rect 2693 28806 2745 28858
rect 2757 28806 2809 28858
rect 2821 28806 2873 28858
rect 2885 28806 2937 28858
rect 5987 28806 6039 28858
rect 6051 28806 6103 28858
rect 6115 28806 6167 28858
rect 6179 28806 6231 28858
rect 6243 28806 6295 28858
rect 9345 28806 9397 28858
rect 9409 28806 9461 28858
rect 9473 28806 9525 28858
rect 9537 28806 9589 28858
rect 9601 28806 9653 28858
rect 12703 28806 12755 28858
rect 12767 28806 12819 28858
rect 12831 28806 12883 28858
rect 12895 28806 12947 28858
rect 12959 28806 13011 28858
rect 1952 28704 2004 28756
rect 12256 28704 12308 28756
rect 13268 28704 13320 28756
rect 10876 28636 10928 28688
rect 7104 28611 7156 28620
rect 7104 28577 7113 28611
rect 7113 28577 7147 28611
rect 7147 28577 7156 28611
rect 7104 28568 7156 28577
rect 11796 28611 11848 28620
rect 11796 28577 11805 28611
rect 11805 28577 11839 28611
rect 11839 28577 11848 28611
rect 11796 28568 11848 28577
rect 15016 28568 15068 28620
rect 756 28500 808 28552
rect 6460 28500 6512 28552
rect 6920 28500 6972 28552
rect 8944 28500 8996 28552
rect 9220 28500 9272 28552
rect 7104 28364 7156 28416
rect 7564 28364 7616 28416
rect 8300 28364 8352 28416
rect 8668 28364 8720 28416
rect 8944 28364 8996 28416
rect 9680 28364 9732 28416
rect 11888 28543 11940 28552
rect 11888 28509 11922 28543
rect 11922 28509 11940 28543
rect 11888 28500 11940 28509
rect 12072 28543 12124 28552
rect 12072 28509 12081 28543
rect 12081 28509 12115 28543
rect 12115 28509 12124 28543
rect 12072 28500 12124 28509
rect 12716 28500 12768 28552
rect 12808 28432 12860 28484
rect 11888 28364 11940 28416
rect 12716 28364 12768 28416
rect 13084 28364 13136 28416
rect 13728 28407 13780 28416
rect 13728 28373 13737 28407
rect 13737 28373 13771 28407
rect 13771 28373 13780 28407
rect 13728 28364 13780 28373
rect 4308 28262 4360 28314
rect 4372 28262 4424 28314
rect 4436 28262 4488 28314
rect 4500 28262 4552 28314
rect 4564 28262 4616 28314
rect 7666 28262 7718 28314
rect 7730 28262 7782 28314
rect 7794 28262 7846 28314
rect 7858 28262 7910 28314
rect 7922 28262 7974 28314
rect 11024 28262 11076 28314
rect 11088 28262 11140 28314
rect 11152 28262 11204 28314
rect 11216 28262 11268 28314
rect 11280 28262 11332 28314
rect 14382 28262 14434 28314
rect 14446 28262 14498 28314
rect 14510 28262 14562 28314
rect 14574 28262 14626 28314
rect 14638 28262 14690 28314
rect 7104 28160 7156 28212
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 11888 28160 11940 28212
rect 8208 28067 8260 28076
rect 8208 28033 8217 28067
rect 8217 28033 8251 28067
rect 8251 28033 8260 28067
rect 8208 28024 8260 28033
rect 7288 27956 7340 28008
rect 7564 27956 7616 28008
rect 7932 27999 7984 28008
rect 7932 27965 7941 27999
rect 7941 27965 7975 27999
rect 7975 27965 7984 27999
rect 7932 27956 7984 27965
rect 8944 27999 8996 28008
rect 8944 27965 8953 27999
rect 8953 27965 8987 27999
rect 8987 27965 8996 27999
rect 8944 27956 8996 27965
rect 9956 28067 10008 28076
rect 9956 28033 9990 28067
rect 9990 28033 10008 28067
rect 9956 28024 10008 28033
rect 10140 28067 10192 28076
rect 10140 28033 10149 28067
rect 10149 28033 10183 28067
rect 10183 28033 10192 28067
rect 10140 28024 10192 28033
rect 10968 28067 11020 28076
rect 10968 28033 10977 28067
rect 10977 28033 11011 28067
rect 11011 28033 11020 28067
rect 10968 28024 11020 28033
rect 11980 28024 12032 28076
rect 13452 28160 13504 28212
rect 14188 28203 14240 28212
rect 14188 28169 14197 28203
rect 14197 28169 14231 28203
rect 14231 28169 14240 28203
rect 14188 28160 14240 28169
rect 9312 27956 9364 28008
rect 1584 27863 1636 27872
rect 1584 27829 1593 27863
rect 1593 27829 1627 27863
rect 1627 27829 1636 27863
rect 1584 27820 1636 27829
rect 8116 27820 8168 27872
rect 8944 27820 8996 27872
rect 10784 27956 10836 28008
rect 10048 27820 10100 27872
rect 10692 27820 10744 27872
rect 10784 27863 10836 27872
rect 10784 27829 10793 27863
rect 10793 27829 10827 27863
rect 10827 27829 10836 27863
rect 10784 27820 10836 27829
rect 11612 27820 11664 27872
rect 12072 27820 12124 27872
rect 13544 28067 13596 28076
rect 13544 28033 13553 28067
rect 13553 28033 13587 28067
rect 13587 28033 13596 28067
rect 13544 28024 13596 28033
rect 12348 27999 12400 28008
rect 12348 27965 12357 27999
rect 12357 27965 12391 27999
rect 12391 27965 12400 27999
rect 12348 27956 12400 27965
rect 12716 27956 12768 28008
rect 13360 27999 13412 28008
rect 13360 27965 13394 27999
rect 13394 27965 13412 27999
rect 13360 27956 13412 27965
rect 13084 27820 13136 27872
rect 2629 27718 2681 27770
rect 2693 27718 2745 27770
rect 2757 27718 2809 27770
rect 2821 27718 2873 27770
rect 2885 27718 2937 27770
rect 5987 27718 6039 27770
rect 6051 27718 6103 27770
rect 6115 27718 6167 27770
rect 6179 27718 6231 27770
rect 6243 27718 6295 27770
rect 9345 27718 9397 27770
rect 9409 27718 9461 27770
rect 9473 27718 9525 27770
rect 9537 27718 9589 27770
rect 9601 27718 9653 27770
rect 12703 27718 12755 27770
rect 12767 27718 12819 27770
rect 12831 27718 12883 27770
rect 12895 27718 12947 27770
rect 12959 27718 13011 27770
rect 6828 27616 6880 27668
rect 3056 27548 3108 27600
rect 3884 27548 3936 27600
rect 7472 27548 7524 27600
rect 1676 27480 1728 27532
rect 7380 27480 7432 27532
rect 1860 27412 1912 27464
rect 2688 27455 2740 27464
rect 2688 27421 2697 27455
rect 2697 27421 2731 27455
rect 2731 27421 2740 27455
rect 2688 27412 2740 27421
rect 6460 27412 6512 27464
rect 8208 27616 8260 27668
rect 8208 27412 8260 27464
rect 10968 27616 11020 27668
rect 11704 27616 11756 27668
rect 9680 27548 9732 27600
rect 9956 27548 10008 27600
rect 10232 27455 10284 27464
rect 10232 27421 10241 27455
rect 10241 27421 10275 27455
rect 10275 27421 10284 27455
rect 10232 27412 10284 27421
rect 11888 27425 11940 27464
rect 7196 27276 7248 27328
rect 8760 27276 8812 27328
rect 9680 27276 9732 27328
rect 10232 27276 10284 27328
rect 11888 27412 11913 27425
rect 11913 27412 11940 27425
rect 12348 27344 12400 27396
rect 13452 27387 13504 27396
rect 13452 27353 13461 27387
rect 13461 27353 13495 27387
rect 13495 27353 13504 27387
rect 13452 27344 13504 27353
rect 11704 27276 11756 27328
rect 12716 27276 12768 27328
rect 4308 27174 4360 27226
rect 4372 27174 4424 27226
rect 4436 27174 4488 27226
rect 4500 27174 4552 27226
rect 4564 27174 4616 27226
rect 7666 27174 7718 27226
rect 7730 27174 7782 27226
rect 7794 27174 7846 27226
rect 7858 27174 7910 27226
rect 7922 27174 7974 27226
rect 11024 27174 11076 27226
rect 11088 27174 11140 27226
rect 11152 27174 11204 27226
rect 11216 27174 11268 27226
rect 11280 27174 11332 27226
rect 14382 27174 14434 27226
rect 14446 27174 14498 27226
rect 14510 27174 14562 27226
rect 14574 27174 14626 27226
rect 14638 27174 14690 27226
rect 1676 27072 1728 27124
rect 2688 27072 2740 27124
rect 7380 27072 7432 27124
rect 5448 27004 5500 27056
rect 6460 27004 6512 27056
rect 8208 27115 8260 27124
rect 8208 27081 8217 27115
rect 8217 27081 8251 27115
rect 8251 27081 8260 27115
rect 8208 27072 8260 27081
rect 10600 27072 10652 27124
rect 11796 27072 11848 27124
rect 756 26936 808 26988
rect 4160 26936 4212 26988
rect 4896 26979 4948 26988
rect 4896 26945 4905 26979
rect 4905 26945 4939 26979
rect 4939 26945 4948 26979
rect 4896 26936 4948 26945
rect 5172 26979 5224 26988
rect 5172 26945 5179 26979
rect 5179 26945 5213 26979
rect 5213 26945 5224 26979
rect 5172 26936 5224 26945
rect 5908 26936 5960 26988
rect 7564 26979 7616 26988
rect 7564 26945 7573 26979
rect 7573 26945 7607 26979
rect 7607 26945 7616 26979
rect 7564 26936 7616 26945
rect 9680 26936 9732 26988
rect 6552 26911 6604 26920
rect 6552 26877 6561 26911
rect 6561 26877 6595 26911
rect 6595 26877 6604 26911
rect 6552 26868 6604 26877
rect 5816 26732 5868 26784
rect 7380 26911 7432 26920
rect 7380 26877 7414 26911
rect 7414 26877 7432 26911
rect 7380 26868 7432 26877
rect 7748 26868 7800 26920
rect 12716 26936 12768 26988
rect 8484 26732 8536 26784
rect 10876 26868 10928 26920
rect 11796 26868 11848 26920
rect 12256 26868 12308 26920
rect 12532 26911 12584 26920
rect 12532 26877 12541 26911
rect 12541 26877 12575 26911
rect 12575 26877 12584 26911
rect 12532 26868 12584 26877
rect 13084 26868 13136 26920
rect 13360 26911 13412 26920
rect 13360 26877 13394 26911
rect 13394 26877 13412 26911
rect 13360 26868 13412 26877
rect 13544 26911 13596 26920
rect 13544 26877 13553 26911
rect 13553 26877 13587 26911
rect 13587 26877 13596 26911
rect 13544 26868 13596 26877
rect 12348 26800 12400 26852
rect 10876 26775 10928 26784
rect 10876 26741 10885 26775
rect 10885 26741 10919 26775
rect 10919 26741 10928 26775
rect 10876 26732 10928 26741
rect 14004 26732 14056 26784
rect 2629 26630 2681 26682
rect 2693 26630 2745 26682
rect 2757 26630 2809 26682
rect 2821 26630 2873 26682
rect 2885 26630 2937 26682
rect 5987 26630 6039 26682
rect 6051 26630 6103 26682
rect 6115 26630 6167 26682
rect 6179 26630 6231 26682
rect 6243 26630 6295 26682
rect 9345 26630 9397 26682
rect 9409 26630 9461 26682
rect 9473 26630 9525 26682
rect 9537 26630 9589 26682
rect 9601 26630 9653 26682
rect 12703 26630 12755 26682
rect 12767 26630 12819 26682
rect 12831 26630 12883 26682
rect 12895 26630 12947 26682
rect 12959 26630 13011 26682
rect 4896 26460 4948 26512
rect 4896 26324 4948 26376
rect 10048 26528 10100 26580
rect 10876 26528 10928 26580
rect 12624 26528 12676 26580
rect 13544 26528 13596 26580
rect 9128 26460 9180 26512
rect 10508 26460 10560 26512
rect 7380 26435 7432 26444
rect 7380 26401 7414 26435
rect 7414 26401 7432 26435
rect 7380 26392 7432 26401
rect 10692 26435 10744 26444
rect 10692 26401 10701 26435
rect 10701 26401 10735 26435
rect 10735 26401 10744 26435
rect 10692 26392 10744 26401
rect 5908 26324 5960 26376
rect 6552 26367 6604 26376
rect 6552 26333 6561 26367
rect 6561 26333 6595 26367
rect 6595 26333 6604 26367
rect 6552 26324 6604 26333
rect 7288 26367 7340 26376
rect 7288 26333 7297 26367
rect 7297 26333 7331 26367
rect 7331 26333 7340 26367
rect 7288 26324 7340 26333
rect 7564 26367 7616 26376
rect 7564 26333 7573 26367
rect 7573 26333 7607 26367
rect 7607 26333 7616 26367
rect 7564 26324 7616 26333
rect 10600 26324 10652 26376
rect 10876 26392 10928 26444
rect 12072 26392 12124 26444
rect 1492 26299 1544 26308
rect 1492 26265 1501 26299
rect 1501 26265 1535 26299
rect 1535 26265 1544 26299
rect 1492 26256 1544 26265
rect 5724 26256 5776 26308
rect 6276 26256 6328 26308
rect 9864 26256 9916 26308
rect 11704 26367 11756 26376
rect 11704 26333 11713 26367
rect 11713 26333 11747 26367
rect 11747 26333 11756 26367
rect 11704 26324 11756 26333
rect 5172 26188 5224 26240
rect 6552 26188 6604 26240
rect 6828 26188 6880 26240
rect 7380 26188 7432 26240
rect 9588 26188 9640 26240
rect 12532 26256 12584 26308
rect 13268 26324 13320 26376
rect 4308 26086 4360 26138
rect 4372 26086 4424 26138
rect 4436 26086 4488 26138
rect 4500 26086 4552 26138
rect 4564 26086 4616 26138
rect 7666 26086 7718 26138
rect 7730 26086 7782 26138
rect 7794 26086 7846 26138
rect 7858 26086 7910 26138
rect 7922 26086 7974 26138
rect 11024 26086 11076 26138
rect 11088 26086 11140 26138
rect 11152 26086 11204 26138
rect 11216 26086 11268 26138
rect 11280 26086 11332 26138
rect 14382 26086 14434 26138
rect 14446 26086 14498 26138
rect 14510 26086 14562 26138
rect 14574 26086 14626 26138
rect 14638 26086 14690 26138
rect 6920 25916 6972 25968
rect 8668 25984 8720 26036
rect 10048 25984 10100 26036
rect 10416 25984 10468 26036
rect 13636 25984 13688 26036
rect 10232 25916 10284 25968
rect 12256 25916 12308 25968
rect 11612 25891 11664 25900
rect 11612 25857 11621 25891
rect 11621 25857 11655 25891
rect 11655 25857 11664 25891
rect 11612 25848 11664 25857
rect 12072 25848 12124 25900
rect 12440 25848 12492 25900
rect 6460 25644 6512 25696
rect 12348 25823 12400 25832
rect 12348 25789 12357 25823
rect 12357 25789 12391 25823
rect 12391 25789 12400 25823
rect 12348 25780 12400 25789
rect 13268 25891 13320 25900
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 13544 25823 13596 25832
rect 13544 25789 13553 25823
rect 13553 25789 13587 25823
rect 13587 25789 13596 25823
rect 13544 25780 13596 25789
rect 8208 25712 8260 25764
rect 7932 25687 7984 25696
rect 7932 25653 7941 25687
rect 7941 25653 7975 25687
rect 7975 25653 7984 25687
rect 7932 25644 7984 25653
rect 9588 25712 9640 25764
rect 9680 25644 9732 25696
rect 11152 25712 11204 25764
rect 12624 25712 12676 25764
rect 10692 25687 10744 25696
rect 10692 25653 10701 25687
rect 10701 25653 10735 25687
rect 10735 25653 10744 25687
rect 10692 25644 10744 25653
rect 11888 25687 11940 25696
rect 11888 25653 11897 25687
rect 11897 25653 11931 25687
rect 11931 25653 11940 25687
rect 11888 25644 11940 25653
rect 12808 25644 12860 25696
rect 13268 25644 13320 25696
rect 2629 25542 2681 25594
rect 2693 25542 2745 25594
rect 2757 25542 2809 25594
rect 2821 25542 2873 25594
rect 2885 25542 2937 25594
rect 5987 25542 6039 25594
rect 6051 25542 6103 25594
rect 6115 25542 6167 25594
rect 6179 25542 6231 25594
rect 6243 25542 6295 25594
rect 9345 25542 9397 25594
rect 9409 25542 9461 25594
rect 9473 25542 9525 25594
rect 9537 25542 9589 25594
rect 9601 25542 9653 25594
rect 12703 25542 12755 25594
rect 12767 25542 12819 25594
rect 12831 25542 12883 25594
rect 12895 25542 12947 25594
rect 12959 25542 13011 25594
rect 7564 25440 7616 25492
rect 7932 25440 7984 25492
rect 11428 25440 11480 25492
rect 11612 25440 11664 25492
rect 12624 25440 12676 25492
rect 14096 25372 14148 25424
rect 4896 25304 4948 25356
rect 6460 25347 6512 25356
rect 6460 25313 6469 25347
rect 6469 25313 6503 25347
rect 6503 25313 6512 25347
rect 6460 25304 6512 25313
rect 7564 25304 7616 25356
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 756 25236 808 25288
rect 5724 25236 5776 25288
rect 8944 25279 8996 25288
rect 8944 25245 8953 25279
rect 8953 25245 8987 25279
rect 8987 25245 8996 25279
rect 8944 25236 8996 25245
rect 9956 25279 10008 25288
rect 10968 25304 11020 25356
rect 11152 25304 11204 25356
rect 9956 25245 9990 25279
rect 9990 25245 10008 25279
rect 9956 25236 10008 25245
rect 10416 25100 10468 25152
rect 14188 25304 14240 25356
rect 11428 25168 11480 25220
rect 11888 25168 11940 25220
rect 12808 25211 12860 25220
rect 12808 25177 12817 25211
rect 12817 25177 12851 25211
rect 12851 25177 12860 25211
rect 12808 25168 12860 25177
rect 13084 25168 13136 25220
rect 11612 25100 11664 25152
rect 13820 25143 13872 25152
rect 13820 25109 13829 25143
rect 13829 25109 13863 25143
rect 13863 25109 13872 25143
rect 13820 25100 13872 25109
rect 4308 24998 4360 25050
rect 4372 24998 4424 25050
rect 4436 24998 4488 25050
rect 4500 24998 4552 25050
rect 4564 24998 4616 25050
rect 7666 24998 7718 25050
rect 7730 24998 7782 25050
rect 7794 24998 7846 25050
rect 7858 24998 7910 25050
rect 7922 24998 7974 25050
rect 11024 24998 11076 25050
rect 11088 24998 11140 25050
rect 11152 24998 11204 25050
rect 11216 24998 11268 25050
rect 11280 24998 11332 25050
rect 14382 24998 14434 25050
rect 14446 24998 14498 25050
rect 14510 24998 14562 25050
rect 14574 24998 14626 25050
rect 14638 24998 14690 25050
rect 7656 24896 7708 24948
rect 8208 24896 8260 24948
rect 8668 24896 8720 24948
rect 9588 24896 9640 24948
rect 13544 24896 13596 24948
rect 756 24760 808 24812
rect 6736 24828 6788 24880
rect 7012 24828 7064 24880
rect 10416 24803 10468 24812
rect 10416 24769 10425 24803
rect 10425 24769 10459 24803
rect 10459 24769 10468 24803
rect 10416 24760 10468 24769
rect 10968 24803 11020 24812
rect 10968 24769 10977 24803
rect 10977 24769 11011 24803
rect 11011 24769 11020 24803
rect 10968 24760 11020 24769
rect 4160 24692 4212 24744
rect 12164 24760 12216 24812
rect 12716 24803 12768 24812
rect 12716 24769 12723 24803
rect 12723 24769 12757 24803
rect 12757 24769 12768 24803
rect 12716 24760 12768 24769
rect 14096 24828 14148 24880
rect 15016 24828 15068 24880
rect 14280 24760 14332 24812
rect 15200 24760 15252 24812
rect 15568 24760 15620 24812
rect 5724 24624 5776 24676
rect 7472 24624 7524 24676
rect 11612 24624 11664 24676
rect 7380 24599 7432 24608
rect 7380 24565 7389 24599
rect 7389 24565 7423 24599
rect 7423 24565 7432 24599
rect 7380 24556 7432 24565
rect 7564 24556 7616 24608
rect 7748 24556 7800 24608
rect 11428 24556 11480 24608
rect 14004 24556 14056 24608
rect 2629 24454 2681 24506
rect 2693 24454 2745 24506
rect 2757 24454 2809 24506
rect 2821 24454 2873 24506
rect 2885 24454 2937 24506
rect 5987 24454 6039 24506
rect 6051 24454 6103 24506
rect 6115 24454 6167 24506
rect 6179 24454 6231 24506
rect 6243 24454 6295 24506
rect 9345 24454 9397 24506
rect 9409 24454 9461 24506
rect 9473 24454 9525 24506
rect 9537 24454 9589 24506
rect 9601 24454 9653 24506
rect 12703 24454 12755 24506
rect 12767 24454 12819 24506
rect 12831 24454 12883 24506
rect 12895 24454 12947 24506
rect 12959 24454 13011 24506
rect 5816 24352 5868 24404
rect 6276 24352 6328 24404
rect 4160 24216 4212 24268
rect 6000 24259 6052 24268
rect 6000 24225 6009 24259
rect 6009 24225 6043 24259
rect 6043 24225 6052 24259
rect 6000 24216 6052 24225
rect 7380 24352 7432 24404
rect 7472 24352 7524 24404
rect 10416 24352 10468 24404
rect 9956 24327 10008 24336
rect 9956 24293 9965 24327
rect 9965 24293 9999 24327
rect 9999 24293 10008 24327
rect 9956 24284 10008 24293
rect 4712 24191 4764 24200
rect 4712 24157 4719 24191
rect 4719 24157 4753 24191
rect 4753 24157 4764 24191
rect 4712 24148 4764 24157
rect 5448 24148 5500 24200
rect 5908 24148 5960 24200
rect 6184 24148 6236 24200
rect 6828 24191 6880 24200
rect 6828 24157 6862 24191
rect 6862 24157 6880 24191
rect 6828 24148 6880 24157
rect 9128 24148 9180 24200
rect 12164 24352 12216 24404
rect 15476 24352 15528 24404
rect 10048 24148 10100 24200
rect 10232 24080 10284 24132
rect 5540 24012 5592 24064
rect 5908 24012 5960 24064
rect 6000 24012 6052 24064
rect 6368 24012 6420 24064
rect 6736 24012 6788 24064
rect 7472 24012 7524 24064
rect 11796 24148 11848 24200
rect 10968 24080 11020 24132
rect 14096 24148 14148 24200
rect 11796 24012 11848 24064
rect 12900 24055 12952 24064
rect 12900 24021 12909 24055
rect 12909 24021 12943 24055
rect 12943 24021 12952 24055
rect 12900 24012 12952 24021
rect 13728 24123 13780 24132
rect 13728 24089 13737 24123
rect 13737 24089 13771 24123
rect 13771 24089 13780 24123
rect 13728 24080 13780 24089
rect 14188 24012 14240 24064
rect 4308 23910 4360 23962
rect 4372 23910 4424 23962
rect 4436 23910 4488 23962
rect 4500 23910 4552 23962
rect 4564 23910 4616 23962
rect 7666 23910 7718 23962
rect 7730 23910 7782 23962
rect 7794 23910 7846 23962
rect 7858 23910 7910 23962
rect 7922 23910 7974 23962
rect 11024 23910 11076 23962
rect 11088 23910 11140 23962
rect 11152 23910 11204 23962
rect 11216 23910 11268 23962
rect 11280 23910 11332 23962
rect 14382 23910 14434 23962
rect 14446 23910 14498 23962
rect 14510 23910 14562 23962
rect 14574 23910 14626 23962
rect 14638 23910 14690 23962
rect 3516 23808 3568 23860
rect 7472 23808 7524 23860
rect 9220 23851 9272 23860
rect 9220 23817 9229 23851
rect 9229 23817 9263 23851
rect 9263 23817 9272 23851
rect 9220 23808 9272 23817
rect 9680 23808 9732 23860
rect 14004 23808 14056 23860
rect 14188 23851 14240 23860
rect 14188 23817 14197 23851
rect 14197 23817 14231 23851
rect 14231 23817 14240 23851
rect 14188 23808 14240 23817
rect 10416 23740 10468 23792
rect 10784 23740 10836 23792
rect 756 23672 808 23724
rect 7564 23715 7616 23724
rect 7564 23681 7573 23715
rect 7573 23681 7607 23715
rect 7607 23681 7616 23715
rect 7564 23672 7616 23681
rect 12256 23672 12308 23724
rect 13452 23672 13504 23724
rect 5172 23604 5224 23656
rect 8300 23647 8352 23656
rect 8300 23613 8309 23647
rect 8309 23613 8343 23647
rect 8343 23613 8352 23647
rect 8300 23604 8352 23613
rect 8484 23604 8536 23656
rect 8760 23604 8812 23656
rect 9680 23604 9732 23656
rect 5080 23536 5132 23588
rect 7840 23536 7892 23588
rect 12900 23604 12952 23656
rect 13268 23647 13320 23656
rect 13268 23613 13277 23647
rect 13277 23613 13311 23647
rect 13311 23613 13320 23647
rect 13268 23604 13320 23613
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 6184 23468 6236 23520
rect 8484 23468 8536 23520
rect 10232 23468 10284 23520
rect 11060 23468 11112 23520
rect 12164 23468 12216 23520
rect 12348 23468 12400 23520
rect 2629 23366 2681 23418
rect 2693 23366 2745 23418
rect 2757 23366 2809 23418
rect 2821 23366 2873 23418
rect 2885 23366 2937 23418
rect 5987 23366 6039 23418
rect 6051 23366 6103 23418
rect 6115 23366 6167 23418
rect 6179 23366 6231 23418
rect 6243 23366 6295 23418
rect 9345 23366 9397 23418
rect 9409 23366 9461 23418
rect 9473 23366 9525 23418
rect 9537 23366 9589 23418
rect 9601 23366 9653 23418
rect 12703 23366 12755 23418
rect 12767 23366 12819 23418
rect 12831 23366 12883 23418
rect 12895 23366 12947 23418
rect 12959 23366 13011 23418
rect 2504 23264 2556 23316
rect 11612 23264 11664 23316
rect 13084 23264 13136 23316
rect 13544 23264 13596 23316
rect 8760 23196 8812 23248
rect 10324 23196 10376 23248
rect 10784 23196 10836 23248
rect 11060 23196 11112 23248
rect 7196 23128 7248 23180
rect 8300 23128 8352 23180
rect 10876 23128 10928 23180
rect 12440 23128 12492 23180
rect 756 22992 808 23044
rect 7472 22992 7524 23044
rect 8208 23060 8260 23112
rect 10508 23060 10560 23112
rect 10600 23103 10652 23112
rect 10600 23069 10609 23103
rect 10609 23069 10643 23103
rect 10643 23069 10652 23103
rect 10600 23060 10652 23069
rect 10324 22992 10376 23044
rect 11796 23103 11848 23112
rect 11796 23069 11805 23103
rect 11805 23069 11839 23103
rect 11839 23069 11848 23103
rect 11796 23060 11848 23069
rect 12348 22992 12400 23044
rect 13176 22992 13228 23044
rect 8392 22924 8444 22976
rect 9036 22924 9088 22976
rect 15200 22924 15252 22976
rect 4308 22822 4360 22874
rect 4372 22822 4424 22874
rect 4436 22822 4488 22874
rect 4500 22822 4552 22874
rect 4564 22822 4616 22874
rect 7666 22822 7718 22874
rect 7730 22822 7782 22874
rect 7794 22822 7846 22874
rect 7858 22822 7910 22874
rect 7922 22822 7974 22874
rect 11024 22822 11076 22874
rect 11088 22822 11140 22874
rect 11152 22822 11204 22874
rect 11216 22822 11268 22874
rect 11280 22822 11332 22874
rect 14382 22822 14434 22874
rect 14446 22822 14498 22874
rect 14510 22822 14562 22874
rect 14574 22822 14626 22874
rect 14638 22822 14690 22874
rect 7196 22720 7248 22772
rect 8024 22720 8076 22772
rect 8392 22720 8444 22772
rect 10784 22720 10836 22772
rect 13360 22720 13412 22772
rect 14924 22720 14976 22772
rect 5540 22584 5592 22636
rect 7196 22584 7248 22636
rect 9680 22652 9732 22704
rect 14004 22652 14056 22704
rect 8668 22584 8720 22636
rect 5816 22380 5868 22432
rect 12624 22584 12676 22636
rect 15384 22584 15436 22636
rect 12256 22516 12308 22568
rect 14924 22516 14976 22568
rect 15292 22516 15344 22568
rect 9772 22423 9824 22432
rect 9772 22389 9781 22423
rect 9781 22389 9815 22423
rect 9815 22389 9824 22423
rect 9772 22380 9824 22389
rect 10232 22380 10284 22432
rect 10600 22380 10652 22432
rect 13820 22448 13872 22500
rect 13452 22423 13504 22432
rect 13452 22389 13461 22423
rect 13461 22389 13495 22423
rect 13495 22389 13504 22423
rect 13452 22380 13504 22389
rect 2629 22278 2681 22330
rect 2693 22278 2745 22330
rect 2757 22278 2809 22330
rect 2821 22278 2873 22330
rect 2885 22278 2937 22330
rect 5987 22278 6039 22330
rect 6051 22278 6103 22330
rect 6115 22278 6167 22330
rect 6179 22278 6231 22330
rect 6243 22278 6295 22330
rect 9345 22278 9397 22330
rect 9409 22278 9461 22330
rect 9473 22278 9525 22330
rect 9537 22278 9589 22330
rect 9601 22278 9653 22330
rect 12703 22278 12755 22330
rect 12767 22278 12819 22330
rect 12831 22278 12883 22330
rect 12895 22278 12947 22330
rect 12959 22278 13011 22330
rect 9864 22176 9916 22228
rect 9772 22108 9824 22160
rect 4896 21972 4948 22024
rect 5540 22015 5592 22024
rect 5540 21981 5549 22015
rect 5549 21981 5583 22015
rect 5583 21981 5592 22015
rect 5540 21972 5592 21981
rect 5816 22015 5868 22024
rect 5816 21981 5825 22015
rect 5825 21981 5868 22015
rect 5816 21972 5868 21981
rect 7012 21972 7064 22024
rect 7104 21972 7156 22024
rect 7380 21972 7432 22024
rect 756 21904 808 21956
rect 8300 21972 8352 22024
rect 8668 21972 8720 22024
rect 9312 21972 9364 22024
rect 9772 22015 9824 22024
rect 9772 21981 9781 22015
rect 9781 21981 9815 22015
rect 9815 21981 9824 22015
rect 9772 21972 9824 21981
rect 10140 22040 10192 22092
rect 12440 22176 12492 22228
rect 13176 22176 13228 22228
rect 13268 22108 13320 22160
rect 11612 22083 11664 22092
rect 11612 22049 11621 22083
rect 11621 22049 11655 22083
rect 11655 22049 11664 22083
rect 11612 22040 11664 22049
rect 13728 22040 13780 22092
rect 7564 21904 7616 21956
rect 9128 21904 9180 21956
rect 10784 22015 10836 22024
rect 10784 21981 10818 22015
rect 10818 21981 10836 22015
rect 10784 21972 10836 21981
rect 10968 22015 11020 22024
rect 10968 21981 10977 22015
rect 10977 21981 11011 22015
rect 11011 21981 11020 22015
rect 10968 21972 11020 21981
rect 11888 21972 11940 22024
rect 11612 21904 11664 21956
rect 12256 21904 12308 21956
rect 13820 21904 13872 21956
rect 2320 21836 2372 21888
rect 4804 21836 4856 21888
rect 6368 21836 6420 21888
rect 8760 21836 8812 21888
rect 9772 21836 9824 21888
rect 10232 21836 10284 21888
rect 10784 21836 10836 21888
rect 12164 21836 12216 21888
rect 12992 21836 13044 21888
rect 13636 21836 13688 21888
rect 15384 21836 15436 21888
rect 4308 21734 4360 21786
rect 4372 21734 4424 21786
rect 4436 21734 4488 21786
rect 4500 21734 4552 21786
rect 4564 21734 4616 21786
rect 7666 21734 7718 21786
rect 7730 21734 7782 21786
rect 7794 21734 7846 21786
rect 7858 21734 7910 21786
rect 7922 21734 7974 21786
rect 11024 21734 11076 21786
rect 11088 21734 11140 21786
rect 11152 21734 11204 21786
rect 11216 21734 11268 21786
rect 11280 21734 11332 21786
rect 14382 21734 14434 21786
rect 14446 21734 14498 21786
rect 14510 21734 14562 21786
rect 14574 21734 14626 21786
rect 14638 21734 14690 21786
rect 5080 21632 5132 21684
rect 4528 21564 4580 21616
rect 756 21496 808 21548
rect 4896 21539 4948 21548
rect 4896 21505 4905 21539
rect 4905 21505 4939 21539
rect 4939 21505 4948 21539
rect 4896 21496 4948 21505
rect 5540 21564 5592 21616
rect 6828 21564 6880 21616
rect 9404 21675 9456 21684
rect 9404 21641 9413 21675
rect 9413 21641 9447 21675
rect 9447 21641 9456 21675
rect 9404 21632 9456 21641
rect 11796 21564 11848 21616
rect 13636 21632 13688 21684
rect 15476 21632 15528 21684
rect 5264 21496 5316 21548
rect 8484 21539 8536 21548
rect 8484 21505 8493 21539
rect 8493 21505 8527 21539
rect 8527 21505 8536 21539
rect 8484 21496 8536 21505
rect 8760 21539 8812 21548
rect 8760 21505 8769 21539
rect 8769 21505 8803 21539
rect 8803 21505 8812 21539
rect 8760 21496 8812 21505
rect 10692 21539 10744 21548
rect 10692 21505 10701 21539
rect 10701 21505 10735 21539
rect 10735 21505 10744 21539
rect 10692 21496 10744 21505
rect 11704 21539 11756 21548
rect 11704 21505 11713 21539
rect 11713 21505 11747 21539
rect 11747 21505 11756 21539
rect 11704 21496 11756 21505
rect 7748 21471 7800 21480
rect 7748 21437 7757 21471
rect 7757 21437 7791 21471
rect 7791 21437 7800 21471
rect 7748 21428 7800 21437
rect 7932 21428 7984 21480
rect 5908 21335 5960 21344
rect 5908 21301 5917 21335
rect 5917 21301 5951 21335
rect 5951 21301 5960 21335
rect 5908 21292 5960 21301
rect 7380 21292 7432 21344
rect 8208 21403 8260 21412
rect 8208 21369 8217 21403
rect 8217 21369 8251 21403
rect 8251 21369 8260 21403
rect 8208 21360 8260 21369
rect 8668 21292 8720 21344
rect 8944 21292 8996 21344
rect 9312 21428 9364 21480
rect 9772 21428 9824 21480
rect 10140 21471 10192 21480
rect 10140 21437 10149 21471
rect 10149 21437 10183 21471
rect 10183 21437 10192 21471
rect 10140 21428 10192 21437
rect 11060 21428 11112 21480
rect 11244 21428 11296 21480
rect 13544 21539 13596 21548
rect 13544 21505 13553 21539
rect 13553 21505 13587 21539
rect 13587 21505 13596 21539
rect 13544 21496 13596 21505
rect 10048 21292 10100 21344
rect 10140 21292 10192 21344
rect 10600 21292 10652 21344
rect 10692 21292 10744 21344
rect 11612 21360 11664 21412
rect 11796 21360 11848 21412
rect 12992 21471 13044 21480
rect 12992 21437 13001 21471
rect 13001 21437 13035 21471
rect 13035 21437 13044 21471
rect 12992 21428 13044 21437
rect 13268 21471 13320 21480
rect 13268 21437 13277 21471
rect 13277 21437 13311 21471
rect 13311 21437 13320 21471
rect 13268 21428 13320 21437
rect 13360 21471 13412 21480
rect 13360 21437 13394 21471
rect 13394 21437 13412 21471
rect 13360 21428 13412 21437
rect 15476 21428 15528 21480
rect 13084 21360 13136 21412
rect 11888 21292 11940 21344
rect 14096 21292 14148 21344
rect 2629 21190 2681 21242
rect 2693 21190 2745 21242
rect 2757 21190 2809 21242
rect 2821 21190 2873 21242
rect 2885 21190 2937 21242
rect 5987 21190 6039 21242
rect 6051 21190 6103 21242
rect 6115 21190 6167 21242
rect 6179 21190 6231 21242
rect 6243 21190 6295 21242
rect 9345 21190 9397 21242
rect 9409 21190 9461 21242
rect 9473 21190 9525 21242
rect 9537 21190 9589 21242
rect 9601 21190 9653 21242
rect 12703 21190 12755 21242
rect 12767 21190 12819 21242
rect 12831 21190 12883 21242
rect 12895 21190 12947 21242
rect 12959 21190 13011 21242
rect 3240 21131 3292 21140
rect 3240 21097 3249 21131
rect 3249 21097 3283 21131
rect 3283 21097 3292 21131
rect 3240 21088 3292 21097
rect 7288 21131 7340 21140
rect 7288 21097 7297 21131
rect 7297 21097 7331 21131
rect 7331 21097 7340 21131
rect 7288 21088 7340 21097
rect 8484 21088 8536 21140
rect 8944 21088 8996 21140
rect 9772 21088 9824 21140
rect 10876 21088 10928 21140
rect 14004 21088 14056 21140
rect 5908 20952 5960 21004
rect 3056 20927 3108 20936
rect 3056 20893 3065 20927
rect 3065 20893 3099 20927
rect 3099 20893 3108 20927
rect 3056 20884 3108 20893
rect 6368 20927 6420 20936
rect 6368 20893 6377 20927
rect 6377 20893 6411 20927
rect 6411 20893 6420 20927
rect 6368 20884 6420 20893
rect 6460 20884 6512 20936
rect 7748 20952 7800 21004
rect 11244 21020 11296 21072
rect 15016 21088 15068 21140
rect 15200 21088 15252 21140
rect 5724 20816 5776 20868
rect 5540 20748 5592 20800
rect 5908 20748 5960 20800
rect 8116 20884 8168 20936
rect 8852 20884 8904 20936
rect 9588 20884 9640 20936
rect 9772 20927 9824 20936
rect 9772 20893 9781 20927
rect 9781 20893 9815 20927
rect 9815 20893 9824 20927
rect 9772 20884 9824 20893
rect 12716 20995 12768 21004
rect 12716 20961 12725 20995
rect 12725 20961 12759 20995
rect 12759 20961 12768 20995
rect 12716 20952 12768 20961
rect 15016 20952 15068 21004
rect 6736 20859 6788 20868
rect 6736 20825 6745 20859
rect 6745 20825 6779 20859
rect 6779 20825 6788 20859
rect 6736 20816 6788 20825
rect 13360 20884 13412 20936
rect 14280 20884 14332 20936
rect 8116 20748 8168 20800
rect 8484 20748 8536 20800
rect 10232 20748 10284 20800
rect 10876 20748 10928 20800
rect 12532 20816 12584 20868
rect 14004 20816 14056 20868
rect 15292 20748 15344 20800
rect 4308 20646 4360 20698
rect 4372 20646 4424 20698
rect 4436 20646 4488 20698
rect 4500 20646 4552 20698
rect 4564 20646 4616 20698
rect 7666 20646 7718 20698
rect 7730 20646 7782 20698
rect 7794 20646 7846 20698
rect 7858 20646 7910 20698
rect 7922 20646 7974 20698
rect 11024 20646 11076 20698
rect 11088 20646 11140 20698
rect 11152 20646 11204 20698
rect 11216 20646 11268 20698
rect 11280 20646 11332 20698
rect 14382 20646 14434 20698
rect 14446 20646 14498 20698
rect 14510 20646 14562 20698
rect 14574 20646 14626 20698
rect 14638 20646 14690 20698
rect 1676 20476 1728 20528
rect 5448 20476 5500 20528
rect 7104 20476 7156 20528
rect 8208 20544 8260 20596
rect 9128 20544 9180 20596
rect 9772 20544 9824 20596
rect 11888 20544 11940 20596
rect 756 20340 808 20392
rect 5172 20408 5224 20460
rect 7932 20408 7984 20460
rect 9128 20408 9180 20460
rect 12164 20481 12216 20528
rect 12164 20476 12189 20481
rect 12189 20476 12216 20481
rect 13728 20544 13780 20596
rect 6920 20340 6972 20392
rect 7012 20383 7064 20392
rect 7012 20349 7021 20383
rect 7021 20349 7055 20383
rect 7055 20349 7064 20383
rect 7012 20340 7064 20349
rect 8760 20340 8812 20392
rect 9680 20340 9732 20392
rect 9128 20272 9180 20324
rect 8300 20204 8352 20256
rect 9036 20204 9088 20256
rect 10968 20272 11020 20324
rect 14188 20408 14240 20460
rect 11888 20383 11940 20392
rect 11888 20349 11897 20383
rect 11897 20349 11931 20383
rect 11931 20349 11940 20383
rect 11888 20340 11940 20349
rect 13268 20340 13320 20392
rect 13728 20340 13780 20392
rect 11612 20247 11664 20256
rect 11612 20213 11621 20247
rect 11621 20213 11655 20247
rect 11655 20213 11664 20247
rect 11612 20204 11664 20213
rect 12624 20204 12676 20256
rect 14188 20204 14240 20256
rect 2629 20102 2681 20154
rect 2693 20102 2745 20154
rect 2757 20102 2809 20154
rect 2821 20102 2873 20154
rect 2885 20102 2937 20154
rect 5987 20102 6039 20154
rect 6051 20102 6103 20154
rect 6115 20102 6167 20154
rect 6179 20102 6231 20154
rect 6243 20102 6295 20154
rect 9345 20102 9397 20154
rect 9409 20102 9461 20154
rect 9473 20102 9525 20154
rect 9537 20102 9589 20154
rect 9601 20102 9653 20154
rect 12703 20102 12755 20154
rect 12767 20102 12819 20154
rect 12831 20102 12883 20154
rect 12895 20102 12947 20154
rect 12959 20102 13011 20154
rect 1676 20000 1728 20052
rect 9864 20000 9916 20052
rect 11612 20000 11664 20052
rect 11980 20000 12032 20052
rect 4160 19796 4212 19848
rect 7288 19932 7340 19984
rect 7472 19932 7524 19984
rect 8944 19907 8996 19916
rect 8944 19873 8953 19907
rect 8953 19873 8987 19907
rect 8987 19873 8996 19907
rect 8944 19864 8996 19873
rect 7472 19839 7524 19848
rect 7472 19805 7481 19839
rect 7481 19805 7515 19839
rect 7515 19805 7524 19839
rect 7472 19796 7524 19805
rect 756 19728 808 19780
rect 4896 19771 4948 19780
rect 4896 19737 4930 19771
rect 4930 19737 4948 19771
rect 4896 19728 4948 19737
rect 6828 19703 6880 19712
rect 6828 19669 6837 19703
rect 6837 19669 6871 19703
rect 6871 19669 6880 19703
rect 6828 19660 6880 19669
rect 8760 19728 8812 19780
rect 8300 19660 8352 19712
rect 8852 19660 8904 19712
rect 9128 19796 9180 19848
rect 10692 19839 10744 19848
rect 10692 19805 10701 19839
rect 10701 19805 10735 19839
rect 10735 19805 10744 19839
rect 10692 19796 10744 19805
rect 10968 19839 11020 19848
rect 10968 19805 10977 19839
rect 10977 19805 11011 19839
rect 11011 19805 11020 19839
rect 10968 19796 11020 19805
rect 12624 19864 12676 19916
rect 12716 19907 12768 19916
rect 12716 19873 12725 19907
rect 12725 19873 12759 19907
rect 12759 19873 12768 19907
rect 12716 19864 12768 19873
rect 13912 20043 13964 20052
rect 13912 20009 13921 20043
rect 13921 20009 13955 20043
rect 13955 20009 13964 20043
rect 13912 20000 13964 20009
rect 13636 19864 13688 19916
rect 12072 19839 12124 19848
rect 12072 19805 12081 19839
rect 12081 19805 12115 19839
rect 12115 19805 12124 19839
rect 12072 19796 12124 19805
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 12256 19796 12308 19805
rect 12992 19839 13044 19848
rect 12992 19805 13001 19839
rect 13001 19805 13035 19839
rect 13035 19805 13044 19839
rect 12992 19796 13044 19805
rect 13268 19839 13320 19848
rect 13268 19805 13277 19839
rect 13277 19805 13311 19839
rect 13311 19805 13320 19839
rect 13268 19796 13320 19805
rect 11336 19728 11388 19780
rect 9864 19660 9916 19712
rect 9956 19703 10008 19712
rect 9956 19669 9965 19703
rect 9965 19669 9999 19703
rect 9999 19669 10008 19703
rect 9956 19660 10008 19669
rect 13820 19660 13872 19712
rect 4308 19558 4360 19610
rect 4372 19558 4424 19610
rect 4436 19558 4488 19610
rect 4500 19558 4552 19610
rect 4564 19558 4616 19610
rect 7666 19558 7718 19610
rect 7730 19558 7782 19610
rect 7794 19558 7846 19610
rect 7858 19558 7910 19610
rect 7922 19558 7974 19610
rect 11024 19558 11076 19610
rect 11088 19558 11140 19610
rect 11152 19558 11204 19610
rect 11216 19558 11268 19610
rect 11280 19558 11332 19610
rect 14382 19558 14434 19610
rect 14446 19558 14498 19610
rect 14510 19558 14562 19610
rect 14574 19558 14626 19610
rect 14638 19558 14690 19610
rect 6828 19456 6880 19508
rect 7472 19456 7524 19508
rect 11888 19456 11940 19508
rect 3700 19320 3752 19372
rect 5172 19320 5224 19372
rect 6368 19363 6420 19372
rect 6368 19329 6377 19363
rect 6377 19329 6411 19363
rect 6411 19329 6420 19363
rect 6368 19320 6420 19329
rect 6644 19363 6696 19372
rect 6644 19329 6651 19363
rect 6651 19329 6685 19363
rect 6685 19329 6696 19363
rect 6644 19320 6696 19329
rect 7012 19320 7064 19372
rect 7288 19320 7340 19372
rect 7472 19320 7524 19372
rect 10324 19388 10376 19440
rect 8944 19320 8996 19372
rect 11612 19320 11664 19372
rect 12256 19456 12308 19508
rect 12440 19388 12492 19440
rect 13268 19456 13320 19508
rect 14096 19499 14148 19508
rect 14096 19465 14105 19499
rect 14105 19465 14139 19499
rect 14139 19465 14148 19499
rect 14096 19456 14148 19465
rect 13268 19320 13320 19372
rect 13544 19320 13596 19372
rect 13636 19320 13688 19372
rect 14096 19320 14148 19372
rect 6828 19116 6880 19168
rect 7656 19252 7708 19304
rect 8760 19295 8812 19304
rect 8760 19261 8769 19295
rect 8769 19261 8803 19295
rect 8803 19261 8812 19295
rect 8760 19252 8812 19261
rect 8852 19252 8904 19304
rect 7472 19184 7524 19236
rect 7564 19116 7616 19168
rect 7748 19116 7800 19168
rect 7840 19159 7892 19168
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 8852 19116 8904 19168
rect 9588 19295 9640 19304
rect 9588 19261 9622 19295
rect 9622 19261 9640 19295
rect 9588 19252 9640 19261
rect 9772 19295 9824 19304
rect 9772 19261 9781 19295
rect 9781 19261 9815 19295
rect 9815 19261 9824 19295
rect 9772 19252 9824 19261
rect 10784 19252 10836 19304
rect 11244 19295 11296 19304
rect 11244 19261 11253 19295
rect 11253 19261 11287 19295
rect 11287 19261 11296 19295
rect 11244 19252 11296 19261
rect 12164 19252 12216 19304
rect 12440 19252 12492 19304
rect 12532 19116 12584 19168
rect 2629 19014 2681 19066
rect 2693 19014 2745 19066
rect 2757 19014 2809 19066
rect 2821 19014 2873 19066
rect 2885 19014 2937 19066
rect 5987 19014 6039 19066
rect 6051 19014 6103 19066
rect 6115 19014 6167 19066
rect 6179 19014 6231 19066
rect 6243 19014 6295 19066
rect 9345 19014 9397 19066
rect 9409 19014 9461 19066
rect 9473 19014 9525 19066
rect 9537 19014 9589 19066
rect 9601 19014 9653 19066
rect 12703 19014 12755 19066
rect 12767 19014 12819 19066
rect 12831 19014 12883 19066
rect 12895 19014 12947 19066
rect 12959 19014 13011 19066
rect 5816 18912 5868 18964
rect 6460 18912 6512 18964
rect 5908 18708 5960 18760
rect 6736 18819 6788 18828
rect 6736 18785 6745 18819
rect 6745 18785 6779 18819
rect 6779 18785 6788 18819
rect 6736 18776 6788 18785
rect 7840 18912 7892 18964
rect 8300 18912 8352 18964
rect 8576 18912 8628 18964
rect 9772 18912 9824 18964
rect 10232 18912 10284 18964
rect 7472 18844 7524 18896
rect 756 18640 808 18692
rect 6920 18708 6972 18760
rect 7012 18751 7064 18760
rect 7012 18717 7021 18751
rect 7021 18717 7055 18751
rect 7055 18717 7064 18751
rect 7012 18708 7064 18717
rect 4804 18572 4856 18624
rect 6092 18572 6144 18624
rect 6184 18615 6236 18624
rect 6184 18581 6193 18615
rect 6193 18581 6227 18615
rect 6227 18581 6236 18615
rect 6184 18572 6236 18581
rect 6368 18572 6420 18624
rect 7012 18572 7064 18624
rect 7288 18615 7340 18624
rect 7288 18581 7297 18615
rect 7297 18581 7331 18615
rect 7331 18581 7340 18615
rect 7288 18572 7340 18581
rect 14004 18912 14056 18964
rect 12348 18844 12400 18896
rect 8852 18776 8904 18828
rect 9864 18776 9916 18828
rect 12440 18751 12492 18760
rect 12440 18717 12449 18751
rect 12449 18717 12483 18751
rect 12483 18717 12492 18751
rect 12440 18708 12492 18717
rect 8208 18572 8260 18624
rect 8300 18572 8352 18624
rect 8668 18572 8720 18624
rect 13452 18708 13504 18760
rect 14372 18708 14424 18760
rect 15568 18708 15620 18760
rect 10232 18572 10284 18624
rect 10508 18572 10560 18624
rect 11520 18572 11572 18624
rect 12532 18572 12584 18624
rect 13544 18572 13596 18624
rect 4308 18470 4360 18522
rect 4372 18470 4424 18522
rect 4436 18470 4488 18522
rect 4500 18470 4552 18522
rect 4564 18470 4616 18522
rect 7666 18470 7718 18522
rect 7730 18470 7782 18522
rect 7794 18470 7846 18522
rect 7858 18470 7910 18522
rect 7922 18470 7974 18522
rect 11024 18470 11076 18522
rect 11088 18470 11140 18522
rect 11152 18470 11204 18522
rect 11216 18470 11268 18522
rect 11280 18470 11332 18522
rect 14382 18470 14434 18522
rect 14446 18470 14498 18522
rect 14510 18470 14562 18522
rect 14574 18470 14626 18522
rect 14638 18470 14690 18522
rect 5908 18411 5960 18420
rect 5908 18377 5917 18411
rect 5917 18377 5951 18411
rect 5951 18377 5960 18411
rect 5908 18368 5960 18377
rect 6736 18368 6788 18420
rect 6920 18411 6972 18420
rect 6920 18377 6929 18411
rect 6929 18377 6963 18411
rect 6963 18377 6972 18411
rect 6920 18368 6972 18377
rect 7012 18368 7064 18420
rect 3700 18300 3752 18352
rect 4988 18300 5040 18352
rect 6184 18300 6236 18352
rect 11980 18368 12032 18420
rect 15016 18368 15068 18420
rect 1492 18275 1544 18284
rect 1492 18241 1501 18275
rect 1501 18241 1535 18275
rect 1535 18241 1544 18275
rect 1492 18232 1544 18241
rect 2964 18232 3016 18284
rect 4804 18275 4856 18284
rect 4804 18241 4827 18275
rect 4827 18241 4856 18275
rect 4804 18232 4856 18241
rect 480 18164 532 18216
rect 4160 18164 4212 18216
rect 6368 18232 6420 18284
rect 7472 18232 7524 18284
rect 7288 18164 7340 18216
rect 8300 18232 8352 18284
rect 10692 18232 10744 18284
rect 9680 18164 9732 18216
rect 11704 18232 11756 18284
rect 12348 18275 12400 18284
rect 12348 18241 12357 18275
rect 12357 18241 12391 18275
rect 12391 18241 12400 18275
rect 12348 18232 12400 18241
rect 13452 18232 13504 18284
rect 13544 18275 13596 18284
rect 13544 18241 13553 18275
rect 13553 18241 13587 18275
rect 13587 18241 13596 18275
rect 13544 18232 13596 18241
rect 11796 18164 11848 18216
rect 12624 18164 12676 18216
rect 13912 18164 13964 18216
rect 4160 18028 4212 18080
rect 5632 18028 5684 18080
rect 6092 18028 6144 18080
rect 9036 18028 9088 18080
rect 10784 18071 10836 18080
rect 10784 18037 10793 18071
rect 10793 18037 10827 18071
rect 10827 18037 10836 18071
rect 10784 18028 10836 18037
rect 11152 18071 11204 18080
rect 11152 18037 11161 18071
rect 11161 18037 11195 18071
rect 11195 18037 11204 18071
rect 11152 18028 11204 18037
rect 12440 18028 12492 18080
rect 2629 17926 2681 17978
rect 2693 17926 2745 17978
rect 2757 17926 2809 17978
rect 2821 17926 2873 17978
rect 2885 17926 2937 17978
rect 5987 17926 6039 17978
rect 6051 17926 6103 17978
rect 6115 17926 6167 17978
rect 6179 17926 6231 17978
rect 6243 17926 6295 17978
rect 9345 17926 9397 17978
rect 9409 17926 9461 17978
rect 9473 17926 9525 17978
rect 9537 17926 9589 17978
rect 9601 17926 9653 17978
rect 12703 17926 12755 17978
rect 12767 17926 12819 17978
rect 12831 17926 12883 17978
rect 12895 17926 12947 17978
rect 12959 17926 13011 17978
rect 6368 17824 6420 17876
rect 8852 17824 8904 17876
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 2044 17620 2096 17672
rect 5356 17663 5408 17672
rect 3056 17552 3108 17604
rect 5356 17629 5363 17663
rect 5363 17629 5397 17663
rect 5397 17629 5408 17663
rect 5356 17620 5408 17629
rect 6460 17663 6512 17672
rect 6460 17629 6469 17663
rect 6469 17629 6503 17663
rect 6503 17629 6512 17663
rect 6460 17620 6512 17629
rect 11152 17756 11204 17808
rect 12072 17824 12124 17876
rect 12624 17824 12676 17876
rect 13084 17756 13136 17808
rect 12624 17688 12676 17740
rect 6920 17552 6972 17604
rect 10876 17620 10928 17672
rect 11428 17620 11480 17672
rect 11704 17663 11756 17672
rect 11704 17629 11713 17663
rect 11713 17629 11747 17663
rect 11747 17629 11756 17663
rect 11704 17620 11756 17629
rect 13084 17663 13136 17672
rect 13084 17629 13093 17663
rect 13093 17629 13127 17663
rect 13127 17629 13136 17663
rect 13084 17620 13136 17629
rect 13176 17620 13228 17672
rect 2412 17527 2464 17536
rect 2412 17493 2421 17527
rect 2421 17493 2455 17527
rect 2455 17493 2464 17527
rect 2412 17484 2464 17493
rect 7472 17527 7524 17536
rect 7472 17493 7481 17527
rect 7481 17493 7515 17527
rect 7515 17493 7524 17527
rect 7472 17484 7524 17493
rect 7932 17484 7984 17536
rect 8484 17484 8536 17536
rect 9680 17484 9732 17536
rect 10784 17484 10836 17536
rect 10876 17527 10928 17536
rect 10876 17493 10885 17527
rect 10885 17493 10919 17527
rect 10919 17493 10928 17527
rect 10876 17484 10928 17493
rect 11428 17484 11480 17536
rect 11704 17484 11756 17536
rect 4308 17382 4360 17434
rect 4372 17382 4424 17434
rect 4436 17382 4488 17434
rect 4500 17382 4552 17434
rect 4564 17382 4616 17434
rect 7666 17382 7718 17434
rect 7730 17382 7782 17434
rect 7794 17382 7846 17434
rect 7858 17382 7910 17434
rect 7922 17382 7974 17434
rect 11024 17382 11076 17434
rect 11088 17382 11140 17434
rect 11152 17382 11204 17434
rect 11216 17382 11268 17434
rect 11280 17382 11332 17434
rect 14382 17382 14434 17434
rect 14446 17382 14498 17434
rect 14510 17382 14562 17434
rect 14574 17382 14626 17434
rect 14638 17382 14690 17434
rect 2412 17280 2464 17332
rect 7840 17280 7892 17332
rect 8484 17280 8536 17332
rect 8668 17323 8720 17332
rect 8668 17289 8677 17323
rect 8677 17289 8711 17323
rect 8711 17289 8720 17323
rect 8668 17280 8720 17289
rect 8852 17280 8904 17332
rect 9772 17280 9824 17332
rect 756 17144 808 17196
rect 1860 17076 1912 17128
rect 2136 17076 2188 17128
rect 7196 17144 7248 17196
rect 7840 17187 7892 17196
rect 7840 17153 7874 17187
rect 7874 17153 7892 17187
rect 7840 17144 7892 17153
rect 5264 17076 5316 17128
rect 1492 16940 1544 16992
rect 7104 17076 7156 17128
rect 7472 17119 7524 17128
rect 7472 17085 7481 17119
rect 7481 17085 7515 17119
rect 7515 17085 7524 17119
rect 7472 17076 7524 17085
rect 7380 17008 7432 17060
rect 8024 17119 8076 17128
rect 8024 17085 8033 17119
rect 8033 17085 8067 17119
rect 8067 17085 8076 17119
rect 8024 17076 8076 17085
rect 8392 17076 8444 17128
rect 9588 17212 9640 17264
rect 9680 17212 9732 17264
rect 11336 17280 11388 17332
rect 13728 17280 13780 17332
rect 8668 17144 8720 17196
rect 10416 17144 10468 17196
rect 10508 17187 10560 17196
rect 10508 17153 10517 17187
rect 10517 17153 10551 17187
rect 10551 17153 10560 17187
rect 10508 17144 10560 17153
rect 10048 17076 10100 17128
rect 9680 16940 9732 16992
rect 9772 16983 9824 16992
rect 9772 16949 9781 16983
rect 9781 16949 9815 16983
rect 9815 16949 9824 16983
rect 9772 16940 9824 16949
rect 11152 17144 11204 17196
rect 11336 17144 11388 17196
rect 11428 17144 11480 17196
rect 13544 17212 13596 17264
rect 14004 17187 14056 17196
rect 14004 17153 14013 17187
rect 14013 17153 14047 17187
rect 14047 17153 14056 17187
rect 14004 17144 14056 17153
rect 10968 17076 11020 17128
rect 12072 17076 12124 17128
rect 12348 17119 12400 17128
rect 12348 17085 12357 17119
rect 12357 17085 12391 17119
rect 12391 17085 12400 17119
rect 12348 17076 12400 17085
rect 12532 17119 12584 17128
rect 12532 17085 12541 17119
rect 12541 17085 12575 17119
rect 12575 17085 12584 17119
rect 12532 17076 12584 17085
rect 13912 17076 13964 17128
rect 15568 17076 15620 17128
rect 11060 16983 11112 16992
rect 11060 16949 11069 16983
rect 11069 16949 11103 16983
rect 11103 16949 11112 16983
rect 11060 16940 11112 16949
rect 11244 16940 11296 16992
rect 12256 16940 12308 16992
rect 12532 16940 12584 16992
rect 12992 16940 13044 16992
rect 13452 16940 13504 16992
rect 2629 16838 2681 16890
rect 2693 16838 2745 16890
rect 2757 16838 2809 16890
rect 2821 16838 2873 16890
rect 2885 16838 2937 16890
rect 5987 16838 6039 16890
rect 6051 16838 6103 16890
rect 6115 16838 6167 16890
rect 6179 16838 6231 16890
rect 6243 16838 6295 16890
rect 9345 16838 9397 16890
rect 9409 16838 9461 16890
rect 9473 16838 9525 16890
rect 9537 16838 9589 16890
rect 9601 16838 9653 16890
rect 12703 16838 12755 16890
rect 12767 16838 12819 16890
rect 12831 16838 12883 16890
rect 12895 16838 12947 16890
rect 12959 16838 13011 16890
rect 6460 16600 6512 16652
rect 8024 16736 8076 16788
rect 8484 16736 8536 16788
rect 3424 16532 3476 16584
rect 4896 16532 4948 16584
rect 756 16464 808 16516
rect 3516 16464 3568 16516
rect 8852 16600 8904 16652
rect 9220 16643 9272 16652
rect 9220 16609 9229 16643
rect 9229 16609 9263 16643
rect 9263 16609 9272 16643
rect 9220 16600 9272 16609
rect 9496 16600 9548 16652
rect 9772 16736 9824 16788
rect 10876 16668 10928 16720
rect 11612 16736 11664 16788
rect 11980 16736 12032 16788
rect 12716 16736 12768 16788
rect 11244 16668 11296 16720
rect 12532 16668 12584 16720
rect 10600 16600 10652 16652
rect 12164 16600 12216 16652
rect 12716 16643 12768 16652
rect 12716 16609 12725 16643
rect 12725 16609 12759 16643
rect 12759 16609 12768 16643
rect 12716 16600 12768 16609
rect 13176 16736 13228 16788
rect 13820 16736 13872 16788
rect 13452 16600 13504 16652
rect 9588 16532 9640 16584
rect 10140 16575 10192 16584
rect 10140 16541 10149 16575
rect 10149 16541 10183 16575
rect 10183 16541 10192 16575
rect 10140 16532 10192 16541
rect 10416 16575 10468 16584
rect 10416 16541 10425 16575
rect 10425 16541 10459 16575
rect 10459 16541 10468 16575
rect 10416 16532 10468 16541
rect 11152 16575 11204 16584
rect 11152 16541 11161 16575
rect 11161 16541 11195 16575
rect 11195 16541 11204 16575
rect 11152 16532 11204 16541
rect 11888 16532 11940 16584
rect 8392 16464 8444 16516
rect 8668 16396 8720 16448
rect 10232 16396 10284 16448
rect 11428 16396 11480 16448
rect 11612 16439 11664 16448
rect 11612 16405 11621 16439
rect 11621 16405 11655 16439
rect 11655 16405 11664 16439
rect 11612 16396 11664 16405
rect 12164 16464 12216 16516
rect 13176 16532 13228 16584
rect 13820 16396 13872 16448
rect 4308 16294 4360 16346
rect 4372 16294 4424 16346
rect 4436 16294 4488 16346
rect 4500 16294 4552 16346
rect 4564 16294 4616 16346
rect 7666 16294 7718 16346
rect 7730 16294 7782 16346
rect 7794 16294 7846 16346
rect 7858 16294 7910 16346
rect 7922 16294 7974 16346
rect 11024 16294 11076 16346
rect 11088 16294 11140 16346
rect 11152 16294 11204 16346
rect 11216 16294 11268 16346
rect 11280 16294 11332 16346
rect 14382 16294 14434 16346
rect 14446 16294 14498 16346
rect 14510 16294 14562 16346
rect 14574 16294 14626 16346
rect 14638 16294 14690 16346
rect 1952 16192 2004 16244
rect 10416 16192 10468 16244
rect 12716 16192 12768 16244
rect 15292 16192 15344 16244
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 7380 16124 7432 16176
rect 8300 16124 8352 16176
rect 6460 16056 6512 16108
rect 7012 16056 7064 16108
rect 2412 15895 2464 15904
rect 2412 15861 2421 15895
rect 2421 15861 2455 15895
rect 2455 15861 2464 15895
rect 2412 15852 2464 15861
rect 2504 15852 2556 15904
rect 5540 15852 5592 15904
rect 9772 16056 9824 16108
rect 10416 16056 10468 16108
rect 11060 16124 11112 16176
rect 11796 16124 11848 16176
rect 15016 16124 15068 16176
rect 15476 16124 15528 16176
rect 15568 16124 15620 16176
rect 12808 16056 12860 16108
rect 8392 15988 8444 16040
rect 11612 15988 11664 16040
rect 11796 16031 11848 16040
rect 11796 15997 11805 16031
rect 11805 15997 11839 16031
rect 11839 15997 11848 16031
rect 11796 15988 11848 15997
rect 15384 15988 15436 16040
rect 15568 15920 15620 15972
rect 8392 15852 8444 15904
rect 10140 15852 10192 15904
rect 2629 15750 2681 15802
rect 2693 15750 2745 15802
rect 2757 15750 2809 15802
rect 2821 15750 2873 15802
rect 2885 15750 2937 15802
rect 5987 15750 6039 15802
rect 6051 15750 6103 15802
rect 6115 15750 6167 15802
rect 6179 15750 6231 15802
rect 6243 15750 6295 15802
rect 9345 15750 9397 15802
rect 9409 15750 9461 15802
rect 9473 15750 9525 15802
rect 9537 15750 9589 15802
rect 9601 15750 9653 15802
rect 12703 15750 12755 15802
rect 12767 15750 12819 15802
rect 12831 15750 12883 15802
rect 12895 15750 12947 15802
rect 12959 15750 13011 15802
rect 6920 15648 6972 15700
rect 7196 15648 7248 15700
rect 7380 15580 7432 15632
rect 9956 15580 10008 15632
rect 6460 15512 6512 15564
rect 11060 15648 11112 15700
rect 11704 15648 11756 15700
rect 13912 15648 13964 15700
rect 11060 15555 11112 15564
rect 11060 15521 11069 15555
rect 11069 15521 11103 15555
rect 11103 15521 11112 15555
rect 11060 15512 11112 15521
rect 11520 15512 11572 15564
rect 11888 15580 11940 15632
rect 7380 15444 7432 15496
rect 8852 15444 8904 15496
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 11152 15487 11204 15496
rect 11152 15453 11186 15487
rect 11186 15453 11204 15487
rect 12072 15555 12124 15564
rect 12072 15521 12081 15555
rect 12081 15521 12115 15555
rect 12115 15521 12124 15555
rect 12072 15512 12124 15521
rect 11152 15444 11204 15453
rect 14648 15444 14700 15496
rect 756 15376 808 15428
rect 5632 15376 5684 15428
rect 9312 15308 9364 15360
rect 10232 15308 10284 15360
rect 11152 15308 11204 15360
rect 12164 15308 12216 15360
rect 12992 15308 13044 15360
rect 13820 15351 13872 15360
rect 13820 15317 13829 15351
rect 13829 15317 13863 15351
rect 13863 15317 13872 15351
rect 13820 15308 13872 15317
rect 4308 15206 4360 15258
rect 4372 15206 4424 15258
rect 4436 15206 4488 15258
rect 4500 15206 4552 15258
rect 4564 15206 4616 15258
rect 7666 15206 7718 15258
rect 7730 15206 7782 15258
rect 7794 15206 7846 15258
rect 7858 15206 7910 15258
rect 7922 15206 7974 15258
rect 11024 15206 11076 15258
rect 11088 15206 11140 15258
rect 11152 15206 11204 15258
rect 11216 15206 11268 15258
rect 11280 15206 11332 15258
rect 14382 15206 14434 15258
rect 14446 15206 14498 15258
rect 14510 15206 14562 15258
rect 14574 15206 14626 15258
rect 14638 15206 14690 15258
rect 1308 15104 1360 15156
rect 1492 15079 1544 15088
rect 1492 15045 1501 15079
rect 1501 15045 1535 15079
rect 1535 15045 1544 15079
rect 1492 15036 1544 15045
rect 2412 15036 2464 15088
rect 1584 14900 1636 14952
rect 5908 15104 5960 15156
rect 6736 15104 6788 15156
rect 7104 15104 7156 15156
rect 10324 15104 10376 15156
rect 10048 15036 10100 15088
rect 15200 15104 15252 15156
rect 7104 14968 7156 15020
rect 8116 15011 8168 15020
rect 8116 14977 8125 15011
rect 8125 14977 8159 15011
rect 8159 14977 8168 15011
rect 8116 14968 8168 14977
rect 9036 15011 9088 15020
rect 9036 14977 9045 15011
rect 9045 14977 9079 15011
rect 9079 14977 9088 15011
rect 9036 14968 9088 14977
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 10324 15011 10376 15020
rect 10324 14977 10333 15011
rect 10333 14977 10376 15011
rect 10324 14968 10376 14977
rect 6368 14943 6420 14952
rect 848 14764 900 14816
rect 1952 14807 2004 14816
rect 1952 14773 1961 14807
rect 1961 14773 1995 14807
rect 1995 14773 2004 14807
rect 1952 14764 2004 14773
rect 6368 14909 6377 14943
rect 6377 14909 6411 14943
rect 6411 14909 6420 14943
rect 6368 14900 6420 14909
rect 8300 14943 8352 14952
rect 8300 14909 8309 14943
rect 8309 14909 8343 14943
rect 8343 14909 8352 14943
rect 8300 14900 8352 14909
rect 8392 14900 8444 14952
rect 5908 14807 5960 14816
rect 5908 14773 5917 14807
rect 5917 14773 5951 14807
rect 5951 14773 5960 14807
rect 5908 14764 5960 14773
rect 6828 14764 6880 14816
rect 8668 14832 8720 14884
rect 9680 14900 9732 14952
rect 12348 15036 12400 15088
rect 11704 15011 11756 15020
rect 11704 14977 11713 15011
rect 11713 14977 11747 15011
rect 11747 14977 11756 15011
rect 11704 14968 11756 14977
rect 12072 15011 12124 15020
rect 12072 14977 12081 15011
rect 12081 14977 12115 15011
rect 12115 14977 12124 15011
rect 12072 14968 12124 14977
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 11060 14900 11112 14952
rect 12440 14900 12492 14952
rect 12992 14943 13044 14952
rect 12992 14909 13001 14943
rect 13001 14909 13035 14943
rect 13035 14909 13044 14943
rect 12992 14900 13044 14909
rect 13360 14943 13412 14952
rect 13360 14909 13394 14943
rect 13394 14909 13412 14943
rect 13360 14900 13412 14909
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 7380 14807 7432 14816
rect 7380 14773 7389 14807
rect 7389 14773 7423 14807
rect 7423 14773 7432 14807
rect 7380 14764 7432 14773
rect 11336 14764 11388 14816
rect 12072 14764 12124 14816
rect 14372 14764 14424 14816
rect 2629 14662 2681 14714
rect 2693 14662 2745 14714
rect 2757 14662 2809 14714
rect 2821 14662 2873 14714
rect 2885 14662 2937 14714
rect 5987 14662 6039 14714
rect 6051 14662 6103 14714
rect 6115 14662 6167 14714
rect 6179 14662 6231 14714
rect 6243 14662 6295 14714
rect 9345 14662 9397 14714
rect 9409 14662 9461 14714
rect 9473 14662 9525 14714
rect 9537 14662 9589 14714
rect 9601 14662 9653 14714
rect 12703 14662 12755 14714
rect 12767 14662 12819 14714
rect 12831 14662 12883 14714
rect 12895 14662 12947 14714
rect 12959 14662 13011 14714
rect 5908 14560 5960 14612
rect 1400 14467 1452 14476
rect 1400 14433 1409 14467
rect 1409 14433 1443 14467
rect 1443 14433 1452 14467
rect 1400 14424 1452 14433
rect 7104 14560 7156 14612
rect 7380 14560 7432 14612
rect 8024 14560 8076 14612
rect 8576 14560 8628 14612
rect 10508 14560 10560 14612
rect 6828 14467 6880 14476
rect 6828 14433 6862 14467
rect 6862 14433 6880 14467
rect 6828 14424 6880 14433
rect 7564 14492 7616 14544
rect 7932 14492 7984 14544
rect 9772 14492 9824 14544
rect 1308 14356 1360 14408
rect 6000 14399 6052 14408
rect 6000 14365 6009 14399
rect 6009 14365 6043 14399
rect 6043 14365 6052 14399
rect 6000 14356 6052 14365
rect 6736 14399 6788 14408
rect 6736 14365 6745 14399
rect 6745 14365 6779 14399
rect 6779 14365 6788 14399
rect 6736 14356 6788 14365
rect 9036 14424 9088 14476
rect 12164 14492 12216 14544
rect 13544 14603 13596 14612
rect 13544 14569 13553 14603
rect 13553 14569 13587 14603
rect 13587 14569 13596 14603
rect 13544 14560 13596 14569
rect 10324 14467 10376 14476
rect 10324 14433 10333 14467
rect 10333 14433 10367 14467
rect 10367 14433 10376 14467
rect 10324 14424 10376 14433
rect 10784 14467 10836 14476
rect 10784 14433 10793 14467
rect 10793 14433 10827 14467
rect 10827 14433 10836 14467
rect 10784 14424 10836 14433
rect 11060 14467 11112 14476
rect 11060 14433 11087 14467
rect 11087 14433 11112 14467
rect 11060 14424 11112 14433
rect 12440 14424 12492 14476
rect 13820 14424 13872 14476
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 6736 14220 6788 14272
rect 7656 14220 7708 14272
rect 10508 14356 10560 14408
rect 11244 14356 11296 14408
rect 11336 14399 11388 14408
rect 11336 14365 11345 14399
rect 11345 14365 11379 14399
rect 11379 14365 11388 14399
rect 11336 14356 11388 14365
rect 8392 14288 8444 14340
rect 8576 14288 8628 14340
rect 9864 14288 9916 14340
rect 11888 14288 11940 14340
rect 12164 14288 12216 14340
rect 12900 14356 12952 14408
rect 15016 14288 15068 14340
rect 10968 14220 11020 14272
rect 4308 14118 4360 14170
rect 4372 14118 4424 14170
rect 4436 14118 4488 14170
rect 4500 14118 4552 14170
rect 4564 14118 4616 14170
rect 7666 14118 7718 14170
rect 7730 14118 7782 14170
rect 7794 14118 7846 14170
rect 7858 14118 7910 14170
rect 7922 14118 7974 14170
rect 11024 14118 11076 14170
rect 11088 14118 11140 14170
rect 11152 14118 11204 14170
rect 11216 14118 11268 14170
rect 11280 14118 11332 14170
rect 14382 14118 14434 14170
rect 14446 14118 14498 14170
rect 14510 14118 14562 14170
rect 14574 14118 14626 14170
rect 14638 14118 14690 14170
rect 1952 14016 2004 14068
rect 7288 14016 7340 14068
rect 9680 13948 9732 14000
rect 1676 13880 1728 13932
rect 1860 13880 1912 13932
rect 5080 13880 5132 13932
rect 7564 13880 7616 13932
rect 5080 13744 5132 13796
rect 5448 13744 5500 13796
rect 1584 13719 1636 13728
rect 1584 13685 1593 13719
rect 1593 13685 1627 13719
rect 1627 13685 1636 13719
rect 1584 13676 1636 13685
rect 7840 13855 7892 13864
rect 7840 13821 7849 13855
rect 7849 13821 7883 13855
rect 7883 13821 7892 13855
rect 7840 13812 7892 13821
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 9864 14016 9916 14068
rect 10784 14016 10836 14068
rect 13360 14016 13412 14068
rect 9864 13880 9916 13932
rect 10692 13880 10744 13932
rect 11796 13923 11848 13932
rect 11796 13889 11803 13923
rect 11803 13889 11837 13923
rect 11837 13889 11848 13923
rect 12348 13948 12400 14000
rect 12440 13948 12492 14000
rect 13912 13991 13964 14000
rect 13912 13957 13921 13991
rect 13921 13957 13955 13991
rect 13955 13957 13964 13991
rect 13912 13948 13964 13957
rect 11796 13880 11848 13889
rect 7656 13744 7708 13796
rect 8300 13812 8352 13864
rect 9496 13855 9548 13864
rect 9496 13821 9505 13855
rect 9505 13821 9539 13855
rect 9539 13821 9548 13855
rect 9496 13812 9548 13821
rect 11520 13855 11572 13864
rect 11520 13821 11529 13855
rect 11529 13821 11563 13855
rect 11563 13821 11572 13855
rect 11520 13812 11572 13821
rect 13084 13812 13136 13864
rect 13360 13880 13412 13932
rect 11796 13676 11848 13728
rect 12440 13676 12492 13728
rect 13360 13676 13412 13728
rect 2629 13574 2681 13626
rect 2693 13574 2745 13626
rect 2757 13574 2809 13626
rect 2821 13574 2873 13626
rect 2885 13574 2937 13626
rect 5987 13574 6039 13626
rect 6051 13574 6103 13626
rect 6115 13574 6167 13626
rect 6179 13574 6231 13626
rect 6243 13574 6295 13626
rect 9345 13574 9397 13626
rect 9409 13574 9461 13626
rect 9473 13574 9525 13626
rect 9537 13574 9589 13626
rect 9601 13574 9653 13626
rect 12703 13574 12755 13626
rect 12767 13574 12819 13626
rect 12831 13574 12883 13626
rect 12895 13574 12947 13626
rect 12959 13574 13011 13626
rect 6368 13472 6420 13524
rect 2412 13268 2464 13320
rect 7840 13472 7892 13524
rect 8300 13472 8352 13524
rect 8852 13472 8904 13524
rect 9404 13472 9456 13524
rect 8944 13379 8996 13388
rect 8944 13345 8953 13379
rect 8953 13345 8987 13379
rect 8987 13345 8996 13379
rect 8944 13336 8996 13345
rect 10140 13472 10192 13524
rect 10324 13472 10376 13524
rect 10876 13472 10928 13524
rect 7104 13268 7156 13320
rect 7656 13268 7708 13320
rect 8208 13268 8260 13320
rect 8484 13268 8536 13320
rect 848 13132 900 13184
rect 6552 13200 6604 13252
rect 6828 13200 6880 13252
rect 8944 13200 8996 13252
rect 9864 13311 9916 13320
rect 9864 13277 9873 13311
rect 9873 13277 9907 13311
rect 9907 13277 9916 13311
rect 9864 13268 9916 13277
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 11888 13379 11940 13388
rect 11888 13345 11897 13379
rect 11897 13345 11931 13379
rect 11931 13345 11940 13379
rect 11888 13336 11940 13345
rect 13452 13472 13504 13524
rect 12348 13336 12400 13388
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 13176 13404 13228 13456
rect 13268 13404 13320 13456
rect 15292 13472 15344 13524
rect 11244 13311 11296 13320
rect 11244 13277 11253 13311
rect 11253 13277 11287 13311
rect 11287 13277 11296 13311
rect 11244 13268 11296 13277
rect 14372 13268 14424 13320
rect 10692 13200 10744 13252
rect 10784 13200 10836 13252
rect 13728 13243 13780 13252
rect 13728 13209 13737 13243
rect 13737 13209 13771 13243
rect 13771 13209 13780 13243
rect 13728 13200 13780 13209
rect 4068 13132 4120 13184
rect 8576 13132 8628 13184
rect 8668 13132 8720 13184
rect 11428 13132 11480 13184
rect 4308 13030 4360 13082
rect 4372 13030 4424 13082
rect 4436 13030 4488 13082
rect 4500 13030 4552 13082
rect 4564 13030 4616 13082
rect 7666 13030 7718 13082
rect 7730 13030 7782 13082
rect 7794 13030 7846 13082
rect 7858 13030 7910 13082
rect 7922 13030 7974 13082
rect 11024 13030 11076 13082
rect 11088 13030 11140 13082
rect 11152 13030 11204 13082
rect 11216 13030 11268 13082
rect 11280 13030 11332 13082
rect 14382 13030 14434 13082
rect 14446 13030 14498 13082
rect 14510 13030 14562 13082
rect 14574 13030 14626 13082
rect 14638 13030 14690 13082
rect 1676 12928 1728 12980
rect 3792 12928 3844 12980
rect 6920 12928 6972 12980
rect 7288 12928 7340 12980
rect 8392 12928 8444 12980
rect 8576 12928 8628 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 7104 12860 7156 12912
rect 8852 12860 8904 12912
rect 9680 12860 9732 12912
rect 10140 12928 10192 12980
rect 10784 12928 10836 12980
rect 7288 12835 7340 12844
rect 7288 12801 7295 12835
rect 7295 12801 7329 12835
rect 7329 12801 7340 12835
rect 7288 12792 7340 12801
rect 8668 12792 8720 12844
rect 10416 12792 10468 12844
rect 14004 12928 14056 12980
rect 15476 12928 15528 12980
rect 12716 12792 12768 12844
rect 8852 12767 8904 12776
rect 8852 12733 8861 12767
rect 8861 12733 8895 12767
rect 8895 12733 8904 12767
rect 8852 12724 8904 12733
rect 9864 12656 9916 12708
rect 10048 12656 10100 12708
rect 11980 12724 12032 12776
rect 12164 12656 12216 12708
rect 2412 12631 2464 12640
rect 2412 12597 2421 12631
rect 2421 12597 2455 12631
rect 2455 12597 2464 12631
rect 2412 12588 2464 12597
rect 5356 12588 5408 12640
rect 8668 12588 8720 12640
rect 8852 12588 8904 12640
rect 8944 12588 8996 12640
rect 11336 12588 11388 12640
rect 11796 12588 11848 12640
rect 12624 12724 12676 12776
rect 13452 12724 13504 12776
rect 13544 12767 13596 12776
rect 13544 12733 13553 12767
rect 13553 12733 13587 12767
rect 13587 12733 13596 12767
rect 13544 12724 13596 12733
rect 12992 12699 13044 12708
rect 12992 12665 13001 12699
rect 13001 12665 13035 12699
rect 13035 12665 13044 12699
rect 12992 12656 13044 12665
rect 12440 12588 12492 12640
rect 12624 12588 12676 12640
rect 2629 12486 2681 12538
rect 2693 12486 2745 12538
rect 2757 12486 2809 12538
rect 2821 12486 2873 12538
rect 2885 12486 2937 12538
rect 5987 12486 6039 12538
rect 6051 12486 6103 12538
rect 6115 12486 6167 12538
rect 6179 12486 6231 12538
rect 6243 12486 6295 12538
rect 9345 12486 9397 12538
rect 9409 12486 9461 12538
rect 9473 12486 9525 12538
rect 9537 12486 9589 12538
rect 9601 12486 9653 12538
rect 12703 12486 12755 12538
rect 12767 12486 12819 12538
rect 12831 12486 12883 12538
rect 12895 12486 12947 12538
rect 12959 12486 13011 12538
rect 4712 12384 4764 12436
rect 7196 12384 7248 12436
rect 11888 12384 11940 12436
rect 13084 12384 13136 12436
rect 6828 12316 6880 12368
rect 7104 12291 7156 12300
rect 7104 12257 7113 12291
rect 7113 12257 7147 12291
rect 7147 12257 7156 12291
rect 7104 12248 7156 12257
rect 9680 12248 9732 12300
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 2412 12180 2464 12232
rect 5632 12180 5684 12232
rect 848 12044 900 12096
rect 4712 12112 4764 12164
rect 7012 12180 7064 12232
rect 7380 12223 7432 12232
rect 7380 12189 7387 12223
rect 7387 12189 7421 12223
rect 7421 12189 7432 12223
rect 7380 12180 7432 12189
rect 9220 12180 9272 12232
rect 5632 12044 5684 12096
rect 7196 12044 7248 12096
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 12072 12248 12124 12300
rect 10140 12112 10192 12164
rect 11612 12112 11664 12164
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 11980 12112 12032 12164
rect 12164 12112 12216 12164
rect 13452 12044 13504 12096
rect 13636 12044 13688 12096
rect 4308 11942 4360 11994
rect 4372 11942 4424 11994
rect 4436 11942 4488 11994
rect 4500 11942 4552 11994
rect 4564 11942 4616 11994
rect 7666 11942 7718 11994
rect 7730 11942 7782 11994
rect 7794 11942 7846 11994
rect 7858 11942 7910 11994
rect 7922 11942 7974 11994
rect 11024 11942 11076 11994
rect 11088 11942 11140 11994
rect 11152 11942 11204 11994
rect 11216 11942 11268 11994
rect 11280 11942 11332 11994
rect 14382 11942 14434 11994
rect 14446 11942 14498 11994
rect 14510 11942 14562 11994
rect 14574 11942 14626 11994
rect 14638 11942 14690 11994
rect 5816 11840 5868 11892
rect 10140 11840 10192 11892
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 4712 11704 4764 11756
rect 5908 11772 5960 11824
rect 7748 11772 7800 11824
rect 5540 11704 5592 11756
rect 6920 11704 6972 11756
rect 7288 11704 7340 11756
rect 8024 11772 8076 11824
rect 8208 11772 8260 11824
rect 7104 11636 7156 11688
rect 12348 11840 12400 11892
rect 13544 11840 13596 11892
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 12072 11772 12124 11824
rect 11796 11704 11848 11756
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 848 11500 900 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 7288 11500 7340 11552
rect 11888 11568 11940 11620
rect 12348 11568 12400 11620
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 11428 11500 11480 11552
rect 2629 11398 2681 11450
rect 2693 11398 2745 11450
rect 2757 11398 2809 11450
rect 2821 11398 2873 11450
rect 2885 11398 2937 11450
rect 5987 11398 6039 11450
rect 6051 11398 6103 11450
rect 6115 11398 6167 11450
rect 6179 11398 6231 11450
rect 6243 11398 6295 11450
rect 9345 11398 9397 11450
rect 9409 11398 9461 11450
rect 9473 11398 9525 11450
rect 9537 11398 9589 11450
rect 9601 11398 9653 11450
rect 12703 11398 12755 11450
rect 12767 11398 12819 11450
rect 12831 11398 12883 11450
rect 12895 11398 12947 11450
rect 12959 11398 13011 11450
rect 6644 11296 6696 11348
rect 10508 11296 10560 11348
rect 11520 11296 11572 11348
rect 5724 11160 5776 11212
rect 6092 11160 6144 11212
rect 7748 11228 7800 11280
rect 8484 11228 8536 11280
rect 10692 11228 10744 11280
rect 8392 11160 8444 11212
rect 13176 11296 13228 11348
rect 5816 11024 5868 11076
rect 6920 11135 6972 11144
rect 6920 11101 6929 11135
rect 6929 11101 6963 11135
rect 6963 11101 6972 11135
rect 6920 11092 6972 11101
rect 7104 11092 7156 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 8852 11092 8904 11144
rect 9036 11092 9088 11144
rect 2136 10956 2188 11008
rect 10508 11135 10560 11144
rect 10508 11101 10517 11135
rect 10517 11101 10551 11135
rect 10551 11101 10560 11135
rect 10508 11092 10560 11101
rect 10876 11092 10928 11144
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 11612 11092 11664 11144
rect 11704 11135 11756 11144
rect 11704 11101 11713 11135
rect 11713 11101 11747 11135
rect 11747 11101 11756 11135
rect 11704 11092 11756 11101
rect 12716 11105 12768 11144
rect 12716 11092 12741 11105
rect 12741 11092 12768 11105
rect 12900 10956 12952 11008
rect 4308 10854 4360 10906
rect 4372 10854 4424 10906
rect 4436 10854 4488 10906
rect 4500 10854 4552 10906
rect 4564 10854 4616 10906
rect 7666 10854 7718 10906
rect 7730 10854 7782 10906
rect 7794 10854 7846 10906
rect 7858 10854 7910 10906
rect 7922 10854 7974 10906
rect 11024 10854 11076 10906
rect 11088 10854 11140 10906
rect 11152 10854 11204 10906
rect 11216 10854 11268 10906
rect 11280 10854 11332 10906
rect 14382 10854 14434 10906
rect 14446 10854 14498 10906
rect 14510 10854 14562 10906
rect 14574 10854 14626 10906
rect 14638 10854 14690 10906
rect 1492 10752 1544 10804
rect 6920 10752 6972 10804
rect 7564 10752 7616 10804
rect 8208 10752 8260 10804
rect 10324 10752 10376 10804
rect 10600 10752 10652 10804
rect 10692 10752 10744 10804
rect 11428 10752 11480 10804
rect 11888 10752 11940 10804
rect 2044 10616 2096 10668
rect 2136 10659 2188 10668
rect 2136 10625 2145 10659
rect 2145 10625 2179 10659
rect 2179 10625 2188 10659
rect 2136 10616 2188 10625
rect 5632 10616 5684 10668
rect 6368 10659 6420 10668
rect 6368 10625 6377 10659
rect 6377 10625 6411 10659
rect 6411 10625 6420 10659
rect 6368 10616 6420 10625
rect 8392 10727 8444 10736
rect 8392 10693 8401 10727
rect 8401 10693 8435 10727
rect 8435 10693 8444 10727
rect 8392 10684 8444 10693
rect 8668 10684 8720 10736
rect 6552 10548 6604 10600
rect 7104 10616 7156 10668
rect 9680 10616 9732 10668
rect 848 10412 900 10464
rect 5724 10412 5776 10464
rect 6736 10455 6788 10464
rect 6736 10421 6745 10455
rect 6745 10421 6779 10455
rect 6779 10421 6788 10455
rect 6736 10412 6788 10421
rect 6920 10412 6972 10464
rect 7656 10412 7708 10464
rect 8116 10412 8168 10464
rect 9404 10455 9456 10464
rect 9404 10421 9413 10455
rect 9413 10421 9447 10455
rect 9447 10421 9456 10455
rect 9404 10412 9456 10421
rect 12256 10795 12308 10804
rect 12256 10761 12265 10795
rect 12265 10761 12299 10795
rect 12299 10761 12308 10795
rect 12256 10752 12308 10761
rect 12348 10752 12400 10804
rect 13084 10752 13136 10804
rect 14280 10752 14332 10804
rect 9864 10548 9916 10600
rect 11060 10480 11112 10532
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 11888 10616 11940 10668
rect 12072 10659 12124 10668
rect 12072 10625 12081 10659
rect 12081 10625 12115 10659
rect 12115 10625 12124 10659
rect 12072 10616 12124 10625
rect 13268 10659 13320 10668
rect 13268 10625 13277 10659
rect 13277 10625 13311 10659
rect 13311 10625 13320 10659
rect 13268 10616 13320 10625
rect 13360 10659 13412 10668
rect 13360 10625 13394 10659
rect 13394 10625 13412 10659
rect 13360 10616 13412 10625
rect 12440 10548 12492 10600
rect 12900 10548 12952 10600
rect 13544 10591 13596 10600
rect 13544 10557 13553 10591
rect 13553 10557 13587 10591
rect 13587 10557 13596 10591
rect 13544 10548 13596 10557
rect 10784 10412 10836 10464
rect 12532 10412 12584 10464
rect 14004 10412 14056 10464
rect 2629 10310 2681 10362
rect 2693 10310 2745 10362
rect 2757 10310 2809 10362
rect 2821 10310 2873 10362
rect 2885 10310 2937 10362
rect 5987 10310 6039 10362
rect 6051 10310 6103 10362
rect 6115 10310 6167 10362
rect 6179 10310 6231 10362
rect 6243 10310 6295 10362
rect 9345 10310 9397 10362
rect 9409 10310 9461 10362
rect 9473 10310 9525 10362
rect 9537 10310 9589 10362
rect 9601 10310 9653 10362
rect 12703 10310 12755 10362
rect 12767 10310 12819 10362
rect 12831 10310 12883 10362
rect 12895 10310 12947 10362
rect 12959 10310 13011 10362
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 6552 10208 6604 10260
rect 6736 10208 6788 10260
rect 10508 10208 10560 10260
rect 11612 10208 11664 10260
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 2780 10047 2832 10056
rect 2780 10013 2789 10047
rect 2789 10013 2823 10047
rect 2823 10013 2832 10047
rect 2780 10004 2832 10013
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 1860 9936 1912 9988
rect 6368 9936 6420 9988
rect 2504 9868 2556 9920
rect 4712 9868 4764 9920
rect 6552 10047 6604 10056
rect 6552 10013 6561 10047
rect 6561 10013 6595 10047
rect 6595 10013 6604 10047
rect 6552 10004 6604 10013
rect 7104 10140 7156 10192
rect 7196 10072 7248 10124
rect 7288 10115 7340 10124
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 9588 10183 9640 10192
rect 9588 10149 9597 10183
rect 9597 10149 9631 10183
rect 9631 10149 9640 10183
rect 9588 10140 9640 10149
rect 8668 10072 8720 10124
rect 9220 10072 9272 10124
rect 9496 10072 9548 10124
rect 7564 10047 7616 10056
rect 7564 10013 7573 10047
rect 7573 10013 7607 10047
rect 7607 10013 7616 10047
rect 7564 10004 7616 10013
rect 7656 10047 7708 10056
rect 7656 10013 7690 10047
rect 7690 10013 7708 10047
rect 7656 10004 7708 10013
rect 8852 10004 8904 10056
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 10784 10072 10836 10124
rect 10140 10047 10192 10056
rect 10140 10013 10149 10047
rect 10149 10013 10183 10047
rect 10183 10013 10192 10047
rect 10140 10004 10192 10013
rect 9588 9868 9640 9920
rect 9864 9868 9916 9920
rect 11612 10072 11664 10124
rect 11060 10047 11112 10056
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 11796 10047 11848 10056
rect 11796 10013 11805 10047
rect 11805 10013 11839 10047
rect 11839 10013 11848 10047
rect 11796 10004 11848 10013
rect 14096 10072 14148 10124
rect 12072 10047 12124 10056
rect 12072 10013 12081 10047
rect 12081 10013 12115 10047
rect 12115 10013 12124 10047
rect 12072 10004 12124 10013
rect 11612 9868 11664 9920
rect 11796 9868 11848 9920
rect 12164 9868 12216 9920
rect 12348 9868 12400 9920
rect 4308 9766 4360 9818
rect 4372 9766 4424 9818
rect 4436 9766 4488 9818
rect 4500 9766 4552 9818
rect 4564 9766 4616 9818
rect 7666 9766 7718 9818
rect 7730 9766 7782 9818
rect 7794 9766 7846 9818
rect 7858 9766 7910 9818
rect 7922 9766 7974 9818
rect 11024 9766 11076 9818
rect 11088 9766 11140 9818
rect 11152 9766 11204 9818
rect 11216 9766 11268 9818
rect 11280 9766 11332 9818
rect 14382 9766 14434 9818
rect 14446 9766 14498 9818
rect 14510 9766 14562 9818
rect 14574 9766 14626 9818
rect 14638 9766 14690 9818
rect 6828 9664 6880 9716
rect 1768 9596 1820 9648
rect 8208 9664 8260 9716
rect 8576 9664 8628 9716
rect 9588 9664 9640 9716
rect 9680 9664 9732 9716
rect 12440 9664 12492 9716
rect 13820 9664 13872 9716
rect 11612 9596 11664 9648
rect 8300 9528 8352 9580
rect 8576 9528 8628 9580
rect 10140 9571 10192 9580
rect 10140 9537 10149 9571
rect 10149 9537 10183 9571
rect 10183 9537 10192 9571
rect 10140 9528 10192 9537
rect 10232 9571 10284 9580
rect 10232 9537 10266 9571
rect 10266 9537 10284 9571
rect 10232 9528 10284 9537
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 1400 9503 1452 9512
rect 1400 9469 1409 9503
rect 1409 9469 1443 9503
rect 1443 9469 1452 9503
rect 1400 9460 1452 9469
rect 9220 9503 9272 9512
rect 9220 9469 9229 9503
rect 9229 9469 9263 9503
rect 9263 9469 9272 9503
rect 9220 9460 9272 9469
rect 9772 9460 9824 9512
rect 9864 9435 9916 9444
rect 9864 9401 9873 9435
rect 9873 9401 9907 9435
rect 9907 9401 9916 9435
rect 9864 9392 9916 9401
rect 10876 9392 10928 9444
rect 11336 9392 11388 9444
rect 14188 9639 14240 9648
rect 14188 9605 14197 9639
rect 14197 9605 14231 9639
rect 14231 9605 14240 9639
rect 14188 9596 14240 9605
rect 12348 9571 12400 9580
rect 12348 9537 12357 9571
rect 12357 9537 12391 9571
rect 12391 9537 12400 9571
rect 12348 9528 12400 9537
rect 12164 9460 12216 9512
rect 12624 9460 12676 9512
rect 13452 9528 13504 9580
rect 13728 9460 13780 9512
rect 2412 9367 2464 9376
rect 2412 9333 2421 9367
rect 2421 9333 2455 9367
rect 2455 9333 2464 9367
rect 2412 9324 2464 9333
rect 7380 9324 7432 9376
rect 9772 9324 9824 9376
rect 12624 9324 12676 9376
rect 13084 9392 13136 9444
rect 14004 9324 14056 9376
rect 2629 9222 2681 9274
rect 2693 9222 2745 9274
rect 2757 9222 2809 9274
rect 2821 9222 2873 9274
rect 2885 9222 2937 9274
rect 5987 9222 6039 9274
rect 6051 9222 6103 9274
rect 6115 9222 6167 9274
rect 6179 9222 6231 9274
rect 6243 9222 6295 9274
rect 9345 9222 9397 9274
rect 9409 9222 9461 9274
rect 9473 9222 9525 9274
rect 9537 9222 9589 9274
rect 9601 9222 9653 9274
rect 12703 9222 12755 9274
rect 12767 9222 12819 9274
rect 12831 9222 12883 9274
rect 12895 9222 12947 9274
rect 12959 9222 13011 9274
rect 1768 9120 1820 9172
rect 2412 9052 2464 9104
rect 2044 8916 2096 8968
rect 9772 8984 9824 9036
rect 9864 8984 9916 9036
rect 10692 9027 10744 9036
rect 10692 8993 10701 9027
rect 10701 8993 10735 9027
rect 10735 8993 10744 9027
rect 10692 8984 10744 8993
rect 2504 8959 2556 8968
rect 2504 8925 2513 8959
rect 2513 8925 2547 8959
rect 2547 8925 2556 8959
rect 2504 8916 2556 8925
rect 2596 8959 2648 8968
rect 2596 8925 2605 8959
rect 2605 8925 2639 8959
rect 2639 8925 2648 8959
rect 2596 8916 2648 8925
rect 4804 8916 4856 8968
rect 7380 8916 7432 8968
rect 848 8780 900 8832
rect 2320 8823 2372 8832
rect 2320 8789 2329 8823
rect 2329 8789 2363 8823
rect 2363 8789 2372 8823
rect 2320 8780 2372 8789
rect 5540 8780 5592 8832
rect 7288 8780 7340 8832
rect 8484 8916 8536 8968
rect 10416 8959 10468 8968
rect 10416 8925 10425 8959
rect 10425 8925 10459 8959
rect 10459 8925 10468 8959
rect 10416 8916 10468 8925
rect 10508 8959 10560 8968
rect 10508 8925 10542 8959
rect 10542 8925 10560 8959
rect 11520 9120 11572 9172
rect 11704 9120 11756 9172
rect 13820 9120 13872 9172
rect 12624 9052 12676 9104
rect 11336 8984 11388 9036
rect 12532 8984 12584 9036
rect 13912 8984 13964 9036
rect 10508 8916 10560 8925
rect 12624 8916 12676 8968
rect 14832 8916 14884 8968
rect 14188 8848 14240 8900
rect 8392 8780 8444 8832
rect 10508 8780 10560 8832
rect 10692 8780 10744 8832
rect 12072 8780 12124 8832
rect 12532 8780 12584 8832
rect 13176 8780 13228 8832
rect 4308 8678 4360 8730
rect 4372 8678 4424 8730
rect 4436 8678 4488 8730
rect 4500 8678 4552 8730
rect 4564 8678 4616 8730
rect 7666 8678 7718 8730
rect 7730 8678 7782 8730
rect 7794 8678 7846 8730
rect 7858 8678 7910 8730
rect 7922 8678 7974 8730
rect 11024 8678 11076 8730
rect 11088 8678 11140 8730
rect 11152 8678 11204 8730
rect 11216 8678 11268 8730
rect 11280 8678 11332 8730
rect 14382 8678 14434 8730
rect 14446 8678 14498 8730
rect 14510 8678 14562 8730
rect 14574 8678 14626 8730
rect 14638 8678 14690 8730
rect 2320 8576 2372 8628
rect 2596 8576 2648 8628
rect 8852 8576 8904 8628
rect 10324 8576 10376 8628
rect 11796 8576 11848 8628
rect 4804 8440 4856 8492
rect 5908 8508 5960 8560
rect 1676 8347 1728 8356
rect 1676 8313 1685 8347
rect 1685 8313 1719 8347
rect 1719 8313 1728 8347
rect 1676 8304 1728 8313
rect 6736 8483 6788 8492
rect 6736 8449 6745 8483
rect 6745 8449 6779 8483
rect 6779 8449 6788 8483
rect 6736 8440 6788 8449
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 8300 8372 8352 8424
rect 8208 8304 8260 8356
rect 11704 8508 11756 8560
rect 11428 8440 11480 8492
rect 12164 8440 12216 8492
rect 10876 8372 10928 8424
rect 11244 8372 11296 8424
rect 11152 8304 11204 8356
rect 12624 8508 12676 8560
rect 13544 8619 13596 8628
rect 13544 8585 13553 8619
rect 13553 8585 13587 8619
rect 13587 8585 13596 8619
rect 13544 8576 13596 8585
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 13636 8440 13688 8492
rect 8116 8236 8168 8288
rect 8392 8236 8444 8288
rect 9956 8279 10008 8288
rect 9956 8245 9965 8279
rect 9965 8245 9999 8279
rect 9999 8245 10008 8279
rect 9956 8236 10008 8245
rect 10600 8236 10652 8288
rect 2629 8134 2681 8186
rect 2693 8134 2745 8186
rect 2757 8134 2809 8186
rect 2821 8134 2873 8186
rect 2885 8134 2937 8186
rect 5987 8134 6039 8186
rect 6051 8134 6103 8186
rect 6115 8134 6167 8186
rect 6179 8134 6231 8186
rect 6243 8134 6295 8186
rect 9345 8134 9397 8186
rect 9409 8134 9461 8186
rect 9473 8134 9525 8186
rect 9537 8134 9589 8186
rect 9601 8134 9653 8186
rect 12703 8134 12755 8186
rect 12767 8134 12819 8186
rect 12831 8134 12883 8186
rect 12895 8134 12947 8186
rect 12959 8134 13011 8186
rect 6736 8032 6788 8084
rect 7196 8032 7248 8084
rect 7932 8032 7984 8084
rect 8944 8032 8996 8084
rect 9128 8032 9180 8084
rect 9588 7964 9640 8016
rect 10140 7964 10192 8016
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 8024 7896 8076 7948
rect 8116 7939 8168 7948
rect 8116 7905 8125 7939
rect 8125 7905 8159 7939
rect 8159 7905 8168 7939
rect 8116 7896 8168 7905
rect 9312 7896 9364 7948
rect 9680 7896 9732 7948
rect 9956 7896 10008 7948
rect 10508 7939 10560 7948
rect 10508 7905 10517 7939
rect 10517 7905 10551 7939
rect 10551 7905 10560 7939
rect 10508 7896 10560 7905
rect 10600 7939 10652 7948
rect 10600 7905 10634 7939
rect 10634 7905 10652 7939
rect 10600 7896 10652 7905
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 5540 7828 5592 7880
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7288 7828 7340 7880
rect 9496 7828 9548 7880
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 10784 7871 10836 7880
rect 10784 7837 10793 7871
rect 10793 7837 10827 7871
rect 10827 7837 10836 7871
rect 10784 7828 10836 7837
rect 11980 8032 12032 8084
rect 13728 8032 13780 8084
rect 12532 7896 12584 7948
rect 11520 7828 11572 7880
rect 11888 7828 11940 7880
rect 13268 7828 13320 7880
rect 13636 7760 13688 7812
rect 10508 7692 10560 7744
rect 10784 7692 10836 7744
rect 13176 7692 13228 7744
rect 13728 7692 13780 7744
rect 4308 7590 4360 7642
rect 4372 7590 4424 7642
rect 4436 7590 4488 7642
rect 4500 7590 4552 7642
rect 4564 7590 4616 7642
rect 7666 7590 7718 7642
rect 7730 7590 7782 7642
rect 7794 7590 7846 7642
rect 7858 7590 7910 7642
rect 7922 7590 7974 7642
rect 11024 7590 11076 7642
rect 11088 7590 11140 7642
rect 11152 7590 11204 7642
rect 11216 7590 11268 7642
rect 11280 7590 11332 7642
rect 14382 7590 14434 7642
rect 14446 7590 14498 7642
rect 14510 7590 14562 7642
rect 14574 7590 14626 7642
rect 14638 7590 14690 7642
rect 2412 7488 2464 7540
rect 6828 7488 6880 7540
rect 9128 7488 9180 7540
rect 11980 7488 12032 7540
rect 12532 7488 12584 7540
rect 13084 7488 13136 7540
rect 13176 7488 13228 7540
rect 14280 7488 14332 7540
rect 8944 7420 8996 7472
rect 7196 7395 7248 7404
rect 7196 7361 7205 7395
rect 7205 7361 7239 7395
rect 7239 7361 7248 7395
rect 7196 7352 7248 7361
rect 848 7148 900 7200
rect 8208 7352 8260 7404
rect 9312 7352 9364 7404
rect 14832 7420 14884 7472
rect 7564 7284 7616 7336
rect 7932 7284 7984 7336
rect 8392 7327 8444 7336
rect 8392 7293 8401 7327
rect 8401 7293 8435 7327
rect 8435 7293 8444 7327
rect 8392 7284 8444 7293
rect 9680 7327 9732 7336
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 10508 7395 10560 7404
rect 10508 7361 10542 7395
rect 10542 7361 10560 7395
rect 10508 7352 10560 7361
rect 11428 7352 11480 7404
rect 13636 7395 13688 7404
rect 13636 7361 13645 7395
rect 13645 7361 13679 7395
rect 13679 7361 13688 7395
rect 13636 7352 13688 7361
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 11980 7327 12032 7336
rect 11980 7293 11989 7327
rect 11989 7293 12023 7327
rect 12023 7293 12032 7327
rect 11980 7284 12032 7293
rect 9588 7216 9640 7268
rect 9772 7216 9824 7268
rect 9956 7216 10008 7268
rect 10140 7259 10192 7268
rect 10140 7225 10149 7259
rect 10149 7225 10183 7259
rect 10183 7225 10192 7259
rect 10140 7216 10192 7225
rect 9680 7148 9732 7200
rect 10048 7148 10100 7200
rect 10600 7148 10652 7200
rect 11612 7148 11664 7200
rect 11888 7148 11940 7200
rect 12256 7148 12308 7200
rect 2629 7046 2681 7098
rect 2693 7046 2745 7098
rect 2757 7046 2809 7098
rect 2821 7046 2873 7098
rect 2885 7046 2937 7098
rect 5987 7046 6039 7098
rect 6051 7046 6103 7098
rect 6115 7046 6167 7098
rect 6179 7046 6231 7098
rect 6243 7046 6295 7098
rect 9345 7046 9397 7098
rect 9409 7046 9461 7098
rect 9473 7046 9525 7098
rect 9537 7046 9589 7098
rect 9601 7046 9653 7098
rect 12703 7046 12755 7098
rect 12767 7046 12819 7098
rect 12831 7046 12883 7098
rect 12895 7046 12947 7098
rect 12959 7046 13011 7098
rect 7564 6944 7616 6996
rect 7932 6944 7984 6996
rect 8300 6944 8352 6996
rect 8668 6808 8720 6860
rect 8852 6808 8904 6860
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 9864 6944 9916 6996
rect 11796 6876 11848 6928
rect 10508 6808 10560 6860
rect 1492 6715 1544 6724
rect 1492 6681 1501 6715
rect 1501 6681 1535 6715
rect 1535 6681 1544 6715
rect 1492 6672 1544 6681
rect 848 6604 900 6656
rect 9956 6783 10008 6792
rect 9956 6749 9990 6783
rect 9990 6749 10008 6783
rect 9956 6740 10008 6749
rect 8208 6672 8260 6724
rect 7380 6604 7432 6656
rect 9036 6604 9088 6656
rect 11244 6783 11296 6792
rect 11244 6749 11251 6783
rect 11251 6749 11285 6783
rect 11285 6749 11296 6783
rect 11244 6740 11296 6749
rect 10876 6672 10928 6724
rect 11796 6672 11848 6724
rect 13360 6672 13412 6724
rect 13452 6672 13504 6724
rect 10784 6647 10836 6656
rect 10784 6613 10793 6647
rect 10793 6613 10827 6647
rect 10827 6613 10836 6647
rect 10784 6604 10836 6613
rect 10968 6604 11020 6656
rect 12624 6604 12676 6656
rect 15016 6604 15068 6656
rect 4308 6502 4360 6554
rect 4372 6502 4424 6554
rect 4436 6502 4488 6554
rect 4500 6502 4552 6554
rect 4564 6502 4616 6554
rect 7666 6502 7718 6554
rect 7730 6502 7782 6554
rect 7794 6502 7846 6554
rect 7858 6502 7910 6554
rect 7922 6502 7974 6554
rect 11024 6502 11076 6554
rect 11088 6502 11140 6554
rect 11152 6502 11204 6554
rect 11216 6502 11268 6554
rect 11280 6502 11332 6554
rect 14382 6502 14434 6554
rect 14446 6502 14498 6554
rect 14510 6502 14562 6554
rect 14574 6502 14626 6554
rect 14638 6502 14690 6554
rect 9772 6400 9824 6452
rect 9956 6400 10008 6452
rect 11888 6400 11940 6452
rect 6460 6332 6512 6384
rect 15108 6400 15160 6452
rect 7380 6264 7432 6316
rect 8576 6264 8628 6316
rect 9680 6264 9732 6316
rect 10324 6307 10376 6316
rect 10324 6273 10358 6307
rect 10358 6273 10376 6307
rect 10324 6264 10376 6273
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 12072 6264 12124 6316
rect 13452 6332 13504 6384
rect 13636 6332 13688 6384
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 9220 6196 9272 6248
rect 2320 6060 2372 6112
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 10876 6196 10928 6248
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 13728 6264 13780 6316
rect 9956 6171 10008 6180
rect 9956 6137 9965 6171
rect 9965 6137 9999 6171
rect 9999 6137 10008 6171
rect 9956 6128 10008 6137
rect 10968 6128 11020 6180
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 12624 6060 12676 6112
rect 2629 5958 2681 6010
rect 2693 5958 2745 6010
rect 2757 5958 2809 6010
rect 2821 5958 2873 6010
rect 2885 5958 2937 6010
rect 5987 5958 6039 6010
rect 6051 5958 6103 6010
rect 6115 5958 6167 6010
rect 6179 5958 6231 6010
rect 6243 5958 6295 6010
rect 9345 5958 9397 6010
rect 9409 5958 9461 6010
rect 9473 5958 9525 6010
rect 9537 5958 9589 6010
rect 9601 5958 9653 6010
rect 12703 5958 12755 6010
rect 12767 5958 12819 6010
rect 12831 5958 12883 6010
rect 12895 5958 12947 6010
rect 12959 5958 13011 6010
rect 1492 5856 1544 5908
rect 2412 5856 2464 5908
rect 7380 5856 7432 5908
rect 8392 5856 8444 5908
rect 8576 5856 8628 5908
rect 12900 5856 12952 5908
rect 8668 5788 8720 5840
rect 10968 5788 11020 5840
rect 13636 5856 13688 5908
rect 2596 5652 2648 5704
rect 10692 5720 10744 5772
rect 11152 5720 11204 5772
rect 11336 5720 11388 5772
rect 11520 5763 11572 5772
rect 11520 5729 11529 5763
rect 11529 5729 11563 5763
rect 11563 5729 11572 5763
rect 11520 5720 11572 5729
rect 11612 5763 11664 5772
rect 11612 5729 11646 5763
rect 11646 5729 11664 5763
rect 11612 5720 11664 5729
rect 12440 5720 12492 5772
rect 8300 5652 8352 5704
rect 8944 5652 8996 5704
rect 11796 5695 11848 5704
rect 11796 5661 11805 5695
rect 11805 5661 11839 5695
rect 11839 5661 11848 5695
rect 11796 5652 11848 5661
rect 1584 5559 1636 5568
rect 1584 5525 1593 5559
rect 1593 5525 1627 5559
rect 1627 5525 1636 5559
rect 1584 5516 1636 5525
rect 12440 5627 12492 5636
rect 12440 5593 12449 5627
rect 12449 5593 12483 5627
rect 12483 5593 12492 5627
rect 12440 5584 12492 5593
rect 12808 5695 12860 5704
rect 12808 5661 12817 5695
rect 12817 5661 12860 5695
rect 12808 5652 12860 5661
rect 13728 5652 13780 5704
rect 12716 5516 12768 5568
rect 4308 5414 4360 5466
rect 4372 5414 4424 5466
rect 4436 5414 4488 5466
rect 4500 5414 4552 5466
rect 4564 5414 4616 5466
rect 7666 5414 7718 5466
rect 7730 5414 7782 5466
rect 7794 5414 7846 5466
rect 7858 5414 7910 5466
rect 7922 5414 7974 5466
rect 11024 5414 11076 5466
rect 11088 5414 11140 5466
rect 11152 5414 11204 5466
rect 11216 5414 11268 5466
rect 11280 5414 11332 5466
rect 14382 5414 14434 5466
rect 14446 5414 14498 5466
rect 14510 5414 14562 5466
rect 14574 5414 14626 5466
rect 14638 5414 14690 5466
rect 8760 5312 8812 5364
rect 4712 5176 4764 5228
rect 7012 5176 7064 5228
rect 10508 5312 10560 5364
rect 11796 5312 11848 5364
rect 13176 5312 13228 5364
rect 7380 5108 7432 5160
rect 8208 5108 8260 5160
rect 10232 5108 10284 5160
rect 8944 5040 8996 5092
rect 848 4972 900 5024
rect 12716 5108 12768 5160
rect 12532 4972 12584 5024
rect 12900 4972 12952 5024
rect 2629 4870 2681 4922
rect 2693 4870 2745 4922
rect 2757 4870 2809 4922
rect 2821 4870 2873 4922
rect 2885 4870 2937 4922
rect 5987 4870 6039 4922
rect 6051 4870 6103 4922
rect 6115 4870 6167 4922
rect 6179 4870 6231 4922
rect 6243 4870 6295 4922
rect 9345 4870 9397 4922
rect 9409 4870 9461 4922
rect 9473 4870 9525 4922
rect 9537 4870 9589 4922
rect 9601 4870 9653 4922
rect 12703 4870 12755 4922
rect 12767 4870 12819 4922
rect 12831 4870 12883 4922
rect 12895 4870 12947 4922
rect 12959 4870 13011 4922
rect 4988 4768 5040 4820
rect 9956 4811 10008 4820
rect 9956 4777 9965 4811
rect 9965 4777 9999 4811
rect 9999 4777 10008 4811
rect 9956 4768 10008 4777
rect 11244 4768 11296 4820
rect 11428 4768 11480 4820
rect 12532 4768 12584 4820
rect 13360 4768 13412 4820
rect 8208 4632 8260 4684
rect 9220 4607 9272 4616
rect 9220 4573 9227 4607
rect 9227 4573 9261 4607
rect 9261 4573 9272 4607
rect 9220 4564 9272 4573
rect 10232 4632 10284 4684
rect 11336 4632 11388 4684
rect 10600 4607 10652 4616
rect 10600 4573 10609 4607
rect 10609 4573 10652 4607
rect 10600 4564 10652 4573
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 12624 4607 12676 4616
rect 12348 4539 12400 4548
rect 12348 4505 12357 4539
rect 12357 4505 12391 4539
rect 12391 4505 12400 4539
rect 12348 4496 12400 4505
rect 9036 4428 9088 4480
rect 12624 4573 12633 4607
rect 12633 4573 12667 4607
rect 12667 4573 12676 4607
rect 12624 4564 12676 4573
rect 12532 4496 12584 4548
rect 13268 4564 13320 4616
rect 4308 4326 4360 4378
rect 4372 4326 4424 4378
rect 4436 4326 4488 4378
rect 4500 4326 4552 4378
rect 4564 4326 4616 4378
rect 7666 4326 7718 4378
rect 7730 4326 7782 4378
rect 7794 4326 7846 4378
rect 7858 4326 7910 4378
rect 7922 4326 7974 4378
rect 11024 4326 11076 4378
rect 11088 4326 11140 4378
rect 11152 4326 11204 4378
rect 11216 4326 11268 4378
rect 11280 4326 11332 4378
rect 14382 4326 14434 4378
rect 14446 4326 14498 4378
rect 14510 4326 14562 4378
rect 14574 4326 14626 4378
rect 14638 4326 14690 4378
rect 9220 4224 9272 4276
rect 12532 4224 12584 4276
rect 10324 4156 10376 4208
rect 12348 4199 12400 4208
rect 12348 4165 12357 4199
rect 12357 4165 12391 4199
rect 12391 4165 12400 4199
rect 12348 4156 12400 4165
rect 13912 4156 13964 4208
rect 15292 4156 15344 4208
rect 756 4088 808 4140
rect 11704 4088 11756 4140
rect 13452 4088 13504 4140
rect 13636 4131 13688 4140
rect 13636 4097 13645 4131
rect 13645 4097 13679 4131
rect 13679 4097 13688 4131
rect 13636 4088 13688 4097
rect 15384 4088 15436 4140
rect 5080 3952 5132 4004
rect 3424 3884 3476 3936
rect 13820 3884 13872 3936
rect 2629 3782 2681 3834
rect 2693 3782 2745 3834
rect 2757 3782 2809 3834
rect 2821 3782 2873 3834
rect 2885 3782 2937 3834
rect 5987 3782 6039 3834
rect 6051 3782 6103 3834
rect 6115 3782 6167 3834
rect 6179 3782 6231 3834
rect 6243 3782 6295 3834
rect 9345 3782 9397 3834
rect 9409 3782 9461 3834
rect 9473 3782 9525 3834
rect 9537 3782 9589 3834
rect 9601 3782 9653 3834
rect 12703 3782 12755 3834
rect 12767 3782 12819 3834
rect 12831 3782 12883 3834
rect 12895 3782 12947 3834
rect 12959 3782 13011 3834
rect 8484 3680 8536 3732
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 4308 3238 4360 3290
rect 4372 3238 4424 3290
rect 4436 3238 4488 3290
rect 4500 3238 4552 3290
rect 4564 3238 4616 3290
rect 7666 3238 7718 3290
rect 7730 3238 7782 3290
rect 7794 3238 7846 3290
rect 7858 3238 7910 3290
rect 7922 3238 7974 3290
rect 11024 3238 11076 3290
rect 11088 3238 11140 3290
rect 11152 3238 11204 3290
rect 11216 3238 11268 3290
rect 11280 3238 11332 3290
rect 14382 3238 14434 3290
rect 14446 3238 14498 3290
rect 14510 3238 14562 3290
rect 14574 3238 14626 3290
rect 14638 3238 14690 3290
rect 13084 2796 13136 2848
rect 13360 2796 13412 2848
rect 2629 2694 2681 2746
rect 2693 2694 2745 2746
rect 2757 2694 2809 2746
rect 2821 2694 2873 2746
rect 2885 2694 2937 2746
rect 5987 2694 6039 2746
rect 6051 2694 6103 2746
rect 6115 2694 6167 2746
rect 6179 2694 6231 2746
rect 6243 2694 6295 2746
rect 9345 2694 9397 2746
rect 9409 2694 9461 2746
rect 9473 2694 9525 2746
rect 9537 2694 9589 2746
rect 9601 2694 9653 2746
rect 12703 2694 12755 2746
rect 12767 2694 12819 2746
rect 12831 2694 12883 2746
rect 12895 2694 12947 2746
rect 12959 2694 13011 2746
rect 4308 2150 4360 2202
rect 4372 2150 4424 2202
rect 4436 2150 4488 2202
rect 4500 2150 4552 2202
rect 4564 2150 4616 2202
rect 7666 2150 7718 2202
rect 7730 2150 7782 2202
rect 7794 2150 7846 2202
rect 7858 2150 7910 2202
rect 7922 2150 7974 2202
rect 11024 2150 11076 2202
rect 11088 2150 11140 2202
rect 11152 2150 11204 2202
rect 11216 2150 11268 2202
rect 11280 2150 11332 2202
rect 14382 2150 14434 2202
rect 14446 2150 14498 2202
rect 14510 2150 14562 2202
rect 14574 2150 14626 2202
rect 14638 2150 14690 2202
rect 6644 2048 6696 2100
rect 7196 2091 7248 2100
rect 7196 2057 7205 2091
rect 7205 2057 7239 2091
rect 7239 2057 7248 2091
rect 7196 2048 7248 2057
rect 7472 2048 7524 2100
rect 8668 2091 8720 2100
rect 8668 2057 8677 2091
rect 8677 2057 8711 2091
rect 8711 2057 8720 2091
rect 8668 2048 8720 2057
rect 9404 2091 9456 2100
rect 9404 2057 9413 2091
rect 9413 2057 9447 2091
rect 9447 2057 9456 2091
rect 9404 2048 9456 2057
rect 10140 2091 10192 2100
rect 10140 2057 10149 2091
rect 10149 2057 10183 2091
rect 10183 2057 10192 2091
rect 10140 2048 10192 2057
rect 10876 2091 10928 2100
rect 10876 2057 10885 2091
rect 10885 2057 10919 2091
rect 10919 2057 10928 2091
rect 10876 2048 10928 2057
rect 13452 2091 13504 2100
rect 13452 2057 13461 2091
rect 13461 2057 13495 2091
rect 13495 2057 13504 2091
rect 13452 2048 13504 2057
rect 9036 1980 9088 2032
rect 2044 1955 2096 1964
rect 2044 1921 2053 1955
rect 2053 1921 2087 1955
rect 2087 1921 2096 1955
rect 2044 1912 2096 1921
rect 6460 1955 6512 1964
rect 6460 1921 6469 1955
rect 6469 1921 6503 1955
rect 6503 1921 6512 1955
rect 6460 1912 6512 1921
rect 7104 1955 7156 1964
rect 7104 1921 7113 1955
rect 7113 1921 7147 1955
rect 7147 1921 7156 1955
rect 7104 1912 7156 1921
rect 7840 1955 7892 1964
rect 7840 1921 7849 1955
rect 7849 1921 7883 1955
rect 7883 1921 7892 1955
rect 7840 1912 7892 1921
rect 8576 1955 8628 1964
rect 8576 1921 8585 1955
rect 8585 1921 8619 1955
rect 8619 1921 8628 1955
rect 8576 1912 8628 1921
rect 9220 1912 9272 1964
rect 10048 1955 10100 1964
rect 10048 1921 10057 1955
rect 10057 1921 10091 1955
rect 10091 1921 10100 1955
rect 10048 1912 10100 1921
rect 10784 1955 10836 1964
rect 10784 1921 10793 1955
rect 10793 1921 10827 1955
rect 10827 1921 10836 1955
rect 10784 1912 10836 1921
rect 11612 1955 11664 1964
rect 11612 1921 11621 1955
rect 11621 1921 11655 1955
rect 11655 1921 11664 1955
rect 11612 1912 11664 1921
rect 12256 1955 12308 1964
rect 12256 1921 12265 1955
rect 12265 1921 12299 1955
rect 12299 1921 12308 1955
rect 12256 1912 12308 1921
rect 13084 1912 13136 1964
rect 13728 1955 13780 1964
rect 13728 1921 13737 1955
rect 13737 1921 13771 1955
rect 13771 1921 13780 1955
rect 13728 1912 13780 1921
rect 14188 1955 14240 1964
rect 14188 1921 14197 1955
rect 14197 1921 14231 1955
rect 14231 1921 14240 1955
rect 14188 1912 14240 1921
rect 4160 1776 4212 1828
rect 14740 1844 14792 1896
rect 15568 1844 15620 1896
rect 14832 1708 14884 1760
rect 2629 1606 2681 1658
rect 2693 1606 2745 1658
rect 2757 1606 2809 1658
rect 2821 1606 2873 1658
rect 2885 1606 2937 1658
rect 5987 1606 6039 1658
rect 6051 1606 6103 1658
rect 6115 1606 6167 1658
rect 6179 1606 6231 1658
rect 6243 1606 6295 1658
rect 9345 1606 9397 1658
rect 9409 1606 9461 1658
rect 9473 1606 9525 1658
rect 9537 1606 9589 1658
rect 9601 1606 9653 1658
rect 12703 1606 12755 1658
rect 12767 1606 12819 1658
rect 12831 1606 12883 1658
rect 12895 1606 12947 1658
rect 12959 1606 13011 1658
rect 6460 1504 6512 1556
rect 7104 1504 7156 1556
rect 7840 1504 7892 1556
rect 8576 1504 8628 1556
rect 9220 1504 9272 1556
rect 10048 1504 10100 1556
rect 10784 1504 10836 1556
rect 11612 1547 11664 1556
rect 11612 1513 11621 1547
rect 11621 1513 11655 1547
rect 11655 1513 11664 1547
rect 11612 1504 11664 1513
rect 12256 1504 12308 1556
rect 13084 1547 13136 1556
rect 13084 1513 13093 1547
rect 13093 1513 13127 1547
rect 13127 1513 13136 1547
rect 13084 1504 13136 1513
rect 13728 1504 13780 1556
rect 9128 1436 9180 1488
rect 1216 1300 1268 1352
rect 2504 1300 2556 1352
rect 2688 1343 2740 1352
rect 2688 1309 2697 1343
rect 2697 1309 2731 1343
rect 2731 1309 2740 1343
rect 2688 1300 2740 1309
rect 2320 1232 2372 1284
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 4620 1343 4672 1352
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 5172 1300 5224 1352
rect 6184 1343 6236 1352
rect 6184 1309 6193 1343
rect 6193 1309 6227 1343
rect 6227 1309 6236 1343
rect 6184 1300 6236 1309
rect 4160 1232 4212 1284
rect 5080 1275 5132 1284
rect 5080 1241 5089 1275
rect 5089 1241 5123 1275
rect 5123 1241 5132 1275
rect 5080 1232 5132 1241
rect 5632 1232 5684 1284
rect 6644 1343 6696 1352
rect 6644 1309 6653 1343
rect 6653 1309 6687 1343
rect 6687 1309 6696 1343
rect 6644 1300 6696 1309
rect 7104 1300 7156 1352
rect 8116 1343 8168 1352
rect 8116 1309 8125 1343
rect 8125 1309 8159 1343
rect 8159 1309 8168 1343
rect 8116 1300 8168 1309
rect 8576 1300 8628 1352
rect 9312 1300 9364 1352
rect 10048 1300 10100 1352
rect 10784 1300 10836 1352
rect 11520 1300 11572 1352
rect 12256 1300 12308 1352
rect 13268 1343 13320 1352
rect 13268 1309 13277 1343
rect 13277 1309 13311 1343
rect 13311 1309 13320 1343
rect 13268 1300 13320 1309
rect 13544 1343 13596 1352
rect 13544 1309 13553 1343
rect 13553 1309 13587 1343
rect 13587 1309 13596 1343
rect 13544 1300 13596 1309
rect 15200 1300 15252 1352
rect 13820 1207 13872 1216
rect 13820 1173 13829 1207
rect 13829 1173 13863 1207
rect 13863 1173 13872 1207
rect 13820 1164 13872 1173
rect 4308 1062 4360 1114
rect 4372 1062 4424 1114
rect 4436 1062 4488 1114
rect 4500 1062 4552 1114
rect 4564 1062 4616 1114
rect 7666 1062 7718 1114
rect 7730 1062 7782 1114
rect 7794 1062 7846 1114
rect 7858 1062 7910 1114
rect 7922 1062 7974 1114
rect 11024 1062 11076 1114
rect 11088 1062 11140 1114
rect 11152 1062 11204 1114
rect 11216 1062 11268 1114
rect 11280 1062 11332 1114
rect 14382 1062 14434 1114
rect 14446 1062 14498 1114
rect 14510 1062 14562 1114
rect 14574 1062 14626 1114
rect 14638 1062 14690 1114
<< metal2 >>
rect 478 44540 534 45000
rect 1214 44540 1270 45000
rect 1950 44540 2006 45000
rect 2686 44540 2742 45000
rect 3422 44540 3478 45000
rect 4158 44540 4214 45000
rect 4894 44540 4950 45000
rect 5630 44540 5686 45000
rect 6366 44540 6422 45000
rect 7102 44540 7158 45000
rect 7838 44540 7894 45000
rect 8574 44540 8630 45000
rect 9310 44540 9366 45000
rect 10046 44540 10102 45000
rect 10782 44540 10838 45000
rect 11518 44540 11574 45000
rect 12254 44540 12310 45000
rect 12990 44540 13046 45000
rect 13726 44540 13782 45000
rect 14462 44540 14518 45000
rect 15198 44540 15254 45000
rect 492 43450 520 44540
rect 480 43444 532 43450
rect 480 43386 532 43392
rect 1228 43058 1256 44540
rect 1768 43308 1820 43314
rect 1768 43250 1820 43256
rect 1400 43104 1452 43110
rect 1228 43052 1400 43058
rect 1228 43046 1452 43052
rect 1228 43030 1440 43046
rect 1400 42628 1452 42634
rect 1400 42570 1452 42576
rect 1412 41449 1440 42570
rect 1398 41440 1454 41449
rect 1398 41375 1454 41384
rect 756 41132 808 41138
rect 756 41074 808 41080
rect 768 40633 796 41074
rect 754 40624 810 40633
rect 754 40559 810 40568
rect 1492 40112 1544 40118
rect 1492 40054 1544 40060
rect 1504 39953 1532 40054
rect 1490 39944 1546 39953
rect 1490 39879 1546 39888
rect 756 39364 808 39370
rect 756 39306 808 39312
rect 768 39001 796 39306
rect 754 38992 810 39001
rect 754 38927 810 38936
rect 756 38344 808 38350
rect 756 38286 808 38292
rect 768 38185 796 38286
rect 754 38176 810 38185
rect 754 38111 810 38120
rect 756 37868 808 37874
rect 756 37810 808 37816
rect 768 37369 796 37810
rect 754 37360 810 37369
rect 754 37295 810 37304
rect 1584 37188 1636 37194
rect 1584 37130 1636 37136
rect 756 36780 808 36786
rect 756 36722 808 36728
rect 768 36553 796 36722
rect 754 36544 810 36553
rect 754 36479 810 36488
rect 1492 36100 1544 36106
rect 1492 36042 1544 36048
rect 1504 35873 1532 36042
rect 1490 35864 1546 35873
rect 1490 35799 1546 35808
rect 756 35080 808 35086
rect 756 35022 808 35028
rect 768 34921 796 35022
rect 754 34912 810 34921
rect 754 34847 810 34856
rect 1400 34604 1452 34610
rect 1400 34546 1452 34552
rect 1412 34513 1440 34546
rect 1398 34504 1454 34513
rect 1398 34439 1454 34448
rect 756 33516 808 33522
rect 756 33458 808 33464
rect 768 33289 796 33458
rect 754 33280 810 33289
rect 754 33215 810 33224
rect 756 32904 808 32910
rect 756 32846 808 32852
rect 768 32473 796 32846
rect 1596 32774 1624 37130
rect 1780 36650 1808 43250
rect 1964 43178 1992 44540
rect 2700 43874 2728 44540
rect 2700 43846 2820 43874
rect 2044 43308 2096 43314
rect 2044 43250 2096 43256
rect 1952 43172 2004 43178
rect 1952 43114 2004 43120
rect 2056 42362 2084 43250
rect 2792 43110 2820 43846
rect 3436 43450 3464 44540
rect 4172 43450 4200 44540
rect 4308 43548 4616 43557
rect 4308 43546 4314 43548
rect 4370 43546 4394 43548
rect 4450 43546 4474 43548
rect 4530 43546 4554 43548
rect 4610 43546 4616 43548
rect 4370 43494 4372 43546
rect 4552 43494 4554 43546
rect 4308 43492 4314 43494
rect 4370 43492 4394 43494
rect 4450 43492 4474 43494
rect 4530 43492 4554 43494
rect 4610 43492 4616 43494
rect 4308 43483 4616 43492
rect 4908 43450 4936 44540
rect 5644 43450 5672 44540
rect 6380 43450 6408 44540
rect 7116 43450 7144 44540
rect 7852 43874 7880 44540
rect 7852 43846 8064 43874
rect 7666 43548 7974 43557
rect 7666 43546 7672 43548
rect 7728 43546 7752 43548
rect 7808 43546 7832 43548
rect 7888 43546 7912 43548
rect 7968 43546 7974 43548
rect 7728 43494 7730 43546
rect 7910 43494 7912 43546
rect 7666 43492 7672 43494
rect 7728 43492 7752 43494
rect 7808 43492 7832 43494
rect 7888 43492 7912 43494
rect 7968 43492 7974 43494
rect 7666 43483 7974 43492
rect 8036 43450 8064 43846
rect 8588 43450 8616 44540
rect 9324 43450 9352 44540
rect 10060 43450 10088 44540
rect 10796 43450 10824 44540
rect 11024 43548 11332 43557
rect 11024 43546 11030 43548
rect 11086 43546 11110 43548
rect 11166 43546 11190 43548
rect 11246 43546 11270 43548
rect 11326 43546 11332 43548
rect 11086 43494 11088 43546
rect 11268 43494 11270 43546
rect 11024 43492 11030 43494
rect 11086 43492 11110 43494
rect 11166 43492 11190 43494
rect 11246 43492 11270 43494
rect 11326 43492 11332 43494
rect 11024 43483 11332 43492
rect 11532 43450 11560 44540
rect 12268 43450 12296 44540
rect 13004 43450 13032 44540
rect 3424 43444 3476 43450
rect 3424 43386 3476 43392
rect 4160 43444 4212 43450
rect 4160 43386 4212 43392
rect 4896 43444 4948 43450
rect 4896 43386 4948 43392
rect 5632 43444 5684 43450
rect 5632 43386 5684 43392
rect 6368 43444 6420 43450
rect 6368 43386 6420 43392
rect 7104 43444 7156 43450
rect 7104 43386 7156 43392
rect 8024 43444 8076 43450
rect 8024 43386 8076 43392
rect 8576 43444 8628 43450
rect 8576 43386 8628 43392
rect 9312 43444 9364 43450
rect 9312 43386 9364 43392
rect 10048 43444 10100 43450
rect 10048 43386 10100 43392
rect 10784 43444 10836 43450
rect 10784 43386 10836 43392
rect 11520 43444 11572 43450
rect 11520 43386 11572 43392
rect 12256 43444 12308 43450
rect 12256 43386 12308 43392
rect 12992 43444 13044 43450
rect 12992 43386 13044 43392
rect 3056 43308 3108 43314
rect 3056 43250 3108 43256
rect 3148 43308 3200 43314
rect 3148 43250 3200 43256
rect 3792 43308 3844 43314
rect 3792 43250 3844 43256
rect 4344 43308 4396 43314
rect 4344 43250 4396 43256
rect 4988 43308 5040 43314
rect 5724 43308 5776 43314
rect 4988 43250 5040 43256
rect 5552 43268 5724 43296
rect 2780 43104 2832 43110
rect 2780 43046 2832 43052
rect 2629 43004 2937 43013
rect 2629 43002 2635 43004
rect 2691 43002 2715 43004
rect 2771 43002 2795 43004
rect 2851 43002 2875 43004
rect 2931 43002 2937 43004
rect 2691 42950 2693 43002
rect 2873 42950 2875 43002
rect 2629 42948 2635 42950
rect 2691 42948 2715 42950
rect 2771 42948 2795 42950
rect 2851 42948 2875 42950
rect 2931 42948 2937 42950
rect 2629 42939 2937 42948
rect 2044 42356 2096 42362
rect 2044 42298 2096 42304
rect 2136 42220 2188 42226
rect 2136 42162 2188 42168
rect 1952 36780 2004 36786
rect 1952 36722 2004 36728
rect 1768 36644 1820 36650
rect 1768 36586 1820 36592
rect 1964 36378 1992 36722
rect 1952 36372 2004 36378
rect 1952 36314 2004 36320
rect 1584 32768 1636 32774
rect 1584 32710 1636 32716
rect 1860 32768 1912 32774
rect 1860 32710 1912 32716
rect 754 32464 810 32473
rect 754 32399 810 32408
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31657 1440 31758
rect 1768 31680 1820 31686
rect 1398 31648 1454 31657
rect 1768 31622 1820 31628
rect 1398 31583 1454 31592
rect 756 31340 808 31346
rect 756 31282 808 31288
rect 768 30841 796 31282
rect 754 30832 810 30841
rect 754 30767 810 30776
rect 756 30252 808 30258
rect 756 30194 808 30200
rect 768 30025 796 30194
rect 754 30016 810 30025
rect 754 29951 810 29960
rect 756 29640 808 29646
rect 756 29582 808 29588
rect 768 29209 796 29582
rect 754 29200 810 29209
rect 754 29135 810 29144
rect 1780 29073 1808 31622
rect 1766 29064 1822 29073
rect 1766 28999 1822 29008
rect 756 28552 808 28558
rect 756 28494 808 28500
rect 1582 28520 1638 28529
rect 768 28393 796 28494
rect 1582 28455 1638 28464
rect 754 28384 810 28393
rect 754 28319 810 28328
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27577 1440 28018
rect 1596 27878 1624 28455
rect 1584 27872 1636 27878
rect 1584 27814 1636 27820
rect 1398 27568 1454 27577
rect 1398 27503 1454 27512
rect 756 26988 808 26994
rect 756 26930 808 26936
rect 768 26761 796 26930
rect 754 26752 810 26761
rect 754 26687 810 26696
rect 1492 26308 1544 26314
rect 1492 26250 1544 26256
rect 1504 26217 1532 26250
rect 1490 26208 1546 26217
rect 1490 26143 1546 26152
rect 1596 25888 1624 27814
rect 1676 27532 1728 27538
rect 1676 27474 1728 27480
rect 1688 27130 1716 27474
rect 1676 27124 1728 27130
rect 1676 27066 1728 27072
rect 1504 25860 1624 25888
rect 756 25288 808 25294
rect 756 25230 808 25236
rect 768 25129 796 25230
rect 754 25120 810 25129
rect 754 25055 810 25064
rect 756 24812 808 24818
rect 756 24754 808 24760
rect 768 24313 796 24754
rect 754 24304 810 24313
rect 754 24239 810 24248
rect 756 23724 808 23730
rect 756 23666 808 23672
rect 768 23497 796 23666
rect 754 23488 810 23497
rect 754 23423 810 23432
rect 756 23044 808 23050
rect 756 22986 808 22992
rect 768 22681 796 22986
rect 754 22672 810 22681
rect 754 22607 810 22616
rect 756 21956 808 21962
rect 756 21898 808 21904
rect 768 21865 796 21898
rect 754 21856 810 21865
rect 754 21791 810 21800
rect 756 21548 808 21554
rect 756 21490 808 21496
rect 768 21049 796 21490
rect 754 21040 810 21049
rect 754 20975 810 20984
rect 756 20392 808 20398
rect 756 20334 808 20340
rect 768 20233 796 20334
rect 754 20224 810 20233
rect 754 20159 810 20168
rect 756 19780 808 19786
rect 756 19722 808 19728
rect 768 19417 796 19722
rect 754 19408 810 19417
rect 754 19343 810 19352
rect 1504 19334 1532 25860
rect 1688 20618 1716 27066
rect 1320 19306 1532 19334
rect 1596 20590 1716 20618
rect 756 18692 808 18698
rect 756 18634 808 18640
rect 768 18601 796 18634
rect 754 18592 810 18601
rect 754 18527 810 18536
rect 480 18216 532 18222
rect 480 18158 532 18164
rect 492 160 520 18158
rect 756 17196 808 17202
rect 756 17138 808 17144
rect 768 16969 796 17138
rect 754 16960 810 16969
rect 754 16895 810 16904
rect 756 16516 808 16522
rect 756 16458 808 16464
rect 768 16153 796 16458
rect 754 16144 810 16153
rect 754 16079 810 16088
rect 756 15428 808 15434
rect 756 15370 808 15376
rect 768 15337 796 15370
rect 754 15328 810 15337
rect 754 15263 810 15272
rect 1320 15162 1348 19306
rect 1492 18284 1544 18290
rect 1492 18226 1544 18232
rect 1504 17921 1532 18226
rect 1490 17912 1546 17921
rect 1490 17847 1546 17856
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1412 16114 1440 17614
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1308 15156 1360 15162
rect 1308 15098 1360 15104
rect 848 14816 900 14822
rect 848 14758 900 14764
rect 860 14521 888 14758
rect 846 14512 902 14521
rect 846 14447 902 14456
rect 1320 14414 1348 15098
rect 1412 14482 1440 16050
rect 1504 15094 1532 16934
rect 1492 15088 1544 15094
rect 1492 15030 1544 15036
rect 1596 14958 1624 20590
rect 1676 20528 1728 20534
rect 1676 20470 1728 20476
rect 1688 20058 1716 20470
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1780 19334 1808 28999
rect 1872 27470 1900 32710
rect 2148 29850 2176 42162
rect 2629 41916 2937 41925
rect 2629 41914 2635 41916
rect 2691 41914 2715 41916
rect 2771 41914 2795 41916
rect 2851 41914 2875 41916
rect 2931 41914 2937 41916
rect 2691 41862 2693 41914
rect 2873 41862 2875 41914
rect 2629 41860 2635 41862
rect 2691 41860 2715 41862
rect 2771 41860 2795 41862
rect 2851 41860 2875 41862
rect 2931 41860 2937 41862
rect 2629 41851 2937 41860
rect 2629 40828 2937 40837
rect 2629 40826 2635 40828
rect 2691 40826 2715 40828
rect 2771 40826 2795 40828
rect 2851 40826 2875 40828
rect 2931 40826 2937 40828
rect 2691 40774 2693 40826
rect 2873 40774 2875 40826
rect 2629 40772 2635 40774
rect 2691 40772 2715 40774
rect 2771 40772 2795 40774
rect 2851 40772 2875 40774
rect 2931 40772 2937 40774
rect 2629 40763 2937 40772
rect 2629 39740 2937 39749
rect 2629 39738 2635 39740
rect 2691 39738 2715 39740
rect 2771 39738 2795 39740
rect 2851 39738 2875 39740
rect 2931 39738 2937 39740
rect 2691 39686 2693 39738
rect 2873 39686 2875 39738
rect 2629 39684 2635 39686
rect 2691 39684 2715 39686
rect 2771 39684 2795 39686
rect 2851 39684 2875 39686
rect 2931 39684 2937 39686
rect 2629 39675 2937 39684
rect 2629 38652 2937 38661
rect 2629 38650 2635 38652
rect 2691 38650 2715 38652
rect 2771 38650 2795 38652
rect 2851 38650 2875 38652
rect 2931 38650 2937 38652
rect 2691 38598 2693 38650
rect 2873 38598 2875 38650
rect 2629 38596 2635 38598
rect 2691 38596 2715 38598
rect 2771 38596 2795 38598
rect 2851 38596 2875 38598
rect 2931 38596 2937 38598
rect 2629 38587 2937 38596
rect 2629 37564 2937 37573
rect 2629 37562 2635 37564
rect 2691 37562 2715 37564
rect 2771 37562 2795 37564
rect 2851 37562 2875 37564
rect 2931 37562 2937 37564
rect 2691 37510 2693 37562
rect 2873 37510 2875 37562
rect 2629 37508 2635 37510
rect 2691 37508 2715 37510
rect 2771 37508 2795 37510
rect 2851 37508 2875 37510
rect 2931 37508 2937 37510
rect 2629 37499 2937 37508
rect 2629 36476 2937 36485
rect 2629 36474 2635 36476
rect 2691 36474 2715 36476
rect 2771 36474 2795 36476
rect 2851 36474 2875 36476
rect 2931 36474 2937 36476
rect 2691 36422 2693 36474
rect 2873 36422 2875 36474
rect 2629 36420 2635 36422
rect 2691 36420 2715 36422
rect 2771 36420 2795 36422
rect 2851 36420 2875 36422
rect 2931 36420 2937 36422
rect 2629 36411 2937 36420
rect 2629 35388 2937 35397
rect 2629 35386 2635 35388
rect 2691 35386 2715 35388
rect 2771 35386 2795 35388
rect 2851 35386 2875 35388
rect 2931 35386 2937 35388
rect 2691 35334 2693 35386
rect 2873 35334 2875 35386
rect 2629 35332 2635 35334
rect 2691 35332 2715 35334
rect 2771 35332 2795 35334
rect 2851 35332 2875 35334
rect 2931 35332 2937 35334
rect 2629 35323 2937 35332
rect 2629 34300 2937 34309
rect 2629 34298 2635 34300
rect 2691 34298 2715 34300
rect 2771 34298 2795 34300
rect 2851 34298 2875 34300
rect 2931 34298 2937 34300
rect 2691 34246 2693 34298
rect 2873 34246 2875 34298
rect 2629 34244 2635 34246
rect 2691 34244 2715 34246
rect 2771 34244 2795 34246
rect 2851 34244 2875 34246
rect 2931 34244 2937 34246
rect 2629 34235 2937 34244
rect 2629 33212 2937 33221
rect 2629 33210 2635 33212
rect 2691 33210 2715 33212
rect 2771 33210 2795 33212
rect 2851 33210 2875 33212
rect 2931 33210 2937 33212
rect 2691 33158 2693 33210
rect 2873 33158 2875 33210
rect 2629 33156 2635 33158
rect 2691 33156 2715 33158
rect 2771 33156 2795 33158
rect 2851 33156 2875 33158
rect 2931 33156 2937 33158
rect 2629 33147 2937 33156
rect 2629 32124 2937 32133
rect 2629 32122 2635 32124
rect 2691 32122 2715 32124
rect 2771 32122 2795 32124
rect 2851 32122 2875 32124
rect 2931 32122 2937 32124
rect 2691 32070 2693 32122
rect 2873 32070 2875 32122
rect 2629 32068 2635 32070
rect 2691 32068 2715 32070
rect 2771 32068 2795 32070
rect 2851 32068 2875 32070
rect 2931 32068 2937 32070
rect 2629 32059 2937 32068
rect 2629 31036 2937 31045
rect 2629 31034 2635 31036
rect 2691 31034 2715 31036
rect 2771 31034 2795 31036
rect 2851 31034 2875 31036
rect 2931 31034 2937 31036
rect 2691 30982 2693 31034
rect 2873 30982 2875 31034
rect 2629 30980 2635 30982
rect 2691 30980 2715 30982
rect 2771 30980 2795 30982
rect 2851 30980 2875 30982
rect 2931 30980 2937 30982
rect 2629 30971 2937 30980
rect 2629 29948 2937 29957
rect 2629 29946 2635 29948
rect 2691 29946 2715 29948
rect 2771 29946 2795 29948
rect 2851 29946 2875 29948
rect 2931 29946 2937 29948
rect 2691 29894 2693 29946
rect 2873 29894 2875 29946
rect 2629 29892 2635 29894
rect 2691 29892 2715 29894
rect 2771 29892 2795 29894
rect 2851 29892 2875 29894
rect 2931 29892 2937 29894
rect 2629 29883 2937 29892
rect 2136 29844 2188 29850
rect 2136 29786 2188 29792
rect 2044 29504 2096 29510
rect 2044 29446 2096 29452
rect 1952 28756 2004 28762
rect 1952 28698 2004 28704
rect 1860 27464 1912 27470
rect 1860 27406 1912 27412
rect 1688 19306 1808 19334
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1400 14476 1452 14482
rect 1400 14418 1452 14424
rect 1308 14408 1360 14414
rect 1308 14350 1360 14356
rect 848 13184 900 13190
rect 848 13126 900 13132
rect 860 12889 888 13126
rect 846 12880 902 12889
rect 1412 12850 1440 14418
rect 1596 13818 1624 14894
rect 1688 13938 1716 19306
rect 1872 17134 1900 27406
rect 1964 17490 1992 28698
rect 2056 17678 2084 29446
rect 2629 28860 2937 28869
rect 2629 28858 2635 28860
rect 2691 28858 2715 28860
rect 2771 28858 2795 28860
rect 2851 28858 2875 28860
rect 2931 28858 2937 28860
rect 2691 28806 2693 28858
rect 2873 28806 2875 28858
rect 2629 28804 2635 28806
rect 2691 28804 2715 28806
rect 2771 28804 2795 28806
rect 2851 28804 2875 28806
rect 2931 28804 2937 28806
rect 2629 28795 2937 28804
rect 2629 27772 2937 27781
rect 2629 27770 2635 27772
rect 2691 27770 2715 27772
rect 2771 27770 2795 27772
rect 2851 27770 2875 27772
rect 2931 27770 2937 27772
rect 2691 27718 2693 27770
rect 2873 27718 2875 27770
rect 2629 27716 2635 27718
rect 2691 27716 2715 27718
rect 2771 27716 2795 27718
rect 2851 27716 2875 27718
rect 2931 27716 2937 27718
rect 2629 27707 2937 27716
rect 3068 27606 3096 43250
rect 3160 42906 3188 43250
rect 3804 42906 3832 43250
rect 4356 42906 4384 43250
rect 5000 42906 5028 43250
rect 3148 42900 3200 42906
rect 3148 42842 3200 42848
rect 3792 42900 3844 42906
rect 3792 42842 3844 42848
rect 4344 42900 4396 42906
rect 4344 42842 4396 42848
rect 4988 42900 5040 42906
rect 4988 42842 5040 42848
rect 3424 42696 3476 42702
rect 3424 42638 3476 42644
rect 4068 42696 4120 42702
rect 4068 42638 4120 42644
rect 4988 42696 5040 42702
rect 4988 42638 5040 42644
rect 3056 27600 3108 27606
rect 3056 27542 3108 27548
rect 2688 27464 2740 27470
rect 2688 27406 2740 27412
rect 2700 27130 2728 27406
rect 2688 27124 2740 27130
rect 2688 27066 2740 27072
rect 2629 26684 2937 26693
rect 2629 26682 2635 26684
rect 2691 26682 2715 26684
rect 2771 26682 2795 26684
rect 2851 26682 2875 26684
rect 2931 26682 2937 26684
rect 2691 26630 2693 26682
rect 2873 26630 2875 26682
rect 2629 26628 2635 26630
rect 2691 26628 2715 26630
rect 2771 26628 2795 26630
rect 2851 26628 2875 26630
rect 2931 26628 2937 26630
rect 2629 26619 2937 26628
rect 2629 25596 2937 25605
rect 2629 25594 2635 25596
rect 2691 25594 2715 25596
rect 2771 25594 2795 25596
rect 2851 25594 2875 25596
rect 2931 25594 2937 25596
rect 2691 25542 2693 25594
rect 2873 25542 2875 25594
rect 2629 25540 2635 25542
rect 2691 25540 2715 25542
rect 2771 25540 2795 25542
rect 2851 25540 2875 25542
rect 2931 25540 2937 25542
rect 2629 25531 2937 25540
rect 2629 24508 2937 24517
rect 2629 24506 2635 24508
rect 2691 24506 2715 24508
rect 2771 24506 2795 24508
rect 2851 24506 2875 24508
rect 2931 24506 2937 24508
rect 2691 24454 2693 24506
rect 2873 24454 2875 24506
rect 2629 24452 2635 24454
rect 2691 24452 2715 24454
rect 2771 24452 2795 24454
rect 2851 24452 2875 24454
rect 2931 24452 2937 24454
rect 2629 24443 2937 24452
rect 2629 23420 2937 23429
rect 2629 23418 2635 23420
rect 2691 23418 2715 23420
rect 2771 23418 2795 23420
rect 2851 23418 2875 23420
rect 2931 23418 2937 23420
rect 2691 23366 2693 23418
rect 2873 23366 2875 23418
rect 2629 23364 2635 23366
rect 2691 23364 2715 23366
rect 2771 23364 2795 23366
rect 2851 23364 2875 23366
rect 2931 23364 2937 23366
rect 2629 23355 2937 23364
rect 2504 23316 2556 23322
rect 2504 23258 2556 23264
rect 2320 21888 2372 21894
rect 2320 21830 2372 21836
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 1964 17462 2084 17490
rect 1860 17128 1912 17134
rect 1860 17070 1912 17076
rect 2056 16946 2084 17462
rect 2136 17128 2188 17134
rect 2136 17070 2188 17076
rect 2332 17082 2360 21830
rect 2412 17536 2464 17542
rect 2412 17478 2464 17484
rect 2424 17338 2452 17478
rect 2412 17332 2464 17338
rect 2412 17274 2464 17280
rect 2410 17096 2466 17105
rect 1964 16918 2084 16946
rect 1964 16250 1992 16918
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 2148 14906 2176 17070
rect 2332 17054 2410 17082
rect 2410 17031 2466 17040
rect 2516 15910 2544 23258
rect 2629 22332 2937 22341
rect 2629 22330 2635 22332
rect 2691 22330 2715 22332
rect 2771 22330 2795 22332
rect 2851 22330 2875 22332
rect 2931 22330 2937 22332
rect 2691 22278 2693 22330
rect 2873 22278 2875 22330
rect 2629 22276 2635 22278
rect 2691 22276 2715 22278
rect 2771 22276 2795 22278
rect 2851 22276 2875 22278
rect 2931 22276 2937 22278
rect 2629 22267 2937 22276
rect 3436 22094 3464 42638
rect 3608 42628 3660 42634
rect 3608 42570 3660 42576
rect 3516 23860 3568 23866
rect 3516 23802 3568 23808
rect 3252 22066 3464 22094
rect 2629 21244 2937 21253
rect 2629 21242 2635 21244
rect 2691 21242 2715 21244
rect 2771 21242 2795 21244
rect 2851 21242 2875 21244
rect 2931 21242 2937 21244
rect 2691 21190 2693 21242
rect 2873 21190 2875 21242
rect 2629 21188 2635 21190
rect 2691 21188 2715 21190
rect 2771 21188 2795 21190
rect 2851 21188 2875 21190
rect 2931 21188 2937 21190
rect 2629 21179 2937 21188
rect 3252 21146 3280 22066
rect 3240 21140 3292 21146
rect 3240 21082 3292 21088
rect 3056 20936 3108 20942
rect 3056 20878 3108 20884
rect 2629 20156 2937 20165
rect 2629 20154 2635 20156
rect 2691 20154 2715 20156
rect 2771 20154 2795 20156
rect 2851 20154 2875 20156
rect 2931 20154 2937 20156
rect 2691 20102 2693 20154
rect 2873 20102 2875 20154
rect 2629 20100 2635 20102
rect 2691 20100 2715 20102
rect 2771 20100 2795 20102
rect 2851 20100 2875 20102
rect 2931 20100 2937 20102
rect 2629 20091 2937 20100
rect 2629 19068 2937 19077
rect 2629 19066 2635 19068
rect 2691 19066 2715 19068
rect 2771 19066 2795 19068
rect 2851 19066 2875 19068
rect 2931 19066 2937 19068
rect 2691 19014 2693 19066
rect 2873 19014 2875 19066
rect 2629 19012 2635 19014
rect 2691 19012 2715 19014
rect 2771 19012 2795 19014
rect 2851 19012 2875 19014
rect 2931 19012 2937 19014
rect 2629 19003 2937 19012
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 2629 17980 2937 17989
rect 2629 17978 2635 17980
rect 2691 17978 2715 17980
rect 2771 17978 2795 17980
rect 2851 17978 2875 17980
rect 2931 17978 2937 17980
rect 2691 17926 2693 17978
rect 2873 17926 2875 17978
rect 2629 17924 2635 17926
rect 2691 17924 2715 17926
rect 2771 17924 2795 17926
rect 2851 17924 2875 17926
rect 2931 17924 2937 17926
rect 2629 17915 2937 17924
rect 2629 16892 2937 16901
rect 2629 16890 2635 16892
rect 2691 16890 2715 16892
rect 2771 16890 2795 16892
rect 2851 16890 2875 16892
rect 2931 16890 2937 16892
rect 2691 16838 2693 16890
rect 2873 16838 2875 16890
rect 2629 16836 2635 16838
rect 2691 16836 2715 16838
rect 2771 16836 2795 16838
rect 2851 16836 2875 16838
rect 2931 16836 2937 16838
rect 2629 16827 2937 16836
rect 2412 15904 2464 15910
rect 2412 15846 2464 15852
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2424 15094 2452 15846
rect 2629 15804 2937 15813
rect 2629 15802 2635 15804
rect 2691 15802 2715 15804
rect 2771 15802 2795 15804
rect 2851 15802 2875 15804
rect 2931 15802 2937 15804
rect 2691 15750 2693 15802
rect 2873 15750 2875 15802
rect 2629 15748 2635 15750
rect 2691 15748 2715 15750
rect 2771 15748 2795 15750
rect 2851 15748 2875 15750
rect 2931 15748 2937 15750
rect 2629 15739 2937 15748
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 1780 14878 2176 14906
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1596 13790 1716 13818
rect 1584 13728 1636 13734
rect 1582 13696 1584 13705
rect 1636 13696 1638 13705
rect 1582 13631 1638 13640
rect 1688 12986 1716 13790
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 846 12815 902 12824
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 848 12096 900 12102
rect 846 12064 848 12073
rect 900 12064 902 12073
rect 846 11999 902 12008
rect 848 11552 900 11558
rect 848 11494 900 11500
rect 860 11257 888 11494
rect 846 11248 902 11257
rect 846 11183 902 11192
rect 848 10464 900 10470
rect 846 10432 848 10441
rect 900 10432 902 10441
rect 846 10367 902 10376
rect 1412 10062 1440 12786
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 10810 1532 11698
rect 1492 10804 1544 10810
rect 1492 10746 1544 10752
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9518 1440 9998
rect 1780 9654 1808 14878
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1964 14074 1992 14758
rect 2629 14716 2937 14725
rect 2629 14714 2635 14716
rect 2691 14714 2715 14716
rect 2771 14714 2795 14716
rect 2851 14714 2875 14716
rect 2931 14714 2937 14716
rect 2691 14662 2693 14714
rect 2873 14662 2875 14714
rect 2629 14660 2635 14662
rect 2691 14660 2715 14662
rect 2771 14660 2795 14662
rect 2851 14660 2875 14662
rect 2931 14660 2937 14662
rect 2629 14651 2937 14660
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1860 13932 1912 13938
rect 1860 13874 1912 13880
rect 1872 10713 1900 13874
rect 2424 13326 2452 14214
rect 2629 13628 2937 13637
rect 2629 13626 2635 13628
rect 2691 13626 2715 13628
rect 2771 13626 2795 13628
rect 2851 13626 2875 13628
rect 2931 13626 2937 13628
rect 2691 13574 2693 13626
rect 2873 13574 2875 13626
rect 2629 13572 2635 13574
rect 2691 13572 2715 13574
rect 2771 13572 2795 13574
rect 2851 13572 2875 13574
rect 2931 13572 2937 13574
rect 2629 13563 2937 13572
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2412 12640 2464 12646
rect 2412 12582 2464 12588
rect 2424 12238 2452 12582
rect 2629 12540 2937 12549
rect 2629 12538 2635 12540
rect 2691 12538 2715 12540
rect 2771 12538 2795 12540
rect 2851 12538 2875 12540
rect 2931 12538 2937 12540
rect 2691 12486 2693 12538
rect 2873 12486 2875 12538
rect 2629 12484 2635 12486
rect 2691 12484 2715 12486
rect 2771 12484 2795 12486
rect 2851 12484 2875 12486
rect 2931 12484 2937 12486
rect 2629 12475 2937 12484
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2629 11452 2937 11461
rect 2629 11450 2635 11452
rect 2691 11450 2715 11452
rect 2771 11450 2795 11452
rect 2851 11450 2875 11452
rect 2931 11450 2937 11452
rect 2691 11398 2693 11450
rect 2873 11398 2875 11450
rect 2629 11396 2635 11398
rect 2691 11396 2715 11398
rect 2771 11396 2795 11398
rect 2851 11396 2875 11398
rect 2931 11396 2937 11398
rect 2629 11387 2937 11396
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 1858 10704 1914 10713
rect 2148 10674 2176 10950
rect 1858 10639 1914 10648
rect 2044 10668 2096 10674
rect 1872 9994 1900 10639
rect 2044 10610 2096 10616
rect 2136 10668 2188 10674
rect 2136 10610 2188 10616
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 1400 9512 1452 9518
rect 1400 9454 1452 9460
rect 848 8832 900 8838
rect 846 8800 848 8809
rect 900 8800 902 8809
rect 846 8735 902 8744
rect 1412 7886 1440 9454
rect 1780 9178 1808 9590
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 2056 8974 2084 10610
rect 2629 10364 2937 10373
rect 2629 10362 2635 10364
rect 2691 10362 2715 10364
rect 2771 10362 2795 10364
rect 2851 10362 2875 10364
rect 2931 10362 2937 10364
rect 2691 10310 2693 10362
rect 2873 10310 2875 10362
rect 2629 10308 2635 10310
rect 2691 10308 2715 10310
rect 2771 10308 2795 10310
rect 2851 10308 2875 10310
rect 2931 10308 2937 10310
rect 2629 10299 2937 10308
rect 2976 10266 3004 18226
rect 3068 17610 3096 20878
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 3424 16584 3476 16590
rect 3424 16526 3476 16532
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2504 9920 2556 9926
rect 2504 9862 2556 9868
rect 2412 9376 2464 9382
rect 2412 9318 2464 9324
rect 2424 9110 2452 9318
rect 2412 9104 2464 9110
rect 2412 9046 2464 9052
rect 2516 8974 2544 9862
rect 2792 9625 2820 9998
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2629 9276 2937 9285
rect 2629 9274 2635 9276
rect 2691 9274 2715 9276
rect 2771 9274 2795 9276
rect 2851 9274 2875 9276
rect 2931 9274 2937 9276
rect 2691 9222 2693 9274
rect 2873 9222 2875 9274
rect 2629 9220 2635 9222
rect 2691 9220 2715 9222
rect 2771 9220 2795 9222
rect 2851 9220 2875 9222
rect 2931 9220 2937 9222
rect 2629 9211 2937 9220
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2596 8968 2648 8974
rect 2596 8910 2648 8916
rect 2320 8832 2372 8838
rect 2320 8774 2372 8780
rect 2332 8634 2360 8774
rect 2608 8634 2636 8910
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 1676 8356 1728 8362
rect 1676 8298 1728 8304
rect 1688 8265 1716 8298
rect 1674 8256 1730 8265
rect 1674 8191 1730 8200
rect 2629 8188 2937 8197
rect 2629 8186 2635 8188
rect 2691 8186 2715 8188
rect 2771 8186 2795 8188
rect 2851 8186 2875 8188
rect 2931 8186 2937 8188
rect 2691 8134 2693 8186
rect 2873 8134 2875 8186
rect 2629 8132 2635 8134
rect 2691 8132 2715 8134
rect 2771 8132 2795 8134
rect 2851 8132 2875 8134
rect 2931 8132 2937 8134
rect 2629 8123 2937 8132
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 848 7200 900 7206
rect 846 7168 848 7177
rect 900 7168 902 7177
rect 846 7103 902 7112
rect 848 6656 900 6662
rect 848 6598 900 6604
rect 860 6361 888 6598
rect 846 6352 902 6361
rect 846 6287 902 6296
rect 1412 6254 1440 7822
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7546 2452 7686
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2629 7100 2937 7109
rect 2629 7098 2635 7100
rect 2691 7098 2715 7100
rect 2771 7098 2795 7100
rect 2851 7098 2875 7100
rect 2931 7098 2937 7100
rect 2691 7046 2693 7098
rect 2873 7046 2875 7098
rect 2629 7044 2635 7046
rect 2691 7044 2715 7046
rect 2771 7044 2795 7046
rect 2851 7044 2875 7046
rect 2931 7044 2937 7046
rect 2629 7035 2937 7044
rect 1492 6724 1544 6730
rect 1492 6666 1544 6672
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1504 5914 1532 6666
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1584 5568 1636 5574
rect 1582 5536 1584 5545
rect 1636 5536 1638 5545
rect 1582 5471 1638 5480
rect 848 5024 900 5030
rect 848 4966 900 4972
rect 860 4729 888 4966
rect 846 4720 902 4729
rect 846 4655 902 4664
rect 756 4140 808 4146
rect 756 4082 808 4088
rect 768 3913 796 4082
rect 754 3904 810 3913
rect 754 3839 810 3848
rect 2044 1964 2096 1970
rect 1964 1924 2044 1952
rect 1216 1352 1268 1358
rect 1216 1294 1268 1300
rect 1228 160 1256 1294
rect 1964 160 1992 1924
rect 2044 1906 2096 1912
rect 2332 1290 2360 6054
rect 2424 5914 2452 6054
rect 2629 6012 2937 6021
rect 2629 6010 2635 6012
rect 2691 6010 2715 6012
rect 2771 6010 2795 6012
rect 2851 6010 2875 6012
rect 2931 6010 2937 6012
rect 2691 5958 2693 6010
rect 2873 5958 2875 6010
rect 2629 5956 2635 5958
rect 2691 5956 2715 5958
rect 2771 5956 2795 5958
rect 2851 5956 2875 5958
rect 2931 5956 2937 5958
rect 2629 5947 2937 5956
rect 2412 5908 2464 5914
rect 2412 5850 2464 5856
rect 2596 5704 2648 5710
rect 2516 5664 2596 5692
rect 2516 1358 2544 5664
rect 2596 5646 2648 5652
rect 2629 4924 2937 4933
rect 2629 4922 2635 4924
rect 2691 4922 2715 4924
rect 2771 4922 2795 4924
rect 2851 4922 2875 4924
rect 2931 4922 2937 4924
rect 2691 4870 2693 4922
rect 2873 4870 2875 4922
rect 2629 4868 2635 4870
rect 2691 4868 2715 4870
rect 2771 4868 2795 4870
rect 2851 4868 2875 4870
rect 2931 4868 2937 4870
rect 2629 4859 2937 4868
rect 3436 3942 3464 16526
rect 3528 16522 3556 23802
rect 3620 18329 3648 42570
rect 4080 42362 4108 42638
rect 4308 42460 4616 42469
rect 4308 42458 4314 42460
rect 4370 42458 4394 42460
rect 4450 42458 4474 42460
rect 4530 42458 4554 42460
rect 4610 42458 4616 42460
rect 4370 42406 4372 42458
rect 4552 42406 4554 42458
rect 4308 42404 4314 42406
rect 4370 42404 4394 42406
rect 4450 42404 4474 42406
rect 4530 42404 4554 42406
rect 4610 42404 4616 42406
rect 4308 42395 4616 42404
rect 5000 42362 5028 42638
rect 4068 42356 4120 42362
rect 4068 42298 4120 42304
rect 4988 42356 5040 42362
rect 4988 42298 5040 42304
rect 3976 42288 4028 42294
rect 3976 42230 4028 42236
rect 3700 36372 3752 36378
rect 3700 36314 3752 36320
rect 3712 19378 3740 36314
rect 3792 31136 3844 31142
rect 3792 31078 3844 31084
rect 3804 29646 3832 31078
rect 3792 29640 3844 29646
rect 3792 29582 3844 29588
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3698 18728 3754 18737
rect 3698 18663 3754 18672
rect 3712 18358 3740 18663
rect 3700 18352 3752 18358
rect 3606 18320 3662 18329
rect 3700 18294 3752 18300
rect 3606 18255 3662 18264
rect 3516 16516 3568 16522
rect 3516 16458 3568 16464
rect 3804 12986 3832 29582
rect 3884 27600 3936 27606
rect 3884 27542 3936 27548
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3896 10577 3924 27542
rect 3988 17105 4016 42230
rect 4252 42220 4304 42226
rect 4252 42162 4304 42168
rect 4896 42220 4948 42226
rect 4896 42162 4948 42168
rect 4264 41585 4292 42162
rect 4250 41576 4306 41585
rect 4250 41511 4306 41520
rect 4908 41449 4936 42162
rect 4894 41440 4950 41449
rect 4308 41372 4616 41381
rect 4894 41375 4950 41384
rect 4308 41370 4314 41372
rect 4370 41370 4394 41372
rect 4450 41370 4474 41372
rect 4530 41370 4554 41372
rect 4610 41370 4616 41372
rect 4370 41318 4372 41370
rect 4552 41318 4554 41370
rect 4308 41316 4314 41318
rect 4370 41316 4394 41318
rect 4450 41316 4474 41318
rect 4530 41316 4554 41318
rect 4610 41316 4616 41318
rect 4308 41307 4616 41316
rect 4308 40284 4616 40293
rect 4308 40282 4314 40284
rect 4370 40282 4394 40284
rect 4450 40282 4474 40284
rect 4530 40282 4554 40284
rect 4610 40282 4616 40284
rect 4370 40230 4372 40282
rect 4552 40230 4554 40282
rect 4308 40228 4314 40230
rect 4370 40228 4394 40230
rect 4450 40228 4474 40230
rect 4530 40228 4554 40230
rect 4610 40228 4616 40230
rect 4308 40219 4616 40228
rect 4712 39908 4764 39914
rect 4712 39850 4764 39856
rect 4724 39438 4752 39850
rect 4712 39432 4764 39438
rect 4712 39374 4764 39380
rect 4308 39196 4616 39205
rect 4308 39194 4314 39196
rect 4370 39194 4394 39196
rect 4450 39194 4474 39196
rect 4530 39194 4554 39196
rect 4610 39194 4616 39196
rect 4370 39142 4372 39194
rect 4552 39142 4554 39194
rect 4308 39140 4314 39142
rect 4370 39140 4394 39142
rect 4450 39140 4474 39142
rect 4530 39140 4554 39142
rect 4610 39140 4616 39142
rect 4308 39131 4616 39140
rect 4308 38108 4616 38117
rect 4308 38106 4314 38108
rect 4370 38106 4394 38108
rect 4450 38106 4474 38108
rect 4530 38106 4554 38108
rect 4610 38106 4616 38108
rect 4370 38054 4372 38106
rect 4552 38054 4554 38106
rect 4308 38052 4314 38054
rect 4370 38052 4394 38054
rect 4450 38052 4474 38054
rect 4530 38052 4554 38054
rect 4610 38052 4616 38054
rect 4308 38043 4616 38052
rect 4308 37020 4616 37029
rect 4308 37018 4314 37020
rect 4370 37018 4394 37020
rect 4450 37018 4474 37020
rect 4530 37018 4554 37020
rect 4610 37018 4616 37020
rect 4370 36966 4372 37018
rect 4552 36966 4554 37018
rect 4308 36964 4314 36966
rect 4370 36964 4394 36966
rect 4450 36964 4474 36966
rect 4530 36964 4554 36966
rect 4610 36964 4616 36966
rect 4308 36955 4616 36964
rect 4308 35932 4616 35941
rect 4308 35930 4314 35932
rect 4370 35930 4394 35932
rect 4450 35930 4474 35932
rect 4530 35930 4554 35932
rect 4610 35930 4616 35932
rect 4370 35878 4372 35930
rect 4552 35878 4554 35930
rect 4308 35876 4314 35878
rect 4370 35876 4394 35878
rect 4450 35876 4474 35878
rect 4530 35876 4554 35878
rect 4610 35876 4616 35878
rect 4308 35867 4616 35876
rect 4308 34844 4616 34853
rect 4308 34842 4314 34844
rect 4370 34842 4394 34844
rect 4450 34842 4474 34844
rect 4530 34842 4554 34844
rect 4610 34842 4616 34844
rect 4370 34790 4372 34842
rect 4552 34790 4554 34842
rect 4308 34788 4314 34790
rect 4370 34788 4394 34790
rect 4450 34788 4474 34790
rect 4530 34788 4554 34790
rect 4610 34788 4616 34790
rect 4308 34779 4616 34788
rect 4308 33756 4616 33765
rect 4308 33754 4314 33756
rect 4370 33754 4394 33756
rect 4450 33754 4474 33756
rect 4530 33754 4554 33756
rect 4610 33754 4616 33756
rect 4370 33702 4372 33754
rect 4552 33702 4554 33754
rect 4308 33700 4314 33702
rect 4370 33700 4394 33702
rect 4450 33700 4474 33702
rect 4530 33700 4554 33702
rect 4610 33700 4616 33702
rect 4308 33691 4616 33700
rect 4308 32668 4616 32677
rect 4308 32666 4314 32668
rect 4370 32666 4394 32668
rect 4450 32666 4474 32668
rect 4530 32666 4554 32668
rect 4610 32666 4616 32668
rect 4370 32614 4372 32666
rect 4552 32614 4554 32666
rect 4308 32612 4314 32614
rect 4370 32612 4394 32614
rect 4450 32612 4474 32614
rect 4530 32612 4554 32614
rect 4610 32612 4616 32614
rect 4308 32603 4616 32612
rect 4308 31580 4616 31589
rect 4308 31578 4314 31580
rect 4370 31578 4394 31580
rect 4450 31578 4474 31580
rect 4530 31578 4554 31580
rect 4610 31578 4616 31580
rect 4370 31526 4372 31578
rect 4552 31526 4554 31578
rect 4308 31524 4314 31526
rect 4370 31524 4394 31526
rect 4450 31524 4474 31526
rect 4530 31524 4554 31526
rect 4610 31524 4616 31526
rect 4308 31515 4616 31524
rect 4308 30492 4616 30501
rect 4308 30490 4314 30492
rect 4370 30490 4394 30492
rect 4450 30490 4474 30492
rect 4530 30490 4554 30492
rect 4610 30490 4616 30492
rect 4370 30438 4372 30490
rect 4552 30438 4554 30490
rect 4308 30436 4314 30438
rect 4370 30436 4394 30438
rect 4450 30436 4474 30438
rect 4530 30436 4554 30438
rect 4610 30436 4616 30438
rect 4308 30427 4616 30436
rect 4308 29404 4616 29413
rect 4308 29402 4314 29404
rect 4370 29402 4394 29404
rect 4450 29402 4474 29404
rect 4530 29402 4554 29404
rect 4610 29402 4616 29404
rect 4370 29350 4372 29402
rect 4552 29350 4554 29402
rect 4308 29348 4314 29350
rect 4370 29348 4394 29350
rect 4450 29348 4474 29350
rect 4530 29348 4554 29350
rect 4610 29348 4616 29350
rect 4308 29339 4616 29348
rect 4308 28316 4616 28325
rect 4308 28314 4314 28316
rect 4370 28314 4394 28316
rect 4450 28314 4474 28316
rect 4530 28314 4554 28316
rect 4610 28314 4616 28316
rect 4370 28262 4372 28314
rect 4552 28262 4554 28314
rect 4308 28260 4314 28262
rect 4370 28260 4394 28262
rect 4450 28260 4474 28262
rect 4530 28260 4554 28262
rect 4610 28260 4616 28262
rect 4308 28251 4616 28260
rect 4066 27976 4122 27985
rect 4066 27911 4122 27920
rect 3974 17096 4030 17105
rect 3974 17031 4030 17040
rect 4080 13190 4108 27911
rect 4308 27228 4616 27237
rect 4308 27226 4314 27228
rect 4370 27226 4394 27228
rect 4450 27226 4474 27228
rect 4530 27226 4554 27228
rect 4610 27226 4616 27228
rect 4370 27174 4372 27226
rect 4552 27174 4554 27226
rect 4308 27172 4314 27174
rect 4370 27172 4394 27174
rect 4450 27172 4474 27174
rect 4530 27172 4554 27174
rect 4610 27172 4616 27174
rect 4308 27163 4616 27172
rect 4160 26988 4212 26994
rect 4160 26930 4212 26936
rect 4172 24750 4200 26930
rect 4308 26140 4616 26149
rect 4308 26138 4314 26140
rect 4370 26138 4394 26140
rect 4450 26138 4474 26140
rect 4530 26138 4554 26140
rect 4610 26138 4616 26140
rect 4370 26086 4372 26138
rect 4552 26086 4554 26138
rect 4308 26084 4314 26086
rect 4370 26084 4394 26086
rect 4450 26084 4474 26086
rect 4530 26084 4554 26086
rect 4610 26084 4616 26086
rect 4308 26075 4616 26084
rect 4308 25052 4616 25061
rect 4308 25050 4314 25052
rect 4370 25050 4394 25052
rect 4450 25050 4474 25052
rect 4530 25050 4554 25052
rect 4610 25050 4616 25052
rect 4370 24998 4372 25050
rect 4552 24998 4554 25050
rect 4308 24996 4314 24998
rect 4370 24996 4394 24998
rect 4450 24996 4474 24998
rect 4530 24996 4554 24998
rect 4610 24996 4616 24998
rect 4308 24987 4616 24996
rect 4160 24744 4212 24750
rect 4160 24686 4212 24692
rect 4172 24274 4200 24686
rect 4160 24268 4212 24274
rect 4160 24210 4212 24216
rect 4724 24206 4752 39374
rect 5552 35290 5580 43268
rect 5724 43250 5776 43256
rect 6460 43308 6512 43314
rect 6460 43250 6512 43256
rect 7196 43308 7248 43314
rect 7196 43250 7248 43256
rect 7932 43308 7984 43314
rect 7932 43250 7984 43256
rect 8944 43308 8996 43314
rect 8944 43250 8996 43256
rect 9220 43308 9272 43314
rect 9220 43250 9272 43256
rect 10140 43308 10192 43314
rect 10140 43250 10192 43256
rect 10968 43308 11020 43314
rect 10968 43250 11020 43256
rect 11612 43308 11664 43314
rect 11612 43250 11664 43256
rect 12440 43308 12492 43314
rect 12440 43250 12492 43256
rect 13084 43308 13136 43314
rect 13084 43250 13136 43256
rect 13544 43308 13596 43314
rect 13544 43250 13596 43256
rect 5987 43004 6295 43013
rect 5987 43002 5993 43004
rect 6049 43002 6073 43004
rect 6129 43002 6153 43004
rect 6209 43002 6233 43004
rect 6289 43002 6295 43004
rect 6049 42950 6051 43002
rect 6231 42950 6233 43002
rect 5987 42948 5993 42950
rect 6049 42948 6073 42950
rect 6129 42948 6153 42950
rect 6209 42948 6233 42950
rect 6289 42948 6295 42950
rect 5987 42939 6295 42948
rect 6472 42906 6500 43250
rect 7208 42906 7236 43250
rect 7944 42906 7972 43250
rect 8956 42906 8984 43250
rect 9232 42906 9260 43250
rect 9345 43004 9653 43013
rect 9345 43002 9351 43004
rect 9407 43002 9431 43004
rect 9487 43002 9511 43004
rect 9567 43002 9591 43004
rect 9647 43002 9653 43004
rect 9407 42950 9409 43002
rect 9589 42950 9591 43002
rect 9345 42948 9351 42950
rect 9407 42948 9431 42950
rect 9487 42948 9511 42950
rect 9567 42948 9591 42950
rect 9647 42948 9653 42950
rect 9345 42939 9653 42948
rect 10152 42906 10180 43250
rect 10980 42906 11008 43250
rect 11624 42906 11652 43250
rect 12452 42906 12480 43250
rect 12703 43004 13011 43013
rect 12703 43002 12709 43004
rect 12765 43002 12789 43004
rect 12845 43002 12869 43004
rect 12925 43002 12949 43004
rect 13005 43002 13011 43004
rect 12765 42950 12767 43002
rect 12947 42950 12949 43002
rect 12703 42948 12709 42950
rect 12765 42948 12789 42950
rect 12845 42948 12869 42950
rect 12925 42948 12949 42950
rect 13005 42948 13011 42950
rect 12703 42939 13011 42948
rect 13096 42906 13124 43250
rect 6460 42900 6512 42906
rect 6460 42842 6512 42848
rect 7196 42900 7248 42906
rect 7196 42842 7248 42848
rect 7932 42900 7984 42906
rect 7932 42842 7984 42848
rect 8944 42900 8996 42906
rect 8944 42842 8996 42848
rect 9220 42900 9272 42906
rect 9220 42842 9272 42848
rect 10140 42900 10192 42906
rect 10140 42842 10192 42848
rect 10968 42900 11020 42906
rect 10968 42842 11020 42848
rect 11612 42900 11664 42906
rect 11612 42842 11664 42848
rect 12440 42900 12492 42906
rect 12440 42842 12492 42848
rect 13084 42900 13136 42906
rect 13084 42842 13136 42848
rect 10046 42800 10102 42809
rect 10046 42735 10102 42744
rect 10060 42702 10088 42735
rect 6460 42696 6512 42702
rect 6460 42638 6512 42644
rect 7196 42696 7248 42702
rect 7932 42696 7984 42702
rect 7196 42638 7248 42644
rect 7930 42664 7932 42673
rect 8668 42696 8720 42702
rect 7984 42664 7986 42673
rect 5632 42356 5684 42362
rect 5632 42298 5684 42304
rect 5540 35284 5592 35290
rect 5540 35226 5592 35232
rect 5356 34672 5408 34678
rect 5356 34614 5408 34620
rect 4988 34196 5040 34202
rect 4988 34138 5040 34144
rect 5000 33318 5028 34138
rect 4988 33312 5040 33318
rect 4988 33254 5040 33260
rect 4804 32292 4856 32298
rect 4804 32234 4856 32240
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4308 23964 4616 23973
rect 4308 23962 4314 23964
rect 4370 23962 4394 23964
rect 4450 23962 4474 23964
rect 4530 23962 4554 23964
rect 4610 23962 4616 23964
rect 4370 23910 4372 23962
rect 4552 23910 4554 23962
rect 4308 23908 4314 23910
rect 4370 23908 4394 23910
rect 4450 23908 4474 23910
rect 4530 23908 4554 23910
rect 4610 23908 4616 23910
rect 4308 23899 4616 23908
rect 4308 22876 4616 22885
rect 4308 22874 4314 22876
rect 4370 22874 4394 22876
rect 4450 22874 4474 22876
rect 4530 22874 4554 22876
rect 4610 22874 4616 22876
rect 4370 22822 4372 22874
rect 4552 22822 4554 22874
rect 4308 22820 4314 22822
rect 4370 22820 4394 22822
rect 4450 22820 4474 22822
rect 4530 22820 4554 22822
rect 4610 22820 4616 22822
rect 4308 22811 4616 22820
rect 4816 21894 4844 32234
rect 4896 26988 4948 26994
rect 4896 26930 4948 26936
rect 4908 26518 4936 26930
rect 4896 26512 4948 26518
rect 4896 26454 4948 26460
rect 4896 26376 4948 26382
rect 4896 26318 4948 26324
rect 4908 25362 4936 26318
rect 4896 25356 4948 25362
rect 4896 25298 4948 25304
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4308 21788 4616 21797
rect 4308 21786 4314 21788
rect 4370 21786 4394 21788
rect 4450 21786 4474 21788
rect 4530 21786 4554 21788
rect 4610 21786 4616 21788
rect 4370 21734 4372 21786
rect 4552 21734 4554 21786
rect 4308 21732 4314 21734
rect 4370 21732 4394 21734
rect 4450 21732 4474 21734
rect 4530 21732 4554 21734
rect 4610 21732 4616 21734
rect 4308 21723 4616 21732
rect 4528 21616 4580 21622
rect 4526 21584 4528 21593
rect 4580 21584 4582 21593
rect 4908 21554 4936 21966
rect 4896 21548 4948 21554
rect 4526 21519 4582 21528
rect 4724 21508 4896 21536
rect 4308 20700 4616 20709
rect 4308 20698 4314 20700
rect 4370 20698 4394 20700
rect 4450 20698 4474 20700
rect 4530 20698 4554 20700
rect 4610 20698 4616 20700
rect 4370 20646 4372 20698
rect 4552 20646 4554 20698
rect 4308 20644 4314 20646
rect 4370 20644 4394 20646
rect 4450 20644 4474 20646
rect 4530 20644 4554 20646
rect 4610 20644 4616 20646
rect 4308 20635 4616 20644
rect 4158 20496 4214 20505
rect 4158 20431 4214 20440
rect 4172 19854 4200 20431
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4172 18222 4200 19790
rect 4308 19612 4616 19621
rect 4308 19610 4314 19612
rect 4370 19610 4394 19612
rect 4450 19610 4474 19612
rect 4530 19610 4554 19612
rect 4610 19610 4616 19612
rect 4370 19558 4372 19610
rect 4552 19558 4554 19610
rect 4308 19556 4314 19558
rect 4370 19556 4394 19558
rect 4450 19556 4474 19558
rect 4530 19556 4554 19558
rect 4610 19556 4616 19558
rect 4308 19547 4616 19556
rect 4308 18524 4616 18533
rect 4308 18522 4314 18524
rect 4370 18522 4394 18524
rect 4450 18522 4474 18524
rect 4530 18522 4554 18524
rect 4610 18522 4616 18524
rect 4370 18470 4372 18522
rect 4552 18470 4554 18522
rect 4308 18468 4314 18470
rect 4370 18468 4394 18470
rect 4450 18468 4474 18470
rect 4530 18468 4554 18470
rect 4610 18468 4616 18470
rect 4308 18459 4616 18468
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 4160 18080 4212 18086
rect 4160 18022 4212 18028
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 3882 10568 3938 10577
rect 3882 10503 3938 10512
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 2629 3836 2937 3845
rect 2629 3834 2635 3836
rect 2691 3834 2715 3836
rect 2771 3834 2795 3836
rect 2851 3834 2875 3836
rect 2931 3834 2937 3836
rect 2691 3782 2693 3834
rect 2873 3782 2875 3834
rect 2629 3780 2635 3782
rect 2691 3780 2715 3782
rect 2771 3780 2795 3782
rect 2851 3780 2875 3782
rect 2931 3780 2937 3782
rect 2629 3771 2937 3780
rect 2629 2748 2937 2757
rect 2629 2746 2635 2748
rect 2691 2746 2715 2748
rect 2771 2746 2795 2748
rect 2851 2746 2875 2748
rect 2931 2746 2937 2748
rect 2691 2694 2693 2746
rect 2873 2694 2875 2746
rect 2629 2692 2635 2694
rect 2691 2692 2715 2694
rect 2771 2692 2795 2694
rect 2851 2692 2875 2694
rect 2931 2692 2937 2694
rect 2629 2683 2937 2692
rect 4172 1834 4200 18022
rect 4308 17436 4616 17445
rect 4308 17434 4314 17436
rect 4370 17434 4394 17436
rect 4450 17434 4474 17436
rect 4530 17434 4554 17436
rect 4610 17434 4616 17436
rect 4370 17382 4372 17434
rect 4552 17382 4554 17434
rect 4308 17380 4314 17382
rect 4370 17380 4394 17382
rect 4450 17380 4474 17382
rect 4530 17380 4554 17382
rect 4610 17380 4616 17382
rect 4308 17371 4616 17380
rect 4308 16348 4616 16357
rect 4308 16346 4314 16348
rect 4370 16346 4394 16348
rect 4450 16346 4474 16348
rect 4530 16346 4554 16348
rect 4610 16346 4616 16348
rect 4370 16294 4372 16346
rect 4552 16294 4554 16346
rect 4308 16292 4314 16294
rect 4370 16292 4394 16294
rect 4450 16292 4474 16294
rect 4530 16292 4554 16294
rect 4610 16292 4616 16294
rect 4308 16283 4616 16292
rect 4308 15260 4616 15269
rect 4308 15258 4314 15260
rect 4370 15258 4394 15260
rect 4450 15258 4474 15260
rect 4530 15258 4554 15260
rect 4610 15258 4616 15260
rect 4370 15206 4372 15258
rect 4552 15206 4554 15258
rect 4308 15204 4314 15206
rect 4370 15204 4394 15206
rect 4450 15204 4474 15206
rect 4530 15204 4554 15206
rect 4610 15204 4616 15206
rect 4308 15195 4616 15204
rect 4308 14172 4616 14181
rect 4308 14170 4314 14172
rect 4370 14170 4394 14172
rect 4450 14170 4474 14172
rect 4530 14170 4554 14172
rect 4610 14170 4616 14172
rect 4370 14118 4372 14170
rect 4552 14118 4554 14170
rect 4308 14116 4314 14118
rect 4370 14116 4394 14118
rect 4450 14116 4474 14118
rect 4530 14116 4554 14118
rect 4610 14116 4616 14118
rect 4308 14107 4616 14116
rect 4308 13084 4616 13093
rect 4308 13082 4314 13084
rect 4370 13082 4394 13084
rect 4450 13082 4474 13084
rect 4530 13082 4554 13084
rect 4610 13082 4616 13084
rect 4370 13030 4372 13082
rect 4552 13030 4554 13082
rect 4308 13028 4314 13030
rect 4370 13028 4394 13030
rect 4450 13028 4474 13030
rect 4530 13028 4554 13030
rect 4610 13028 4616 13030
rect 4308 13019 4616 13028
rect 4724 12442 4752 21508
rect 4896 21490 4948 21496
rect 4896 19780 4948 19786
rect 4896 19722 4948 19728
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4816 18290 4844 18566
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4908 16590 4936 19722
rect 5000 18873 5028 33254
rect 5172 26988 5224 26994
rect 5172 26930 5224 26936
rect 5184 26246 5212 26930
rect 5172 26240 5224 26246
rect 5172 26182 5224 26188
rect 5172 23656 5224 23662
rect 5172 23598 5224 23604
rect 5080 23588 5132 23594
rect 5080 23530 5132 23536
rect 5092 21690 5120 23530
rect 5080 21684 5132 21690
rect 5080 21626 5132 21632
rect 5184 20618 5212 23598
rect 5264 21548 5316 21554
rect 5264 21490 5316 21496
rect 5092 20590 5212 20618
rect 4986 18864 5042 18873
rect 4986 18799 5042 18808
rect 4988 18352 5040 18358
rect 4988 18294 5040 18300
rect 4896 16584 4948 16590
rect 4896 16526 4948 16532
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4724 12170 4752 12378
rect 4712 12164 4764 12170
rect 4712 12106 4764 12112
rect 4308 11996 4616 12005
rect 4308 11994 4314 11996
rect 4370 11994 4394 11996
rect 4450 11994 4474 11996
rect 4530 11994 4554 11996
rect 4610 11994 4616 11996
rect 4370 11942 4372 11994
rect 4552 11942 4554 11994
rect 4308 11940 4314 11942
rect 4370 11940 4394 11942
rect 4450 11940 4474 11942
rect 4530 11940 4554 11942
rect 4610 11940 4616 11942
rect 4308 11931 4616 11940
rect 4724 11762 4752 12106
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4308 10908 4616 10917
rect 4308 10906 4314 10908
rect 4370 10906 4394 10908
rect 4450 10906 4474 10908
rect 4530 10906 4554 10908
rect 4610 10906 4616 10908
rect 4370 10854 4372 10906
rect 4552 10854 4554 10906
rect 4308 10852 4314 10854
rect 4370 10852 4394 10854
rect 4450 10852 4474 10854
rect 4530 10852 4554 10854
rect 4610 10852 4616 10854
rect 4308 10843 4616 10852
rect 4724 10010 4752 11698
rect 4724 9982 4844 10010
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4308 9820 4616 9829
rect 4308 9818 4314 9820
rect 4370 9818 4394 9820
rect 4450 9818 4474 9820
rect 4530 9818 4554 9820
rect 4610 9818 4616 9820
rect 4370 9766 4372 9818
rect 4552 9766 4554 9818
rect 4308 9764 4314 9766
rect 4370 9764 4394 9766
rect 4450 9764 4474 9766
rect 4530 9764 4554 9766
rect 4610 9764 4616 9766
rect 4308 9755 4616 9764
rect 4308 8732 4616 8741
rect 4308 8730 4314 8732
rect 4370 8730 4394 8732
rect 4450 8730 4474 8732
rect 4530 8730 4554 8732
rect 4610 8730 4616 8732
rect 4370 8678 4372 8730
rect 4552 8678 4554 8730
rect 4308 8676 4314 8678
rect 4370 8676 4394 8678
rect 4450 8676 4474 8678
rect 4530 8676 4554 8678
rect 4610 8676 4616 8678
rect 4308 8667 4616 8676
rect 4308 7644 4616 7653
rect 4308 7642 4314 7644
rect 4370 7642 4394 7644
rect 4450 7642 4474 7644
rect 4530 7642 4554 7644
rect 4610 7642 4616 7644
rect 4370 7590 4372 7642
rect 4552 7590 4554 7642
rect 4308 7588 4314 7590
rect 4370 7588 4394 7590
rect 4450 7588 4474 7590
rect 4530 7588 4554 7590
rect 4610 7588 4616 7590
rect 4308 7579 4616 7588
rect 4308 6556 4616 6565
rect 4308 6554 4314 6556
rect 4370 6554 4394 6556
rect 4450 6554 4474 6556
rect 4530 6554 4554 6556
rect 4610 6554 4616 6556
rect 4370 6502 4372 6554
rect 4552 6502 4554 6554
rect 4308 6500 4314 6502
rect 4370 6500 4394 6502
rect 4450 6500 4474 6502
rect 4530 6500 4554 6502
rect 4610 6500 4616 6502
rect 4308 6491 4616 6500
rect 4308 5468 4616 5477
rect 4308 5466 4314 5468
rect 4370 5466 4394 5468
rect 4450 5466 4474 5468
rect 4530 5466 4554 5468
rect 4610 5466 4616 5468
rect 4370 5414 4372 5466
rect 4552 5414 4554 5466
rect 4308 5412 4314 5414
rect 4370 5412 4394 5414
rect 4450 5412 4474 5414
rect 4530 5412 4554 5414
rect 4610 5412 4616 5414
rect 4308 5403 4616 5412
rect 4724 5234 4752 9862
rect 4816 8974 4844 9982
rect 4804 8968 4856 8974
rect 4804 8910 4856 8916
rect 4816 8498 4844 8910
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 5000 4826 5028 18294
rect 5092 13938 5120 20590
rect 5172 20460 5224 20466
rect 5172 20402 5224 20408
rect 5184 19378 5212 20402
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5080 13796 5132 13802
rect 5080 13738 5132 13744
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4308 4380 4616 4389
rect 4308 4378 4314 4380
rect 4370 4378 4394 4380
rect 4450 4378 4474 4380
rect 4530 4378 4554 4380
rect 4610 4378 4616 4380
rect 4370 4326 4372 4378
rect 4552 4326 4554 4378
rect 4308 4324 4314 4326
rect 4370 4324 4394 4326
rect 4450 4324 4474 4326
rect 4530 4324 4554 4326
rect 4610 4324 4616 4326
rect 4308 4315 4616 4324
rect 5092 4010 5120 13738
rect 5184 12832 5212 19314
rect 5276 17134 5304 21490
rect 5368 17678 5396 34614
rect 5540 33448 5592 33454
rect 5540 33390 5592 33396
rect 5552 30054 5580 33390
rect 5540 30048 5592 30054
rect 5540 29990 5592 29996
rect 5552 29050 5580 29990
rect 5460 29022 5580 29050
rect 5460 27062 5488 29022
rect 5540 28960 5592 28966
rect 5540 28902 5592 28908
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5460 20534 5488 24142
rect 5552 24070 5580 28902
rect 5540 24064 5592 24070
rect 5540 24006 5592 24012
rect 5540 22636 5592 22642
rect 5540 22578 5592 22584
rect 5552 22030 5580 22578
rect 5540 22024 5592 22030
rect 5540 21966 5592 21972
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5552 20806 5580 21558
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5448 20528 5500 20534
rect 5448 20470 5500 20476
rect 5446 20360 5502 20369
rect 5446 20295 5502 20304
rect 5356 17672 5408 17678
rect 5356 17614 5408 17620
rect 5264 17128 5316 17134
rect 5264 17070 5316 17076
rect 5184 12804 5304 12832
rect 5276 9674 5304 12804
rect 5368 12646 5396 17614
rect 5460 13802 5488 20295
rect 5644 18086 5672 42298
rect 5987 41916 6295 41925
rect 5987 41914 5993 41916
rect 6049 41914 6073 41916
rect 6129 41914 6153 41916
rect 6209 41914 6233 41916
rect 6289 41914 6295 41916
rect 6049 41862 6051 41914
rect 6231 41862 6233 41914
rect 5987 41860 5993 41862
rect 6049 41860 6073 41862
rect 6129 41860 6153 41862
rect 6209 41860 6233 41862
rect 6289 41860 6295 41862
rect 5987 41851 6295 41860
rect 6472 41449 6500 42638
rect 7208 41721 7236 42638
rect 8668 42638 8720 42644
rect 10048 42696 10100 42702
rect 10048 42638 10100 42644
rect 12348 42696 12400 42702
rect 12348 42638 12400 42644
rect 7930 42599 7986 42608
rect 7666 42460 7974 42469
rect 7666 42458 7672 42460
rect 7728 42458 7752 42460
rect 7808 42458 7832 42460
rect 7888 42458 7912 42460
rect 7968 42458 7974 42460
rect 7728 42406 7730 42458
rect 7910 42406 7912 42458
rect 7666 42404 7672 42406
rect 7728 42404 7752 42406
rect 7808 42404 7832 42406
rect 7888 42404 7912 42406
rect 7968 42404 7974 42406
rect 7666 42395 7974 42404
rect 8680 42129 8708 42638
rect 10324 42560 10376 42566
rect 10324 42502 10376 42508
rect 10336 42294 10364 42502
rect 11024 42460 11332 42469
rect 11024 42458 11030 42460
rect 11086 42458 11110 42460
rect 11166 42458 11190 42460
rect 11246 42458 11270 42460
rect 11326 42458 11332 42460
rect 11086 42406 11088 42458
rect 11268 42406 11270 42458
rect 11024 42404 11030 42406
rect 11086 42404 11110 42406
rect 11166 42404 11190 42406
rect 11246 42404 11270 42406
rect 11326 42404 11332 42406
rect 11024 42395 11332 42404
rect 12360 42362 12388 42638
rect 13176 42628 13228 42634
rect 13176 42570 13228 42576
rect 12348 42356 12400 42362
rect 12348 42298 12400 42304
rect 10324 42288 10376 42294
rect 10324 42230 10376 42236
rect 8666 42120 8722 42129
rect 8666 42055 8722 42064
rect 9345 41916 9653 41925
rect 9345 41914 9351 41916
rect 9407 41914 9431 41916
rect 9487 41914 9511 41916
rect 9567 41914 9591 41916
rect 9647 41914 9653 41916
rect 9407 41862 9409 41914
rect 9589 41862 9591 41914
rect 9345 41860 9351 41862
rect 9407 41860 9431 41862
rect 9487 41860 9511 41862
rect 9567 41860 9591 41862
rect 9647 41860 9653 41862
rect 9345 41851 9653 41860
rect 12703 41916 13011 41925
rect 12703 41914 12709 41916
rect 12765 41914 12789 41916
rect 12845 41914 12869 41916
rect 12925 41914 12949 41916
rect 13005 41914 13011 41916
rect 12765 41862 12767 41914
rect 12947 41862 12949 41914
rect 12703 41860 12709 41862
rect 12765 41860 12789 41862
rect 12845 41860 12869 41862
rect 12925 41860 12949 41862
rect 13005 41860 13011 41862
rect 12703 41851 13011 41860
rect 13188 41818 13216 42570
rect 13556 42362 13584 43250
rect 13740 42362 13768 44540
rect 14476 43738 14504 44540
rect 14292 43710 14504 43738
rect 14292 42770 14320 43710
rect 14382 43548 14690 43557
rect 14382 43546 14388 43548
rect 14444 43546 14468 43548
rect 14524 43546 14548 43548
rect 14604 43546 14628 43548
rect 14684 43546 14690 43548
rect 14444 43494 14446 43546
rect 14626 43494 14628 43546
rect 14382 43492 14388 43494
rect 14444 43492 14468 43494
rect 14524 43492 14548 43494
rect 14604 43492 14628 43494
rect 14684 43492 14690 43494
rect 14382 43483 14690 43492
rect 15212 43450 15240 44540
rect 15200 43444 15252 43450
rect 15200 43386 15252 43392
rect 14280 42764 14332 42770
rect 14280 42706 14332 42712
rect 13820 42696 13872 42702
rect 13820 42638 13872 42644
rect 13544 42356 13596 42362
rect 13544 42298 13596 42304
rect 13728 42356 13780 42362
rect 13728 42298 13780 42304
rect 13728 42220 13780 42226
rect 13728 42162 13780 42168
rect 13740 41818 13768 42162
rect 13176 41812 13228 41818
rect 13176 41754 13228 41760
rect 13728 41812 13780 41818
rect 13728 41754 13780 41760
rect 7194 41712 7250 41721
rect 7194 41647 7250 41656
rect 13832 41585 13860 42638
rect 15568 42560 15620 42566
rect 15568 42502 15620 42508
rect 14382 42460 14690 42469
rect 14382 42458 14388 42460
rect 14444 42458 14468 42460
rect 14524 42458 14548 42460
rect 14604 42458 14628 42460
rect 14684 42458 14690 42460
rect 14444 42406 14446 42458
rect 14626 42406 14628 42458
rect 14382 42404 14388 42406
rect 14444 42404 14468 42406
rect 14524 42404 14548 42406
rect 14604 42404 14628 42406
rect 14684 42404 14690 42406
rect 14382 42395 14690 42404
rect 15476 42084 15528 42090
rect 15476 42026 15528 42032
rect 14740 41608 14792 41614
rect 13818 41576 13874 41585
rect 14740 41550 14792 41556
rect 13818 41511 13874 41520
rect 14004 41540 14056 41546
rect 14004 41482 14056 41488
rect 6458 41440 6514 41449
rect 6458 41375 6514 41384
rect 7666 41372 7974 41381
rect 7666 41370 7672 41372
rect 7728 41370 7752 41372
rect 7808 41370 7832 41372
rect 7888 41370 7912 41372
rect 7968 41370 7974 41372
rect 7728 41318 7730 41370
rect 7910 41318 7912 41370
rect 7666 41316 7672 41318
rect 7728 41316 7752 41318
rect 7808 41316 7832 41318
rect 7888 41316 7912 41318
rect 7968 41316 7974 41318
rect 7666 41307 7974 41316
rect 11024 41372 11332 41381
rect 11024 41370 11030 41372
rect 11086 41370 11110 41372
rect 11166 41370 11190 41372
rect 11246 41370 11270 41372
rect 11326 41370 11332 41372
rect 11086 41318 11088 41370
rect 11268 41318 11270 41370
rect 11024 41316 11030 41318
rect 11086 41316 11110 41318
rect 11166 41316 11190 41318
rect 11246 41316 11270 41318
rect 11326 41316 11332 41318
rect 11024 41307 11332 41316
rect 6368 40928 6420 40934
rect 6368 40870 6420 40876
rect 5987 40828 6295 40837
rect 5987 40826 5993 40828
rect 6049 40826 6073 40828
rect 6129 40826 6153 40828
rect 6209 40826 6233 40828
rect 6289 40826 6295 40828
rect 6049 40774 6051 40826
rect 6231 40774 6233 40826
rect 5987 40772 5993 40774
rect 6049 40772 6073 40774
rect 6129 40772 6153 40774
rect 6209 40772 6233 40774
rect 6289 40772 6295 40774
rect 5987 40763 6295 40772
rect 5987 39740 6295 39749
rect 5987 39738 5993 39740
rect 6049 39738 6073 39740
rect 6129 39738 6153 39740
rect 6209 39738 6233 39740
rect 6289 39738 6295 39740
rect 6049 39686 6051 39738
rect 6231 39686 6233 39738
rect 5987 39684 5993 39686
rect 6049 39684 6073 39686
rect 6129 39684 6153 39686
rect 6209 39684 6233 39686
rect 6289 39684 6295 39686
rect 5987 39675 6295 39684
rect 6380 39642 6408 40870
rect 9345 40828 9653 40837
rect 9345 40826 9351 40828
rect 9407 40826 9431 40828
rect 9487 40826 9511 40828
rect 9567 40826 9591 40828
rect 9647 40826 9653 40828
rect 9407 40774 9409 40826
rect 9589 40774 9591 40826
rect 9345 40772 9351 40774
rect 9407 40772 9431 40774
rect 9487 40772 9511 40774
rect 9567 40772 9591 40774
rect 9647 40772 9653 40774
rect 9345 40763 9653 40772
rect 12703 40828 13011 40837
rect 12703 40826 12709 40828
rect 12765 40826 12789 40828
rect 12845 40826 12869 40828
rect 12925 40826 12949 40828
rect 13005 40826 13011 40828
rect 12765 40774 12767 40826
rect 12947 40774 12949 40826
rect 12703 40772 12709 40774
rect 12765 40772 12789 40774
rect 12845 40772 12869 40774
rect 12925 40772 12949 40774
rect 13005 40772 13011 40774
rect 12703 40763 13011 40772
rect 7666 40284 7974 40293
rect 7666 40282 7672 40284
rect 7728 40282 7752 40284
rect 7808 40282 7832 40284
rect 7888 40282 7912 40284
rect 7968 40282 7974 40284
rect 7728 40230 7730 40282
rect 7910 40230 7912 40282
rect 7666 40228 7672 40230
rect 7728 40228 7752 40230
rect 7808 40228 7832 40230
rect 7888 40228 7912 40230
rect 7968 40228 7974 40230
rect 7666 40219 7974 40228
rect 11024 40284 11332 40293
rect 11024 40282 11030 40284
rect 11086 40282 11110 40284
rect 11166 40282 11190 40284
rect 11246 40282 11270 40284
rect 11326 40282 11332 40284
rect 11086 40230 11088 40282
rect 11268 40230 11270 40282
rect 11024 40228 11030 40230
rect 11086 40228 11110 40230
rect 11166 40228 11190 40230
rect 11246 40228 11270 40230
rect 11326 40228 11332 40230
rect 11024 40219 11332 40228
rect 7472 40044 7524 40050
rect 7472 39986 7524 39992
rect 13820 40044 13872 40050
rect 13820 39986 13872 39992
rect 6368 39636 6420 39642
rect 6368 39578 6420 39584
rect 6736 39636 6788 39642
rect 6736 39578 6788 39584
rect 5987 38652 6295 38661
rect 5987 38650 5993 38652
rect 6049 38650 6073 38652
rect 6129 38650 6153 38652
rect 6209 38650 6233 38652
rect 6289 38650 6295 38652
rect 6049 38598 6051 38650
rect 6231 38598 6233 38650
rect 6748 38654 6776 39578
rect 7484 39370 7512 39986
rect 13268 39840 13320 39846
rect 13268 39782 13320 39788
rect 9345 39740 9653 39749
rect 9345 39738 9351 39740
rect 9407 39738 9431 39740
rect 9487 39738 9511 39740
rect 9567 39738 9591 39740
rect 9647 39738 9653 39740
rect 9407 39686 9409 39738
rect 9589 39686 9591 39738
rect 9345 39684 9351 39686
rect 9407 39684 9431 39686
rect 9487 39684 9511 39686
rect 9567 39684 9591 39686
rect 9647 39684 9653 39686
rect 9345 39675 9653 39684
rect 12703 39740 13011 39749
rect 12703 39738 12709 39740
rect 12765 39738 12789 39740
rect 12845 39738 12869 39740
rect 12925 39738 12949 39740
rect 13005 39738 13011 39740
rect 12765 39686 12767 39738
rect 12947 39686 12949 39738
rect 12703 39684 12709 39686
rect 12765 39684 12789 39686
rect 12845 39684 12869 39686
rect 12925 39684 12949 39686
rect 13005 39684 13011 39686
rect 12703 39675 13011 39684
rect 12900 39432 12952 39438
rect 12900 39374 12952 39380
rect 7472 39364 7524 39370
rect 7472 39306 7524 39312
rect 6748 38626 6868 38654
rect 5987 38596 5993 38598
rect 6049 38596 6073 38598
rect 6129 38596 6153 38598
rect 6209 38596 6233 38598
rect 6289 38596 6295 38598
rect 5987 38587 6295 38596
rect 5987 37564 6295 37573
rect 5987 37562 5993 37564
rect 6049 37562 6073 37564
rect 6129 37562 6153 37564
rect 6209 37562 6233 37564
rect 6289 37562 6295 37564
rect 6049 37510 6051 37562
rect 6231 37510 6233 37562
rect 5987 37508 5993 37510
rect 6049 37508 6073 37510
rect 6129 37508 6153 37510
rect 6209 37508 6233 37510
rect 6289 37508 6295 37510
rect 5987 37499 6295 37508
rect 5987 36476 6295 36485
rect 5987 36474 5993 36476
rect 6049 36474 6073 36476
rect 6129 36474 6153 36476
rect 6209 36474 6233 36476
rect 6289 36474 6295 36476
rect 6049 36422 6051 36474
rect 6231 36422 6233 36474
rect 5987 36420 5993 36422
rect 6049 36420 6073 36422
rect 6129 36420 6153 36422
rect 6209 36420 6233 36422
rect 6289 36420 6295 36422
rect 5987 36411 6295 36420
rect 6458 35592 6514 35601
rect 6458 35527 6514 35536
rect 5987 35388 6295 35397
rect 5987 35386 5993 35388
rect 6049 35386 6073 35388
rect 6129 35386 6153 35388
rect 6209 35386 6233 35388
rect 6289 35386 6295 35388
rect 6049 35334 6051 35386
rect 6231 35334 6233 35386
rect 5987 35332 5993 35334
rect 6049 35332 6073 35334
rect 6129 35332 6153 35334
rect 6209 35332 6233 35334
rect 6289 35332 6295 35334
rect 5987 35323 6295 35332
rect 5724 35080 5776 35086
rect 5724 35022 5776 35028
rect 5736 34746 5764 35022
rect 6472 34950 6500 35527
rect 6460 34944 6512 34950
rect 6460 34886 6512 34892
rect 5724 34740 5776 34746
rect 5724 34682 5776 34688
rect 5722 34640 5778 34649
rect 5722 34575 5724 34584
rect 5776 34575 5778 34584
rect 5724 34546 5776 34552
rect 5987 34300 6295 34309
rect 5987 34298 5993 34300
rect 6049 34298 6073 34300
rect 6129 34298 6153 34300
rect 6209 34298 6233 34300
rect 6289 34298 6295 34300
rect 6049 34246 6051 34298
rect 6231 34246 6233 34298
rect 5987 34244 5993 34246
rect 6049 34244 6073 34246
rect 6129 34244 6153 34246
rect 6209 34244 6233 34246
rect 6289 34244 6295 34246
rect 5987 34235 6295 34244
rect 5987 33212 6295 33221
rect 5987 33210 5993 33212
rect 6049 33210 6073 33212
rect 6129 33210 6153 33212
rect 6209 33210 6233 33212
rect 6289 33210 6295 33212
rect 6049 33158 6051 33210
rect 6231 33158 6233 33210
rect 5987 33156 5993 33158
rect 6049 33156 6073 33158
rect 6129 33156 6153 33158
rect 6209 33156 6233 33158
rect 6289 33156 6295 33158
rect 5987 33147 6295 33156
rect 5987 32124 6295 32133
rect 5987 32122 5993 32124
rect 6049 32122 6073 32124
rect 6129 32122 6153 32124
rect 6209 32122 6233 32124
rect 6289 32122 6295 32124
rect 6049 32070 6051 32122
rect 6231 32070 6233 32122
rect 5987 32068 5993 32070
rect 6049 32068 6073 32070
rect 6129 32068 6153 32070
rect 6209 32068 6233 32070
rect 6289 32068 6295 32070
rect 5987 32059 6295 32068
rect 6472 31464 6500 34886
rect 6840 31498 6868 38626
rect 7484 36258 7512 39306
rect 7666 39196 7974 39205
rect 7666 39194 7672 39196
rect 7728 39194 7752 39196
rect 7808 39194 7832 39196
rect 7888 39194 7912 39196
rect 7968 39194 7974 39196
rect 7728 39142 7730 39194
rect 7910 39142 7912 39194
rect 7666 39140 7672 39142
rect 7728 39140 7752 39142
rect 7808 39140 7832 39142
rect 7888 39140 7912 39142
rect 7968 39140 7974 39142
rect 7666 39131 7974 39140
rect 11024 39196 11332 39205
rect 11024 39194 11030 39196
rect 11086 39194 11110 39196
rect 11166 39194 11190 39196
rect 11246 39194 11270 39196
rect 11326 39194 11332 39196
rect 11086 39142 11088 39194
rect 11268 39142 11270 39194
rect 11024 39140 11030 39142
rect 11086 39140 11110 39142
rect 11166 39140 11190 39142
rect 11246 39140 11270 39142
rect 11326 39140 11332 39142
rect 11024 39131 11332 39140
rect 12912 39098 12940 39374
rect 13280 39098 13308 39782
rect 13832 39642 13860 39986
rect 13820 39636 13872 39642
rect 13820 39578 13872 39584
rect 12900 39092 12952 39098
rect 12900 39034 12952 39040
rect 13268 39092 13320 39098
rect 13268 39034 13320 39040
rect 13636 38956 13688 38962
rect 13636 38898 13688 38904
rect 12256 38888 12308 38894
rect 12256 38830 12308 38836
rect 9345 38652 9653 38661
rect 9345 38650 9351 38652
rect 9407 38650 9431 38652
rect 9487 38650 9511 38652
rect 9567 38650 9591 38652
rect 9647 38650 9653 38652
rect 9407 38598 9409 38650
rect 9589 38598 9591 38650
rect 9345 38596 9351 38598
rect 9407 38596 9431 38598
rect 9487 38596 9511 38598
rect 9567 38596 9591 38598
rect 9647 38596 9653 38598
rect 9345 38587 9653 38596
rect 12164 38480 12216 38486
rect 12164 38422 12216 38428
rect 11796 38344 11848 38350
rect 11796 38286 11848 38292
rect 7666 38108 7974 38117
rect 7666 38106 7672 38108
rect 7728 38106 7752 38108
rect 7808 38106 7832 38108
rect 7888 38106 7912 38108
rect 7968 38106 7974 38108
rect 7728 38054 7730 38106
rect 7910 38054 7912 38106
rect 7666 38052 7672 38054
rect 7728 38052 7752 38054
rect 7808 38052 7832 38054
rect 7888 38052 7912 38054
rect 7968 38052 7974 38054
rect 7666 38043 7974 38052
rect 11024 38108 11332 38117
rect 11024 38106 11030 38108
rect 11086 38106 11110 38108
rect 11166 38106 11190 38108
rect 11246 38106 11270 38108
rect 11326 38106 11332 38108
rect 11086 38054 11088 38106
rect 11268 38054 11270 38106
rect 11024 38052 11030 38054
rect 11086 38052 11110 38054
rect 11166 38052 11190 38054
rect 11246 38052 11270 38054
rect 11326 38052 11332 38054
rect 11024 38043 11332 38052
rect 10324 37868 10376 37874
rect 10324 37810 10376 37816
rect 9345 37564 9653 37573
rect 9345 37562 9351 37564
rect 9407 37562 9431 37564
rect 9487 37562 9511 37564
rect 9567 37562 9591 37564
rect 9647 37562 9653 37564
rect 9407 37510 9409 37562
rect 9589 37510 9591 37562
rect 9345 37508 9351 37510
rect 9407 37508 9431 37510
rect 9487 37508 9511 37510
rect 9567 37508 9591 37510
rect 9647 37508 9653 37510
rect 9345 37499 9653 37508
rect 10336 37466 10364 37810
rect 10416 37800 10468 37806
rect 10416 37742 10468 37748
rect 10324 37460 10376 37466
rect 10324 37402 10376 37408
rect 10428 37369 10456 37742
rect 10508 37460 10560 37466
rect 10508 37402 10560 37408
rect 10414 37360 10470 37369
rect 10414 37295 10470 37304
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 7666 37020 7974 37029
rect 7666 37018 7672 37020
rect 7728 37018 7752 37020
rect 7808 37018 7832 37020
rect 7888 37018 7912 37020
rect 7968 37018 7974 37020
rect 7728 36966 7730 37018
rect 7910 36966 7912 37018
rect 7666 36964 7672 36966
rect 7728 36964 7752 36966
rect 7808 36964 7832 36966
rect 7888 36964 7912 36966
rect 7968 36964 7974 36966
rect 7666 36955 7974 36964
rect 8312 36922 8340 37198
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 7300 36230 7512 36258
rect 6920 32836 6972 32842
rect 6920 32778 6972 32784
rect 6748 31470 6868 31498
rect 6472 31436 6684 31464
rect 6552 31340 6604 31346
rect 6552 31282 6604 31288
rect 5987 31036 6295 31045
rect 5987 31034 5993 31036
rect 6049 31034 6073 31036
rect 6129 31034 6153 31036
rect 6209 31034 6233 31036
rect 6289 31034 6295 31036
rect 6049 30982 6051 31034
rect 6231 30982 6233 31034
rect 5987 30980 5993 30982
rect 6049 30980 6073 30982
rect 6129 30980 6153 30982
rect 6209 30980 6233 30982
rect 6289 30980 6295 30982
rect 5987 30971 6295 30980
rect 5987 29948 6295 29957
rect 5987 29946 5993 29948
rect 6049 29946 6073 29948
rect 6129 29946 6153 29948
rect 6209 29946 6233 29948
rect 6289 29946 6295 29948
rect 6049 29894 6051 29946
rect 6231 29894 6233 29946
rect 5987 29892 5993 29894
rect 6049 29892 6073 29894
rect 6129 29892 6153 29894
rect 6209 29892 6233 29894
rect 6289 29892 6295 29894
rect 5987 29883 6295 29892
rect 5987 28860 6295 28869
rect 5987 28858 5993 28860
rect 6049 28858 6073 28860
rect 6129 28858 6153 28860
rect 6209 28858 6233 28860
rect 6289 28858 6295 28860
rect 6049 28806 6051 28858
rect 6231 28806 6233 28858
rect 5987 28804 5993 28806
rect 6049 28804 6073 28806
rect 6129 28804 6153 28806
rect 6209 28804 6233 28806
rect 6289 28804 6295 28806
rect 5987 28795 6295 28804
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 5987 27772 6295 27781
rect 5987 27770 5993 27772
rect 6049 27770 6073 27772
rect 6129 27770 6153 27772
rect 6209 27770 6233 27772
rect 6289 27770 6295 27772
rect 6049 27718 6051 27770
rect 6231 27718 6233 27770
rect 5987 27716 5993 27718
rect 6049 27716 6073 27718
rect 6129 27716 6153 27718
rect 6209 27716 6233 27718
rect 6289 27716 6295 27718
rect 5987 27707 6295 27716
rect 6472 27470 6500 28494
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6472 27062 6500 27406
rect 6460 27056 6512 27062
rect 6460 26998 6512 27004
rect 5908 26988 5960 26994
rect 5908 26930 5960 26936
rect 5816 26784 5868 26790
rect 5816 26726 5868 26732
rect 5724 26308 5776 26314
rect 5724 26250 5776 26256
rect 5736 25294 5764 26250
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5724 24676 5776 24682
rect 5724 24618 5776 24624
rect 5736 24290 5764 24618
rect 5828 24410 5856 26726
rect 5920 26382 5948 26930
rect 5987 26684 6295 26693
rect 5987 26682 5993 26684
rect 6049 26682 6073 26684
rect 6129 26682 6153 26684
rect 6209 26682 6233 26684
rect 6289 26682 6295 26684
rect 6049 26630 6051 26682
rect 6231 26630 6233 26682
rect 5987 26628 5993 26630
rect 6049 26628 6073 26630
rect 6129 26628 6153 26630
rect 6209 26628 6233 26630
rect 6289 26628 6295 26630
rect 5987 26619 6295 26628
rect 5908 26376 5960 26382
rect 5908 26318 5960 26324
rect 5816 24404 5868 24410
rect 5816 24346 5868 24352
rect 5736 24262 5856 24290
rect 5828 22438 5856 24262
rect 5920 24206 5948 26318
rect 6276 26308 6328 26314
rect 6328 26268 6408 26296
rect 6276 26250 6328 26256
rect 5987 25596 6295 25605
rect 5987 25594 5993 25596
rect 6049 25594 6073 25596
rect 6129 25594 6153 25596
rect 6209 25594 6233 25596
rect 6289 25594 6295 25596
rect 6049 25542 6051 25594
rect 6231 25542 6233 25594
rect 5987 25540 5993 25542
rect 6049 25540 6073 25542
rect 6129 25540 6153 25542
rect 6209 25540 6233 25542
rect 6289 25540 6295 25542
rect 5987 25531 6295 25540
rect 5987 24508 6295 24517
rect 5987 24506 5993 24508
rect 6049 24506 6073 24508
rect 6129 24506 6153 24508
rect 6209 24506 6233 24508
rect 6289 24506 6295 24508
rect 6049 24454 6051 24506
rect 6231 24454 6233 24506
rect 5987 24452 5993 24454
rect 6049 24452 6073 24454
rect 6129 24452 6153 24454
rect 6209 24452 6233 24454
rect 6289 24452 6295 24454
rect 5987 24443 6295 24452
rect 6276 24404 6328 24410
rect 6276 24346 6328 24352
rect 6000 24268 6052 24274
rect 6000 24210 6052 24216
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 6012 24070 6040 24210
rect 6184 24200 6236 24206
rect 6184 24142 6236 24148
rect 5908 24064 5960 24070
rect 5908 24006 5960 24012
rect 6000 24064 6052 24070
rect 6000 24006 6052 24012
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 5828 22030 5856 22374
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5920 21434 5948 24006
rect 6196 23526 6224 24142
rect 6288 23882 6316 24346
rect 6380 24070 6408 26268
rect 6472 25702 6500 26998
rect 6564 26926 6592 31282
rect 6552 26920 6604 26926
rect 6552 26862 6604 26868
rect 6564 26382 6592 26862
rect 6552 26376 6604 26382
rect 6552 26318 6604 26324
rect 6552 26240 6604 26246
rect 6552 26182 6604 26188
rect 6460 25696 6512 25702
rect 6460 25638 6512 25644
rect 6472 25362 6500 25638
rect 6460 25356 6512 25362
rect 6460 25298 6512 25304
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6288 23854 6408 23882
rect 6184 23520 6236 23526
rect 6184 23462 6236 23468
rect 5987 23420 6295 23429
rect 5987 23418 5993 23420
rect 6049 23418 6073 23420
rect 6129 23418 6153 23420
rect 6209 23418 6233 23420
rect 6289 23418 6295 23420
rect 6049 23366 6051 23418
rect 6231 23366 6233 23418
rect 5987 23364 5993 23366
rect 6049 23364 6073 23366
rect 6129 23364 6153 23366
rect 6209 23364 6233 23366
rect 6289 23364 6295 23366
rect 5987 23355 6295 23364
rect 5987 22332 6295 22341
rect 5987 22330 5993 22332
rect 6049 22330 6073 22332
rect 6129 22330 6153 22332
rect 6209 22330 6233 22332
rect 6289 22330 6295 22332
rect 6049 22278 6051 22330
rect 6231 22278 6233 22330
rect 5987 22276 5993 22278
rect 6049 22276 6073 22278
rect 6129 22276 6153 22278
rect 6209 22276 6233 22278
rect 6289 22276 6295 22278
rect 5987 22267 6295 22276
rect 6380 21978 6408 23854
rect 6380 21950 6500 21978
rect 6368 21888 6420 21894
rect 6368 21830 6420 21836
rect 5828 21406 5948 21434
rect 5724 20868 5776 20874
rect 5724 20810 5776 20816
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5540 15904 5592 15910
rect 5540 15846 5592 15852
rect 5448 13796 5500 13802
rect 5448 13738 5500 13744
rect 5356 12640 5408 12646
rect 5356 12582 5408 12588
rect 5552 11762 5580 15846
rect 5632 15428 5684 15434
rect 5632 15370 5684 15376
rect 5644 12238 5672 15370
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5632 12096 5684 12102
rect 5632 12038 5684 12044
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5644 10674 5672 12038
rect 5736 11218 5764 20810
rect 5828 18970 5856 21406
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5920 21010 5948 21286
rect 5987 21244 6295 21253
rect 5987 21242 5993 21244
rect 6049 21242 6073 21244
rect 6129 21242 6153 21244
rect 6209 21242 6233 21244
rect 6289 21242 6295 21244
rect 6049 21190 6051 21242
rect 6231 21190 6233 21242
rect 5987 21188 5993 21190
rect 6049 21188 6073 21190
rect 6129 21188 6153 21190
rect 6209 21188 6233 21190
rect 6289 21188 6295 21190
rect 5987 21179 6295 21188
rect 5908 21004 5960 21010
rect 5908 20946 5960 20952
rect 6380 20942 6408 21830
rect 6472 20942 6500 21950
rect 6368 20936 6420 20942
rect 6368 20878 6420 20884
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 5908 20800 5960 20806
rect 5908 20742 5960 20748
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5828 11898 5856 18906
rect 5920 18850 5948 20742
rect 5987 20156 6295 20165
rect 5987 20154 5993 20156
rect 6049 20154 6073 20156
rect 6129 20154 6153 20156
rect 6209 20154 6233 20156
rect 6289 20154 6295 20156
rect 6049 20102 6051 20154
rect 6231 20102 6233 20154
rect 5987 20100 5993 20102
rect 6049 20100 6073 20102
rect 6129 20100 6153 20102
rect 6209 20100 6233 20102
rect 6289 20100 6295 20102
rect 5987 20091 6295 20100
rect 6368 19372 6420 19378
rect 6368 19314 6420 19320
rect 5987 19068 6295 19077
rect 5987 19066 5993 19068
rect 6049 19066 6073 19068
rect 6129 19066 6153 19068
rect 6209 19066 6233 19068
rect 6289 19066 6295 19068
rect 6049 19014 6051 19066
rect 6231 19014 6233 19066
rect 5987 19012 5993 19014
rect 6049 19012 6073 19014
rect 6129 19012 6153 19014
rect 6209 19012 6233 19014
rect 6289 19012 6295 19014
rect 5987 19003 6295 19012
rect 5920 18822 6040 18850
rect 5908 18760 5960 18766
rect 5908 18702 5960 18708
rect 5920 18426 5948 18702
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 6012 18136 6040 18822
rect 6380 18714 6408 19314
rect 6472 18970 6500 20878
rect 6460 18964 6512 18970
rect 6460 18906 6512 18912
rect 6380 18686 6500 18714
rect 6092 18624 6144 18630
rect 6092 18566 6144 18572
rect 6184 18624 6236 18630
rect 6184 18566 6236 18572
rect 6368 18624 6420 18630
rect 6368 18566 6420 18572
rect 5920 18108 6040 18136
rect 5920 15162 5948 18108
rect 6104 18086 6132 18566
rect 6196 18358 6224 18566
rect 6184 18352 6236 18358
rect 6184 18294 6236 18300
rect 6380 18290 6408 18566
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6092 18080 6144 18086
rect 6092 18022 6144 18028
rect 5987 17980 6295 17989
rect 5987 17978 5993 17980
rect 6049 17978 6073 17980
rect 6129 17978 6153 17980
rect 6209 17978 6233 17980
rect 6289 17978 6295 17980
rect 6049 17926 6051 17978
rect 6231 17926 6233 17978
rect 5987 17924 5993 17926
rect 6049 17924 6073 17926
rect 6129 17924 6153 17926
rect 6209 17924 6233 17926
rect 6289 17924 6295 17926
rect 5987 17915 6295 17924
rect 6380 17882 6408 18226
rect 6368 17876 6420 17882
rect 6368 17818 6420 17824
rect 6472 17678 6500 18686
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 5987 16892 6295 16901
rect 5987 16890 5993 16892
rect 6049 16890 6073 16892
rect 6129 16890 6153 16892
rect 6209 16890 6233 16892
rect 6289 16890 6295 16892
rect 6049 16838 6051 16890
rect 6231 16838 6233 16890
rect 5987 16836 5993 16838
rect 6049 16836 6073 16838
rect 6129 16836 6153 16838
rect 6209 16836 6233 16838
rect 6289 16836 6295 16838
rect 5987 16827 6295 16836
rect 6472 16658 6500 17614
rect 6460 16652 6512 16658
rect 6460 16594 6512 16600
rect 6472 16114 6500 16594
rect 6460 16108 6512 16114
rect 6460 16050 6512 16056
rect 5987 15804 6295 15813
rect 5987 15802 5993 15804
rect 6049 15802 6073 15804
rect 6129 15802 6153 15804
rect 6209 15802 6233 15804
rect 6289 15802 6295 15804
rect 6049 15750 6051 15802
rect 6231 15750 6233 15802
rect 5987 15748 5993 15750
rect 6049 15748 6073 15750
rect 6129 15748 6153 15750
rect 6209 15748 6233 15750
rect 6289 15748 6295 15750
rect 5987 15739 6295 15748
rect 6472 15570 6500 16050
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 5908 14816 5960 14822
rect 5908 14758 5960 14764
rect 5920 14618 5948 14758
rect 5987 14716 6295 14725
rect 5987 14714 5993 14716
rect 6049 14714 6073 14716
rect 6129 14714 6153 14716
rect 6209 14714 6233 14716
rect 6289 14714 6295 14716
rect 6049 14662 6051 14714
rect 6231 14662 6233 14714
rect 5987 14660 5993 14662
rect 6049 14660 6073 14662
rect 6129 14660 6153 14662
rect 6209 14660 6233 14662
rect 6289 14660 6295 14662
rect 5987 14651 6295 14660
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6012 13716 6040 14350
rect 5920 13688 6040 13716
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5920 11830 5948 13688
rect 5987 13628 6295 13637
rect 5987 13626 5993 13628
rect 6049 13626 6073 13628
rect 6129 13626 6153 13628
rect 6209 13626 6233 13628
rect 6289 13626 6295 13628
rect 6049 13574 6051 13626
rect 6231 13574 6233 13626
rect 5987 13572 5993 13574
rect 6049 13572 6073 13574
rect 6129 13572 6153 13574
rect 6209 13572 6233 13574
rect 6289 13572 6295 13574
rect 5987 13563 6295 13572
rect 6380 13530 6408 14894
rect 6368 13524 6420 13530
rect 6368 13466 6420 13472
rect 6564 13258 6592 26182
rect 6656 19378 6684 31436
rect 6748 24886 6776 31470
rect 6828 29504 6880 29510
rect 6828 29446 6880 29452
rect 6840 29306 6868 29446
rect 6828 29300 6880 29306
rect 6828 29242 6880 29248
rect 6932 29073 6960 32778
rect 7196 31816 7248 31822
rect 7196 31758 7248 31764
rect 7012 31476 7064 31482
rect 7012 31418 7064 31424
rect 6918 29064 6974 29073
rect 6918 28999 6974 29008
rect 6932 28558 6960 28999
rect 6920 28552 6972 28558
rect 6826 28520 6882 28529
rect 6920 28494 6972 28500
rect 6826 28455 6882 28464
rect 6840 27674 6868 28455
rect 6828 27668 6880 27674
rect 6828 27610 6880 27616
rect 6828 26240 6880 26246
rect 6828 26182 6880 26188
rect 6736 24880 6788 24886
rect 6736 24822 6788 24828
rect 6840 24206 6868 26182
rect 6920 25968 6972 25974
rect 6920 25910 6972 25916
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6736 24064 6788 24070
rect 6736 24006 6788 24012
rect 6748 21468 6776 24006
rect 6840 21622 6868 24142
rect 6828 21616 6880 21622
rect 6828 21558 6880 21564
rect 6748 21440 6868 21468
rect 6736 20868 6788 20874
rect 6736 20810 6788 20816
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6552 13252 6604 13258
rect 6552 13194 6604 13200
rect 5987 12540 6295 12549
rect 5987 12538 5993 12540
rect 6049 12538 6073 12540
rect 6129 12538 6153 12540
rect 6209 12538 6233 12540
rect 6289 12538 6295 12540
rect 6049 12486 6051 12538
rect 6231 12486 6233 12538
rect 5987 12484 5993 12486
rect 6049 12484 6073 12486
rect 6129 12484 6153 12486
rect 6209 12484 6233 12486
rect 6289 12484 6295 12486
rect 5987 12475 6295 12484
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5920 11642 5948 11766
rect 6656 11642 6684 19314
rect 6748 18986 6776 20810
rect 6840 20244 6868 21440
rect 6932 20777 6960 25910
rect 7024 24970 7052 31418
rect 7104 29844 7156 29850
rect 7104 29786 7156 29792
rect 7116 29170 7144 29786
rect 7104 29164 7156 29170
rect 7104 29106 7156 29112
rect 7116 28626 7144 29106
rect 7104 28620 7156 28626
rect 7104 28562 7156 28568
rect 7208 28529 7236 31758
rect 7300 29850 7328 36230
rect 7380 36168 7432 36174
rect 7380 36110 7432 36116
rect 7392 32366 7420 36110
rect 7666 35932 7974 35941
rect 7666 35930 7672 35932
rect 7728 35930 7752 35932
rect 7808 35930 7832 35932
rect 7888 35930 7912 35932
rect 7968 35930 7974 35932
rect 7728 35878 7730 35930
rect 7910 35878 7912 35930
rect 7666 35876 7672 35878
rect 7728 35876 7752 35878
rect 7808 35876 7832 35878
rect 7888 35876 7912 35878
rect 7968 35876 7974 35878
rect 7666 35867 7974 35876
rect 8116 35080 8168 35086
rect 8116 35022 8168 35028
rect 7666 34844 7974 34853
rect 7666 34842 7672 34844
rect 7728 34842 7752 34844
rect 7808 34842 7832 34844
rect 7888 34842 7912 34844
rect 7968 34842 7974 34844
rect 7728 34790 7730 34842
rect 7910 34790 7912 34842
rect 7666 34788 7672 34790
rect 7728 34788 7752 34790
rect 7808 34788 7832 34790
rect 7888 34788 7912 34790
rect 7968 34788 7974 34790
rect 7666 34779 7974 34788
rect 7666 33756 7974 33765
rect 7666 33754 7672 33756
rect 7728 33754 7752 33756
rect 7808 33754 7832 33756
rect 7888 33754 7912 33756
rect 7968 33754 7974 33756
rect 7728 33702 7730 33754
rect 7910 33702 7912 33754
rect 7666 33700 7672 33702
rect 7728 33700 7752 33702
rect 7808 33700 7832 33702
rect 7888 33700 7912 33702
rect 7968 33700 7974 33702
rect 7666 33691 7974 33700
rect 7666 32668 7974 32677
rect 7666 32666 7672 32668
rect 7728 32666 7752 32668
rect 7808 32666 7832 32668
rect 7888 32666 7912 32668
rect 7968 32666 7974 32668
rect 7728 32614 7730 32666
rect 7910 32614 7912 32666
rect 7666 32612 7672 32614
rect 7728 32612 7752 32614
rect 7808 32612 7832 32614
rect 7888 32612 7912 32614
rect 7968 32612 7974 32614
rect 7666 32603 7974 32612
rect 7380 32360 7432 32366
rect 7380 32302 7432 32308
rect 7392 31890 7420 32302
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7392 30938 7420 31826
rect 7666 31580 7974 31589
rect 7666 31578 7672 31580
rect 7728 31578 7752 31580
rect 7808 31578 7832 31580
rect 7888 31578 7912 31580
rect 7968 31578 7974 31580
rect 7728 31526 7730 31578
rect 7910 31526 7912 31578
rect 7666 31524 7672 31526
rect 7728 31524 7752 31526
rect 7808 31524 7832 31526
rect 7888 31524 7912 31526
rect 7968 31524 7974 31526
rect 7666 31515 7974 31524
rect 8024 31272 8076 31278
rect 8024 31214 8076 31220
rect 7380 30932 7432 30938
rect 7432 30892 7512 30920
rect 7380 30874 7432 30880
rect 7380 30592 7432 30598
rect 7380 30534 7432 30540
rect 7288 29844 7340 29850
rect 7288 29786 7340 29792
rect 7288 29640 7340 29646
rect 7288 29582 7340 29588
rect 7194 28520 7250 28529
rect 7194 28455 7250 28464
rect 7104 28416 7156 28422
rect 7104 28358 7156 28364
rect 7116 28218 7144 28358
rect 7104 28212 7156 28218
rect 7104 28154 7156 28160
rect 7300 28098 7328 29582
rect 7116 28070 7328 28098
rect 7116 25106 7144 28070
rect 7288 28008 7340 28014
rect 7288 27950 7340 27956
rect 7196 27328 7248 27334
rect 7196 27270 7248 27276
rect 7208 26194 7236 27270
rect 7300 26382 7328 27950
rect 7392 27538 7420 30534
rect 7484 29646 7512 30892
rect 7666 30492 7974 30501
rect 7666 30490 7672 30492
rect 7728 30490 7752 30492
rect 7808 30490 7832 30492
rect 7888 30490 7912 30492
rect 7968 30490 7974 30492
rect 7728 30438 7730 30490
rect 7910 30438 7912 30490
rect 7666 30436 7672 30438
rect 7728 30436 7752 30438
rect 7808 30436 7832 30438
rect 7888 30436 7912 30438
rect 7968 30436 7974 30438
rect 7666 30427 7974 30436
rect 7472 29640 7524 29646
rect 7472 29582 7524 29588
rect 7472 29504 7524 29510
rect 7472 29446 7524 29452
rect 7484 27860 7512 29446
rect 7666 29404 7974 29413
rect 7666 29402 7672 29404
rect 7728 29402 7752 29404
rect 7808 29402 7832 29404
rect 7888 29402 7912 29404
rect 7968 29402 7974 29404
rect 7728 29350 7730 29402
rect 7910 29350 7912 29402
rect 7666 29348 7672 29350
rect 7728 29348 7752 29350
rect 7808 29348 7832 29350
rect 7888 29348 7912 29350
rect 7968 29348 7974 29350
rect 7666 29339 7974 29348
rect 7564 28416 7616 28422
rect 7564 28358 7616 28364
rect 7576 28014 7604 28358
rect 7666 28316 7974 28325
rect 7666 28314 7672 28316
rect 7728 28314 7752 28316
rect 7808 28314 7832 28316
rect 7888 28314 7912 28316
rect 7968 28314 7974 28316
rect 7728 28262 7730 28314
rect 7910 28262 7912 28314
rect 7666 28260 7672 28262
rect 7728 28260 7752 28262
rect 7808 28260 7832 28262
rect 7888 28260 7912 28262
rect 7968 28260 7974 28262
rect 7666 28251 7974 28260
rect 7564 28008 7616 28014
rect 7564 27950 7616 27956
rect 7932 28008 7984 28014
rect 7932 27950 7984 27956
rect 7484 27832 7604 27860
rect 7944 27849 7972 27950
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7380 27532 7432 27538
rect 7380 27474 7432 27480
rect 7392 27130 7420 27474
rect 7380 27124 7432 27130
rect 7380 27066 7432 27072
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7484 26874 7512 27542
rect 7576 26994 7604 27832
rect 7930 27840 7986 27849
rect 7930 27775 7986 27784
rect 7666 27228 7974 27237
rect 7666 27226 7672 27228
rect 7728 27226 7752 27228
rect 7808 27226 7832 27228
rect 7888 27226 7912 27228
rect 7968 27226 7974 27228
rect 7728 27174 7730 27226
rect 7910 27174 7912 27226
rect 7666 27172 7672 27174
rect 7728 27172 7752 27174
rect 7808 27172 7832 27174
rect 7888 27172 7912 27174
rect 7968 27172 7974 27174
rect 7666 27163 7974 27172
rect 7564 26988 7616 26994
rect 7564 26930 7616 26936
rect 7748 26920 7800 26926
rect 7484 26868 7748 26874
rect 7484 26862 7800 26868
rect 7392 26450 7420 26862
rect 7484 26846 7788 26862
rect 7380 26444 7432 26450
rect 7380 26386 7432 26392
rect 7288 26376 7340 26382
rect 7286 26344 7288 26353
rect 7340 26344 7342 26353
rect 7286 26279 7342 26288
rect 7392 26246 7420 26386
rect 7564 26376 7616 26382
rect 7564 26318 7616 26324
rect 7380 26240 7432 26246
rect 7208 26166 7328 26194
rect 7380 26182 7432 26188
rect 7116 25078 7236 25106
rect 7024 24942 7144 24970
rect 7012 24880 7064 24886
rect 7012 24822 7064 24828
rect 7024 22030 7052 24822
rect 7116 22658 7144 24942
rect 7208 23186 7236 25078
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 7208 22778 7236 23122
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7116 22642 7236 22658
rect 7116 22636 7248 22642
rect 7116 22630 7196 22636
rect 7196 22578 7248 22584
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 7116 21876 7144 21966
rect 7024 21848 7144 21876
rect 6918 20768 6974 20777
rect 6918 20703 6974 20712
rect 6918 20496 6974 20505
rect 6918 20431 6974 20440
rect 6932 20398 6960 20431
rect 7024 20398 7052 21848
rect 7104 20528 7156 20534
rect 7104 20470 7156 20476
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 6840 20216 6960 20244
rect 6828 19712 6880 19718
rect 6828 19654 6880 19660
rect 6840 19514 6868 19654
rect 6828 19508 6880 19514
rect 6828 19450 6880 19456
rect 6932 19360 6960 20216
rect 7024 19961 7052 20334
rect 7010 19952 7066 19961
rect 7010 19887 7066 19896
rect 7012 19372 7064 19378
rect 6932 19332 7012 19360
rect 7012 19314 7064 19320
rect 7010 19272 7066 19281
rect 7010 19207 7066 19216
rect 6828 19168 6880 19174
rect 6826 19136 6828 19145
rect 6880 19136 6882 19145
rect 6826 19071 6882 19080
rect 6748 18958 6868 18986
rect 6736 18828 6788 18834
rect 6736 18770 6788 18776
rect 6748 18426 6776 18770
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6736 15156 6788 15162
rect 6736 15098 6788 15104
rect 6748 14414 6776 15098
rect 6840 14822 6868 18958
rect 7024 18766 7052 19207
rect 6920 18760 6972 18766
rect 6920 18702 6972 18708
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6932 18426 6960 18702
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 7024 18426 7052 18566
rect 6920 18420 6972 18426
rect 6920 18362 6972 18368
rect 7012 18420 7064 18426
rect 7012 18362 7064 18368
rect 6918 17640 6974 17649
rect 6918 17575 6920 17584
rect 6972 17575 6974 17584
rect 6920 17546 6972 17552
rect 6932 15706 6960 17546
rect 7116 17354 7144 20470
rect 7208 19258 7236 22578
rect 7300 21146 7328 26166
rect 7576 25498 7604 26318
rect 7666 26140 7974 26149
rect 7666 26138 7672 26140
rect 7728 26138 7752 26140
rect 7808 26138 7832 26140
rect 7888 26138 7912 26140
rect 7968 26138 7974 26140
rect 7728 26086 7730 26138
rect 7910 26086 7912 26138
rect 7666 26084 7672 26086
rect 7728 26084 7752 26086
rect 7808 26084 7832 26086
rect 7888 26084 7912 26086
rect 7968 26084 7974 26086
rect 7666 26075 7974 26084
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7944 25498 7972 25638
rect 7564 25492 7616 25498
rect 7564 25434 7616 25440
rect 7932 25492 7984 25498
rect 7932 25434 7984 25440
rect 7564 25356 7616 25362
rect 7564 25298 7616 25304
rect 7472 24676 7524 24682
rect 7472 24618 7524 24624
rect 7380 24608 7432 24614
rect 7380 24550 7432 24556
rect 7392 24410 7420 24550
rect 7484 24410 7512 24618
rect 7576 24614 7604 25298
rect 7666 25052 7974 25061
rect 7666 25050 7672 25052
rect 7728 25050 7752 25052
rect 7808 25050 7832 25052
rect 7888 25050 7912 25052
rect 7968 25050 7974 25052
rect 7728 24998 7730 25050
rect 7910 24998 7912 25050
rect 7666 24996 7672 24998
rect 7728 24996 7752 24998
rect 7808 24996 7832 24998
rect 7888 24996 7912 24998
rect 7968 24996 7974 24998
rect 7666 24987 7974 24996
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7564 24608 7616 24614
rect 7564 24550 7616 24556
rect 7380 24404 7432 24410
rect 7380 24346 7432 24352
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7668 24290 7696 24890
rect 7748 24608 7800 24614
rect 7748 24550 7800 24556
rect 7392 24262 7696 24290
rect 7392 22030 7420 24262
rect 7760 24154 7788 24550
rect 7576 24126 7788 24154
rect 7472 24064 7524 24070
rect 7472 24006 7524 24012
rect 7484 23866 7512 24006
rect 7472 23860 7524 23866
rect 7472 23802 7524 23808
rect 7576 23730 7604 24126
rect 7666 23964 7974 23973
rect 7666 23962 7672 23964
rect 7728 23962 7752 23964
rect 7808 23962 7832 23964
rect 7888 23962 7912 23964
rect 7968 23962 7974 23964
rect 7728 23910 7730 23962
rect 7910 23910 7912 23962
rect 7666 23908 7672 23910
rect 7728 23908 7752 23910
rect 7808 23908 7832 23910
rect 7888 23908 7912 23910
rect 7968 23908 7974 23910
rect 7666 23899 7974 23908
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7576 23633 7604 23666
rect 7562 23624 7618 23633
rect 7562 23559 7618 23568
rect 7840 23588 7892 23594
rect 7840 23530 7892 23536
rect 7472 23044 7524 23050
rect 7472 22986 7524 22992
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 7378 21856 7434 21865
rect 7378 21791 7434 21800
rect 7392 21350 7420 21791
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7288 21140 7340 21146
rect 7288 21082 7340 21088
rect 7392 21026 7420 21286
rect 7300 20998 7420 21026
rect 7300 20074 7328 20998
rect 7300 20046 7420 20074
rect 7288 19984 7340 19990
rect 7288 19926 7340 19932
rect 7300 19378 7328 19926
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7208 19230 7328 19258
rect 7300 18714 7328 19230
rect 7024 17326 7144 17354
rect 7208 18686 7328 18714
rect 7024 16114 7052 17326
rect 7208 17202 7236 18686
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 7300 18222 7328 18566
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7196 17196 7248 17202
rect 7248 17156 7328 17184
rect 7196 17138 7248 17144
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 6920 15700 6972 15706
rect 6920 15642 6972 15648
rect 6828 14816 6880 14822
rect 6828 14758 6880 14764
rect 6840 14482 6868 14758
rect 6828 14476 6880 14482
rect 6828 14418 6880 14424
rect 6736 14408 6788 14414
rect 6736 14350 6788 14356
rect 6748 14278 6776 14350
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 6828 13252 6880 13258
rect 6828 13194 6880 13200
rect 6840 12434 6868 13194
rect 6920 12980 6972 12986
rect 6920 12922 6972 12928
rect 5828 11614 5948 11642
rect 6380 11614 6684 11642
rect 6748 12406 6868 12434
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5828 11082 5856 11614
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11200 5948 11494
rect 5987 11452 6295 11461
rect 5987 11450 5993 11452
rect 6049 11450 6073 11452
rect 6129 11450 6153 11452
rect 6209 11450 6233 11452
rect 6289 11450 6295 11452
rect 6049 11398 6051 11450
rect 6231 11398 6233 11450
rect 5987 11396 5993 11398
rect 6049 11396 6073 11398
rect 6129 11396 6153 11398
rect 6209 11396 6233 11398
rect 6289 11396 6295 11398
rect 5987 11387 6295 11396
rect 6092 11212 6144 11218
rect 5920 11172 6092 11200
rect 6092 11154 6144 11160
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 6380 10996 6408 11614
rect 6748 11506 6776 12406
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6840 11642 6868 12310
rect 6932 11762 6960 12922
rect 7024 12238 7052 16050
rect 7116 15162 7144 17070
rect 7196 15700 7248 15706
rect 7196 15642 7248 15648
rect 7104 15156 7156 15162
rect 7104 15098 7156 15104
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14618 7144 14962
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7116 12918 7144 13262
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7208 12442 7236 15642
rect 7300 14074 7328 17156
rect 7392 17066 7420 20046
rect 7484 19990 7512 22986
rect 7852 22964 7880 23530
rect 8036 23032 8064 31214
rect 8128 29714 8156 35022
rect 8208 34604 8260 34610
rect 8208 34546 8260 34552
rect 8220 31822 8248 34546
rect 8208 31816 8260 31822
rect 8208 31758 8260 31764
rect 8208 30388 8260 30394
rect 8208 30330 8260 30336
rect 8116 29708 8168 29714
rect 8116 29650 8168 29656
rect 8116 28960 8168 28966
rect 8116 28902 8168 28908
rect 8128 27878 8156 28902
rect 8220 28200 8248 30330
rect 8312 28422 8340 36858
rect 9772 36780 9824 36786
rect 9772 36722 9824 36728
rect 9345 36476 9653 36485
rect 9345 36474 9351 36476
rect 9407 36474 9431 36476
rect 9487 36474 9511 36476
rect 9567 36474 9591 36476
rect 9647 36474 9653 36476
rect 9407 36422 9409 36474
rect 9589 36422 9591 36474
rect 9345 36420 9351 36422
rect 9407 36420 9431 36422
rect 9487 36420 9511 36422
rect 9567 36420 9591 36422
rect 9647 36420 9653 36422
rect 9345 36411 9653 36420
rect 8944 35692 8996 35698
rect 8944 35634 8996 35640
rect 8956 35290 8984 35634
rect 9345 35388 9653 35397
rect 9345 35386 9351 35388
rect 9407 35386 9431 35388
rect 9487 35386 9511 35388
rect 9567 35386 9591 35388
rect 9647 35386 9653 35388
rect 9407 35334 9409 35386
rect 9589 35334 9591 35386
rect 9345 35332 9351 35334
rect 9407 35332 9431 35334
rect 9487 35332 9511 35334
rect 9567 35332 9591 35334
rect 9647 35332 9653 35334
rect 9345 35323 9653 35332
rect 8944 35284 8996 35290
rect 8944 35226 8996 35232
rect 9680 35080 9732 35086
rect 9680 35022 9732 35028
rect 9345 34300 9653 34309
rect 9345 34298 9351 34300
rect 9407 34298 9431 34300
rect 9487 34298 9511 34300
rect 9567 34298 9591 34300
rect 9647 34298 9653 34300
rect 9407 34246 9409 34298
rect 9589 34246 9591 34298
rect 9345 34244 9351 34246
rect 9407 34244 9431 34246
rect 9487 34244 9511 34246
rect 9567 34244 9591 34246
rect 9647 34244 9653 34246
rect 9345 34235 9653 34244
rect 9692 33454 9720 35022
rect 9784 34678 9812 36722
rect 10232 36712 10284 36718
rect 10232 36654 10284 36660
rect 10244 35834 10272 36654
rect 10520 36378 10548 37402
rect 11808 37369 11836 38286
rect 11888 38276 11940 38282
rect 11888 38218 11940 38224
rect 11900 38010 11928 38218
rect 11888 38004 11940 38010
rect 11888 37946 11940 37952
rect 11794 37360 11850 37369
rect 11794 37295 11850 37304
rect 11888 37256 11940 37262
rect 11702 37224 11758 37233
rect 11940 37204 12112 37210
rect 11888 37198 12112 37204
rect 11900 37182 12112 37198
rect 11702 37159 11758 37168
rect 11716 37126 11744 37159
rect 12084 37126 12112 37182
rect 11704 37120 11756 37126
rect 11704 37062 11756 37068
rect 11980 37120 12032 37126
rect 11980 37062 12032 37068
rect 12072 37120 12124 37126
rect 12072 37062 12124 37068
rect 11024 37020 11332 37029
rect 11024 37018 11030 37020
rect 11086 37018 11110 37020
rect 11166 37018 11190 37020
rect 11246 37018 11270 37020
rect 11326 37018 11332 37020
rect 11086 36966 11088 37018
rect 11268 36966 11270 37018
rect 11024 36964 11030 36966
rect 11086 36964 11110 36966
rect 11166 36964 11190 36966
rect 11246 36964 11270 36966
rect 11326 36964 11332 36966
rect 11024 36955 11332 36964
rect 11426 36952 11482 36961
rect 11426 36887 11482 36896
rect 10600 36848 10652 36854
rect 10600 36790 10652 36796
rect 10508 36372 10560 36378
rect 10508 36314 10560 36320
rect 10508 36236 10560 36242
rect 10508 36178 10560 36184
rect 10232 35828 10284 35834
rect 10232 35770 10284 35776
rect 10416 35692 10468 35698
rect 10416 35634 10468 35640
rect 10428 35290 10456 35634
rect 10416 35284 10468 35290
rect 10416 35226 10468 35232
rect 9864 35216 9916 35222
rect 9864 35158 9916 35164
rect 9772 34672 9824 34678
rect 9772 34614 9824 34620
rect 9772 34400 9824 34406
rect 9772 34342 9824 34348
rect 9680 33448 9732 33454
rect 9680 33390 9732 33396
rect 9345 33212 9653 33221
rect 9345 33210 9351 33212
rect 9407 33210 9431 33212
rect 9487 33210 9511 33212
rect 9567 33210 9591 33212
rect 9647 33210 9653 33212
rect 9407 33158 9409 33210
rect 9589 33158 9591 33210
rect 9345 33156 9351 33158
rect 9407 33156 9431 33158
rect 9487 33156 9511 33158
rect 9567 33156 9591 33158
rect 9647 33156 9653 33158
rect 9345 33147 9653 33156
rect 8760 33040 8812 33046
rect 8760 32982 8812 32988
rect 8576 32428 8628 32434
rect 8576 32370 8628 32376
rect 8484 30048 8536 30054
rect 8484 29990 8536 29996
rect 8392 29164 8444 29170
rect 8392 29106 8444 29112
rect 8300 28416 8352 28422
rect 8300 28358 8352 28364
rect 8220 28172 8340 28200
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8116 27872 8168 27878
rect 8116 27814 8168 27820
rect 8220 27674 8248 28018
rect 8208 27668 8260 27674
rect 8208 27610 8260 27616
rect 8208 27464 8260 27470
rect 8208 27406 8260 27412
rect 8220 27130 8248 27406
rect 8208 27124 8260 27130
rect 8208 27066 8260 27072
rect 8208 25764 8260 25770
rect 8208 25706 8260 25712
rect 8220 24954 8248 25706
rect 8208 24948 8260 24954
rect 8208 24890 8260 24896
rect 8312 23746 8340 28172
rect 8404 28121 8432 29106
rect 8390 28112 8446 28121
rect 8390 28047 8446 28056
rect 8496 26790 8524 29990
rect 8484 26784 8536 26790
rect 8484 26726 8536 26732
rect 8220 23718 8340 23746
rect 8220 23118 8248 23718
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8484 23656 8536 23662
rect 8484 23598 8536 23604
rect 8312 23186 8340 23598
rect 8496 23526 8524 23598
rect 8484 23520 8536 23526
rect 8484 23462 8536 23468
rect 8300 23180 8352 23186
rect 8352 23140 8524 23168
rect 8300 23122 8352 23128
rect 8208 23112 8260 23118
rect 8208 23054 8260 23060
rect 8036 23004 8156 23032
rect 7852 22936 8064 22964
rect 7666 22876 7974 22885
rect 7666 22874 7672 22876
rect 7728 22874 7752 22876
rect 7808 22874 7832 22876
rect 7888 22874 7912 22876
rect 7968 22874 7974 22876
rect 7728 22822 7730 22874
rect 7910 22822 7912 22874
rect 7666 22820 7672 22822
rect 7728 22820 7752 22822
rect 7808 22820 7832 22822
rect 7888 22820 7912 22822
rect 7968 22820 7974 22822
rect 7666 22811 7974 22820
rect 8036 22778 8064 22936
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 7564 21956 7616 21962
rect 7564 21898 7616 21904
rect 7472 19984 7524 19990
rect 7472 19926 7524 19932
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7484 19514 7512 19790
rect 7472 19508 7524 19514
rect 7472 19450 7524 19456
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7484 19281 7512 19314
rect 7470 19272 7526 19281
rect 7470 19207 7472 19216
rect 7524 19207 7526 19216
rect 7472 19178 7524 19184
rect 7576 19174 7604 21898
rect 7666 21788 7974 21797
rect 7666 21786 7672 21788
rect 7728 21786 7752 21788
rect 7808 21786 7832 21788
rect 7888 21786 7912 21788
rect 7968 21786 7974 21788
rect 7728 21734 7730 21786
rect 7910 21734 7912 21786
rect 7666 21732 7672 21734
rect 7728 21732 7752 21734
rect 7808 21732 7832 21734
rect 7888 21732 7912 21734
rect 7968 21732 7974 21734
rect 7666 21723 7974 21732
rect 7748 21480 7800 21486
rect 7748 21422 7800 21428
rect 7932 21480 7984 21486
rect 7984 21440 8064 21468
rect 7932 21422 7984 21428
rect 7760 21010 7788 21422
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7666 20700 7974 20709
rect 7666 20698 7672 20700
rect 7728 20698 7752 20700
rect 7808 20698 7832 20700
rect 7888 20698 7912 20700
rect 7968 20698 7974 20700
rect 7728 20646 7730 20698
rect 7910 20646 7912 20698
rect 7666 20644 7672 20646
rect 7728 20644 7752 20646
rect 7808 20644 7832 20646
rect 7888 20644 7912 20646
rect 7968 20644 7974 20646
rect 7666 20635 7974 20644
rect 7930 20496 7986 20505
rect 7930 20431 7932 20440
rect 7984 20431 7986 20440
rect 7932 20402 7984 20408
rect 7666 19612 7974 19621
rect 7666 19610 7672 19612
rect 7728 19610 7752 19612
rect 7808 19610 7832 19612
rect 7888 19610 7912 19612
rect 7968 19610 7974 19612
rect 7728 19558 7730 19610
rect 7910 19558 7912 19610
rect 7666 19556 7672 19558
rect 7728 19556 7752 19558
rect 7808 19556 7832 19558
rect 7888 19556 7912 19558
rect 7968 19556 7974 19558
rect 7666 19547 7974 19556
rect 7656 19304 7708 19310
rect 7656 19246 7708 19252
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7472 18896 7524 18902
rect 7472 18838 7524 18844
rect 7484 18290 7512 18838
rect 7562 18728 7618 18737
rect 7668 18714 7696 19246
rect 7748 19168 7800 19174
rect 7748 19110 7800 19116
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7618 18686 7696 18714
rect 7562 18663 7618 18672
rect 7760 18612 7788 19110
rect 7852 18970 7880 19110
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 7576 18584 7788 18612
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7484 17134 7512 17478
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7380 17060 7432 17066
rect 7380 17002 7432 17008
rect 7576 16640 7604 18584
rect 7666 18524 7974 18533
rect 7666 18522 7672 18524
rect 7728 18522 7752 18524
rect 7808 18522 7832 18524
rect 7888 18522 7912 18524
rect 7968 18522 7974 18524
rect 7728 18470 7730 18522
rect 7910 18470 7912 18522
rect 7666 18468 7672 18470
rect 7728 18468 7752 18470
rect 7808 18468 7832 18470
rect 7888 18468 7912 18470
rect 7968 18468 7974 18470
rect 7666 18459 7974 18468
rect 8036 18136 8064 21440
rect 8128 20942 8156 23004
rect 8392 22976 8444 22982
rect 8392 22918 8444 22924
rect 8404 22778 8432 22918
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8208 21412 8260 21418
rect 8208 21354 8260 21360
rect 8116 20936 8168 20942
rect 8116 20878 8168 20884
rect 8116 20800 8168 20806
rect 8116 20742 8168 20748
rect 7944 18108 8064 18136
rect 7944 17542 7972 18108
rect 8022 18048 8078 18057
rect 8022 17983 8078 17992
rect 7932 17536 7984 17542
rect 7932 17478 7984 17484
rect 7666 17436 7974 17445
rect 7666 17434 7672 17436
rect 7728 17434 7752 17436
rect 7808 17434 7832 17436
rect 7888 17434 7912 17436
rect 7968 17434 7974 17436
rect 7728 17382 7730 17434
rect 7910 17382 7912 17434
rect 7666 17380 7672 17382
rect 7728 17380 7752 17382
rect 7808 17380 7832 17382
rect 7888 17380 7912 17382
rect 7968 17380 7974 17382
rect 7666 17371 7974 17380
rect 7840 17332 7892 17338
rect 7840 17274 7892 17280
rect 7852 17202 7880 17274
rect 8036 17218 8064 17983
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7944 17190 8064 17218
rect 7484 16612 7604 16640
rect 7380 16176 7432 16182
rect 7380 16118 7432 16124
rect 7392 15638 7420 16118
rect 7380 15632 7432 15638
rect 7380 15574 7432 15580
rect 7380 15496 7432 15502
rect 7484 15484 7512 16612
rect 7944 16538 7972 17190
rect 8024 17128 8076 17134
rect 8024 17070 8076 17076
rect 8036 16794 8064 17070
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7944 16510 8064 16538
rect 7666 16348 7974 16357
rect 7666 16346 7672 16348
rect 7728 16346 7752 16348
rect 7808 16346 7832 16348
rect 7888 16346 7912 16348
rect 7968 16346 7974 16348
rect 7728 16294 7730 16346
rect 7910 16294 7912 16346
rect 7666 16292 7672 16294
rect 7728 16292 7752 16294
rect 7808 16292 7832 16294
rect 7888 16292 7912 16294
rect 7968 16292 7974 16294
rect 7666 16283 7974 16292
rect 7562 15872 7618 15881
rect 7562 15807 7618 15816
rect 7432 15456 7512 15484
rect 7380 15438 7432 15444
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 14618 7420 14758
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7576 14550 7604 15807
rect 7666 15260 7974 15269
rect 7666 15258 7672 15260
rect 7728 15258 7752 15260
rect 7808 15258 7832 15260
rect 7888 15258 7912 15260
rect 7968 15258 7974 15260
rect 7728 15206 7730 15258
rect 7910 15206 7912 15258
rect 7666 15204 7672 15206
rect 7728 15204 7752 15206
rect 7808 15204 7832 15206
rect 7888 15204 7912 15206
rect 7968 15204 7974 15206
rect 7666 15195 7974 15204
rect 8036 14618 8064 16510
rect 8128 15026 8156 20742
rect 8220 20602 8248 21354
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8312 20482 8340 21966
rect 8496 21554 8524 23140
rect 8588 21593 8616 32370
rect 8668 31204 8720 31210
rect 8668 31146 8720 31152
rect 8680 30938 8708 31146
rect 8668 30932 8720 30938
rect 8668 30874 8720 30880
rect 8668 30116 8720 30122
rect 8668 30058 8720 30064
rect 8680 29170 8708 30058
rect 8668 29164 8720 29170
rect 8668 29106 8720 29112
rect 8668 28416 8720 28422
rect 8668 28358 8720 28364
rect 8680 26042 8708 28358
rect 8772 27334 8800 32982
rect 9404 32904 9456 32910
rect 9404 32846 9456 32852
rect 9416 32434 9444 32846
rect 9404 32428 9456 32434
rect 9404 32370 9456 32376
rect 9345 32124 9653 32133
rect 9345 32122 9351 32124
rect 9407 32122 9431 32124
rect 9487 32122 9511 32124
rect 9567 32122 9591 32124
rect 9647 32122 9653 32124
rect 9407 32070 9409 32122
rect 9589 32070 9591 32122
rect 9345 32068 9351 32070
rect 9407 32068 9431 32070
rect 9487 32068 9511 32070
rect 9567 32068 9591 32070
rect 9647 32068 9653 32070
rect 9345 32059 9653 32068
rect 8852 31816 8904 31822
rect 8852 31758 8904 31764
rect 8864 30666 8892 31758
rect 9220 31680 9272 31686
rect 9220 31622 9272 31628
rect 9680 31680 9732 31686
rect 9680 31622 9732 31628
rect 9232 31346 9260 31622
rect 8944 31340 8996 31346
rect 8944 31282 8996 31288
rect 9220 31340 9272 31346
rect 9220 31282 9272 31288
rect 8852 30660 8904 30666
rect 8852 30602 8904 30608
rect 8760 27328 8812 27334
rect 8760 27270 8812 27276
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 8680 24954 8708 25978
rect 8668 24948 8720 24954
rect 8668 24890 8720 24896
rect 8760 23656 8812 23662
rect 8666 23624 8722 23633
rect 8760 23598 8812 23604
rect 8666 23559 8722 23568
rect 8680 22642 8708 23559
rect 8772 23254 8800 23598
rect 8760 23248 8812 23254
rect 8760 23190 8812 23196
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8680 22030 8708 22578
rect 8668 22024 8720 22030
rect 8668 21966 8720 21972
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8574 21584 8630 21593
rect 8484 21548 8536 21554
rect 8772 21554 8800 21830
rect 8574 21519 8630 21528
rect 8760 21548 8812 21554
rect 8484 21490 8536 21496
rect 8496 21146 8524 21490
rect 8484 21140 8536 21146
rect 8484 21082 8536 21088
rect 8484 20800 8536 20806
rect 8484 20742 8536 20748
rect 8220 20454 8340 20482
rect 8220 18850 8248 20454
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 19718 8340 20198
rect 8300 19712 8352 19718
rect 8300 19654 8352 19660
rect 8298 19408 8354 19417
rect 8298 19343 8354 19352
rect 8312 18970 8340 19343
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8220 18822 8340 18850
rect 8312 18748 8340 18822
rect 8206 18728 8262 18737
rect 8312 18720 8432 18748
rect 8206 18663 8262 18672
rect 8220 18630 8248 18663
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 7944 14328 7972 14486
rect 7944 14300 8064 14328
rect 7656 14272 7708 14278
rect 7576 14232 7656 14260
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7300 13138 7328 14010
rect 7576 13938 7604 14232
rect 7656 14214 7708 14220
rect 7666 14172 7974 14181
rect 7666 14170 7672 14172
rect 7728 14170 7752 14172
rect 7808 14170 7832 14172
rect 7888 14170 7912 14172
rect 7968 14170 7974 14172
rect 7728 14118 7730 14170
rect 7910 14118 7912 14170
rect 7666 14116 7672 14118
rect 7728 14116 7752 14118
rect 7808 14116 7832 14118
rect 7888 14116 7912 14118
rect 7968 14116 7974 14118
rect 7666 14107 7974 14116
rect 7654 13968 7710 13977
rect 7564 13932 7616 13938
rect 7654 13903 7710 13912
rect 7564 13874 7616 13880
rect 7668 13802 7696 13903
rect 7840 13864 7892 13870
rect 7840 13806 7892 13812
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7562 13696 7618 13705
rect 7618 13654 7696 13682
rect 7562 13631 7618 13640
rect 7668 13326 7696 13654
rect 7852 13530 7880 13806
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 7656 13320 7708 13326
rect 7576 13280 7656 13308
rect 7300 13110 7420 13138
rect 7288 12980 7340 12986
rect 7288 12922 7340 12928
rect 7300 12850 7328 12922
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7012 12232 7064 12238
rect 7012 12174 7064 12180
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 7116 11694 7144 12242
rect 7392 12238 7420 13110
rect 7380 12232 7432 12238
rect 7576 12186 7604 13280
rect 7656 13262 7708 13268
rect 7666 13084 7974 13093
rect 7666 13082 7672 13084
rect 7728 13082 7752 13084
rect 7808 13082 7832 13084
rect 7888 13082 7912 13084
rect 7968 13082 7974 13084
rect 7728 13030 7730 13082
rect 7910 13030 7912 13082
rect 7666 13028 7672 13030
rect 7728 13028 7752 13030
rect 7808 13028 7832 13030
rect 7888 13028 7912 13030
rect 7968 13028 7974 13030
rect 7666 13019 7974 13028
rect 7380 12174 7432 12180
rect 7484 12158 7604 12186
rect 7196 12096 7248 12102
rect 7196 12038 7248 12044
rect 7104 11688 7156 11694
rect 6840 11614 7052 11642
rect 7104 11630 7156 11636
rect 5920 10968 6408 10996
rect 6472 11478 6776 11506
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5644 10062 5672 10610
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5736 10266 5764 10406
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5184 9646 5304 9674
rect 5184 7313 5212 9646
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5552 7886 5580 8774
rect 5920 8566 5948 10968
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 5987 10364 6295 10373
rect 5987 10362 5993 10364
rect 6049 10362 6073 10364
rect 6129 10362 6153 10364
rect 6209 10362 6233 10364
rect 6289 10362 6295 10364
rect 6049 10310 6051 10362
rect 6231 10310 6233 10362
rect 5987 10308 5993 10310
rect 6049 10308 6073 10310
rect 6129 10308 6153 10310
rect 6209 10308 6233 10310
rect 6289 10308 6295 10310
rect 5987 10299 6295 10308
rect 6380 9994 6408 10610
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 5987 9276 6295 9285
rect 5987 9274 5993 9276
rect 6049 9274 6073 9276
rect 6129 9274 6153 9276
rect 6209 9274 6233 9276
rect 6289 9274 6295 9276
rect 6049 9222 6051 9274
rect 6231 9222 6233 9274
rect 5987 9220 5993 9222
rect 6049 9220 6073 9222
rect 6129 9220 6153 9222
rect 6209 9220 6233 9222
rect 6289 9220 6295 9222
rect 5987 9211 6295 9220
rect 5908 8560 5960 8566
rect 5906 8528 5908 8537
rect 5960 8528 5962 8537
rect 5906 8463 5962 8472
rect 5987 8188 6295 8197
rect 5987 8186 5993 8188
rect 6049 8186 6073 8188
rect 6129 8186 6153 8188
rect 6209 8186 6233 8188
rect 6289 8186 6295 8188
rect 6049 8134 6051 8186
rect 6231 8134 6233 8186
rect 5987 8132 5993 8134
rect 6049 8132 6073 8134
rect 6129 8132 6153 8134
rect 6209 8132 6233 8134
rect 6289 8132 6295 8134
rect 5987 8123 6295 8132
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5170 7304 5226 7313
rect 5170 7239 5226 7248
rect 5987 7100 6295 7109
rect 5987 7098 5993 7100
rect 6049 7098 6073 7100
rect 6129 7098 6153 7100
rect 6209 7098 6233 7100
rect 6289 7098 6295 7100
rect 6049 7046 6051 7098
rect 6231 7046 6233 7098
rect 5987 7044 5993 7046
rect 6049 7044 6073 7046
rect 6129 7044 6153 7046
rect 6209 7044 6233 7046
rect 6289 7044 6295 7046
rect 5987 7035 6295 7044
rect 6472 6390 6500 11478
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6564 10266 6592 10542
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6656 10146 6684 11290
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6932 10810 6960 11086
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6736 10464 6788 10470
rect 6736 10406 6788 10412
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6748 10266 6776 10406
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6564 10118 6684 10146
rect 6828 10124 6880 10130
rect 6564 10062 6592 10118
rect 6828 10066 6880 10072
rect 6552 10056 6604 10062
rect 6552 9998 6604 10004
rect 6840 9722 6868 10066
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6736 8492 6788 8498
rect 6736 8434 6788 8440
rect 6748 8090 6776 8434
rect 6736 8084 6788 8090
rect 6736 8026 6788 8032
rect 6932 7954 6960 10406
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7880 6880 7886
rect 6828 7822 6880 7828
rect 6840 7546 6868 7822
rect 6828 7540 6880 7546
rect 6828 7482 6880 7488
rect 6460 6384 6512 6390
rect 6460 6326 6512 6332
rect 5987 6012 6295 6021
rect 5987 6010 5993 6012
rect 6049 6010 6073 6012
rect 6129 6010 6153 6012
rect 6209 6010 6233 6012
rect 6289 6010 6295 6012
rect 6049 5958 6051 6010
rect 6231 5958 6233 6010
rect 5987 5956 5993 5958
rect 6049 5956 6073 5958
rect 6129 5956 6153 5958
rect 6209 5956 6233 5958
rect 6289 5956 6295 5958
rect 5987 5947 6295 5956
rect 7024 5234 7052 11614
rect 7208 11150 7236 12038
rect 7288 11756 7340 11762
rect 7340 11716 7420 11744
rect 7288 11698 7340 11704
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7104 11144 7156 11150
rect 7104 11086 7156 11092
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7116 10674 7144 11086
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7104 10192 7156 10198
rect 7104 10134 7156 10140
rect 7116 7993 7144 10134
rect 7208 10130 7236 11086
rect 7300 10130 7328 11494
rect 7196 10124 7248 10130
rect 7196 10066 7248 10072
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7392 9674 7420 11716
rect 7484 11200 7512 12158
rect 7666 11996 7974 12005
rect 7666 11994 7672 11996
rect 7728 11994 7752 11996
rect 7808 11994 7832 11996
rect 7888 11994 7912 11996
rect 7968 11994 7974 11996
rect 7728 11942 7730 11994
rect 7910 11942 7912 11994
rect 7666 11940 7672 11942
rect 7728 11940 7752 11942
rect 7808 11940 7832 11942
rect 7888 11940 7912 11942
rect 7968 11940 7974 11942
rect 7666 11931 7974 11940
rect 8036 11830 8064 14300
rect 8128 12434 8156 14962
rect 8220 13326 8248 18566
rect 8312 18290 8340 18566
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8404 18170 8432 18720
rect 8312 18142 8432 18170
rect 8312 16182 8340 18142
rect 8496 18057 8524 20742
rect 8588 18970 8616 21519
rect 8760 21490 8812 21496
rect 8864 21400 8892 30602
rect 8956 30054 8984 31282
rect 9128 31136 9180 31142
rect 9128 31078 9180 31084
rect 9220 31136 9272 31142
rect 9220 31078 9272 31084
rect 9036 30932 9088 30938
rect 9036 30874 9088 30880
rect 9048 30598 9076 30874
rect 9036 30592 9088 30598
rect 9036 30534 9088 30540
rect 9140 30190 9168 31078
rect 9232 30682 9260 31078
rect 9345 31036 9653 31045
rect 9345 31034 9351 31036
rect 9407 31034 9431 31036
rect 9487 31034 9511 31036
rect 9567 31034 9591 31036
rect 9647 31034 9653 31036
rect 9407 30982 9409 31034
rect 9589 30982 9591 31034
rect 9345 30980 9351 30982
rect 9407 30980 9431 30982
rect 9487 30980 9511 30982
rect 9567 30980 9591 30982
rect 9647 30980 9653 30982
rect 9345 30971 9653 30980
rect 9692 30734 9720 31622
rect 9784 31278 9812 34342
rect 9876 34202 9904 35158
rect 10416 35012 10468 35018
rect 10416 34954 10468 34960
rect 10428 34202 10456 34954
rect 9864 34196 9916 34202
rect 9864 34138 9916 34144
rect 10416 34196 10468 34202
rect 10416 34138 10468 34144
rect 9956 34060 10008 34066
rect 9956 34002 10008 34008
rect 10060 34054 10180 34082
rect 9864 33992 9916 33998
rect 9862 33960 9864 33969
rect 9916 33960 9918 33969
rect 9862 33895 9918 33904
rect 9864 33856 9916 33862
rect 9864 33798 9916 33804
rect 9876 33658 9904 33798
rect 9864 33652 9916 33658
rect 9864 33594 9916 33600
rect 9864 32360 9916 32366
rect 9864 32302 9916 32308
rect 9876 31482 9904 32302
rect 9864 31476 9916 31482
rect 9864 31418 9916 31424
rect 9772 31272 9824 31278
rect 9772 31214 9824 31220
rect 9968 30938 9996 34002
rect 9956 30932 10008 30938
rect 9956 30874 10008 30880
rect 9680 30728 9732 30734
rect 9232 30654 9352 30682
rect 9680 30670 9732 30676
rect 9220 30592 9272 30598
rect 9220 30534 9272 30540
rect 9036 30184 9088 30190
rect 9036 30126 9088 30132
rect 9128 30184 9180 30190
rect 9128 30126 9180 30132
rect 8944 30048 8996 30054
rect 8944 29990 8996 29996
rect 8944 29572 8996 29578
rect 8944 29514 8996 29520
rect 8956 28558 8984 29514
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 8944 28416 8996 28422
rect 8944 28358 8996 28364
rect 8956 28121 8984 28358
rect 8942 28112 8998 28121
rect 8942 28047 8998 28056
rect 8956 28014 8984 28047
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 8944 27872 8996 27878
rect 8942 27840 8944 27849
rect 8996 27840 8998 27849
rect 8942 27775 8998 27784
rect 8956 27554 8984 27775
rect 9048 27713 9076 30126
rect 9140 29073 9168 30126
rect 9126 29064 9182 29073
rect 9126 28999 9182 29008
rect 9232 28948 9260 30534
rect 9324 30122 9352 30654
rect 9588 30592 9640 30598
rect 9588 30534 9640 30540
rect 9600 30190 9628 30534
rect 9588 30184 9640 30190
rect 9588 30126 9640 30132
rect 9312 30116 9364 30122
rect 9312 30058 9364 30064
rect 9345 29948 9653 29957
rect 9345 29946 9351 29948
rect 9407 29946 9431 29948
rect 9487 29946 9511 29948
rect 9567 29946 9591 29948
rect 9647 29946 9653 29948
rect 9407 29894 9409 29946
rect 9589 29894 9591 29946
rect 9345 29892 9351 29894
rect 9407 29892 9431 29894
rect 9487 29892 9511 29894
rect 9567 29892 9591 29894
rect 9647 29892 9653 29894
rect 9345 29883 9653 29892
rect 9692 29646 9720 30670
rect 10060 30274 10088 34054
rect 10152 33998 10180 34054
rect 10140 33992 10192 33998
rect 10140 33934 10192 33940
rect 10324 32904 10376 32910
rect 10324 32846 10376 32852
rect 10140 32768 10192 32774
rect 10140 32710 10192 32716
rect 10152 32570 10180 32710
rect 10140 32564 10192 32570
rect 10140 32506 10192 32512
rect 10140 32224 10192 32230
rect 10192 32184 10272 32212
rect 10140 32166 10192 32172
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 9876 30246 10088 30274
rect 9680 29640 9732 29646
rect 9680 29582 9732 29588
rect 9692 29510 9720 29582
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9772 29504 9824 29510
rect 9772 29446 9824 29452
rect 9692 29102 9720 29446
rect 9784 29170 9812 29446
rect 9772 29164 9824 29170
rect 9772 29106 9824 29112
rect 9680 29096 9732 29102
rect 9680 29038 9732 29044
rect 9140 28920 9260 28948
rect 9034 27704 9090 27713
rect 9034 27639 9090 27648
rect 8956 27526 9076 27554
rect 8944 25288 8996 25294
rect 8944 25230 8996 25236
rect 8772 21372 8892 21400
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8680 18714 8708 21286
rect 8772 20398 8800 21372
rect 8956 21350 8984 25230
rect 9048 24018 9076 27526
rect 9140 26518 9168 28920
rect 9345 28860 9653 28869
rect 9345 28858 9351 28860
rect 9407 28858 9431 28860
rect 9487 28858 9511 28860
rect 9567 28858 9591 28860
rect 9647 28858 9653 28860
rect 9407 28806 9409 28858
rect 9589 28806 9591 28858
rect 9345 28804 9351 28806
rect 9407 28804 9431 28806
rect 9487 28804 9511 28806
rect 9567 28804 9591 28806
rect 9647 28804 9653 28806
rect 9345 28795 9653 28804
rect 9220 28552 9272 28558
rect 9220 28494 9272 28500
rect 9128 26512 9180 26518
rect 9128 26454 9180 26460
rect 9140 24206 9168 26454
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9048 23990 9168 24018
rect 9036 22976 9088 22982
rect 9036 22918 9088 22924
rect 9048 22545 9076 22918
rect 9034 22536 9090 22545
rect 9034 22471 9090 22480
rect 9140 22094 9168 23990
rect 9232 23866 9260 28494
rect 9680 28416 9732 28422
rect 9680 28358 9732 28364
rect 9312 28008 9364 28014
rect 9692 27985 9720 28358
rect 9312 27950 9364 27956
rect 9678 27976 9734 27985
rect 9324 27860 9352 27950
rect 9678 27911 9734 27920
rect 9324 27832 9720 27860
rect 9345 27772 9653 27781
rect 9345 27770 9351 27772
rect 9407 27770 9431 27772
rect 9487 27770 9511 27772
rect 9567 27770 9591 27772
rect 9647 27770 9653 27772
rect 9407 27718 9409 27770
rect 9589 27718 9591 27770
rect 9345 27716 9351 27718
rect 9407 27716 9431 27718
rect 9487 27716 9511 27718
rect 9567 27716 9591 27718
rect 9647 27716 9653 27718
rect 9345 27707 9653 27716
rect 9692 27606 9720 27832
rect 9680 27600 9732 27606
rect 9680 27542 9732 27548
rect 9680 27328 9732 27334
rect 9680 27270 9732 27276
rect 9692 26994 9720 27270
rect 9680 26988 9732 26994
rect 9680 26930 9732 26936
rect 9345 26684 9653 26693
rect 9345 26682 9351 26684
rect 9407 26682 9431 26684
rect 9487 26682 9511 26684
rect 9567 26682 9591 26684
rect 9647 26682 9653 26684
rect 9407 26630 9409 26682
rect 9589 26630 9591 26682
rect 9345 26628 9351 26630
rect 9407 26628 9431 26630
rect 9487 26628 9511 26630
rect 9567 26628 9591 26630
rect 9647 26628 9653 26630
rect 9345 26619 9653 26628
rect 9692 26568 9720 26930
rect 9600 26540 9720 26568
rect 9600 26246 9628 26540
rect 9588 26240 9640 26246
rect 9588 26182 9640 26188
rect 9600 25770 9628 26182
rect 9588 25764 9640 25770
rect 9588 25706 9640 25712
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9345 25596 9653 25605
rect 9345 25594 9351 25596
rect 9407 25594 9431 25596
rect 9487 25594 9511 25596
rect 9567 25594 9591 25596
rect 9647 25594 9653 25596
rect 9407 25542 9409 25594
rect 9589 25542 9591 25594
rect 9345 25540 9351 25542
rect 9407 25540 9431 25542
rect 9487 25540 9511 25542
rect 9567 25540 9591 25542
rect 9647 25540 9653 25542
rect 9345 25531 9653 25540
rect 9692 25265 9720 25638
rect 9678 25256 9734 25265
rect 9678 25191 9734 25200
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9600 24834 9628 24890
rect 9600 24806 9720 24834
rect 9345 24508 9653 24517
rect 9345 24506 9351 24508
rect 9407 24506 9431 24508
rect 9487 24506 9511 24508
rect 9567 24506 9591 24508
rect 9647 24506 9653 24508
rect 9407 24454 9409 24506
rect 9589 24454 9591 24506
rect 9345 24452 9351 24454
rect 9407 24452 9431 24454
rect 9487 24452 9511 24454
rect 9567 24452 9591 24454
rect 9647 24452 9653 24454
rect 9345 24443 9653 24452
rect 9692 23866 9720 24806
rect 9220 23860 9272 23866
rect 9220 23802 9272 23808
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9680 23656 9732 23662
rect 9678 23624 9680 23633
rect 9732 23624 9734 23633
rect 9678 23559 9734 23568
rect 9345 23420 9653 23429
rect 9345 23418 9351 23420
rect 9407 23418 9431 23420
rect 9487 23418 9511 23420
rect 9567 23418 9591 23420
rect 9647 23418 9653 23420
rect 9407 23366 9409 23418
rect 9589 23366 9591 23418
rect 9345 23364 9351 23366
rect 9407 23364 9431 23366
rect 9487 23364 9511 23366
rect 9567 23364 9591 23366
rect 9647 23364 9653 23366
rect 9345 23355 9653 23364
rect 9680 22704 9732 22710
rect 9680 22646 9732 22652
rect 9345 22332 9653 22341
rect 9345 22330 9351 22332
rect 9407 22330 9431 22332
rect 9487 22330 9511 22332
rect 9567 22330 9591 22332
rect 9647 22330 9653 22332
rect 9407 22278 9409 22330
rect 9589 22278 9591 22330
rect 9345 22276 9351 22278
rect 9407 22276 9431 22278
rect 9487 22276 9511 22278
rect 9567 22276 9591 22278
rect 9647 22276 9653 22278
rect 9345 22267 9653 22276
rect 9048 22066 9168 22094
rect 8944 21344 8996 21350
rect 8944 21286 8996 21292
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 8852 20936 8904 20942
rect 8852 20878 8904 20884
rect 8760 20392 8812 20398
rect 8760 20334 8812 20340
rect 8772 19786 8800 20334
rect 8864 19802 8892 20878
rect 8956 20074 8984 21082
rect 9048 20262 9076 22066
rect 9312 22024 9364 22030
rect 9312 21966 9364 21972
rect 9402 21992 9458 22001
rect 9128 21956 9180 21962
rect 9128 21898 9180 21904
rect 9140 20602 9168 21898
rect 9324 21486 9352 21966
rect 9402 21927 9458 21936
rect 9416 21690 9444 21927
rect 9404 21684 9456 21690
rect 9404 21626 9456 21632
rect 9312 21480 9364 21486
rect 9232 21440 9312 21468
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 9140 20466 9168 20538
rect 9128 20460 9180 20466
rect 9128 20402 9180 20408
rect 9128 20324 9180 20330
rect 9128 20266 9180 20272
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 8956 20046 9076 20074
rect 8942 19952 8998 19961
rect 8942 19887 8944 19896
rect 8996 19887 8998 19896
rect 8944 19858 8996 19864
rect 8760 19780 8812 19786
rect 8864 19774 8984 19802
rect 8760 19722 8812 19728
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8864 19310 8892 19654
rect 8956 19378 8984 19774
rect 8944 19372 8996 19378
rect 8944 19314 8996 19320
rect 8760 19304 8812 19310
rect 8760 19246 8812 19252
rect 8852 19304 8904 19310
rect 8852 19246 8904 19252
rect 8588 18686 8708 18714
rect 8482 18048 8538 18057
rect 8482 17983 8538 17992
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8496 17338 8524 17478
rect 8484 17332 8536 17338
rect 8484 17274 8536 17280
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8404 16522 8432 17070
rect 8496 16794 8524 17274
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8392 16516 8444 16522
rect 8392 16458 8444 16464
rect 8300 16176 8352 16182
rect 8300 16118 8352 16124
rect 8404 16046 8432 16458
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8392 15904 8444 15910
rect 8392 15846 8444 15852
rect 8404 14958 8432 15846
rect 8300 14952 8352 14958
rect 8300 14894 8352 14900
rect 8392 14952 8444 14958
rect 8392 14894 8444 14900
rect 8312 14328 8340 14894
rect 8588 14618 8616 18686
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8680 17338 8708 18566
rect 8772 18193 8800 19246
rect 8852 19168 8904 19174
rect 8850 19136 8852 19145
rect 8904 19136 8906 19145
rect 8850 19071 8906 19080
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8758 18184 8814 18193
rect 8758 18119 8814 18128
rect 8864 17882 8892 18770
rect 8852 17876 8904 17882
rect 8852 17818 8904 17824
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8668 17196 8720 17202
rect 8668 17138 8720 17144
rect 8680 16454 8708 17138
rect 8864 16658 8892 17274
rect 8852 16652 8904 16658
rect 8852 16594 8904 16600
rect 8668 16448 8720 16454
rect 8720 16396 8800 16402
rect 8668 16390 8800 16396
rect 8680 16374 8800 16390
rect 8668 14884 8720 14890
rect 8668 14826 8720 14832
rect 8576 14612 8628 14618
rect 8496 14572 8576 14600
rect 8392 14340 8444 14346
rect 8312 14300 8392 14328
rect 8392 14282 8444 14288
rect 8496 14056 8524 14572
rect 8576 14554 8628 14560
rect 8576 14340 8628 14346
rect 8576 14282 8628 14288
rect 8312 14028 8524 14056
rect 8312 13870 8340 14028
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8208 13320 8260 13326
rect 8208 13262 8260 13268
rect 8128 12406 8248 12434
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 7760 11286 7788 11766
rect 7748 11280 7800 11286
rect 7748 11222 7800 11228
rect 7484 11172 7696 11200
rect 7668 11132 7696 11172
rect 7470 11112 7526 11121
rect 7668 11104 8064 11132
rect 7470 11047 7526 11056
rect 7300 9646 7420 9674
rect 7300 8838 7328 9646
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 8974 7420 9318
rect 7380 8968 7432 8974
rect 7380 8910 7432 8916
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7208 8090 7236 8434
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7102 7984 7158 7993
rect 7102 7919 7158 7928
rect 7116 7886 7144 7919
rect 7104 7880 7156 7886
rect 7288 7880 7340 7886
rect 7104 7822 7156 7828
rect 7194 7848 7250 7857
rect 7288 7822 7340 7828
rect 7194 7783 7250 7792
rect 7208 7410 7236 7783
rect 7300 7449 7328 7822
rect 7286 7440 7342 7449
rect 7196 7404 7248 7410
rect 7286 7375 7342 7384
rect 7196 7346 7248 7352
rect 7392 6662 7420 8910
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6322 7420 6598
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7392 5914 7420 6258
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 7392 5166 7420 5850
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 5987 4924 6295 4933
rect 5987 4922 5993 4924
rect 6049 4922 6073 4924
rect 6129 4922 6153 4924
rect 6209 4922 6233 4924
rect 6289 4922 6295 4924
rect 6049 4870 6051 4922
rect 6231 4870 6233 4922
rect 5987 4868 5993 4870
rect 6049 4868 6073 4870
rect 6129 4868 6153 4870
rect 6209 4868 6233 4870
rect 6289 4868 6295 4870
rect 5987 4859 6295 4868
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5987 3836 6295 3845
rect 5987 3834 5993 3836
rect 6049 3834 6073 3836
rect 6129 3834 6153 3836
rect 6209 3834 6233 3836
rect 6289 3834 6295 3836
rect 6049 3782 6051 3834
rect 6231 3782 6233 3834
rect 5987 3780 5993 3782
rect 6049 3780 6073 3782
rect 6129 3780 6153 3782
rect 6209 3780 6233 3782
rect 6289 3780 6295 3782
rect 5987 3771 6295 3780
rect 4308 3292 4616 3301
rect 4308 3290 4314 3292
rect 4370 3290 4394 3292
rect 4450 3290 4474 3292
rect 4530 3290 4554 3292
rect 4610 3290 4616 3292
rect 4370 3238 4372 3290
rect 4552 3238 4554 3290
rect 4308 3236 4314 3238
rect 4370 3236 4394 3238
rect 4450 3236 4474 3238
rect 4530 3236 4554 3238
rect 4610 3236 4616 3238
rect 4308 3227 4616 3236
rect 5987 2748 6295 2757
rect 5987 2746 5993 2748
rect 6049 2746 6073 2748
rect 6129 2746 6153 2748
rect 6209 2746 6233 2748
rect 6289 2746 6295 2748
rect 6049 2694 6051 2746
rect 6231 2694 6233 2746
rect 5987 2692 5993 2694
rect 6049 2692 6073 2694
rect 6129 2692 6153 2694
rect 6209 2692 6233 2694
rect 6289 2692 6295 2694
rect 5987 2683 6295 2692
rect 6642 2680 6698 2689
rect 6642 2615 6698 2624
rect 4308 2204 4616 2213
rect 4308 2202 4314 2204
rect 4370 2202 4394 2204
rect 4450 2202 4474 2204
rect 4530 2202 4554 2204
rect 4610 2202 4616 2204
rect 4370 2150 4372 2202
rect 4552 2150 4554 2202
rect 4308 2148 4314 2150
rect 4370 2148 4394 2150
rect 4450 2148 4474 2150
rect 4530 2148 4554 2150
rect 4610 2148 4616 2150
rect 4308 2139 4616 2148
rect 6656 2106 6684 2615
rect 7194 2544 7250 2553
rect 7194 2479 7250 2488
rect 7208 2106 7236 2479
rect 7484 2106 7512 11047
rect 7666 10908 7974 10917
rect 7666 10906 7672 10908
rect 7728 10906 7752 10908
rect 7808 10906 7832 10908
rect 7888 10906 7912 10908
rect 7968 10906 7974 10908
rect 7728 10854 7730 10906
rect 7910 10854 7912 10906
rect 7666 10852 7672 10854
rect 7728 10852 7752 10854
rect 7808 10852 7832 10854
rect 7888 10852 7912 10854
rect 7968 10852 7974 10854
rect 7666 10843 7974 10852
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7576 10062 7604 10746
rect 7656 10464 7708 10470
rect 7656 10406 7708 10412
rect 7668 10062 7696 10406
rect 7564 10056 7616 10062
rect 7564 9998 7616 10004
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7576 8616 7604 9998
rect 7666 9820 7974 9829
rect 7666 9818 7672 9820
rect 7728 9818 7752 9820
rect 7808 9818 7832 9820
rect 7888 9818 7912 9820
rect 7968 9818 7974 9820
rect 7728 9766 7730 9818
rect 7910 9766 7912 9818
rect 7666 9764 7672 9766
rect 7728 9764 7752 9766
rect 7808 9764 7832 9766
rect 7888 9764 7912 9766
rect 7968 9764 7974 9766
rect 7666 9755 7974 9764
rect 7666 8732 7974 8741
rect 7666 8730 7672 8732
rect 7728 8730 7752 8732
rect 7808 8730 7832 8732
rect 7888 8730 7912 8732
rect 7968 8730 7974 8732
rect 7728 8678 7730 8730
rect 7910 8678 7912 8730
rect 7666 8676 7672 8678
rect 7728 8676 7752 8678
rect 7808 8676 7832 8678
rect 7888 8676 7912 8678
rect 7968 8676 7974 8678
rect 7666 8667 7974 8676
rect 7576 8588 7696 8616
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7576 7342 7604 7890
rect 7668 7857 7696 8588
rect 8036 8129 8064 11104
rect 8128 10470 8156 12038
rect 8220 11830 8248 12406
rect 8208 11824 8260 11830
rect 8208 11766 8260 11772
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8220 10713 8248 10746
rect 8206 10704 8262 10713
rect 8206 10639 8262 10648
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8220 9466 8248 9658
rect 8312 9586 8340 13466
rect 8404 12986 8432 13874
rect 8484 13320 8536 13326
rect 8588 13297 8616 14282
rect 8484 13262 8536 13268
rect 8574 13288 8630 13297
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 8496 11370 8524 13262
rect 8574 13223 8630 13232
rect 8680 13190 8708 14826
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8588 12986 8616 13126
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8680 12646 8708 12786
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8496 11342 8616 11370
rect 8484 11280 8536 11286
rect 8484 11222 8536 11228
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8404 10742 8432 11154
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8300 9580 8352 9586
rect 8300 9522 8352 9528
rect 8220 9438 8340 9466
rect 8312 8650 8340 9438
rect 8404 8838 8432 10678
rect 8496 8974 8524 11222
rect 8588 9722 8616 11342
rect 8680 10742 8708 11494
rect 8668 10736 8720 10742
rect 8668 10678 8720 10684
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8576 9716 8628 9722
rect 8576 9658 8628 9664
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8392 8832 8444 8838
rect 8496 8809 8524 8910
rect 8392 8774 8444 8780
rect 8482 8800 8538 8809
rect 8482 8735 8538 8744
rect 8312 8622 8524 8650
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8208 8356 8260 8362
rect 8208 8298 8260 8304
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8022 8120 8078 8129
rect 7932 8084 7984 8090
rect 8022 8055 8078 8064
rect 7932 8026 7984 8032
rect 7840 7948 7892 7954
rect 7944 7936 7972 8026
rect 8128 7954 8156 8230
rect 8024 7948 8076 7954
rect 7944 7908 8024 7936
rect 7840 7890 7892 7896
rect 8024 7890 8076 7896
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 7654 7848 7710 7857
rect 7852 7834 7880 7890
rect 7852 7806 8064 7834
rect 7654 7783 7710 7792
rect 7666 7644 7974 7653
rect 7666 7642 7672 7644
rect 7728 7642 7752 7644
rect 7808 7642 7832 7644
rect 7888 7642 7912 7644
rect 7968 7642 7974 7644
rect 7728 7590 7730 7642
rect 7910 7590 7912 7642
rect 7666 7588 7672 7590
rect 7728 7588 7752 7590
rect 7808 7588 7832 7590
rect 7888 7588 7912 7590
rect 7968 7588 7974 7590
rect 7666 7579 7974 7588
rect 8036 7562 8064 7806
rect 8114 7576 8170 7585
rect 8036 7534 8114 7562
rect 8114 7511 8170 7520
rect 8220 7410 8248 8298
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 7564 7336 7616 7342
rect 7564 7278 7616 7284
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7576 7002 7604 7278
rect 7944 7002 7972 7278
rect 8312 7002 8340 8366
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 7342 8432 8230
rect 8392 7336 8444 7342
rect 8392 7278 8444 7284
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 7666 6556 7974 6565
rect 7666 6554 7672 6556
rect 7728 6554 7752 6556
rect 7808 6554 7832 6556
rect 7888 6554 7912 6556
rect 7968 6554 7974 6556
rect 7728 6502 7730 6554
rect 7910 6502 7912 6554
rect 7666 6500 7672 6502
rect 7728 6500 7752 6502
rect 7808 6500 7832 6502
rect 7888 6500 7912 6502
rect 7968 6500 7974 6502
rect 7666 6491 7974 6500
rect 8220 6225 8248 6666
rect 8206 6216 8262 6225
rect 8206 6151 8262 6160
rect 8404 5914 8432 7278
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8300 5704 8352 5710
rect 8298 5672 8300 5681
rect 8352 5672 8354 5681
rect 8298 5607 8354 5616
rect 7666 5468 7974 5477
rect 7666 5466 7672 5468
rect 7728 5466 7752 5468
rect 7808 5466 7832 5468
rect 7888 5466 7912 5468
rect 7968 5466 7974 5468
rect 7728 5414 7730 5466
rect 7910 5414 7912 5466
rect 7666 5412 7672 5414
rect 7728 5412 7752 5414
rect 7808 5412 7832 5414
rect 7888 5412 7912 5414
rect 7968 5412 7974 5414
rect 7666 5403 7974 5412
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8220 4690 8248 5102
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 7666 4380 7974 4389
rect 7666 4378 7672 4380
rect 7728 4378 7752 4380
rect 7808 4378 7832 4380
rect 7888 4378 7912 4380
rect 7968 4378 7974 4380
rect 7728 4326 7730 4378
rect 7910 4326 7912 4378
rect 7666 4324 7672 4326
rect 7728 4324 7752 4326
rect 7808 4324 7832 4326
rect 7888 4324 7912 4326
rect 7968 4324 7974 4326
rect 7666 4315 7974 4324
rect 8496 3738 8524 8622
rect 8588 6322 8616 9522
rect 8680 6866 8708 10066
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8588 5914 8616 6258
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8680 5846 8708 6802
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8772 5370 8800 16374
rect 8852 15496 8904 15502
rect 8852 15438 8904 15444
rect 8864 13530 8892 15438
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8956 13512 8984 19314
rect 9048 18086 9076 20046
rect 9140 19854 9168 20266
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9036 18080 9088 18086
rect 9036 18022 9088 18028
rect 9232 16658 9260 21440
rect 9312 21422 9364 21428
rect 9345 21244 9653 21253
rect 9345 21242 9351 21244
rect 9407 21242 9431 21244
rect 9487 21242 9511 21244
rect 9567 21242 9591 21244
rect 9647 21242 9653 21244
rect 9407 21190 9409 21242
rect 9589 21190 9591 21242
rect 9345 21188 9351 21190
rect 9407 21188 9431 21190
rect 9487 21188 9511 21190
rect 9567 21188 9591 21190
rect 9647 21188 9653 21190
rect 9345 21179 9653 21188
rect 9692 21026 9720 22646
rect 9784 22545 9812 29106
rect 9876 26489 9904 30246
rect 10048 30184 10100 30190
rect 10048 30126 10100 30132
rect 10060 28121 10088 30126
rect 10152 29170 10180 31758
rect 10244 30258 10272 32184
rect 10336 30938 10364 32846
rect 10520 32842 10548 36178
rect 10612 35834 10640 36790
rect 10876 36168 10928 36174
rect 10876 36110 10928 36116
rect 10888 35834 10916 36110
rect 11024 35932 11332 35941
rect 11024 35930 11030 35932
rect 11086 35930 11110 35932
rect 11166 35930 11190 35932
rect 11246 35930 11270 35932
rect 11326 35930 11332 35932
rect 11086 35878 11088 35930
rect 11268 35878 11270 35930
rect 11024 35876 11030 35878
rect 11086 35876 11110 35878
rect 11166 35876 11190 35878
rect 11246 35876 11270 35878
rect 11326 35876 11332 35878
rect 11024 35867 11332 35876
rect 11440 35834 11468 36887
rect 11992 36786 12020 37062
rect 11980 36780 12032 36786
rect 11980 36722 12032 36728
rect 12176 36582 12204 38422
rect 12268 37398 12296 38830
rect 12440 38820 12492 38826
rect 12440 38762 12492 38768
rect 12452 38026 12480 38762
rect 13084 38752 13136 38758
rect 13084 38694 13136 38700
rect 13360 38752 13412 38758
rect 13360 38694 13412 38700
rect 12703 38652 13011 38661
rect 12703 38650 12709 38652
rect 12765 38650 12789 38652
rect 12845 38650 12869 38652
rect 12925 38650 12949 38652
rect 13005 38650 13011 38652
rect 12765 38598 12767 38650
rect 12947 38598 12949 38650
rect 12703 38596 12709 38598
rect 12765 38596 12789 38598
rect 12845 38596 12869 38598
rect 12925 38596 12949 38598
rect 13005 38596 13011 38598
rect 12703 38587 13011 38596
rect 12624 38344 12676 38350
rect 12360 38010 12480 38026
rect 12348 38004 12480 38010
rect 12400 37998 12480 38004
rect 12544 38292 12624 38298
rect 12544 38286 12676 38292
rect 12544 38270 12664 38286
rect 12348 37946 12400 37952
rect 12256 37392 12308 37398
rect 12256 37334 12308 37340
rect 12544 37346 12572 38270
rect 12624 38208 12676 38214
rect 12624 38150 12676 38156
rect 12636 38010 12664 38150
rect 12624 38004 12676 38010
rect 12624 37946 12676 37952
rect 13096 37942 13124 38694
rect 13372 38457 13400 38694
rect 13648 38554 13676 38898
rect 13912 38752 13964 38758
rect 13910 38720 13912 38729
rect 13964 38720 13966 38729
rect 13910 38655 13966 38664
rect 13636 38548 13688 38554
rect 13636 38490 13688 38496
rect 13452 38480 13504 38486
rect 13358 38448 13414 38457
rect 13452 38422 13504 38428
rect 13358 38383 13414 38392
rect 13360 38276 13412 38282
rect 13360 38218 13412 38224
rect 13372 38010 13400 38218
rect 13464 38010 13492 38422
rect 13360 38004 13412 38010
rect 13360 37946 13412 37952
rect 13452 38004 13504 38010
rect 13452 37946 13504 37952
rect 13084 37936 13136 37942
rect 13084 37878 13136 37884
rect 12624 37868 12676 37874
rect 12624 37810 12676 37816
rect 12636 37466 12664 37810
rect 13728 37664 13780 37670
rect 13728 37606 13780 37612
rect 12703 37564 13011 37573
rect 12703 37562 12709 37564
rect 12765 37562 12789 37564
rect 12845 37562 12869 37564
rect 12925 37562 12949 37564
rect 13005 37562 13011 37564
rect 12765 37510 12767 37562
rect 12947 37510 12949 37562
rect 12703 37508 12709 37510
rect 12765 37508 12789 37510
rect 12845 37508 12869 37510
rect 12925 37508 12949 37510
rect 13005 37508 13011 37510
rect 12703 37499 13011 37508
rect 12624 37460 12676 37466
rect 12624 37402 12676 37408
rect 12348 37324 12400 37330
rect 12544 37318 12848 37346
rect 12348 37266 12400 37272
rect 12360 37233 12388 37266
rect 12624 37256 12676 37262
rect 12346 37224 12402 37233
rect 12624 37198 12676 37204
rect 12716 37256 12768 37262
rect 12716 37198 12768 37204
rect 12346 37159 12402 37168
rect 12440 36780 12492 36786
rect 12440 36722 12492 36728
rect 12532 36780 12584 36786
rect 12532 36722 12584 36728
rect 12164 36576 12216 36582
rect 12164 36518 12216 36524
rect 12452 36378 12480 36722
rect 12440 36372 12492 36378
rect 12440 36314 12492 36320
rect 12256 36100 12308 36106
rect 12256 36042 12308 36048
rect 11796 36032 11848 36038
rect 11796 35974 11848 35980
rect 11888 36032 11940 36038
rect 11888 35974 11940 35980
rect 10600 35828 10652 35834
rect 10600 35770 10652 35776
rect 10876 35828 10928 35834
rect 10876 35770 10928 35776
rect 11244 35828 11296 35834
rect 11244 35770 11296 35776
rect 11428 35828 11480 35834
rect 11428 35770 11480 35776
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10876 35488 10928 35494
rect 10876 35430 10928 35436
rect 10600 35080 10652 35086
rect 10600 35022 10652 35028
rect 10612 34746 10640 35022
rect 10600 34740 10652 34746
rect 10600 34682 10652 34688
rect 10888 33998 10916 35430
rect 10980 35290 11008 35566
rect 10968 35284 11020 35290
rect 10968 35226 11020 35232
rect 11256 35222 11284 35770
rect 11704 35760 11756 35766
rect 11532 35708 11704 35714
rect 11532 35702 11756 35708
rect 11428 35692 11480 35698
rect 11428 35634 11480 35640
rect 11532 35686 11744 35702
rect 11808 35698 11836 35974
rect 11796 35692 11848 35698
rect 11244 35216 11296 35222
rect 11244 35158 11296 35164
rect 11024 34844 11332 34853
rect 11024 34842 11030 34844
rect 11086 34842 11110 34844
rect 11166 34842 11190 34844
rect 11246 34842 11270 34844
rect 11326 34842 11332 34844
rect 11086 34790 11088 34842
rect 11268 34790 11270 34842
rect 11024 34788 11030 34790
rect 11086 34788 11110 34790
rect 11166 34788 11190 34790
rect 11246 34788 11270 34790
rect 11326 34788 11332 34790
rect 11024 34779 11332 34788
rect 11244 34672 11296 34678
rect 11244 34614 11296 34620
rect 10968 34604 11020 34610
rect 10968 34546 11020 34552
rect 10980 34202 11008 34546
rect 11256 34202 11284 34614
rect 11440 34610 11468 35634
rect 11532 35562 11560 35686
rect 11796 35634 11848 35640
rect 11520 35556 11572 35562
rect 11520 35498 11572 35504
rect 11520 35080 11572 35086
rect 11520 35022 11572 35028
rect 11336 34604 11388 34610
rect 11336 34546 11388 34552
rect 11428 34604 11480 34610
rect 11428 34546 11480 34552
rect 10968 34196 11020 34202
rect 10968 34138 11020 34144
rect 11244 34196 11296 34202
rect 11244 34138 11296 34144
rect 11348 34105 11376 34546
rect 11532 34542 11560 35022
rect 11900 34950 11928 35974
rect 12164 35828 12216 35834
rect 12164 35770 12216 35776
rect 12072 35692 12124 35698
rect 12072 35634 12124 35640
rect 11888 34944 11940 34950
rect 11888 34886 11940 34892
rect 11520 34536 11572 34542
rect 11520 34478 11572 34484
rect 11334 34096 11390 34105
rect 11334 34031 11390 34040
rect 10876 33992 10928 33998
rect 10876 33934 10928 33940
rect 11428 33856 11480 33862
rect 11428 33798 11480 33804
rect 11024 33756 11332 33765
rect 11024 33754 11030 33756
rect 11086 33754 11110 33756
rect 11166 33754 11190 33756
rect 11246 33754 11270 33756
rect 11326 33754 11332 33756
rect 11086 33702 11088 33754
rect 11268 33702 11270 33754
rect 11024 33700 11030 33702
rect 11086 33700 11110 33702
rect 11166 33700 11190 33702
rect 11246 33700 11270 33702
rect 11326 33700 11332 33702
rect 11024 33691 11332 33700
rect 11440 33522 11468 33798
rect 10692 33516 10744 33522
rect 10612 33476 10692 33504
rect 10508 32836 10560 32842
rect 10508 32778 10560 32784
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10416 31272 10468 31278
rect 10416 31214 10468 31220
rect 10324 30932 10376 30938
rect 10324 30874 10376 30880
rect 10322 30832 10378 30841
rect 10322 30767 10378 30776
rect 10232 30252 10284 30258
rect 10232 30194 10284 30200
rect 10232 29232 10284 29238
rect 10232 29174 10284 29180
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 10140 28960 10192 28966
rect 10140 28902 10192 28908
rect 10046 28112 10102 28121
rect 9956 28076 10008 28082
rect 10152 28082 10180 28902
rect 10046 28047 10102 28056
rect 10140 28076 10192 28082
rect 9956 28018 10008 28024
rect 10140 28018 10192 28024
rect 9968 27606 9996 28018
rect 10244 27962 10272 29174
rect 10152 27934 10272 27962
rect 10048 27872 10100 27878
rect 10048 27814 10100 27820
rect 9956 27600 10008 27606
rect 9956 27542 10008 27548
rect 9862 26480 9918 26489
rect 9862 26415 9918 26424
rect 9864 26308 9916 26314
rect 9864 26250 9916 26256
rect 9876 25362 9904 26250
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9968 25294 9996 27542
rect 10060 26586 10088 27814
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 10048 26036 10100 26042
rect 10048 25978 10100 25984
rect 10060 25945 10088 25978
rect 10046 25936 10102 25945
rect 10046 25871 10102 25880
rect 9956 25288 10008 25294
rect 9956 25230 10008 25236
rect 9968 25140 9996 25230
rect 9876 25112 9996 25140
rect 9876 22964 9904 25112
rect 9956 24336 10008 24342
rect 9956 24278 10008 24284
rect 9968 23066 9996 24278
rect 10060 24206 10088 25871
rect 10048 24200 10100 24206
rect 10046 24168 10048 24177
rect 10100 24168 10102 24177
rect 10046 24103 10102 24112
rect 9968 23038 10088 23066
rect 9876 22936 9996 22964
rect 9770 22536 9826 22545
rect 9770 22471 9826 22480
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9784 22166 9812 22374
rect 9864 22228 9916 22234
rect 9864 22170 9916 22176
rect 9772 22160 9824 22166
rect 9772 22102 9824 22108
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9784 21894 9812 21966
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9772 21480 9824 21486
rect 9772 21422 9824 21428
rect 9784 21146 9812 21422
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9692 20998 9812 21026
rect 9784 20942 9812 20998
rect 9588 20936 9640 20942
rect 9772 20936 9824 20942
rect 9678 20904 9734 20913
rect 9640 20884 9678 20890
rect 9588 20878 9678 20884
rect 9600 20862 9678 20878
rect 9772 20878 9824 20884
rect 9678 20839 9734 20848
rect 9772 20596 9824 20602
rect 9772 20538 9824 20544
rect 9680 20392 9732 20398
rect 9680 20334 9732 20340
rect 9345 20156 9653 20165
rect 9345 20154 9351 20156
rect 9407 20154 9431 20156
rect 9487 20154 9511 20156
rect 9567 20154 9591 20156
rect 9647 20154 9653 20156
rect 9407 20102 9409 20154
rect 9589 20102 9591 20154
rect 9345 20100 9351 20102
rect 9407 20100 9431 20102
rect 9487 20100 9511 20102
rect 9567 20100 9591 20102
rect 9647 20100 9653 20102
rect 9345 20091 9653 20100
rect 9588 19304 9640 19310
rect 9416 19281 9588 19292
rect 9402 19272 9588 19281
rect 9458 19264 9588 19272
rect 9588 19246 9640 19252
rect 9402 19207 9458 19216
rect 9345 19068 9653 19077
rect 9345 19066 9351 19068
rect 9407 19066 9431 19068
rect 9487 19066 9511 19068
rect 9567 19066 9591 19068
rect 9647 19066 9653 19068
rect 9407 19014 9409 19066
rect 9589 19014 9591 19066
rect 9345 19012 9351 19014
rect 9407 19012 9431 19014
rect 9487 19012 9511 19014
rect 9567 19012 9591 19014
rect 9647 19012 9653 19014
rect 9345 19003 9653 19012
rect 9692 18222 9720 20334
rect 9784 19417 9812 20538
rect 9876 20058 9904 22170
rect 9968 21162 9996 22936
rect 10060 21468 10088 23038
rect 10152 22098 10180 27934
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10244 27334 10272 27406
rect 10232 27328 10284 27334
rect 10232 27270 10284 27276
rect 10232 25968 10284 25974
rect 10232 25910 10284 25916
rect 10244 24138 10272 25910
rect 10232 24132 10284 24138
rect 10232 24074 10284 24080
rect 10244 23633 10272 24074
rect 10230 23624 10286 23633
rect 10230 23559 10286 23568
rect 10232 23520 10284 23526
rect 10232 23462 10284 23468
rect 10244 22438 10272 23462
rect 10336 23254 10364 30767
rect 10428 26042 10456 31214
rect 10520 29646 10548 31758
rect 10612 30734 10640 33476
rect 10692 33458 10744 33464
rect 11336 33516 11388 33522
rect 11336 33458 11388 33464
rect 11428 33516 11480 33522
rect 11428 33458 11480 33464
rect 11152 33040 11204 33046
rect 11152 32982 11204 32988
rect 10968 32904 11020 32910
rect 10966 32872 10968 32881
rect 11020 32872 11022 32881
rect 10784 32836 10836 32842
rect 11164 32842 11192 32982
rect 11242 32872 11298 32881
rect 10966 32807 11022 32816
rect 11152 32836 11204 32842
rect 10784 32778 10836 32784
rect 11242 32807 11298 32816
rect 11152 32778 11204 32784
rect 10692 32428 10744 32434
rect 10692 32370 10744 32376
rect 10704 32026 10732 32370
rect 10796 32026 10824 32778
rect 11256 32774 11284 32807
rect 11244 32768 11296 32774
rect 11348 32756 11376 33458
rect 11532 33454 11560 34478
rect 11796 33924 11848 33930
rect 11796 33866 11848 33872
rect 11612 33856 11664 33862
rect 11612 33798 11664 33804
rect 11624 33590 11652 33798
rect 11612 33584 11664 33590
rect 11612 33526 11664 33532
rect 11520 33448 11572 33454
rect 11520 33390 11572 33396
rect 11532 32978 11560 33390
rect 11520 32972 11572 32978
rect 11520 32914 11572 32920
rect 11348 32728 11468 32756
rect 11244 32710 11296 32716
rect 11024 32668 11332 32677
rect 11024 32666 11030 32668
rect 11086 32666 11110 32668
rect 11166 32666 11190 32668
rect 11246 32666 11270 32668
rect 11326 32666 11332 32668
rect 11086 32614 11088 32666
rect 11268 32614 11270 32666
rect 11024 32612 11030 32614
rect 11086 32612 11110 32614
rect 11166 32612 11190 32614
rect 11246 32612 11270 32614
rect 11326 32612 11332 32614
rect 11024 32603 11332 32612
rect 11440 32552 11468 32728
rect 11256 32524 11468 32552
rect 11152 32428 11204 32434
rect 11152 32370 11204 32376
rect 11060 32360 11112 32366
rect 10888 32320 11060 32348
rect 10692 32020 10744 32026
rect 10692 31962 10744 31968
rect 10784 32020 10836 32026
rect 10784 31962 10836 31968
rect 10784 31816 10836 31822
rect 10784 31758 10836 31764
rect 10796 31482 10824 31758
rect 10888 31754 10916 32320
rect 11060 32302 11112 32308
rect 11164 32298 11192 32370
rect 11152 32292 11204 32298
rect 11152 32234 11204 32240
rect 11256 31958 11284 32524
rect 11532 32366 11560 32914
rect 11520 32360 11572 32366
rect 11520 32302 11572 32308
rect 11808 31958 11836 33866
rect 11244 31952 11296 31958
rect 11244 31894 11296 31900
rect 11796 31952 11848 31958
rect 11796 31894 11848 31900
rect 11336 31816 11388 31822
rect 11704 31816 11756 31822
rect 11388 31764 11468 31770
rect 11336 31758 11468 31764
rect 11704 31758 11756 31764
rect 10876 31748 10928 31754
rect 11348 31742 11468 31758
rect 10876 31690 10928 31696
rect 11024 31580 11332 31589
rect 11024 31578 11030 31580
rect 11086 31578 11110 31580
rect 11166 31578 11190 31580
rect 11246 31578 11270 31580
rect 11326 31578 11332 31580
rect 11086 31526 11088 31578
rect 11268 31526 11270 31578
rect 11024 31524 11030 31526
rect 11086 31524 11110 31526
rect 11166 31524 11190 31526
rect 11246 31524 11270 31526
rect 11326 31524 11332 31526
rect 11024 31515 11332 31524
rect 10784 31476 10836 31482
rect 10784 31418 10836 31424
rect 10692 31340 10744 31346
rect 10692 31282 10744 31288
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10704 30394 10732 31282
rect 11440 31210 11468 31742
rect 11520 31272 11572 31278
rect 11520 31214 11572 31220
rect 11428 31204 11480 31210
rect 11428 31146 11480 31152
rect 11152 31136 11204 31142
rect 11152 31078 11204 31084
rect 11164 30938 11192 31078
rect 11152 30932 11204 30938
rect 11152 30874 11204 30880
rect 11024 30492 11332 30501
rect 11024 30490 11030 30492
rect 11086 30490 11110 30492
rect 11166 30490 11190 30492
rect 11246 30490 11270 30492
rect 11326 30490 11332 30492
rect 11086 30438 11088 30490
rect 11268 30438 11270 30490
rect 11024 30436 11030 30438
rect 11086 30436 11110 30438
rect 11166 30436 11190 30438
rect 11246 30436 11270 30438
rect 11326 30436 11332 30438
rect 11024 30427 11332 30436
rect 10692 30388 10744 30394
rect 10692 30330 10744 30336
rect 10692 30116 10744 30122
rect 10692 30058 10744 30064
rect 10508 29640 10560 29646
rect 10508 29582 10560 29588
rect 10520 29238 10548 29582
rect 10704 29510 10732 30058
rect 11428 29572 11480 29578
rect 11428 29514 11480 29520
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 11024 29404 11332 29413
rect 11024 29402 11030 29404
rect 11086 29402 11110 29404
rect 11166 29402 11190 29404
rect 11246 29402 11270 29404
rect 11326 29402 11332 29404
rect 11086 29350 11088 29402
rect 11268 29350 11270 29402
rect 11024 29348 11030 29350
rect 11086 29348 11110 29350
rect 11166 29348 11190 29350
rect 11246 29348 11270 29350
rect 11326 29348 11332 29350
rect 11024 29339 11332 29348
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 10784 29232 10836 29238
rect 10784 29174 10836 29180
rect 11058 29200 11114 29209
rect 10690 28520 10746 28529
rect 10690 28455 10746 28464
rect 10704 27878 10732 28455
rect 10796 28014 10824 29174
rect 11058 29135 11060 29144
rect 11112 29135 11114 29144
rect 11060 29106 11112 29112
rect 10876 28960 10928 28966
rect 10876 28902 10928 28908
rect 10888 28694 10916 28902
rect 10876 28688 10928 28694
rect 10876 28630 10928 28636
rect 11072 28404 11100 29106
rect 11336 29028 11388 29034
rect 11336 28970 11388 28976
rect 10888 28376 11100 28404
rect 11348 28404 11376 28970
rect 11440 28665 11468 29514
rect 11426 28656 11482 28665
rect 11426 28591 11482 28600
rect 11348 28376 11468 28404
rect 10784 28008 10836 28014
rect 10784 27950 10836 27956
rect 10692 27872 10744 27878
rect 10692 27814 10744 27820
rect 10784 27872 10836 27878
rect 10784 27814 10836 27820
rect 10690 27568 10746 27577
rect 10690 27503 10746 27512
rect 10600 27124 10652 27130
rect 10600 27066 10652 27072
rect 10508 26512 10560 26518
rect 10508 26454 10560 26460
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 10428 25158 10456 25978
rect 10416 25152 10468 25158
rect 10416 25094 10468 25100
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 10428 24410 10456 24754
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10416 23792 10468 23798
rect 10416 23734 10468 23740
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10232 22432 10284 22438
rect 10232 22374 10284 22380
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 10232 21888 10284 21894
rect 10232 21830 10284 21836
rect 10140 21480 10192 21486
rect 10060 21440 10140 21468
rect 10140 21422 10192 21428
rect 10048 21344 10100 21350
rect 10046 21312 10048 21321
rect 10140 21344 10192 21350
rect 10100 21312 10102 21321
rect 10140 21286 10192 21292
rect 10046 21247 10102 21256
rect 9968 21134 10088 21162
rect 9864 20052 9916 20058
rect 9864 19994 9916 20000
rect 9864 19712 9916 19718
rect 9864 19654 9916 19660
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 9770 19408 9826 19417
rect 9770 19343 9826 19352
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9784 18970 9812 19246
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9876 18834 9904 19654
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9876 18329 9904 18770
rect 9862 18320 9918 18329
rect 9862 18255 9918 18264
rect 9680 18216 9732 18222
rect 9680 18158 9732 18164
rect 9862 18184 9918 18193
rect 9345 17980 9653 17989
rect 9345 17978 9351 17980
rect 9407 17978 9431 17980
rect 9487 17978 9511 17980
rect 9567 17978 9591 17980
rect 9647 17978 9653 17980
rect 9407 17926 9409 17978
rect 9589 17926 9591 17978
rect 9345 17924 9351 17926
rect 9407 17924 9431 17926
rect 9487 17924 9511 17926
rect 9567 17924 9591 17926
rect 9647 17924 9653 17926
rect 9345 17915 9653 17924
rect 9692 17864 9720 18158
rect 9862 18119 9918 18128
rect 9600 17836 9720 17864
rect 9770 17912 9826 17921
rect 9770 17847 9826 17856
rect 9600 17270 9628 17836
rect 9680 17536 9732 17542
rect 9680 17478 9732 17484
rect 9692 17270 9720 17478
rect 9784 17338 9812 17847
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9588 17264 9640 17270
rect 9588 17206 9640 17212
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9345 16892 9653 16901
rect 9345 16890 9351 16892
rect 9407 16890 9431 16892
rect 9487 16890 9511 16892
rect 9567 16890 9591 16892
rect 9647 16890 9653 16892
rect 9407 16838 9409 16890
rect 9589 16838 9591 16890
rect 9345 16836 9351 16838
rect 9407 16836 9431 16838
rect 9487 16836 9511 16838
rect 9567 16836 9591 16838
rect 9647 16836 9653 16838
rect 9345 16827 9653 16836
rect 9692 16674 9720 16934
rect 9784 16794 9812 16934
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9496 16652 9548 16658
rect 9692 16646 9812 16674
rect 9496 16594 9548 16600
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9048 14482 9076 14962
rect 9036 14476 9088 14482
rect 9036 14418 9088 14424
rect 8956 13484 9134 13512
rect 8956 13394 8984 13484
rect 9106 13410 9134 13484
rect 8944 13388 8996 13394
rect 9106 13382 9168 13410
rect 8944 13330 8996 13336
rect 9034 13288 9090 13297
rect 8944 13252 8996 13258
rect 9034 13223 9090 13232
rect 8944 13194 8996 13200
rect 8852 12912 8904 12918
rect 8852 12854 8904 12860
rect 8864 12782 8892 12854
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8956 12646 8984 13194
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8864 11257 8892 12582
rect 8850 11248 8906 11257
rect 8850 11183 8906 11192
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 8864 10062 8892 11086
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8864 8634 8892 9998
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8864 6866 8892 8570
rect 8956 8090 8984 12582
rect 9048 11150 9076 13223
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9034 10976 9090 10985
rect 9034 10911 9090 10920
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8956 7478 8984 8026
rect 8944 7472 8996 7478
rect 8944 7414 8996 7420
rect 8852 6860 8904 6866
rect 8852 6802 8904 6808
rect 9048 6746 9076 10911
rect 9140 8090 9168 13382
rect 9232 12238 9260 16594
rect 9508 15892 9536 16594
rect 9588 16584 9640 16590
rect 9678 16552 9734 16561
rect 9640 16532 9678 16538
rect 9588 16526 9678 16532
rect 9600 16510 9678 16526
rect 9678 16487 9734 16496
rect 9692 15994 9720 16487
rect 9784 16114 9812 16646
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9692 15966 9812 15994
rect 9508 15864 9720 15892
rect 9345 15804 9653 15813
rect 9345 15802 9351 15804
rect 9407 15802 9431 15804
rect 9487 15802 9511 15804
rect 9567 15802 9591 15804
rect 9647 15802 9653 15804
rect 9407 15750 9409 15802
rect 9589 15750 9591 15802
rect 9345 15748 9351 15750
rect 9407 15748 9431 15750
rect 9487 15748 9511 15750
rect 9567 15748 9591 15750
rect 9647 15748 9653 15750
rect 9345 15739 9653 15748
rect 9692 15609 9720 15864
rect 9678 15600 9734 15609
rect 9678 15535 9734 15544
rect 9312 15360 9364 15366
rect 9312 15302 9364 15308
rect 9324 15026 9352 15302
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9680 14952 9732 14958
rect 9784 14940 9812 15966
rect 9876 15065 9904 18119
rect 9968 15638 9996 19654
rect 10060 17134 10088 21134
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10152 16590 10180 21286
rect 10244 20806 10272 21830
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10336 20618 10364 22986
rect 10244 20590 10364 20618
rect 10244 18970 10272 20590
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 10152 15910 10180 16526
rect 10244 16454 10272 18566
rect 10232 16448 10284 16454
rect 10232 16390 10284 16396
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 9956 15632 10008 15638
rect 9956 15574 10008 15580
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10048 15088 10100 15094
rect 9862 15056 9918 15065
rect 10048 15030 10100 15036
rect 9862 14991 9918 15000
rect 9784 14912 9996 14940
rect 9680 14894 9732 14900
rect 9345 14716 9653 14725
rect 9345 14714 9351 14716
rect 9407 14714 9431 14716
rect 9487 14714 9511 14716
rect 9567 14714 9591 14716
rect 9647 14714 9653 14716
rect 9407 14662 9409 14714
rect 9589 14662 9591 14714
rect 9345 14660 9351 14662
rect 9407 14660 9431 14662
rect 9487 14660 9511 14662
rect 9567 14660 9591 14662
rect 9647 14660 9653 14662
rect 9345 14651 9653 14660
rect 9692 14498 9720 14894
rect 9770 14784 9826 14793
rect 9770 14719 9826 14728
rect 9784 14550 9812 14719
rect 9508 14470 9720 14498
rect 9772 14544 9824 14550
rect 9772 14486 9824 14492
rect 9508 13870 9536 14470
rect 9692 14396 9720 14470
rect 9692 14368 9812 14396
rect 9678 14240 9734 14249
rect 9678 14175 9734 14184
rect 9692 14006 9720 14175
rect 9680 14000 9732 14006
rect 9680 13942 9732 13948
rect 9496 13864 9548 13870
rect 9496 13806 9548 13812
rect 9345 13628 9653 13637
rect 9345 13626 9351 13628
rect 9407 13626 9431 13628
rect 9487 13626 9511 13628
rect 9567 13626 9591 13628
rect 9647 13626 9653 13628
rect 9407 13574 9409 13626
rect 9589 13574 9591 13626
rect 9345 13572 9351 13574
rect 9407 13572 9431 13574
rect 9487 13572 9511 13574
rect 9567 13572 9591 13574
rect 9647 13572 9653 13574
rect 9345 13563 9653 13572
rect 9404 13524 9456 13530
rect 9404 13466 9456 13472
rect 9416 13433 9444 13466
rect 9402 13424 9458 13433
rect 9402 13359 9458 13368
rect 9680 12912 9732 12918
rect 9784 12900 9812 14368
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 9876 14074 9904 14282
rect 9864 14068 9916 14074
rect 9864 14010 9916 14016
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9876 13326 9904 13874
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9732 12872 9812 12900
rect 9680 12854 9732 12860
rect 9345 12540 9653 12549
rect 9345 12538 9351 12540
rect 9407 12538 9431 12540
rect 9487 12538 9511 12540
rect 9567 12538 9591 12540
rect 9647 12538 9653 12540
rect 9407 12486 9409 12538
rect 9589 12486 9591 12538
rect 9345 12484 9351 12486
rect 9407 12484 9431 12486
rect 9487 12484 9511 12486
rect 9567 12484 9591 12486
rect 9647 12484 9653 12486
rect 9345 12475 9653 12484
rect 9402 12336 9458 12345
rect 9692 12306 9720 12854
rect 9864 12708 9916 12714
rect 9864 12650 9916 12656
rect 9402 12271 9458 12280
rect 9680 12300 9732 12306
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9416 11642 9444 12271
rect 9680 12242 9732 12248
rect 9232 11614 9444 11642
rect 9232 10130 9260 11614
rect 9345 11452 9653 11461
rect 9345 11450 9351 11452
rect 9407 11450 9431 11452
rect 9487 11450 9511 11452
rect 9567 11450 9591 11452
rect 9647 11450 9653 11452
rect 9407 11398 9409 11450
rect 9589 11398 9591 11450
rect 9345 11396 9351 11398
rect 9407 11396 9431 11398
rect 9487 11396 9511 11398
rect 9567 11396 9591 11398
rect 9647 11396 9653 11398
rect 9345 11387 9653 11396
rect 9876 10690 9904 12650
rect 9968 12594 9996 14912
rect 10060 12714 10088 15030
rect 10152 13530 10180 15438
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10152 12986 10180 13262
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 9968 12566 10088 12594
rect 9680 10668 9732 10674
rect 9876 10662 9996 10690
rect 9680 10610 9732 10616
rect 9402 10568 9458 10577
rect 9402 10503 9458 10512
rect 9416 10470 9444 10503
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9345 10364 9653 10373
rect 9345 10362 9351 10364
rect 9407 10362 9431 10364
rect 9487 10362 9511 10364
rect 9567 10362 9591 10364
rect 9647 10362 9653 10364
rect 9407 10310 9409 10362
rect 9589 10310 9591 10362
rect 9345 10308 9351 10310
rect 9407 10308 9431 10310
rect 9487 10308 9511 10310
rect 9567 10308 9591 10310
rect 9647 10308 9653 10310
rect 9345 10299 9653 10308
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9220 10124 9272 10130
rect 9220 10066 9272 10072
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9508 9704 9536 10066
rect 9600 9926 9628 10134
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9692 9722 9720 10610
rect 9864 10600 9916 10606
rect 9784 10560 9864 10588
rect 9588 9716 9640 9722
rect 9508 9676 9588 9704
rect 9588 9658 9640 9664
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9220 9512 9272 9518
rect 9600 9489 9628 9658
rect 9220 9454 9272 9460
rect 9586 9480 9642 9489
rect 9232 8344 9260 9454
rect 9586 9415 9642 9424
rect 9345 9276 9653 9285
rect 9345 9274 9351 9276
rect 9407 9274 9431 9276
rect 9487 9274 9511 9276
rect 9567 9274 9591 9276
rect 9647 9274 9653 9276
rect 9407 9222 9409 9274
rect 9589 9222 9591 9274
rect 9345 9220 9351 9222
rect 9407 9220 9431 9222
rect 9487 9220 9511 9222
rect 9567 9220 9591 9222
rect 9647 9220 9653 9222
rect 9345 9211 9653 9220
rect 9230 8316 9260 8344
rect 9128 8084 9180 8090
rect 9230 8072 9258 8316
rect 9345 8188 9653 8197
rect 9345 8186 9351 8188
rect 9407 8186 9431 8188
rect 9487 8186 9511 8188
rect 9567 8186 9591 8188
rect 9647 8186 9653 8188
rect 9407 8134 9409 8186
rect 9589 8134 9591 8186
rect 9345 8132 9351 8134
rect 9407 8132 9431 8134
rect 9487 8132 9511 8134
rect 9567 8132 9591 8134
rect 9647 8132 9653 8134
rect 9345 8123 9653 8132
rect 9230 8044 9260 8072
rect 9128 8026 9180 8032
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 8956 6718 9076 6746
rect 8956 5710 8984 6718
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8760 5364 8812 5370
rect 8760 5306 8812 5312
rect 8956 5098 8984 5646
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 9048 4486 9076 6598
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 7666 3292 7974 3301
rect 7666 3290 7672 3292
rect 7728 3290 7752 3292
rect 7808 3290 7832 3292
rect 7888 3290 7912 3292
rect 7968 3290 7974 3292
rect 7728 3238 7730 3290
rect 7910 3238 7912 3290
rect 7666 3236 7672 3238
rect 7728 3236 7752 3238
rect 7808 3236 7832 3238
rect 7888 3236 7912 3238
rect 7968 3236 7974 3238
rect 7666 3227 7974 3236
rect 8666 2408 8722 2417
rect 8666 2343 8722 2352
rect 7666 2204 7974 2213
rect 7666 2202 7672 2204
rect 7728 2202 7752 2204
rect 7808 2202 7832 2204
rect 7888 2202 7912 2204
rect 7968 2202 7974 2204
rect 7728 2150 7730 2202
rect 7910 2150 7912 2202
rect 7666 2148 7672 2150
rect 7728 2148 7752 2150
rect 7808 2148 7832 2150
rect 7888 2148 7912 2150
rect 7968 2148 7974 2150
rect 7666 2139 7974 2148
rect 8680 2106 8708 2343
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7472 2100 7524 2106
rect 7472 2042 7524 2048
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 9048 2038 9076 4422
rect 9036 2032 9088 2038
rect 9036 1974 9088 1980
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 7104 1964 7156 1970
rect 7104 1906 7156 1912
rect 7840 1964 7892 1970
rect 7840 1906 7892 1912
rect 8576 1964 8628 1970
rect 8576 1906 8628 1912
rect 4160 1828 4212 1834
rect 4160 1770 4212 1776
rect 2629 1660 2937 1669
rect 2629 1658 2635 1660
rect 2691 1658 2715 1660
rect 2771 1658 2795 1660
rect 2851 1658 2875 1660
rect 2931 1658 2937 1660
rect 2691 1606 2693 1658
rect 2873 1606 2875 1658
rect 2629 1604 2635 1606
rect 2691 1604 2715 1606
rect 2771 1604 2795 1606
rect 2851 1604 2875 1606
rect 2931 1604 2937 1606
rect 2629 1595 2937 1604
rect 5987 1660 6295 1669
rect 5987 1658 5993 1660
rect 6049 1658 6073 1660
rect 6129 1658 6153 1660
rect 6209 1658 6233 1660
rect 6289 1658 6295 1660
rect 6049 1606 6051 1658
rect 6231 1606 6233 1658
rect 5987 1604 5993 1606
rect 6049 1604 6073 1606
rect 6129 1604 6153 1606
rect 6209 1604 6233 1606
rect 6289 1604 6295 1606
rect 5987 1595 6295 1604
rect 6472 1562 6500 1906
rect 7116 1562 7144 1906
rect 7852 1562 7880 1906
rect 8588 1562 8616 1906
rect 6460 1556 6512 1562
rect 6460 1498 6512 1504
rect 7104 1556 7156 1562
rect 7104 1498 7156 1504
rect 7840 1556 7892 1562
rect 7840 1498 7892 1504
rect 8576 1556 8628 1562
rect 8576 1498 8628 1504
rect 9140 1494 9168 7482
rect 9232 6254 9260 8044
rect 9588 8016 9640 8022
rect 9588 7958 9640 7964
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 9324 7585 9352 7890
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9508 7721 9536 7822
rect 9600 7732 9628 7958
rect 9692 7954 9720 9658
rect 9784 9518 9812 10560
rect 9864 10542 9916 10548
rect 9864 10056 9916 10062
rect 9968 10044 9996 10662
rect 9916 10016 9996 10044
rect 9864 9998 9916 10004
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9876 9450 9904 9862
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 9784 9042 9812 9318
rect 9876 9042 9904 9386
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9864 9036 9916 9042
rect 9864 8978 9916 8984
rect 9680 7948 9732 7954
rect 9680 7890 9732 7896
rect 9784 7886 9812 8978
rect 9876 8673 9904 8978
rect 9862 8664 9918 8673
rect 9862 8599 9918 8608
rect 9968 8294 9996 10016
rect 9956 8288 10008 8294
rect 9956 8230 10008 8236
rect 9968 8072 9996 8230
rect 9876 8044 9996 8072
rect 9876 7993 9904 8044
rect 9862 7984 9918 7993
rect 9862 7919 9918 7928
rect 9956 7948 10008 7954
rect 9772 7880 9824 7886
rect 9678 7848 9734 7857
rect 9734 7828 9772 7834
rect 9734 7822 9824 7828
rect 9734 7806 9812 7822
rect 9678 7783 9734 7792
rect 9494 7712 9550 7721
rect 9600 7704 9812 7732
rect 9494 7647 9550 7656
rect 9310 7576 9366 7585
rect 9310 7511 9366 7520
rect 9632 7474 9688 7483
rect 9508 7449 9632 7460
rect 9494 7440 9632 7449
rect 9312 7404 9364 7410
rect 9550 7432 9632 7440
rect 9784 7449 9812 7704
rect 9632 7409 9688 7418
rect 9770 7440 9826 7449
rect 9494 7375 9550 7384
rect 9770 7375 9826 7384
rect 9312 7346 9364 7352
rect 9324 7256 9352 7346
rect 9680 7336 9732 7342
rect 9678 7304 9680 7313
rect 9732 7304 9734 7313
rect 9588 7268 9640 7274
rect 9324 7228 9588 7256
rect 9678 7239 9734 7248
rect 9772 7268 9824 7274
rect 9588 7210 9640 7216
rect 9772 7210 9824 7216
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9345 7100 9653 7109
rect 9345 7098 9351 7100
rect 9407 7098 9431 7100
rect 9487 7098 9511 7100
rect 9567 7098 9591 7100
rect 9647 7098 9653 7100
rect 9407 7046 9409 7098
rect 9589 7046 9591 7098
rect 9345 7044 9351 7046
rect 9407 7044 9431 7046
rect 9487 7044 9511 7046
rect 9567 7044 9591 7046
rect 9647 7044 9653 7046
rect 9345 7035 9653 7044
rect 9310 6896 9366 6905
rect 9310 6831 9366 6840
rect 9588 6860 9640 6866
rect 9220 6248 9272 6254
rect 9220 6190 9272 6196
rect 9324 6100 9352 6831
rect 9588 6802 9640 6808
rect 9600 6202 9628 6802
rect 9692 6322 9720 7142
rect 9784 7041 9812 7210
rect 9770 7032 9826 7041
rect 9876 7002 9904 7919
rect 9956 7890 10008 7896
rect 9968 7274 9996 7890
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 10060 7206 10088 12566
rect 10244 12345 10272 15302
rect 10336 15162 10364 19382
rect 10428 17202 10456 23734
rect 10520 23118 10548 26454
rect 10612 26382 10640 27066
rect 10704 26450 10732 27503
rect 10692 26444 10744 26450
rect 10692 26386 10744 26392
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10612 23118 10640 26318
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 10508 23112 10560 23118
rect 10508 23054 10560 23060
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10612 22545 10640 23054
rect 10598 22536 10654 22545
rect 10598 22471 10654 22480
rect 10600 22432 10652 22438
rect 10600 22374 10652 22380
rect 10612 21536 10640 22374
rect 10704 21554 10732 25638
rect 10796 23798 10824 27814
rect 10888 26926 10916 28376
rect 11024 28316 11332 28325
rect 11024 28314 11030 28316
rect 11086 28314 11110 28316
rect 11166 28314 11190 28316
rect 11246 28314 11270 28316
rect 11326 28314 11332 28316
rect 11086 28262 11088 28314
rect 11268 28262 11270 28314
rect 11024 28260 11030 28262
rect 11086 28260 11110 28262
rect 11166 28260 11190 28262
rect 11246 28260 11270 28262
rect 11326 28260 11332 28262
rect 11024 28251 11332 28260
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 10980 27674 11008 28018
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 11024 27228 11332 27237
rect 11024 27226 11030 27228
rect 11086 27226 11110 27228
rect 11166 27226 11190 27228
rect 11246 27226 11270 27228
rect 11326 27226 11332 27228
rect 11086 27174 11088 27226
rect 11268 27174 11270 27226
rect 11024 27172 11030 27174
rect 11086 27172 11110 27174
rect 11166 27172 11190 27174
rect 11246 27172 11270 27174
rect 11326 27172 11332 27174
rect 11024 27163 11332 27172
rect 10876 26920 10928 26926
rect 10876 26862 10928 26868
rect 10876 26784 10928 26790
rect 10876 26726 10928 26732
rect 10888 26586 10916 26726
rect 10876 26580 10928 26586
rect 10876 26522 10928 26528
rect 10876 26444 10928 26450
rect 10876 26386 10928 26392
rect 10784 23792 10836 23798
rect 10784 23734 10836 23740
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 10796 22778 10824 23190
rect 10888 23186 10916 26386
rect 11024 26140 11332 26149
rect 11024 26138 11030 26140
rect 11086 26138 11110 26140
rect 11166 26138 11190 26140
rect 11246 26138 11270 26140
rect 11326 26138 11332 26140
rect 11086 26086 11088 26138
rect 11268 26086 11270 26138
rect 11024 26084 11030 26086
rect 11086 26084 11110 26086
rect 11166 26084 11190 26086
rect 11246 26084 11270 26086
rect 11326 26084 11332 26086
rect 11024 26075 11332 26084
rect 11152 25764 11204 25770
rect 11152 25706 11204 25712
rect 11164 25362 11192 25706
rect 11440 25498 11468 28376
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 11426 25392 11482 25401
rect 10968 25356 11020 25362
rect 10968 25298 11020 25304
rect 11152 25356 11204 25362
rect 11426 25327 11482 25336
rect 11152 25298 11204 25304
rect 10980 25265 11008 25298
rect 10966 25256 11022 25265
rect 11440 25226 11468 25327
rect 10966 25191 11022 25200
rect 11428 25220 11480 25226
rect 11428 25162 11480 25168
rect 11024 25052 11332 25061
rect 11024 25050 11030 25052
rect 11086 25050 11110 25052
rect 11166 25050 11190 25052
rect 11246 25050 11270 25052
rect 11326 25050 11332 25052
rect 11086 24998 11088 25050
rect 11268 24998 11270 25050
rect 11024 24996 11030 24998
rect 11086 24996 11110 24998
rect 11166 24996 11190 24998
rect 11246 24996 11270 24998
rect 11326 24996 11332 24998
rect 11024 24987 11332 24996
rect 10968 24812 11020 24818
rect 10968 24754 11020 24760
rect 10980 24138 11008 24754
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11440 24177 11468 24550
rect 11426 24168 11482 24177
rect 10968 24132 11020 24138
rect 11426 24103 11482 24112
rect 10968 24074 11020 24080
rect 11024 23964 11332 23973
rect 11024 23962 11030 23964
rect 11086 23962 11110 23964
rect 11166 23962 11190 23964
rect 11246 23962 11270 23964
rect 11326 23962 11332 23964
rect 11086 23910 11088 23962
rect 11268 23910 11270 23962
rect 11024 23908 11030 23910
rect 11086 23908 11110 23910
rect 11166 23908 11190 23910
rect 11246 23908 11270 23910
rect 11326 23908 11332 23910
rect 11024 23899 11332 23908
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 11072 23254 11100 23462
rect 11060 23248 11112 23254
rect 11060 23190 11112 23196
rect 10876 23180 10928 23186
rect 10876 23122 10928 23128
rect 11024 22876 11332 22885
rect 11024 22874 11030 22876
rect 11086 22874 11110 22876
rect 11166 22874 11190 22876
rect 11246 22874 11270 22876
rect 11326 22874 11332 22876
rect 11086 22822 11088 22874
rect 11268 22822 11270 22874
rect 11024 22820 11030 22822
rect 11086 22820 11110 22822
rect 11166 22820 11190 22822
rect 11246 22820 11270 22822
rect 11326 22820 11332 22822
rect 11024 22811 11332 22820
rect 10784 22772 10836 22778
rect 10784 22714 10836 22720
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 10968 22024 11020 22030
rect 10968 21966 11020 21972
rect 10796 21894 10824 21966
rect 10784 21888 10836 21894
rect 10980 21876 11008 21966
rect 10784 21830 10836 21836
rect 10888 21848 11008 21876
rect 10520 21508 10640 21536
rect 10692 21548 10744 21554
rect 10520 18630 10548 21508
rect 10692 21490 10744 21496
rect 10796 21434 10824 21830
rect 10612 21406 10824 21434
rect 10612 21350 10640 21406
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10692 21344 10744 21350
rect 10692 21286 10744 21292
rect 10704 19854 10732 21286
rect 10888 21146 10916 21848
rect 11024 21788 11332 21797
rect 11024 21786 11030 21788
rect 11086 21786 11110 21788
rect 11166 21786 11190 21788
rect 11246 21786 11270 21788
rect 11326 21786 11332 21788
rect 11086 21734 11088 21786
rect 11268 21734 11270 21786
rect 11024 21732 11030 21734
rect 11086 21732 11110 21734
rect 11166 21732 11190 21734
rect 11246 21732 11270 21734
rect 11326 21732 11332 21734
rect 11024 21723 11332 21732
rect 11060 21480 11112 21486
rect 10980 21440 11060 21468
rect 10876 21140 10928 21146
rect 10876 21082 10928 21088
rect 10980 21026 11008 21440
rect 11060 21422 11112 21428
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11256 21078 11284 21422
rect 10888 20998 11008 21026
rect 11244 21072 11296 21078
rect 11244 21014 11296 21020
rect 10888 20806 10916 20998
rect 10876 20800 10928 20806
rect 10876 20742 10928 20748
rect 10692 19848 10744 19854
rect 10692 19790 10744 19796
rect 10888 19666 10916 20742
rect 11024 20700 11332 20709
rect 11024 20698 11030 20700
rect 11086 20698 11110 20700
rect 11166 20698 11190 20700
rect 11246 20698 11270 20700
rect 11326 20698 11332 20700
rect 11086 20646 11088 20698
rect 11268 20646 11270 20698
rect 11024 20644 11030 20646
rect 11086 20644 11110 20646
rect 11166 20644 11190 20646
rect 11246 20644 11270 20646
rect 11326 20644 11332 20646
rect 11024 20635 11332 20644
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 10980 19854 11008 20266
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 11348 19786 11468 19802
rect 11336 19780 11468 19786
rect 11388 19774 11468 19780
rect 11336 19722 11388 19728
rect 10612 19638 10916 19666
rect 10508 18624 10560 18630
rect 10508 18566 10560 18572
rect 10506 17776 10562 17785
rect 10506 17711 10562 17720
rect 10520 17202 10548 17711
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10612 16658 10640 19638
rect 11024 19612 11332 19621
rect 11024 19610 11030 19612
rect 11086 19610 11110 19612
rect 11166 19610 11190 19612
rect 11246 19610 11270 19612
rect 11326 19610 11332 19612
rect 11086 19558 11088 19610
rect 11268 19558 11270 19610
rect 11024 19556 11030 19558
rect 11086 19556 11110 19558
rect 11166 19556 11190 19558
rect 11246 19556 11270 19558
rect 11326 19556 11332 19558
rect 11024 19547 11332 19556
rect 11242 19408 11298 19417
rect 11242 19343 11298 19352
rect 11256 19310 11284 19343
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 10690 18864 10746 18873
rect 10690 18799 10746 18808
rect 10704 18290 10732 18799
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10796 18170 10824 19246
rect 11024 18524 11332 18533
rect 11024 18522 11030 18524
rect 11086 18522 11110 18524
rect 11166 18522 11190 18524
rect 11246 18522 11270 18524
rect 11326 18522 11332 18524
rect 11086 18470 11088 18522
rect 11268 18470 11270 18522
rect 11024 18468 11030 18470
rect 11086 18468 11110 18470
rect 11166 18468 11190 18470
rect 11246 18468 11270 18470
rect 11326 18468 11332 18470
rect 11024 18459 11332 18468
rect 10704 18142 10824 18170
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10428 16250 10456 16526
rect 10416 16244 10468 16250
rect 10416 16186 10468 16192
rect 10416 16108 10468 16114
rect 10416 16050 10468 16056
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10336 14793 10364 14962
rect 10322 14784 10378 14793
rect 10322 14719 10378 14728
rect 10322 14648 10378 14657
rect 10322 14583 10378 14592
rect 10336 14482 10364 14583
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10230 12336 10286 12345
rect 10230 12271 10286 12280
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10152 11898 10180 12106
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10336 11200 10364 13466
rect 10428 12850 10456 16050
rect 10508 14612 10560 14618
rect 10560 14572 10640 14600
rect 10508 14554 10560 14560
rect 10612 14521 10640 14572
rect 10598 14512 10654 14521
rect 10598 14447 10654 14456
rect 10508 14408 10560 14414
rect 10560 14356 10640 14362
rect 10508 14350 10640 14356
rect 10520 14334 10640 14350
rect 10416 12844 10468 12850
rect 10416 12786 10468 12792
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10520 11354 10548 12242
rect 10508 11348 10560 11354
rect 10508 11290 10560 11296
rect 10244 11172 10364 11200
rect 10244 10248 10272 11172
rect 10508 11144 10560 11150
rect 10322 11112 10378 11121
rect 10508 11086 10560 11092
rect 10322 11047 10378 11056
rect 10336 10810 10364 11047
rect 10324 10804 10376 10810
rect 10324 10746 10376 10752
rect 10520 10266 10548 11086
rect 10612 10810 10640 14334
rect 10704 13938 10732 18142
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 10796 17542 10824 18022
rect 11164 17814 11192 18022
rect 11152 17808 11204 17814
rect 11152 17750 11204 17756
rect 11440 17678 11468 19774
rect 11532 19530 11560 31214
rect 11612 31136 11664 31142
rect 11612 31078 11664 31084
rect 11624 29209 11652 31078
rect 11716 30326 11744 31758
rect 11796 31748 11848 31754
rect 11900 31736 11928 34886
rect 12084 33969 12112 35634
rect 12070 33960 12126 33969
rect 12070 33895 12126 33904
rect 12176 33522 12204 35770
rect 12268 35630 12296 36042
rect 12544 35850 12572 36722
rect 12636 36258 12664 37198
rect 12728 36961 12756 37198
rect 12714 36952 12770 36961
rect 12714 36887 12770 36896
rect 12820 36650 12848 37318
rect 13360 37188 13412 37194
rect 13360 37130 13412 37136
rect 13544 37188 13596 37194
rect 13544 37130 13596 37136
rect 13372 37097 13400 37130
rect 13358 37088 13414 37097
rect 13358 37023 13414 37032
rect 13556 36922 13584 37130
rect 13636 37120 13688 37126
rect 13636 37062 13688 37068
rect 13544 36916 13596 36922
rect 13544 36858 13596 36864
rect 12808 36644 12860 36650
rect 12808 36586 12860 36592
rect 13544 36576 13596 36582
rect 13648 36553 13676 37062
rect 13740 36825 13768 37606
rect 13726 36816 13782 36825
rect 13726 36751 13782 36760
rect 13544 36518 13596 36524
rect 13634 36544 13690 36553
rect 12703 36476 13011 36485
rect 12703 36474 12709 36476
rect 12765 36474 12789 36476
rect 12845 36474 12869 36476
rect 12925 36474 12949 36476
rect 13005 36474 13011 36476
rect 12765 36422 12767 36474
rect 12947 36422 12949 36474
rect 12703 36420 12709 36422
rect 12765 36420 12789 36422
rect 12845 36420 12869 36422
rect 12925 36420 12949 36422
rect 13005 36420 13011 36422
rect 12703 36411 13011 36420
rect 12636 36230 12756 36258
rect 12624 36100 12676 36106
rect 12624 36042 12676 36048
rect 12452 35822 12572 35850
rect 12348 35760 12400 35766
rect 12348 35702 12400 35708
rect 12256 35624 12308 35630
rect 12256 35566 12308 35572
rect 12360 34202 12388 35702
rect 12452 35698 12480 35822
rect 12636 35737 12664 36042
rect 12622 35728 12678 35737
rect 12440 35692 12492 35698
rect 12440 35634 12492 35640
rect 12532 35692 12584 35698
rect 12622 35663 12678 35672
rect 12532 35634 12584 35640
rect 12440 34944 12492 34950
rect 12440 34886 12492 34892
rect 12348 34196 12400 34202
rect 12348 34138 12400 34144
rect 12452 33946 12480 34886
rect 12544 34134 12572 35634
rect 12728 35601 12756 36230
rect 13176 36100 13228 36106
rect 13176 36042 13228 36048
rect 13360 36100 13412 36106
rect 13360 36042 13412 36048
rect 12714 35592 12770 35601
rect 12714 35527 12770 35536
rect 13188 35465 13216 36042
rect 13268 35488 13320 35494
rect 13174 35456 13230 35465
rect 13268 35430 13320 35436
rect 12703 35388 13011 35397
rect 13174 35391 13230 35400
rect 12703 35386 12709 35388
rect 12765 35386 12789 35388
rect 12845 35386 12869 35388
rect 12925 35386 12949 35388
rect 13005 35386 13011 35388
rect 12765 35334 12767 35386
rect 12947 35334 12949 35386
rect 12703 35332 12709 35334
rect 12765 35332 12789 35334
rect 12845 35332 12869 35334
rect 12925 35332 12949 35334
rect 13005 35332 13011 35334
rect 12703 35323 13011 35332
rect 13084 35080 13136 35086
rect 13084 35022 13136 35028
rect 12624 34944 12676 34950
rect 12624 34886 12676 34892
rect 12532 34128 12584 34134
rect 12532 34070 12584 34076
rect 12636 34066 12664 34886
rect 12992 34740 13044 34746
rect 12992 34682 13044 34688
rect 13004 34490 13032 34682
rect 13096 34649 13124 35022
rect 13176 35012 13228 35018
rect 13176 34954 13228 34960
rect 13082 34640 13138 34649
rect 13082 34575 13138 34584
rect 13004 34462 13124 34490
rect 12703 34300 13011 34309
rect 12703 34298 12709 34300
rect 12765 34298 12789 34300
rect 12845 34298 12869 34300
rect 12925 34298 12949 34300
rect 13005 34298 13011 34300
rect 12765 34246 12767 34298
rect 12947 34246 12949 34298
rect 12703 34244 12709 34246
rect 12765 34244 12789 34246
rect 12845 34244 12869 34246
rect 12925 34244 12949 34246
rect 13005 34244 13011 34246
rect 12703 34235 13011 34244
rect 12624 34060 12676 34066
rect 12624 34002 12676 34008
rect 12256 33924 12308 33930
rect 12452 33918 12664 33946
rect 12256 33866 12308 33872
rect 12164 33516 12216 33522
rect 12164 33458 12216 33464
rect 11980 33312 12032 33318
rect 11980 33254 12032 33260
rect 11992 32026 12020 33254
rect 11980 32020 12032 32026
rect 11980 31962 12032 31968
rect 12072 31884 12124 31890
rect 12072 31826 12124 31832
rect 11900 31708 12020 31736
rect 11796 31690 11848 31696
rect 11808 30977 11836 31690
rect 11888 31272 11940 31278
rect 11888 31214 11940 31220
rect 11794 30968 11850 30977
rect 11794 30903 11850 30912
rect 11900 30734 11928 31214
rect 11796 30728 11848 30734
rect 11794 30696 11796 30705
rect 11888 30728 11940 30734
rect 11848 30696 11850 30705
rect 11888 30670 11940 30676
rect 11794 30631 11850 30640
rect 11900 30433 11928 30670
rect 11886 30424 11942 30433
rect 11886 30359 11942 30368
rect 11704 30320 11756 30326
rect 11992 30308 12020 31708
rect 11704 30262 11756 30268
rect 11900 30280 12020 30308
rect 11796 29708 11848 29714
rect 11796 29650 11848 29656
rect 11704 29572 11756 29578
rect 11704 29514 11756 29520
rect 11610 29200 11666 29209
rect 11610 29135 11666 29144
rect 11612 29096 11664 29102
rect 11612 29038 11664 29044
rect 11624 28540 11652 29038
rect 11716 29034 11744 29514
rect 11808 29102 11836 29650
rect 11900 29306 11928 30280
rect 11980 30184 12032 30190
rect 11980 30126 12032 30132
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11796 29096 11848 29102
rect 11796 29038 11848 29044
rect 11704 29028 11756 29034
rect 11704 28970 11756 28976
rect 11992 28801 12020 30126
rect 12084 29850 12112 31826
rect 12176 30716 12204 33458
rect 12268 32337 12296 33866
rect 12532 33856 12584 33862
rect 12532 33798 12584 33804
rect 12544 33402 12572 33798
rect 12452 33374 12572 33402
rect 12452 33046 12480 33374
rect 12532 33312 12584 33318
rect 12532 33254 12584 33260
rect 12440 33040 12492 33046
rect 12346 33008 12402 33017
rect 12440 32982 12492 32988
rect 12346 32943 12402 32952
rect 12360 32434 12388 32943
rect 12544 32824 12572 33254
rect 12452 32796 12572 32824
rect 12348 32428 12400 32434
rect 12348 32370 12400 32376
rect 12254 32328 12310 32337
rect 12254 32263 12310 32272
rect 12256 32224 12308 32230
rect 12256 32166 12308 32172
rect 12268 32026 12296 32166
rect 12256 32020 12308 32026
rect 12256 31962 12308 31968
rect 12256 31816 12308 31822
rect 12256 31758 12308 31764
rect 12268 30841 12296 31758
rect 12452 31498 12480 32796
rect 12532 32224 12584 32230
rect 12532 32166 12584 32172
rect 12360 31470 12480 31498
rect 12360 31278 12388 31470
rect 12544 31396 12572 32166
rect 12636 31754 12664 33918
rect 12703 33212 13011 33221
rect 12703 33210 12709 33212
rect 12765 33210 12789 33212
rect 12845 33210 12869 33212
rect 12925 33210 12949 33212
rect 13005 33210 13011 33212
rect 12765 33158 12767 33210
rect 12947 33158 12949 33210
rect 12703 33156 12709 33158
rect 12765 33156 12789 33158
rect 12845 33156 12869 33158
rect 12925 33156 12949 33158
rect 13005 33156 13011 33158
rect 12703 33147 13011 33156
rect 12900 33040 12952 33046
rect 12900 32982 12952 32988
rect 12808 32768 12860 32774
rect 12808 32710 12860 32716
rect 12820 32212 12848 32710
rect 12912 32473 12940 32982
rect 13096 32858 13124 34462
rect 13188 33658 13216 34954
rect 13280 34241 13308 35430
rect 13372 35290 13400 36042
rect 13452 35488 13504 35494
rect 13452 35430 13504 35436
rect 13360 35284 13412 35290
rect 13360 35226 13412 35232
rect 13360 34400 13412 34406
rect 13464 34377 13492 35430
rect 13556 34649 13584 36518
rect 13634 36479 13690 36488
rect 14016 36122 14044 41482
rect 14382 41372 14690 41381
rect 14382 41370 14388 41372
rect 14444 41370 14468 41372
rect 14524 41370 14548 41372
rect 14604 41370 14628 41372
rect 14684 41370 14690 41372
rect 14444 41318 14446 41370
rect 14626 41318 14628 41370
rect 14382 41316 14388 41318
rect 14444 41316 14468 41318
rect 14524 41316 14548 41318
rect 14604 41316 14628 41318
rect 14684 41316 14690 41318
rect 14382 41307 14690 41316
rect 14382 40284 14690 40293
rect 14382 40282 14388 40284
rect 14444 40282 14468 40284
rect 14524 40282 14548 40284
rect 14604 40282 14628 40284
rect 14684 40282 14690 40284
rect 14444 40230 14446 40282
rect 14626 40230 14628 40282
rect 14382 40228 14388 40230
rect 14444 40228 14468 40230
rect 14524 40228 14548 40230
rect 14604 40228 14628 40230
rect 14684 40228 14690 40230
rect 14382 40219 14690 40228
rect 14096 39840 14148 39846
rect 14096 39782 14148 39788
rect 14108 39545 14136 39782
rect 14094 39536 14150 39545
rect 14094 39471 14150 39480
rect 14280 39296 14332 39302
rect 14280 39238 14332 39244
rect 14292 39001 14320 39238
rect 14382 39196 14690 39205
rect 14382 39194 14388 39196
rect 14444 39194 14468 39196
rect 14524 39194 14548 39196
rect 14604 39194 14628 39196
rect 14684 39194 14690 39196
rect 14444 39142 14446 39194
rect 14626 39142 14628 39194
rect 14382 39140 14388 39142
rect 14444 39140 14468 39142
rect 14524 39140 14548 39142
rect 14604 39140 14628 39142
rect 14684 39140 14690 39142
rect 14382 39131 14690 39140
rect 14278 38992 14334 39001
rect 14278 38927 14334 38936
rect 14280 38208 14332 38214
rect 14280 38150 14332 38156
rect 14292 37913 14320 38150
rect 14382 38108 14690 38117
rect 14382 38106 14388 38108
rect 14444 38106 14468 38108
rect 14524 38106 14548 38108
rect 14604 38106 14628 38108
rect 14684 38106 14690 38108
rect 14444 38054 14446 38106
rect 14626 38054 14628 38106
rect 14382 38052 14388 38054
rect 14444 38052 14468 38054
rect 14524 38052 14548 38054
rect 14604 38052 14628 38054
rect 14684 38052 14690 38054
rect 14382 38043 14690 38052
rect 14278 37904 14334 37913
rect 14278 37839 14334 37848
rect 14372 37800 14424 37806
rect 14372 37742 14424 37748
rect 14188 37732 14240 37738
rect 14188 37674 14240 37680
rect 14200 37369 14228 37674
rect 14384 37641 14412 37742
rect 14370 37632 14426 37641
rect 14370 37567 14426 37576
rect 14186 37360 14242 37369
rect 14186 37295 14242 37304
rect 14382 37020 14690 37029
rect 14382 37018 14388 37020
rect 14444 37018 14468 37020
rect 14524 37018 14548 37020
rect 14604 37018 14628 37020
rect 14684 37018 14690 37020
rect 14444 36966 14446 37018
rect 14626 36966 14628 37018
rect 14382 36964 14388 36966
rect 14444 36964 14468 36966
rect 14524 36964 14548 36966
rect 14604 36964 14628 36966
rect 14684 36964 14690 36966
rect 14382 36955 14690 36964
rect 14188 36644 14240 36650
rect 14188 36586 14240 36592
rect 14200 36281 14228 36586
rect 14752 36530 14780 41550
rect 15488 41414 15516 42026
rect 15304 41386 15516 41414
rect 14832 39364 14884 39370
rect 14832 39306 14884 39312
rect 14844 39273 14872 39306
rect 14830 39264 14886 39273
rect 14830 39199 14886 39208
rect 14832 38276 14884 38282
rect 14832 38218 14884 38224
rect 14844 38185 14872 38218
rect 14830 38176 14886 38185
rect 14830 38111 14886 38120
rect 15016 36780 15068 36786
rect 15016 36722 15068 36728
rect 14752 36502 14872 36530
rect 14186 36272 14242 36281
rect 14186 36207 14242 36216
rect 13728 36100 13780 36106
rect 14016 36094 14780 36122
rect 13728 36042 13780 36048
rect 13740 35057 13768 36042
rect 14382 35932 14690 35941
rect 14382 35930 14388 35932
rect 14444 35930 14468 35932
rect 14524 35930 14548 35932
rect 14604 35930 14628 35932
rect 14684 35930 14690 35932
rect 14444 35878 14446 35930
rect 14626 35878 14628 35930
rect 14382 35876 14388 35878
rect 14444 35876 14468 35878
rect 14524 35876 14548 35878
rect 14604 35876 14628 35878
rect 14684 35876 14690 35878
rect 14382 35867 14690 35876
rect 13820 35692 13872 35698
rect 13820 35634 13872 35640
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 13726 35048 13782 35057
rect 13726 34983 13782 34992
rect 13636 34944 13688 34950
rect 13636 34886 13688 34892
rect 13542 34640 13598 34649
rect 13542 34575 13598 34584
rect 13544 34536 13596 34542
rect 13544 34478 13596 34484
rect 13360 34342 13412 34348
rect 13450 34368 13506 34377
rect 13266 34232 13322 34241
rect 13266 34167 13322 34176
rect 13268 33924 13320 33930
rect 13268 33866 13320 33872
rect 13176 33652 13228 33658
rect 13176 33594 13228 33600
rect 13176 33516 13228 33522
rect 13176 33458 13228 33464
rect 13004 32830 13124 32858
rect 12898 32464 12954 32473
rect 13004 32450 13032 32830
rect 13188 32570 13216 33458
rect 13176 32564 13228 32570
rect 13176 32506 13228 32512
rect 13280 32502 13308 33866
rect 13372 33153 13400 34342
rect 13450 34303 13506 34312
rect 13556 34082 13584 34478
rect 13464 34054 13584 34082
rect 13358 33144 13414 33153
rect 13464 33130 13492 34054
rect 13544 33924 13596 33930
rect 13544 33866 13596 33872
rect 13556 33386 13584 33866
rect 13648 33561 13676 34886
rect 13832 34746 13860 35634
rect 14004 35556 14056 35562
rect 14004 35498 14056 35504
rect 14016 35193 14044 35498
rect 14002 35184 14058 35193
rect 14002 35119 14058 35128
rect 13820 34740 13872 34746
rect 13820 34682 13872 34688
rect 13820 34604 13872 34610
rect 13820 34546 13872 34552
rect 13726 34232 13782 34241
rect 13726 34167 13782 34176
rect 13740 33969 13768 34167
rect 13726 33960 13782 33969
rect 13726 33895 13782 33904
rect 13728 33856 13780 33862
rect 13728 33798 13780 33804
rect 13740 33658 13768 33798
rect 13728 33652 13780 33658
rect 13728 33594 13780 33600
rect 13634 33552 13690 33561
rect 13634 33487 13690 33496
rect 13728 33516 13780 33522
rect 13728 33458 13780 33464
rect 13636 33448 13688 33454
rect 13636 33390 13688 33396
rect 13544 33380 13596 33386
rect 13544 33322 13596 33328
rect 13464 33114 13584 33130
rect 13464 33108 13596 33114
rect 13464 33102 13544 33108
rect 13358 33079 13414 33088
rect 13544 33050 13596 33056
rect 13544 32972 13596 32978
rect 13544 32914 13596 32920
rect 13450 32872 13506 32881
rect 13360 32836 13412 32842
rect 13450 32807 13506 32816
rect 13360 32778 13412 32784
rect 13268 32496 13320 32502
rect 13004 32422 13216 32450
rect 13268 32438 13320 32444
rect 12898 32399 12954 32408
rect 12820 32184 13124 32212
rect 12703 32124 13011 32133
rect 12703 32122 12709 32124
rect 12765 32122 12789 32124
rect 12845 32122 12869 32124
rect 12925 32122 12949 32124
rect 13005 32122 13011 32124
rect 12765 32070 12767 32122
rect 12947 32070 12949 32122
rect 12703 32068 12709 32070
rect 12765 32068 12789 32070
rect 12845 32068 12869 32070
rect 12925 32068 12949 32070
rect 13005 32068 13011 32070
rect 12703 32059 13011 32068
rect 12636 31726 12940 31754
rect 12716 31476 12768 31482
rect 12716 31418 12768 31424
rect 12452 31368 12572 31396
rect 12348 31272 12400 31278
rect 12348 31214 12400 31220
rect 12452 30870 12480 31368
rect 12624 31272 12676 31278
rect 12624 31214 12676 31220
rect 12530 30968 12586 30977
rect 12530 30903 12586 30912
rect 12440 30864 12492 30870
rect 12254 30832 12310 30841
rect 12440 30806 12492 30812
rect 12254 30767 12310 30776
rect 12176 30688 12388 30716
rect 12256 30592 12308 30598
rect 12256 30534 12308 30540
rect 12268 30190 12296 30534
rect 12164 30184 12216 30190
rect 12164 30126 12216 30132
rect 12256 30184 12308 30190
rect 12256 30126 12308 30132
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 12072 29504 12124 29510
rect 12072 29446 12124 29452
rect 11978 28792 12034 28801
rect 11978 28727 12034 28736
rect 11808 28626 12020 28642
rect 11796 28620 12020 28626
rect 11848 28614 12020 28620
rect 11796 28562 11848 28568
rect 11888 28552 11940 28558
rect 11624 28512 11744 28540
rect 11612 27872 11664 27878
rect 11612 27814 11664 27820
rect 11624 26897 11652 27814
rect 11716 27674 11744 28512
rect 11882 28506 11888 28540
rect 11826 28500 11888 28506
rect 11826 28494 11940 28500
rect 11826 28478 11910 28494
rect 11826 28472 11854 28478
rect 11808 28444 11854 28472
rect 11704 27668 11756 27674
rect 11704 27610 11756 27616
rect 11704 27328 11756 27334
rect 11704 27270 11756 27276
rect 11610 26888 11666 26897
rect 11610 26823 11666 26832
rect 11610 26752 11666 26761
rect 11610 26687 11666 26696
rect 11624 26194 11652 26687
rect 11716 26382 11744 27270
rect 11808 27130 11836 28444
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11900 28218 11928 28358
rect 11888 28212 11940 28218
rect 11888 28154 11940 28160
rect 11992 28082 12020 28614
rect 12084 28558 12112 29446
rect 12072 28552 12124 28558
rect 12072 28494 12124 28500
rect 11980 28076 12032 28082
rect 11980 28018 12032 28024
rect 12072 27872 12124 27878
rect 11978 27840 12034 27849
rect 12072 27814 12124 27820
rect 11978 27775 12034 27784
rect 11888 27464 11940 27470
rect 11886 27432 11888 27441
rect 11940 27432 11942 27441
rect 11886 27367 11942 27376
rect 11796 27124 11848 27130
rect 11796 27066 11848 27072
rect 11796 26920 11848 26926
rect 11796 26862 11848 26868
rect 11704 26376 11756 26382
rect 11704 26318 11756 26324
rect 11624 26166 11744 26194
rect 11612 25900 11664 25906
rect 11612 25842 11664 25848
rect 11624 25498 11652 25842
rect 11612 25492 11664 25498
rect 11612 25434 11664 25440
rect 11612 25152 11664 25158
rect 11612 25094 11664 25100
rect 11624 24682 11652 25094
rect 11612 24676 11664 24682
rect 11612 24618 11664 24624
rect 11612 23316 11664 23322
rect 11612 23258 11664 23264
rect 11624 23225 11652 23258
rect 11610 23216 11666 23225
rect 11610 23151 11666 23160
rect 11610 23080 11666 23089
rect 11610 23015 11666 23024
rect 11624 22098 11652 23015
rect 11612 22092 11664 22098
rect 11612 22034 11664 22040
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 11624 21418 11652 21898
rect 11716 21554 11744 26166
rect 11808 24206 11836 26862
rect 11888 25696 11940 25702
rect 11888 25638 11940 25644
rect 11900 25401 11928 25638
rect 11886 25392 11942 25401
rect 11886 25327 11942 25336
rect 11888 25220 11940 25226
rect 11888 25162 11940 25168
rect 11796 24200 11848 24206
rect 11796 24142 11848 24148
rect 11796 24064 11848 24070
rect 11796 24006 11848 24012
rect 11808 23118 11836 24006
rect 11796 23112 11848 23118
rect 11796 23054 11848 23060
rect 11900 22030 11928 25162
rect 11888 22024 11940 22030
rect 11808 21984 11888 22012
rect 11808 21622 11836 21984
rect 11888 21966 11940 21972
rect 11796 21616 11848 21622
rect 11796 21558 11848 21564
rect 11704 21548 11756 21554
rect 11704 21490 11756 21496
rect 11612 21412 11664 21418
rect 11612 21354 11664 21360
rect 11716 20754 11744 21490
rect 11796 21412 11848 21418
rect 11796 21354 11848 21360
rect 11624 20726 11744 20754
rect 11624 20369 11652 20726
rect 11808 20380 11836 21354
rect 11888 21344 11940 21350
rect 11888 21286 11940 21292
rect 11900 20602 11928 21286
rect 11888 20596 11940 20602
rect 11888 20538 11940 20544
rect 11888 20392 11940 20398
rect 11610 20360 11666 20369
rect 11808 20352 11888 20380
rect 11888 20334 11940 20340
rect 11610 20295 11666 20304
rect 11612 20256 11664 20262
rect 11612 20198 11664 20204
rect 11624 20058 11652 20198
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11532 19502 11744 19530
rect 11900 19514 11928 20334
rect 11992 20058 12020 27775
rect 12084 27033 12112 27814
rect 12070 27024 12126 27033
rect 12070 26959 12126 26968
rect 12072 26444 12124 26450
rect 12072 26386 12124 26392
rect 12084 25906 12112 26386
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 12176 24936 12204 30126
rect 12360 29510 12388 30688
rect 12440 30388 12492 30394
rect 12440 30330 12492 30336
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 12348 29504 12400 29510
rect 12348 29446 12400 29452
rect 12268 29050 12296 29446
rect 12268 29022 12388 29050
rect 12256 28960 12308 28966
rect 12254 28928 12256 28937
rect 12308 28928 12310 28937
rect 12254 28863 12310 28872
rect 12254 28792 12310 28801
rect 12254 28727 12256 28736
rect 12308 28727 12310 28736
rect 12256 28698 12308 28704
rect 12360 28121 12388 29022
rect 12346 28112 12402 28121
rect 12346 28047 12402 28056
rect 12348 28008 12400 28014
rect 12348 27950 12400 27956
rect 12360 27713 12388 27950
rect 12346 27704 12402 27713
rect 12346 27639 12402 27648
rect 12452 27554 12480 30330
rect 12544 29617 12572 30903
rect 12636 30716 12664 31214
rect 12728 31142 12756 31418
rect 12912 31346 12940 31726
rect 12992 31680 13044 31686
rect 12992 31622 13044 31628
rect 12900 31340 12952 31346
rect 12900 31282 12952 31288
rect 13004 31249 13032 31622
rect 12990 31240 13046 31249
rect 12990 31175 13046 31184
rect 12716 31136 12768 31142
rect 12716 31078 12768 31084
rect 12703 31036 13011 31045
rect 12703 31034 12709 31036
rect 12765 31034 12789 31036
rect 12845 31034 12869 31036
rect 12925 31034 12949 31036
rect 13005 31034 13011 31036
rect 12765 30982 12767 31034
rect 12947 30982 12949 31034
rect 12703 30980 12709 30982
rect 12765 30980 12789 30982
rect 12845 30980 12869 30982
rect 12925 30980 12949 30982
rect 13005 30980 13011 30982
rect 12703 30971 13011 30980
rect 13096 30818 13124 32184
rect 13004 30790 13124 30818
rect 13004 30734 13032 30790
rect 12716 30728 12768 30734
rect 12636 30688 12716 30716
rect 12716 30670 12768 30676
rect 12808 30728 12860 30734
rect 12808 30670 12860 30676
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 12728 30190 12756 30670
rect 12820 30394 12848 30670
rect 12808 30388 12860 30394
rect 12808 30330 12860 30336
rect 13188 30258 13216 32422
rect 13268 32224 13320 32230
rect 13268 32166 13320 32172
rect 13280 31385 13308 32166
rect 13372 31482 13400 32778
rect 13464 31929 13492 32807
rect 13450 31920 13506 31929
rect 13450 31855 13506 31864
rect 13556 31686 13584 32914
rect 13648 31929 13676 33390
rect 13634 31920 13690 31929
rect 13634 31855 13690 31864
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13544 31680 13596 31686
rect 13544 31622 13596 31628
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13266 31376 13322 31385
rect 13266 31311 13322 31320
rect 13648 31260 13676 31758
rect 13464 31232 13676 31260
rect 13268 31136 13320 31142
rect 13268 31078 13320 31084
rect 13176 30252 13228 30258
rect 13176 30194 13228 30200
rect 12716 30184 12768 30190
rect 12636 30144 12716 30172
rect 12530 29608 12586 29617
rect 12530 29543 12586 29552
rect 12532 29504 12584 29510
rect 12532 29446 12584 29452
rect 12544 28801 12572 29446
rect 12636 29238 12664 30144
rect 12716 30126 12768 30132
rect 12992 30184 13044 30190
rect 13044 30144 13124 30172
rect 12992 30126 13044 30132
rect 12703 29948 13011 29957
rect 12703 29946 12709 29948
rect 12765 29946 12789 29948
rect 12845 29946 12869 29948
rect 12925 29946 12949 29948
rect 13005 29946 13011 29948
rect 12765 29894 12767 29946
rect 12947 29894 12949 29946
rect 12703 29892 12709 29894
rect 12765 29892 12789 29894
rect 12845 29892 12869 29894
rect 12925 29892 12949 29894
rect 13005 29892 13011 29894
rect 12703 29883 13011 29892
rect 12624 29232 12676 29238
rect 12624 29174 12676 29180
rect 13096 29050 13124 30144
rect 13176 29572 13228 29578
rect 13176 29514 13228 29520
rect 13004 29022 13124 29050
rect 12716 28960 12768 28966
rect 13004 28948 13032 29022
rect 12768 28920 13032 28948
rect 13084 28960 13136 28966
rect 12716 28902 12768 28908
rect 13084 28902 13136 28908
rect 12703 28860 13011 28869
rect 12703 28858 12709 28860
rect 12765 28858 12789 28860
rect 12845 28858 12869 28860
rect 12925 28858 12949 28860
rect 13005 28858 13011 28860
rect 12765 28806 12767 28858
rect 12947 28806 12949 28858
rect 12703 28804 12709 28806
rect 12765 28804 12789 28806
rect 12845 28804 12869 28806
rect 12925 28804 12949 28806
rect 13005 28804 13011 28806
rect 12530 28792 12586 28801
rect 12703 28795 13011 28804
rect 12530 28727 12586 28736
rect 12268 27526 12480 27554
rect 12268 26926 12296 27526
rect 12544 27441 12572 28727
rect 12716 28552 12768 28558
rect 12714 28520 12716 28529
rect 12768 28520 12770 28529
rect 12714 28455 12770 28464
rect 12808 28484 12860 28490
rect 12808 28426 12860 28432
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 12728 28014 12756 28358
rect 12716 28008 12768 28014
rect 12716 27950 12768 27956
rect 12820 27860 12848 28426
rect 13096 28422 13124 28902
rect 13084 28416 13136 28422
rect 13084 28358 13136 28364
rect 12636 27832 12848 27860
rect 13084 27872 13136 27878
rect 12530 27432 12586 27441
rect 12348 27396 12400 27402
rect 12530 27367 12586 27376
rect 12348 27338 12400 27344
rect 12256 26920 12308 26926
rect 12256 26862 12308 26868
rect 12268 25974 12296 26862
rect 12360 26858 12388 27338
rect 12532 26920 12584 26926
rect 12532 26862 12584 26868
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 12544 26432 12572 26862
rect 12636 26586 12664 27832
rect 13084 27814 13136 27820
rect 12703 27772 13011 27781
rect 12703 27770 12709 27772
rect 12765 27770 12789 27772
rect 12845 27770 12869 27772
rect 12925 27770 12949 27772
rect 13005 27770 13011 27772
rect 12765 27718 12767 27770
rect 12947 27718 12949 27770
rect 12703 27716 12709 27718
rect 12765 27716 12789 27718
rect 12845 27716 12869 27718
rect 12925 27716 12949 27718
rect 13005 27716 13011 27718
rect 12703 27707 13011 27716
rect 12716 27328 12768 27334
rect 12716 27270 12768 27276
rect 12728 26994 12756 27270
rect 12716 26988 12768 26994
rect 12716 26930 12768 26936
rect 13096 26926 13124 27814
rect 13084 26920 13136 26926
rect 13084 26862 13136 26868
rect 12703 26684 13011 26693
rect 12703 26682 12709 26684
rect 12765 26682 12789 26684
rect 12845 26682 12869 26684
rect 12925 26682 12949 26684
rect 13005 26682 13011 26684
rect 12765 26630 12767 26682
rect 12947 26630 12949 26682
rect 12703 26628 12709 26630
rect 12765 26628 12789 26630
rect 12845 26628 12869 26630
rect 12925 26628 12949 26630
rect 13005 26628 13011 26630
rect 12703 26619 13011 26628
rect 12624 26580 12676 26586
rect 13096 26568 13124 26862
rect 12624 26522 12676 26528
rect 12820 26540 13124 26568
rect 12360 26404 12572 26432
rect 12256 25968 12308 25974
rect 12256 25910 12308 25916
rect 12084 24908 12204 24936
rect 11980 20052 12032 20058
rect 11980 19994 12032 20000
rect 12084 19854 12112 24908
rect 12164 24812 12216 24818
rect 12164 24754 12216 24760
rect 12176 24410 12204 24754
rect 12164 24404 12216 24410
rect 12164 24346 12216 24352
rect 12268 23730 12296 25910
rect 12360 25838 12388 26404
rect 12532 26308 12584 26314
rect 12532 26250 12584 26256
rect 12438 25936 12494 25945
rect 12438 25871 12440 25880
rect 12492 25871 12494 25880
rect 12440 25842 12492 25848
rect 12348 25832 12400 25838
rect 12348 25774 12400 25780
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 12254 23624 12310 23633
rect 12254 23559 12310 23568
rect 12164 23520 12216 23526
rect 12164 23462 12216 23468
rect 12176 21894 12204 23462
rect 12268 23032 12296 23559
rect 12360 23526 12388 25774
rect 12348 23520 12400 23526
rect 12348 23462 12400 23468
rect 12452 23186 12480 25842
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12348 23044 12400 23050
rect 12268 23004 12348 23032
rect 12348 22986 12400 22992
rect 12256 22568 12308 22574
rect 12360 22556 12388 22986
rect 12308 22528 12388 22556
rect 12256 22510 12308 22516
rect 12268 21962 12296 22510
rect 12452 22234 12480 23122
rect 12440 22228 12492 22234
rect 12440 22170 12492 22176
rect 12544 22094 12572 26250
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 12636 25498 12664 25706
rect 12820 25702 12848 26540
rect 12898 26480 12954 26489
rect 12954 26438 13124 26466
rect 12898 26415 12954 26424
rect 12808 25696 12860 25702
rect 12808 25638 12860 25644
rect 12703 25596 13011 25605
rect 12703 25594 12709 25596
rect 12765 25594 12789 25596
rect 12845 25594 12869 25596
rect 12925 25594 12949 25596
rect 13005 25594 13011 25596
rect 12765 25542 12767 25594
rect 12947 25542 12949 25594
rect 12703 25540 12709 25542
rect 12765 25540 12789 25542
rect 12845 25540 12869 25542
rect 12925 25540 12949 25542
rect 13005 25540 13011 25542
rect 12703 25531 13011 25540
rect 12624 25492 12676 25498
rect 12624 25434 12676 25440
rect 13096 25378 13124 26438
rect 13004 25350 13124 25378
rect 12808 25220 12860 25226
rect 12808 25162 12860 25168
rect 12820 24993 12848 25162
rect 12806 24984 12862 24993
rect 12806 24919 12862 24928
rect 12716 24812 12768 24818
rect 12636 24772 12716 24800
rect 12636 22642 12664 24772
rect 13004 24800 13032 25350
rect 13084 25220 13136 25226
rect 13084 25162 13136 25168
rect 12768 24772 13032 24800
rect 12716 24754 12768 24760
rect 12703 24508 13011 24517
rect 12703 24506 12709 24508
rect 12765 24506 12789 24508
rect 12845 24506 12869 24508
rect 12925 24506 12949 24508
rect 13005 24506 13011 24508
rect 12765 24454 12767 24506
rect 12947 24454 12949 24506
rect 12703 24452 12709 24454
rect 12765 24452 12789 24454
rect 12845 24452 12869 24454
rect 12925 24452 12949 24454
rect 13005 24452 13011 24454
rect 12703 24443 13011 24452
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12912 23662 12940 24006
rect 12900 23656 12952 23662
rect 12900 23598 12952 23604
rect 12703 23420 13011 23429
rect 12703 23418 12709 23420
rect 12765 23418 12789 23420
rect 12845 23418 12869 23420
rect 12925 23418 12949 23420
rect 13005 23418 13011 23420
rect 12765 23366 12767 23418
rect 12947 23366 12949 23418
rect 12703 23364 12709 23366
rect 12765 23364 12789 23366
rect 12845 23364 12869 23366
rect 12925 23364 12949 23366
rect 13005 23364 13011 23366
rect 12703 23355 13011 23364
rect 13096 23322 13124 25162
rect 13084 23316 13136 23322
rect 13084 23258 13136 23264
rect 13188 23225 13216 29514
rect 13280 28762 13308 31078
rect 13360 29300 13412 29306
rect 13360 29242 13412 29248
rect 13268 28756 13320 28762
rect 13268 28698 13320 28704
rect 13372 28642 13400 29242
rect 13280 28614 13400 28642
rect 13280 26382 13308 28614
rect 13464 28529 13492 31232
rect 13636 31136 13688 31142
rect 13636 31078 13688 31084
rect 13648 30172 13676 31078
rect 13740 30870 13768 33458
rect 13728 30864 13780 30870
rect 13728 30806 13780 30812
rect 13832 30326 13860 34546
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 13924 33017 13952 34002
rect 14108 33289 14136 35634
rect 14382 34844 14690 34853
rect 14382 34842 14388 34844
rect 14444 34842 14468 34844
rect 14524 34842 14548 34844
rect 14604 34842 14628 34844
rect 14684 34842 14690 34844
rect 14444 34790 14446 34842
rect 14626 34790 14628 34842
rect 14382 34788 14388 34790
rect 14444 34788 14468 34790
rect 14524 34788 14548 34790
rect 14604 34788 14628 34790
rect 14684 34788 14690 34790
rect 14382 34779 14690 34788
rect 14382 33756 14690 33765
rect 14382 33754 14388 33756
rect 14444 33754 14468 33756
rect 14524 33754 14548 33756
rect 14604 33754 14628 33756
rect 14684 33754 14690 33756
rect 14444 33702 14446 33754
rect 14626 33702 14628 33754
rect 14382 33700 14388 33702
rect 14444 33700 14468 33702
rect 14524 33700 14548 33702
rect 14604 33700 14628 33702
rect 14684 33700 14690 33702
rect 14382 33691 14690 33700
rect 14188 33380 14240 33386
rect 14188 33322 14240 33328
rect 14094 33280 14150 33289
rect 14094 33215 14150 33224
rect 13910 33008 13966 33017
rect 13910 32943 13966 32952
rect 13912 32360 13964 32366
rect 13912 32302 13964 32308
rect 13820 30320 13872 30326
rect 13820 30262 13872 30268
rect 13648 30144 13860 30172
rect 13544 29504 13596 29510
rect 13544 29446 13596 29452
rect 13450 28520 13506 28529
rect 13450 28455 13506 28464
rect 13452 28212 13504 28218
rect 13452 28154 13504 28160
rect 13360 28008 13412 28014
rect 13360 27950 13412 27956
rect 13372 26926 13400 27950
rect 13464 27713 13492 28154
rect 13556 28082 13584 29446
rect 13832 29186 13860 30144
rect 13924 30122 13952 32302
rect 14200 32065 14228 33322
rect 14280 32836 14332 32842
rect 14280 32778 14332 32784
rect 14186 32056 14242 32065
rect 14186 31991 14242 32000
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 13636 29164 13688 29170
rect 13832 29158 13952 29186
rect 13636 29106 13688 29112
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13450 27704 13506 27713
rect 13450 27639 13506 27648
rect 13452 27396 13504 27402
rect 13452 27338 13504 27344
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 13268 26376 13320 26382
rect 13268 26318 13320 26324
rect 13268 25900 13320 25906
rect 13372 25888 13400 26862
rect 13320 25860 13400 25888
rect 13268 25842 13320 25848
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13280 23662 13308 25638
rect 13372 24460 13400 25860
rect 13464 24585 13492 27338
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13556 26586 13584 26862
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13648 26042 13676 29106
rect 13820 29028 13872 29034
rect 13820 28970 13872 28976
rect 13728 28416 13780 28422
rect 13728 28358 13780 28364
rect 13636 26036 13688 26042
rect 13636 25978 13688 25984
rect 13740 25945 13768 28358
rect 13726 25936 13782 25945
rect 13726 25871 13782 25880
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 13556 24954 13584 25774
rect 13832 25673 13860 28970
rect 13924 27577 13952 29158
rect 13910 27568 13966 27577
rect 13910 27503 13966 27512
rect 14016 26874 14044 31826
rect 14292 31754 14320 32778
rect 14382 32668 14690 32677
rect 14382 32666 14388 32668
rect 14444 32666 14468 32668
rect 14524 32666 14548 32668
rect 14604 32666 14628 32668
rect 14684 32666 14690 32668
rect 14444 32614 14446 32666
rect 14626 32614 14628 32666
rect 14382 32612 14388 32614
rect 14444 32612 14468 32614
rect 14524 32612 14548 32614
rect 14604 32612 14628 32614
rect 14684 32612 14690 32614
rect 14382 32603 14690 32612
rect 14200 31726 14320 31754
rect 14200 31634 14228 31726
rect 14108 31606 14228 31634
rect 14280 31680 14332 31686
rect 14280 31622 14332 31628
rect 14108 30297 14136 31606
rect 14188 31340 14240 31346
rect 14188 31282 14240 31288
rect 14094 30288 14150 30297
rect 14094 30223 14150 30232
rect 14200 28218 14228 31282
rect 14292 31226 14320 31622
rect 14382 31580 14690 31589
rect 14382 31578 14388 31580
rect 14444 31578 14468 31580
rect 14524 31578 14548 31580
rect 14604 31578 14628 31580
rect 14684 31578 14690 31580
rect 14444 31526 14446 31578
rect 14626 31526 14628 31578
rect 14382 31524 14388 31526
rect 14444 31524 14468 31526
rect 14524 31524 14548 31526
rect 14604 31524 14628 31526
rect 14684 31524 14690 31526
rect 14382 31515 14690 31524
rect 14292 31198 14412 31226
rect 14280 31136 14332 31142
rect 14280 31078 14332 31084
rect 14188 28212 14240 28218
rect 14188 28154 14240 28160
rect 14292 28121 14320 31078
rect 14384 30666 14412 31198
rect 14372 30660 14424 30666
rect 14372 30602 14424 30608
rect 14382 30492 14690 30501
rect 14382 30490 14388 30492
rect 14444 30490 14468 30492
rect 14524 30490 14548 30492
rect 14604 30490 14628 30492
rect 14684 30490 14690 30492
rect 14444 30438 14446 30490
rect 14626 30438 14628 30490
rect 14382 30436 14388 30438
rect 14444 30436 14468 30438
rect 14524 30436 14548 30438
rect 14604 30436 14628 30438
rect 14684 30436 14690 30438
rect 14382 30427 14690 30436
rect 14382 29404 14690 29413
rect 14382 29402 14388 29404
rect 14444 29402 14468 29404
rect 14524 29402 14548 29404
rect 14604 29402 14628 29404
rect 14684 29402 14690 29404
rect 14444 29350 14446 29402
rect 14626 29350 14628 29402
rect 14382 29348 14388 29350
rect 14444 29348 14468 29350
rect 14524 29348 14548 29350
rect 14604 29348 14628 29350
rect 14684 29348 14690 29350
rect 14382 29339 14690 29348
rect 14382 28316 14690 28325
rect 14382 28314 14388 28316
rect 14444 28314 14468 28316
rect 14524 28314 14548 28316
rect 14604 28314 14628 28316
rect 14684 28314 14690 28316
rect 14444 28262 14446 28314
rect 14626 28262 14628 28314
rect 14382 28260 14388 28262
rect 14444 28260 14468 28262
rect 14524 28260 14548 28262
rect 14604 28260 14628 28262
rect 14684 28260 14690 28262
rect 14382 28251 14690 28260
rect 14278 28112 14334 28121
rect 14278 28047 14334 28056
rect 14382 27228 14690 27237
rect 14382 27226 14388 27228
rect 14444 27226 14468 27228
rect 14524 27226 14548 27228
rect 14604 27226 14628 27228
rect 14684 27226 14690 27228
rect 14444 27174 14446 27226
rect 14626 27174 14628 27226
rect 14382 27172 14388 27174
rect 14444 27172 14468 27174
rect 14524 27172 14548 27174
rect 14604 27172 14628 27174
rect 14684 27172 14690 27174
rect 14382 27163 14690 27172
rect 13924 26846 14044 26874
rect 13818 25664 13874 25673
rect 13818 25599 13874 25608
rect 13820 25152 13872 25158
rect 13820 25094 13872 25100
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 13450 24576 13506 24585
rect 13450 24511 13506 24520
rect 13372 24432 13676 24460
rect 13648 23746 13676 24432
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13464 23730 13676 23746
rect 13452 23724 13676 23730
rect 13504 23718 13676 23724
rect 13452 23666 13504 23672
rect 13268 23656 13320 23662
rect 13268 23598 13320 23604
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13174 23216 13230 23225
rect 13174 23151 13230 23160
rect 13188 23050 13216 23151
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 12703 22332 13011 22341
rect 12703 22330 12709 22332
rect 12765 22330 12789 22332
rect 12845 22330 12869 22332
rect 12925 22330 12949 22332
rect 13005 22330 13011 22332
rect 12765 22278 12767 22330
rect 12947 22278 12949 22330
rect 12703 22276 12709 22278
rect 12765 22276 12789 22278
rect 12845 22276 12869 22278
rect 12925 22276 12949 22278
rect 13005 22276 13011 22278
rect 12703 22267 13011 22276
rect 13176 22228 13228 22234
rect 13176 22170 13228 22176
rect 12452 22066 12572 22094
rect 12256 21956 12308 21962
rect 12256 21898 12308 21904
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 12254 21312 12310 21321
rect 12254 21247 12310 21256
rect 12162 20632 12218 20641
rect 12162 20567 12218 20576
rect 12176 20534 12204 20567
rect 12164 20528 12216 20534
rect 12164 20470 12216 20476
rect 12268 20482 12296 21247
rect 12268 20454 12388 20482
rect 12072 19848 12124 19854
rect 12256 19848 12308 19854
rect 12072 19790 12124 19796
rect 12162 19816 12218 19825
rect 11612 19372 11664 19378
rect 11612 19314 11664 19320
rect 11520 18624 11572 18630
rect 11520 18566 11572 18572
rect 10876 17672 10928 17678
rect 10874 17640 10876 17649
rect 11428 17672 11480 17678
rect 10928 17640 10930 17649
rect 11428 17614 11480 17620
rect 10874 17575 10930 17584
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10876 17536 10928 17542
rect 10876 17478 10928 17484
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 10782 17368 10838 17377
rect 10782 17303 10838 17312
rect 10796 16980 10824 17303
rect 10888 17116 10916 17478
rect 11024 17436 11332 17445
rect 11024 17434 11030 17436
rect 11086 17434 11110 17436
rect 11166 17434 11190 17436
rect 11246 17434 11270 17436
rect 11326 17434 11332 17436
rect 11086 17382 11088 17434
rect 11268 17382 11270 17434
rect 11024 17380 11030 17382
rect 11086 17380 11110 17382
rect 11166 17380 11190 17382
rect 11246 17380 11270 17382
rect 11326 17380 11332 17382
rect 11024 17371 11332 17380
rect 11336 17332 11388 17338
rect 11336 17274 11388 17280
rect 11348 17202 11376 17274
rect 11440 17202 11468 17478
rect 11152 17196 11204 17202
rect 11152 17138 11204 17144
rect 11336 17196 11388 17202
rect 11336 17138 11388 17144
rect 11428 17196 11480 17202
rect 11428 17138 11480 17144
rect 10968 17128 11020 17134
rect 10888 17088 10968 17116
rect 11164 17105 11192 17138
rect 10968 17070 11020 17076
rect 11150 17096 11206 17105
rect 11150 17031 11206 17040
rect 11060 16992 11112 16998
rect 10796 16952 11060 16980
rect 11060 16934 11112 16940
rect 11244 16992 11296 16998
rect 11244 16934 11296 16940
rect 11256 16726 11284 16934
rect 10876 16720 10928 16726
rect 11244 16720 11296 16726
rect 10876 16662 10928 16668
rect 11150 16688 11206 16697
rect 10888 15144 10916 16662
rect 11244 16662 11296 16668
rect 11150 16623 11206 16632
rect 11164 16590 11192 16623
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11024 16348 11332 16357
rect 11024 16346 11030 16348
rect 11086 16346 11110 16348
rect 11166 16346 11190 16348
rect 11246 16346 11270 16348
rect 11326 16346 11332 16348
rect 11086 16294 11088 16346
rect 11268 16294 11270 16346
rect 11024 16292 11030 16294
rect 11086 16292 11110 16294
rect 11166 16292 11190 16294
rect 11246 16292 11270 16294
rect 11326 16292 11332 16294
rect 11024 16283 11332 16292
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11072 15706 11100 16118
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11058 15600 11114 15609
rect 11058 15535 11060 15544
rect 11112 15535 11114 15544
rect 11060 15506 11112 15512
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11164 15366 11192 15438
rect 11152 15360 11204 15366
rect 11152 15302 11204 15308
rect 11024 15260 11332 15269
rect 11024 15258 11030 15260
rect 11086 15258 11110 15260
rect 11166 15258 11190 15260
rect 11246 15258 11270 15260
rect 11326 15258 11332 15260
rect 11086 15206 11088 15258
rect 11268 15206 11270 15258
rect 11024 15204 11030 15206
rect 11086 15204 11110 15206
rect 11166 15204 11190 15206
rect 11246 15204 11270 15206
rect 11326 15204 11332 15206
rect 11024 15195 11332 15204
rect 10888 15116 11008 15144
rect 10782 14920 10838 14929
rect 10838 14878 10916 14906
rect 10782 14855 10838 14864
rect 10784 14476 10836 14482
rect 10784 14418 10836 14424
rect 10796 14074 10824 14418
rect 10784 14068 10836 14074
rect 10784 14010 10836 14016
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10888 13530 10916 14878
rect 10980 14278 11008 15116
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 11072 14657 11100 14894
rect 11336 14816 11388 14822
rect 11336 14758 11388 14764
rect 11058 14648 11114 14657
rect 11058 14583 11114 14592
rect 11150 14512 11206 14521
rect 11060 14476 11112 14482
rect 11150 14447 11206 14456
rect 11060 14418 11112 14424
rect 10968 14272 11020 14278
rect 11072 14260 11100 14418
rect 11164 14396 11192 14447
rect 11348 14414 11376 14758
rect 11244 14408 11296 14414
rect 11164 14368 11244 14396
rect 11244 14350 11296 14356
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11440 14260 11468 16390
rect 11532 15570 11560 18566
rect 11624 16794 11652 19314
rect 11716 18290 11744 19502
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 12084 18986 12112 19790
rect 12256 19790 12308 19796
rect 12162 19751 12218 19760
rect 12176 19310 12204 19751
rect 12268 19514 12296 19790
rect 12256 19508 12308 19514
rect 12256 19450 12308 19456
rect 12360 19394 12388 20454
rect 12452 19446 12480 22066
rect 12992 21888 13044 21894
rect 12992 21830 13044 21836
rect 13004 21486 13032 21830
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 13084 21412 13136 21418
rect 13084 21354 13136 21360
rect 12703 21244 13011 21253
rect 12703 21242 12709 21244
rect 12765 21242 12789 21244
rect 12845 21242 12869 21244
rect 12925 21242 12949 21244
rect 13005 21242 13011 21244
rect 12765 21190 12767 21242
rect 12947 21190 12949 21242
rect 12703 21188 12709 21190
rect 12765 21188 12789 21190
rect 12845 21188 12869 21190
rect 12925 21188 12949 21190
rect 13005 21188 13011 21190
rect 12703 21179 13011 21188
rect 12716 21004 12768 21010
rect 12716 20946 12768 20952
rect 12532 20868 12584 20874
rect 12532 20810 12584 20816
rect 12268 19366 12388 19394
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12084 18958 12204 18986
rect 12070 18864 12126 18873
rect 12070 18799 12126 18808
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11704 17672 11756 17678
rect 11702 17640 11704 17649
rect 11756 17640 11758 17649
rect 11702 17575 11758 17584
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11716 17241 11744 17478
rect 11702 17232 11758 17241
rect 11702 17167 11758 17176
rect 11612 16788 11664 16794
rect 11612 16730 11664 16736
rect 11612 16448 11664 16454
rect 11610 16416 11612 16425
rect 11664 16416 11666 16425
rect 11610 16351 11666 16360
rect 11612 16040 11664 16046
rect 11612 15982 11664 15988
rect 11520 15564 11572 15570
rect 11520 15506 11572 15512
rect 11072 14232 11468 14260
rect 10968 14214 11020 14220
rect 11024 14172 11332 14181
rect 11024 14170 11030 14172
rect 11086 14170 11110 14172
rect 11166 14170 11190 14172
rect 11246 14170 11270 14172
rect 11326 14170 11332 14172
rect 11086 14118 11088 14170
rect 11268 14118 11270 14170
rect 11024 14116 11030 14118
rect 11086 14116 11110 14118
rect 11166 14116 11190 14118
rect 11246 14116 11270 14118
rect 11326 14116 11332 14118
rect 11024 14107 11332 14116
rect 11334 13968 11390 13977
rect 11440 13954 11468 14232
rect 11390 13926 11468 13954
rect 11334 13903 11390 13912
rect 11520 13864 11572 13870
rect 11624 13852 11652 15982
rect 11716 15706 11744 17167
rect 11808 16182 11836 18158
rect 11886 17232 11942 17241
rect 11886 17167 11942 17176
rect 11900 16590 11928 17167
rect 11992 16794 12020 18362
rect 12084 17882 12112 18799
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 12070 17640 12126 17649
rect 12070 17575 12126 17584
rect 12084 17134 12112 17575
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 11980 16788 12032 16794
rect 11980 16730 12032 16736
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11796 16176 11848 16182
rect 11796 16118 11848 16124
rect 11796 16040 11848 16046
rect 12084 16028 12112 17070
rect 12176 16658 12204 18958
rect 12268 16998 12296 19366
rect 12440 19304 12492 19310
rect 12440 19246 12492 19252
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12360 18612 12388 18838
rect 12452 18766 12480 19246
rect 12544 19174 12572 20810
rect 12728 20641 12756 20946
rect 12714 20632 12770 20641
rect 12714 20567 12770 20576
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12636 20040 12664 20198
rect 12703 20156 13011 20165
rect 12703 20154 12709 20156
rect 12765 20154 12789 20156
rect 12845 20154 12869 20156
rect 12925 20154 12949 20156
rect 13005 20154 13011 20156
rect 12765 20102 12767 20154
rect 12947 20102 12949 20154
rect 12703 20100 12709 20102
rect 12765 20100 12789 20102
rect 12845 20100 12869 20102
rect 12925 20100 12949 20102
rect 13005 20100 13011 20102
rect 12703 20091 13011 20100
rect 12636 20012 12756 20040
rect 12622 19952 12678 19961
rect 12728 19922 12756 20012
rect 13096 19938 13124 21354
rect 12622 19887 12624 19896
rect 12676 19887 12678 19896
rect 12716 19916 12768 19922
rect 12624 19858 12676 19864
rect 12716 19858 12768 19864
rect 12912 19910 13124 19938
rect 12912 19334 12940 19910
rect 12992 19848 13044 19854
rect 13188 19836 13216 22170
rect 13280 22166 13308 23598
rect 13556 23322 13584 23598
rect 13544 23316 13596 23322
rect 13544 23258 13596 23264
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13268 22160 13320 22166
rect 13268 22102 13320 22108
rect 13372 22094 13400 22714
rect 13452 22432 13504 22438
rect 13452 22374 13504 22380
rect 13464 22250 13492 22374
rect 13464 22222 13584 22250
rect 13372 22066 13492 22094
rect 13268 21480 13320 21486
rect 13360 21480 13412 21486
rect 13268 21422 13320 21428
rect 13358 21448 13360 21457
rect 13412 21448 13414 21457
rect 13280 21049 13308 21422
rect 13358 21383 13414 21392
rect 13266 21040 13322 21049
rect 13266 20975 13322 20984
rect 13280 20398 13308 20975
rect 13360 20936 13412 20942
rect 13360 20878 13412 20884
rect 13268 20392 13320 20398
rect 13268 20334 13320 20340
rect 13044 19808 13216 19836
rect 12992 19790 13044 19796
rect 12912 19306 13124 19334
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12703 19068 13011 19077
rect 12703 19066 12709 19068
rect 12765 19066 12789 19068
rect 12845 19066 12869 19068
rect 12925 19066 12949 19068
rect 13005 19066 13011 19068
rect 12765 19014 12767 19066
rect 12947 19014 12949 19066
rect 12703 19012 12709 19014
rect 12765 19012 12789 19014
rect 12845 19012 12869 19014
rect 12925 19012 12949 19014
rect 13005 19012 13011 19014
rect 12703 19003 13011 19012
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12532 18624 12584 18630
rect 12360 18584 12480 18612
rect 12346 18320 12402 18329
rect 12346 18255 12348 18264
rect 12400 18255 12402 18264
rect 12348 18226 12400 18232
rect 12346 18184 12402 18193
rect 12346 18119 12402 18128
rect 12360 17134 12388 18119
rect 12452 18086 12480 18584
rect 12532 18566 12584 18572
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12348 17128 12400 17134
rect 12348 17070 12400 17076
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12268 16708 12296 16934
rect 12268 16680 12388 16708
rect 12164 16652 12216 16658
rect 12216 16612 12296 16640
rect 12164 16594 12216 16600
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 11848 16000 12112 16028
rect 11796 15982 11848 15988
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11888 15632 11940 15638
rect 11888 15574 11940 15580
rect 12070 15600 12126 15609
rect 11702 15464 11758 15473
rect 11758 15422 11836 15450
rect 11702 15399 11758 15408
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11716 14249 11744 14962
rect 11702 14240 11758 14249
rect 11702 14175 11758 14184
rect 11808 13938 11836 15422
rect 11900 14657 11928 15574
rect 12070 15535 12072 15544
rect 12124 15535 12126 15544
rect 12072 15506 12124 15512
rect 12176 15366 12204 16458
rect 12164 15360 12216 15366
rect 12164 15302 12216 15308
rect 12162 15192 12218 15201
rect 12162 15127 12218 15136
rect 12072 15020 12124 15026
rect 12072 14962 12124 14968
rect 12084 14822 12112 14962
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11886 14648 11942 14657
rect 11886 14583 11942 14592
rect 11900 14346 11928 14583
rect 12176 14550 12204 15127
rect 12164 14544 12216 14550
rect 11978 14512 12034 14521
rect 12164 14486 12216 14492
rect 11978 14447 12034 14456
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11796 13932 11848 13938
rect 11796 13874 11848 13880
rect 11572 13824 11652 13852
rect 11808 13818 11836 13874
rect 11520 13806 11572 13812
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 11244 13320 11296 13326
rect 11242 13288 11244 13297
rect 11296 13288 11298 13297
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10784 13252 10836 13258
rect 11242 13223 11298 13232
rect 10784 13194 10836 13200
rect 10704 12050 10732 13194
rect 10796 12986 10824 13194
rect 11428 13184 11480 13190
rect 11428 13126 11480 13132
rect 11024 13084 11332 13093
rect 11024 13082 11030 13084
rect 11086 13082 11110 13084
rect 11166 13082 11190 13084
rect 11246 13082 11270 13084
rect 11326 13082 11332 13084
rect 11086 13030 11088 13082
rect 11268 13030 11270 13082
rect 11024 13028 11030 13030
rect 11086 13028 11110 13030
rect 11166 13028 11190 13030
rect 11246 13028 11270 13030
rect 11326 13028 11332 13030
rect 11024 13019 11332 13028
rect 10784 12980 10836 12986
rect 10784 12922 10836 12928
rect 11336 12640 11388 12646
rect 11334 12608 11336 12617
rect 11388 12608 11390 12617
rect 11334 12543 11390 12552
rect 10704 12022 10824 12050
rect 10796 11762 10824 12022
rect 11024 11996 11332 12005
rect 11024 11994 11030 11996
rect 11086 11994 11110 11996
rect 11166 11994 11190 11996
rect 11246 11994 11270 11996
rect 11326 11994 11332 11996
rect 11086 11942 11088 11994
rect 11268 11942 11270 11994
rect 11024 11940 11030 11942
rect 11086 11940 11110 11942
rect 11166 11940 11190 11942
rect 11246 11940 11270 11942
rect 11326 11940 11332 11942
rect 11024 11931 11332 11940
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 11440 11558 11468 13126
rect 11428 11552 11480 11558
rect 11428 11494 11480 11500
rect 11532 11354 11560 13806
rect 11716 13790 11836 13818
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11624 12073 11652 12106
rect 11610 12064 11666 12073
rect 11610 11999 11666 12008
rect 11716 11744 11744 13790
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 12646 11836 13670
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11808 12152 11836 12582
rect 11900 12442 11928 13330
rect 11992 12782 12020 14447
rect 12164 14340 12216 14346
rect 12164 14282 12216 14288
rect 12176 13274 12204 14282
rect 12084 13246 12204 13274
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 12084 12306 12112 13246
rect 12164 12708 12216 12714
rect 12164 12650 12216 12656
rect 12176 12345 12204 12650
rect 12162 12336 12218 12345
rect 12072 12300 12124 12306
rect 12162 12271 12218 12280
rect 12072 12242 12124 12248
rect 11980 12164 12032 12170
rect 11808 12124 11980 12152
rect 11980 12106 12032 12112
rect 12084 11914 12112 12242
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 11992 11886 12112 11914
rect 11796 11756 11848 11762
rect 11716 11716 11796 11744
rect 11796 11698 11848 11704
rect 11992 11642 12020 11886
rect 12072 11824 12124 11830
rect 12070 11792 12072 11801
rect 12124 11792 12126 11801
rect 12070 11727 12126 11736
rect 11900 11626 12020 11642
rect 11888 11620 12020 11626
rect 11940 11614 12020 11620
rect 12070 11656 12126 11665
rect 12070 11591 12126 11600
rect 11888 11562 11940 11568
rect 11886 11520 11942 11529
rect 11886 11455 11942 11464
rect 11520 11348 11572 11354
rect 11520 11290 11572 11296
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 11794 11248 11850 11257
rect 10704 10810 10732 11222
rect 11794 11183 11850 11192
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 11428 11144 11480 11150
rect 11612 11144 11664 11150
rect 11480 11104 11560 11132
rect 11428 11086 11480 11092
rect 10600 10804 10652 10810
rect 10600 10746 10652 10752
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10508 10260 10560 10266
rect 10244 10220 10318 10248
rect 10290 10146 10318 10220
rect 10508 10202 10560 10208
rect 10269 10118 10318 10146
rect 10796 10130 10824 10406
rect 10784 10124 10836 10130
rect 10140 10056 10192 10062
rect 10138 10024 10140 10033
rect 10269 10044 10297 10118
rect 10784 10066 10836 10072
rect 10192 10024 10194 10033
rect 10138 9959 10194 9968
rect 10244 10016 10297 10044
rect 10414 10024 10470 10033
rect 10244 9586 10272 10016
rect 10414 9959 10470 9968
rect 10428 9586 10456 9959
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10416 9580 10468 9586
rect 10468 9540 10640 9568
rect 10416 9522 10468 9528
rect 10152 9353 10180 9522
rect 10138 9344 10194 9353
rect 10138 9279 10194 9288
rect 10152 8022 10180 9279
rect 10140 8016 10192 8022
rect 10140 7958 10192 7964
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10048 7200 10100 7206
rect 10048 7142 10100 7148
rect 9770 6967 9826 6976
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9956 6792 10008 6798
rect 9770 6760 9826 6769
rect 9956 6734 10008 6740
rect 9770 6695 9826 6704
rect 9784 6458 9812 6695
rect 9968 6458 9996 6734
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9600 6174 9812 6202
rect 9784 6168 9812 6174
rect 9956 6180 10008 6186
rect 9784 6140 9956 6168
rect 10152 6168 10180 7210
rect 10244 6304 10272 9522
rect 10506 9344 10562 9353
rect 10428 9302 10506 9330
rect 10428 8974 10456 9302
rect 10506 9279 10562 9288
rect 10612 9024 10640 9540
rect 10888 9450 10916 11086
rect 11024 10908 11332 10917
rect 11024 10906 11030 10908
rect 11086 10906 11110 10908
rect 11166 10906 11190 10908
rect 11246 10906 11270 10908
rect 11326 10906 11332 10908
rect 11086 10854 11088 10906
rect 11268 10854 11270 10906
rect 11024 10852 11030 10854
rect 11086 10852 11110 10854
rect 11166 10852 11190 10854
rect 11246 10852 11270 10854
rect 11326 10852 11332 10854
rect 11024 10843 11332 10852
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11060 10532 11112 10538
rect 11060 10474 11112 10480
rect 11072 10062 11100 10474
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11024 9820 11332 9829
rect 11024 9818 11030 9820
rect 11086 9818 11110 9820
rect 11166 9818 11190 9820
rect 11246 9818 11270 9820
rect 11326 9818 11332 9820
rect 11086 9766 11088 9818
rect 11268 9766 11270 9818
rect 11024 9764 11030 9766
rect 11086 9764 11110 9766
rect 11166 9764 11190 9766
rect 11246 9764 11270 9766
rect 11326 9764 11332 9766
rect 11024 9755 11332 9764
rect 10876 9444 10928 9450
rect 10876 9386 10928 9392
rect 11336 9444 11388 9450
rect 11336 9386 11388 9392
rect 11242 9072 11298 9081
rect 10692 9036 10744 9042
rect 10612 8996 10692 9024
rect 11348 9042 11376 9386
rect 11440 9353 11468 10746
rect 11426 9344 11482 9353
rect 11426 9279 11482 9288
rect 11532 9178 11560 11104
rect 11612 11086 11664 11092
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11624 10266 11652 11086
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11610 10160 11666 10169
rect 11610 10095 11612 10104
rect 11664 10095 11666 10104
rect 11612 10066 11664 10072
rect 11612 9920 11664 9926
rect 11612 9862 11664 9868
rect 11624 9654 11652 9862
rect 11612 9648 11664 9654
rect 11612 9590 11664 9596
rect 11610 9480 11666 9489
rect 11610 9415 11666 9424
rect 11520 9172 11572 9178
rect 11520 9114 11572 9120
rect 11242 9007 11298 9016
rect 11336 9036 11388 9042
rect 10692 8978 10744 8984
rect 10416 8968 10468 8974
rect 10416 8910 10468 8916
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10336 7392 10364 8570
rect 10428 7936 10456 8910
rect 10520 8838 10548 8910
rect 10704 8838 10732 8978
rect 11256 8922 11284 9007
rect 11336 8978 11388 8984
rect 11256 8894 11468 8922
rect 10508 8832 10560 8838
rect 10692 8832 10744 8838
rect 10560 8792 10640 8820
rect 10508 8774 10560 8780
rect 10612 8294 10640 8792
rect 10692 8774 10744 8780
rect 11024 8732 11332 8741
rect 11024 8730 11030 8732
rect 11086 8730 11110 8732
rect 11166 8730 11190 8732
rect 11246 8730 11270 8732
rect 11326 8730 11332 8732
rect 11086 8678 11088 8730
rect 11268 8678 11270 8730
rect 11024 8676 11030 8678
rect 11086 8676 11110 8678
rect 11166 8676 11190 8678
rect 11246 8676 11270 8678
rect 11326 8676 11332 8678
rect 11024 8667 11332 8676
rect 11334 8528 11390 8537
rect 11440 8498 11468 8894
rect 11334 8463 11390 8472
rect 11428 8492 11480 8498
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10612 7954 10640 8230
rect 10508 7948 10560 7954
rect 10428 7908 10508 7936
rect 10508 7890 10560 7896
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10784 7880 10836 7886
rect 10704 7840 10784 7868
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10520 7410 10548 7686
rect 10416 7404 10468 7410
rect 10336 7364 10416 7392
rect 10416 7346 10468 7352
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10704 7342 10732 7840
rect 10784 7822 10836 7828
rect 10784 7744 10836 7750
rect 10782 7712 10784 7721
rect 10836 7712 10838 7721
rect 10782 7647 10838 7656
rect 10782 7440 10838 7449
rect 10782 7375 10838 7384
rect 10692 7336 10744 7342
rect 10520 7284 10692 7290
rect 10520 7278 10744 7284
rect 10520 7262 10732 7278
rect 10520 6866 10548 7262
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10322 6352 10378 6361
rect 10520 6322 10548 6802
rect 10244 6296 10322 6304
rect 10244 6276 10324 6296
rect 10376 6287 10378 6296
rect 10508 6316 10560 6322
rect 10324 6258 10376 6264
rect 10508 6258 10560 6264
rect 10008 6140 10180 6168
rect 9956 6122 10008 6128
rect 9232 6072 9352 6100
rect 9232 4622 9260 6072
rect 9345 6012 9653 6021
rect 9345 6010 9351 6012
rect 9407 6010 9431 6012
rect 9487 6010 9511 6012
rect 9567 6010 9591 6012
rect 9647 6010 9653 6012
rect 9407 5958 9409 6010
rect 9589 5958 9591 6010
rect 9345 5956 9351 5958
rect 9407 5956 9431 5958
rect 9487 5956 9511 5958
rect 9567 5956 9591 5958
rect 9647 5956 9653 5958
rect 9345 5947 9653 5956
rect 9345 4924 9653 4933
rect 9345 4922 9351 4924
rect 9407 4922 9431 4924
rect 9487 4922 9511 4924
rect 9567 4922 9591 4924
rect 9647 4922 9653 4924
rect 9407 4870 9409 4922
rect 9589 4870 9591 4922
rect 9345 4868 9351 4870
rect 9407 4868 9431 4870
rect 9487 4868 9511 4870
rect 9567 4868 9591 4870
rect 9647 4868 9653 4870
rect 9345 4859 9653 4868
rect 9968 4826 9996 6122
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 9956 4820 10008 4826
rect 9956 4762 10008 4768
rect 10244 4690 10272 5102
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9232 4282 9260 4558
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 10336 4214 10364 6258
rect 10520 5370 10548 6258
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10612 4622 10640 7142
rect 10796 6746 10824 7375
rect 10888 6882 10916 8366
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 7857 11192 8298
rect 11256 7993 11284 8366
rect 11242 7984 11298 7993
rect 11242 7919 11298 7928
rect 11150 7848 11206 7857
rect 11150 7783 11206 7792
rect 11348 7732 11376 8463
rect 11428 8434 11480 8440
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 11348 7704 11468 7732
rect 11024 7644 11332 7653
rect 11024 7642 11030 7644
rect 11086 7642 11110 7644
rect 11166 7642 11190 7644
rect 11246 7642 11270 7644
rect 11326 7642 11332 7644
rect 11086 7590 11088 7642
rect 11268 7590 11270 7642
rect 11024 7588 11030 7590
rect 11086 7588 11110 7590
rect 11166 7588 11190 7590
rect 11246 7588 11270 7590
rect 11326 7588 11332 7590
rect 11024 7579 11332 7588
rect 11440 7410 11468 7704
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 10888 6854 11008 6882
rect 10796 6730 10916 6746
rect 10796 6724 10928 6730
rect 10796 6718 10876 6724
rect 10876 6666 10928 6672
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10692 5772 10744 5778
rect 10796 5760 10824 6598
rect 10888 6254 10916 6666
rect 10980 6662 11008 6854
rect 11244 6792 11296 6798
rect 11440 6780 11468 7346
rect 11296 6752 11468 6780
rect 11244 6734 11296 6740
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 11024 6556 11332 6565
rect 11024 6554 11030 6556
rect 11086 6554 11110 6556
rect 11166 6554 11190 6556
rect 11246 6554 11270 6556
rect 11326 6554 11332 6556
rect 11086 6502 11088 6554
rect 11268 6502 11270 6554
rect 11024 6500 11030 6502
rect 11086 6500 11110 6502
rect 11166 6500 11190 6502
rect 11246 6500 11270 6502
rect 11326 6500 11332 6502
rect 11024 6491 11332 6500
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 10968 6180 11020 6186
rect 10968 6122 11020 6128
rect 10980 5846 11008 6122
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 10968 5840 11020 5846
rect 10968 5782 11020 5788
rect 11164 5778 11192 6054
rect 11532 5778 11560 7822
rect 11624 7290 11652 9415
rect 11716 9178 11744 11086
rect 11808 10674 11836 11183
rect 11900 10810 11928 11455
rect 11978 10976 12034 10985
rect 11978 10911 12034 10920
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11886 10704 11942 10713
rect 11796 10668 11848 10674
rect 11886 10639 11888 10648
rect 11796 10610 11848 10616
rect 11940 10639 11942 10648
rect 11888 10610 11940 10616
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11808 9926 11836 9998
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11808 8634 11836 9862
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11716 7449 11744 8502
rect 11900 7886 11928 10610
rect 11992 8090 12020 10911
rect 12084 10674 12112 11591
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12072 10056 12124 10062
rect 12072 9998 12124 10004
rect 12084 8838 12112 9998
rect 12176 9926 12204 12106
rect 12268 10810 12296 16612
rect 12360 15094 12388 16680
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12452 14958 12480 18022
rect 12544 17134 12572 18566
rect 12624 18216 12676 18222
rect 12624 18158 12676 18164
rect 12636 17882 12664 18158
rect 12703 17980 13011 17989
rect 12703 17978 12709 17980
rect 12765 17978 12789 17980
rect 12845 17978 12869 17980
rect 12925 17978 12949 17980
rect 13005 17978 13011 17980
rect 12765 17926 12767 17978
rect 12947 17926 12949 17978
rect 12703 17924 12709 17926
rect 12765 17924 12789 17926
rect 12845 17924 12869 17926
rect 12925 17924 12949 17926
rect 13005 17924 13011 17926
rect 12703 17915 13011 17924
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 13096 17814 13124 19306
rect 13084 17808 13136 17814
rect 13084 17750 13136 17756
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12532 17128 12584 17134
rect 12532 17070 12584 17076
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12544 16726 12572 16934
rect 12532 16720 12584 16726
rect 12532 16662 12584 16668
rect 12530 15056 12586 15065
rect 12530 14991 12532 15000
rect 12584 14991 12586 15000
rect 12532 14962 12584 14968
rect 12440 14952 12492 14958
rect 12492 14900 12572 14906
rect 12440 14894 12572 14900
rect 12452 14878 12572 14894
rect 12438 14648 12494 14657
rect 12438 14583 12494 14592
rect 12452 14482 12480 14583
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12348 14000 12400 14006
rect 12440 14000 12492 14006
rect 12348 13942 12400 13948
rect 12438 13968 12440 13977
rect 12492 13968 12494 13977
rect 12360 13394 12388 13942
rect 12438 13903 12494 13912
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13394 12480 13670
rect 12348 13388 12400 13394
rect 12348 13330 12400 13336
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12544 13274 12572 14878
rect 12452 13246 12572 13274
rect 12346 12880 12402 12889
rect 12346 12815 12402 12824
rect 12360 11898 12388 12815
rect 12452 12646 12480 13246
rect 12636 12782 12664 17682
rect 13188 17678 13216 19808
rect 13268 19848 13320 19854
rect 13268 19790 13320 19796
rect 13280 19514 13308 19790
rect 13268 19508 13320 19514
rect 13268 19450 13320 19456
rect 13268 19372 13320 19378
rect 13268 19314 13320 19320
rect 13084 17672 13136 17678
rect 13084 17614 13136 17620
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 12990 17504 13046 17513
rect 12990 17439 13046 17448
rect 13004 16998 13032 17439
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 12703 16892 13011 16901
rect 12703 16890 12709 16892
rect 12765 16890 12789 16892
rect 12845 16890 12869 16892
rect 12925 16890 12949 16892
rect 13005 16890 13011 16892
rect 12765 16838 12767 16890
rect 12947 16838 12949 16890
rect 12703 16836 12709 16838
rect 12765 16836 12789 16838
rect 12845 16836 12869 16838
rect 12925 16836 12949 16838
rect 13005 16836 13011 16838
rect 12703 16827 13011 16836
rect 12716 16788 12768 16794
rect 12768 16748 12848 16776
rect 12716 16730 12768 16736
rect 12716 16652 12768 16658
rect 12716 16594 12768 16600
rect 12728 16250 12756 16594
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12820 16114 12848 16748
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 13096 15881 13124 17614
rect 13188 16794 13216 17614
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13176 16584 13228 16590
rect 13280 16572 13308 19314
rect 13228 16544 13308 16572
rect 13176 16526 13228 16532
rect 13082 15872 13138 15881
rect 12703 15804 13011 15813
rect 13082 15807 13138 15816
rect 12703 15802 12709 15804
rect 12765 15802 12789 15804
rect 12845 15802 12869 15804
rect 12925 15802 12949 15804
rect 13005 15802 13011 15804
rect 12765 15750 12767 15802
rect 12947 15750 12949 15802
rect 12703 15748 12709 15750
rect 12765 15748 12789 15750
rect 12845 15748 12869 15750
rect 12925 15748 12949 15750
rect 13005 15748 13011 15750
rect 12703 15739 13011 15748
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 14958 13032 15302
rect 12992 14952 13044 14958
rect 12992 14894 13044 14900
rect 12703 14716 13011 14725
rect 12703 14714 12709 14716
rect 12765 14714 12789 14716
rect 12845 14714 12869 14716
rect 12925 14714 12949 14716
rect 13005 14714 13011 14716
rect 12765 14662 12767 14714
rect 12947 14662 12949 14714
rect 12703 14660 12709 14662
rect 12765 14660 12789 14662
rect 12845 14660 12869 14662
rect 12925 14660 12949 14662
rect 13005 14660 13011 14662
rect 12703 14651 13011 14660
rect 12990 14512 13046 14521
rect 12912 14470 12990 14498
rect 12912 14414 12940 14470
rect 12990 14447 13046 14456
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 12703 13628 13011 13637
rect 12703 13626 12709 13628
rect 12765 13626 12789 13628
rect 12845 13626 12869 13628
rect 12925 13626 12949 13628
rect 13005 13626 13011 13628
rect 12765 13574 12767 13626
rect 12947 13574 12949 13626
rect 12703 13572 12709 13574
rect 12765 13572 12789 13574
rect 12845 13572 12869 13574
rect 12925 13572 12949 13574
rect 13005 13572 13011 13574
rect 12703 13563 13011 13572
rect 13096 13297 13124 13806
rect 13280 13462 13308 16544
rect 13372 15042 13400 20878
rect 13464 18766 13492 22066
rect 13556 21554 13584 22222
rect 13648 21894 13676 23718
rect 13740 23225 13768 24074
rect 13832 23497 13860 25094
rect 13818 23488 13874 23497
rect 13818 23423 13874 23432
rect 13726 23216 13782 23225
rect 13726 23151 13782 23160
rect 13820 22500 13872 22506
rect 13820 22442 13872 22448
rect 13726 22264 13782 22273
rect 13726 22199 13782 22208
rect 13740 22098 13768 22199
rect 13832 22137 13860 22442
rect 13818 22128 13874 22137
rect 13728 22092 13780 22098
rect 13818 22063 13874 22072
rect 13728 22034 13780 22040
rect 13924 22001 13952 26846
rect 14004 26784 14056 26790
rect 14004 26726 14056 26732
rect 14016 26489 14044 26726
rect 14002 26480 14058 26489
rect 14002 26415 14058 26424
rect 14382 26140 14690 26149
rect 14382 26138 14388 26140
rect 14444 26138 14468 26140
rect 14524 26138 14548 26140
rect 14604 26138 14628 26140
rect 14684 26138 14690 26140
rect 14444 26086 14446 26138
rect 14626 26086 14628 26138
rect 14382 26084 14388 26086
rect 14444 26084 14468 26086
rect 14524 26084 14548 26086
rect 14604 26084 14628 26086
rect 14684 26084 14690 26086
rect 14382 26075 14690 26084
rect 14096 25424 14148 25430
rect 14096 25366 14148 25372
rect 14108 24886 14136 25366
rect 14188 25356 14240 25362
rect 14188 25298 14240 25304
rect 14200 25265 14228 25298
rect 14186 25256 14242 25265
rect 14186 25191 14242 25200
rect 14382 25052 14690 25061
rect 14382 25050 14388 25052
rect 14444 25050 14468 25052
rect 14524 25050 14548 25052
rect 14604 25050 14628 25052
rect 14684 25050 14690 25052
rect 14444 24998 14446 25050
rect 14626 24998 14628 25050
rect 14382 24996 14388 24998
rect 14444 24996 14468 24998
rect 14524 24996 14548 24998
rect 14604 24996 14628 24998
rect 14684 24996 14690 24998
rect 14382 24987 14690 24996
rect 14096 24880 14148 24886
rect 14002 24848 14058 24857
rect 14096 24822 14148 24828
rect 14002 24783 14058 24792
rect 14280 24812 14332 24818
rect 14016 24614 14044 24783
rect 14280 24754 14332 24760
rect 14004 24608 14056 24614
rect 14004 24550 14056 24556
rect 14002 24304 14058 24313
rect 14002 24239 14058 24248
rect 14016 23866 14044 24239
rect 14096 24200 14148 24206
rect 14096 24142 14148 24148
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 14108 23066 14136 24142
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14200 23866 14228 24006
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14292 23769 14320 24754
rect 14382 23964 14690 23973
rect 14382 23962 14388 23964
rect 14444 23962 14468 23964
rect 14524 23962 14548 23964
rect 14604 23962 14628 23964
rect 14684 23962 14690 23964
rect 14444 23910 14446 23962
rect 14626 23910 14628 23962
rect 14382 23908 14388 23910
rect 14444 23908 14468 23910
rect 14524 23908 14548 23910
rect 14604 23908 14628 23910
rect 14684 23908 14690 23910
rect 14382 23899 14690 23908
rect 14278 23760 14334 23769
rect 14278 23695 14334 23704
rect 14108 23038 14228 23066
rect 14004 22704 14056 22710
rect 14004 22646 14056 22652
rect 13910 21992 13966 22001
rect 13820 21956 13872 21962
rect 13910 21927 13966 21936
rect 13820 21898 13872 21904
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 13544 21548 13596 21554
rect 13544 21490 13596 21496
rect 13648 20482 13676 21626
rect 13726 21584 13782 21593
rect 13726 21519 13782 21528
rect 13740 20602 13768 21519
rect 13832 20777 13860 21898
rect 14016 21434 14044 22646
rect 13924 21406 14044 21434
rect 13818 20768 13874 20777
rect 13818 20703 13874 20712
rect 13728 20596 13780 20602
rect 13728 20538 13780 20544
rect 13648 20454 13860 20482
rect 13728 20392 13780 20398
rect 13728 20334 13780 20340
rect 13636 19916 13688 19922
rect 13556 19876 13636 19904
rect 13556 19378 13584 19876
rect 13636 19858 13688 19864
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13464 18465 13492 18702
rect 13544 18624 13596 18630
rect 13544 18566 13596 18572
rect 13450 18456 13506 18465
rect 13450 18391 13506 18400
rect 13450 18320 13506 18329
rect 13556 18290 13584 18566
rect 13450 18255 13452 18264
rect 13504 18255 13506 18264
rect 13544 18284 13596 18290
rect 13452 18226 13504 18232
rect 13544 18226 13596 18232
rect 13542 17368 13598 17377
rect 13542 17303 13598 17312
rect 13556 17270 13584 17303
rect 13544 17264 13596 17270
rect 13544 17206 13596 17212
rect 13452 16992 13504 16998
rect 13452 16934 13504 16940
rect 13464 16658 13492 16934
rect 13452 16652 13504 16658
rect 13648 16640 13676 19314
rect 13740 17338 13768 20334
rect 13832 19802 13860 20454
rect 13924 20058 13952 21406
rect 14096 21344 14148 21350
rect 14002 21312 14058 21321
rect 14096 21286 14148 21292
rect 14002 21247 14058 21256
rect 14016 21146 14044 21247
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 14108 21049 14136 21286
rect 14094 21040 14150 21049
rect 14094 20975 14150 20984
rect 14004 20868 14056 20874
rect 14004 20810 14056 20816
rect 14016 20346 14044 20810
rect 14200 20466 14228 23038
rect 14382 22876 14690 22885
rect 14382 22874 14388 22876
rect 14444 22874 14468 22876
rect 14524 22874 14548 22876
rect 14604 22874 14628 22876
rect 14684 22874 14690 22876
rect 14444 22822 14446 22874
rect 14626 22822 14628 22874
rect 14382 22820 14388 22822
rect 14444 22820 14468 22822
rect 14524 22820 14548 22822
rect 14604 22820 14628 22822
rect 14684 22820 14690 22822
rect 14382 22811 14690 22820
rect 14278 22672 14334 22681
rect 14278 22607 14334 22616
rect 14292 20942 14320 22607
rect 14382 21788 14690 21797
rect 14382 21786 14388 21788
rect 14444 21786 14468 21788
rect 14524 21786 14548 21788
rect 14604 21786 14628 21788
rect 14684 21786 14690 21788
rect 14444 21734 14446 21786
rect 14626 21734 14628 21786
rect 14382 21732 14388 21734
rect 14444 21732 14468 21734
rect 14524 21732 14548 21734
rect 14604 21732 14628 21734
rect 14684 21732 14690 21734
rect 14382 21723 14690 21732
rect 14280 20936 14332 20942
rect 14280 20878 14332 20884
rect 14382 20700 14690 20709
rect 14382 20698 14388 20700
rect 14444 20698 14468 20700
rect 14524 20698 14548 20700
rect 14604 20698 14628 20700
rect 14684 20698 14690 20700
rect 14444 20646 14446 20698
rect 14626 20646 14628 20698
rect 14382 20644 14388 20646
rect 14444 20644 14468 20646
rect 14524 20644 14548 20646
rect 14604 20644 14628 20646
rect 14684 20644 14690 20646
rect 14382 20635 14690 20644
rect 14188 20460 14240 20466
rect 14188 20402 14240 20408
rect 14016 20318 14320 20346
rect 14188 20256 14240 20262
rect 14094 20224 14150 20233
rect 14188 20198 14240 20204
rect 14094 20159 14150 20168
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 13832 19774 13952 19802
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13832 16794 13860 19654
rect 13924 18222 13952 19774
rect 14108 19514 14136 20159
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14096 19372 14148 19378
rect 14096 19314 14148 19320
rect 14002 19136 14058 19145
rect 14002 19071 14058 19080
rect 14016 18970 14044 19071
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 13912 18216 13964 18222
rect 13912 18158 13964 18164
rect 14004 17196 14056 17202
rect 14004 17138 14056 17144
rect 13912 17128 13964 17134
rect 13912 17070 13964 17076
rect 13820 16788 13872 16794
rect 13820 16730 13872 16736
rect 13648 16612 13768 16640
rect 13452 16594 13504 16600
rect 13634 16552 13690 16561
rect 13634 16487 13690 16496
rect 13372 15014 13492 15042
rect 13360 14952 13412 14958
rect 13360 14894 13412 14900
rect 13372 14074 13400 14894
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13372 13734 13400 13874
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13176 13456 13228 13462
rect 13176 13398 13228 13404
rect 13268 13456 13320 13462
rect 13268 13398 13320 13404
rect 13082 13288 13138 13297
rect 13188 13274 13216 13398
rect 13188 13246 13308 13274
rect 13082 13223 13138 13232
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12624 12776 12676 12782
rect 12544 12736 12624 12764
rect 12440 12640 12492 12646
rect 12440 12582 12492 12588
rect 12438 12472 12494 12481
rect 12438 12407 12494 12416
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12360 10810 12388 11562
rect 12452 11370 12480 12407
rect 12544 11529 12572 12736
rect 12728 12753 12756 12786
rect 12624 12718 12676 12724
rect 12714 12744 12770 12753
rect 12714 12679 12770 12688
rect 12992 12708 13044 12714
rect 13044 12668 13124 12696
rect 12992 12650 13044 12656
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12530 11520 12586 11529
rect 12530 11455 12586 11464
rect 12452 11342 12572 11370
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12346 10704 12402 10713
rect 12268 10662 12346 10690
rect 12164 9920 12216 9926
rect 12164 9862 12216 9868
rect 12164 9512 12216 9518
rect 12164 9454 12216 9460
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12176 8498 12204 9454
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11702 7440 11758 7449
rect 11702 7375 11758 7384
rect 11992 7342 12020 7482
rect 11980 7336 12032 7342
rect 11624 7262 11744 7290
rect 11980 7278 12032 7284
rect 12070 7304 12126 7313
rect 11612 7200 11664 7206
rect 11716 7188 11744 7262
rect 12070 7239 12126 7248
rect 11888 7200 11940 7206
rect 11716 7160 11888 7188
rect 11612 7142 11664 7148
rect 11888 7142 11940 7148
rect 11624 5778 11652 7142
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11702 6760 11758 6769
rect 11808 6730 11836 6870
rect 11702 6695 11758 6704
rect 11796 6724 11848 6730
rect 10744 5732 10824 5760
rect 11152 5772 11204 5778
rect 10692 5714 10744 5720
rect 11152 5714 11204 5720
rect 11336 5772 11388 5778
rect 11520 5772 11572 5778
rect 11388 5732 11468 5760
rect 11336 5714 11388 5720
rect 11024 5468 11332 5477
rect 11024 5466 11030 5468
rect 11086 5466 11110 5468
rect 11166 5466 11190 5468
rect 11246 5466 11270 5468
rect 11326 5466 11332 5468
rect 11086 5414 11088 5466
rect 11268 5414 11270 5466
rect 11024 5412 11030 5414
rect 11086 5412 11110 5414
rect 11166 5412 11190 5414
rect 11246 5412 11270 5414
rect 11326 5412 11332 5414
rect 11024 5403 11332 5412
rect 11440 4826 11468 5732
rect 11520 5714 11572 5720
rect 11612 5772 11664 5778
rect 11612 5714 11664 5720
rect 11244 4820 11296 4826
rect 11428 4820 11480 4826
rect 11296 4780 11376 4808
rect 11244 4762 11296 4768
rect 11348 4690 11376 4780
rect 11428 4762 11480 4768
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 10600 4616 10652 4622
rect 10600 4558 10652 4564
rect 11024 4380 11332 4389
rect 11024 4378 11030 4380
rect 11086 4378 11110 4380
rect 11166 4378 11190 4380
rect 11246 4378 11270 4380
rect 11326 4378 11332 4380
rect 11086 4326 11088 4378
rect 11268 4326 11270 4378
rect 11024 4324 11030 4326
rect 11086 4324 11110 4326
rect 11166 4324 11190 4326
rect 11246 4324 11270 4326
rect 11326 4324 11332 4326
rect 11024 4315 11332 4324
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 11716 4146 11744 6695
rect 11796 6666 11848 6672
rect 11900 6458 11928 7142
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 12084 6322 12112 7239
rect 12268 7206 12296 10662
rect 12346 10639 12402 10648
rect 12440 10600 12492 10606
rect 12346 10568 12402 10577
rect 12440 10542 12492 10548
rect 12346 10503 12402 10512
rect 12360 9926 12388 10503
rect 12452 10169 12480 10542
rect 12544 10470 12572 11342
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12438 10160 12494 10169
rect 12438 10095 12494 10104
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12360 9586 12388 9862
rect 12452 9722 12480 10095
rect 12440 9716 12492 9722
rect 12440 9658 12492 9664
rect 12438 9616 12494 9625
rect 12348 9580 12400 9586
rect 12438 9551 12494 9560
rect 12348 9522 12400 9528
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12254 6352 12310 6361
rect 12072 6316 12124 6322
rect 12254 6287 12310 6296
rect 12072 6258 12124 6264
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11808 5370 11836 5646
rect 11796 5364 11848 5370
rect 11796 5306 11848 5312
rect 11978 5128 12034 5137
rect 11978 5063 12034 5072
rect 11992 4622 12020 5063
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 12268 4434 12296 6287
rect 12346 5808 12402 5817
rect 12452 5778 12480 9551
rect 12544 9042 12572 10406
rect 12636 9518 12664 12582
rect 12703 12540 13011 12549
rect 12703 12538 12709 12540
rect 12765 12538 12789 12540
rect 12845 12538 12869 12540
rect 12925 12538 12949 12540
rect 13005 12538 13011 12540
rect 12765 12486 12767 12538
rect 12947 12486 12949 12538
rect 12703 12484 12709 12486
rect 12765 12484 12789 12486
rect 12845 12484 12869 12486
rect 12925 12484 12949 12486
rect 13005 12484 13011 12486
rect 12703 12475 13011 12484
rect 13096 12442 13124 12668
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 12703 11452 13011 11461
rect 12703 11450 12709 11452
rect 12765 11450 12789 11452
rect 12845 11450 12869 11452
rect 12925 11450 12949 11452
rect 13005 11450 13011 11452
rect 12765 11398 12767 11450
rect 12947 11398 12949 11450
rect 12703 11396 12709 11398
rect 12765 11396 12789 11398
rect 12845 11396 12869 11398
rect 12925 11396 12949 11398
rect 13005 11396 13011 11398
rect 12703 11387 13011 11396
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12716 11144 12768 11150
rect 12714 11112 12716 11121
rect 12768 11112 12770 11121
rect 12714 11047 12770 11056
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10606 12940 10950
rect 13084 10804 13136 10810
rect 13084 10746 13136 10752
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12703 10364 13011 10373
rect 12703 10362 12709 10364
rect 12765 10362 12789 10364
rect 12845 10362 12869 10364
rect 12925 10362 12949 10364
rect 13005 10362 13011 10364
rect 12765 10310 12767 10362
rect 12947 10310 12949 10362
rect 12703 10308 12709 10310
rect 12765 10308 12789 10310
rect 12845 10308 12869 10310
rect 12925 10308 12949 10310
rect 13005 10308 13011 10310
rect 12703 10299 13011 10308
rect 13096 9625 13124 10746
rect 13082 9616 13138 9625
rect 13082 9551 13138 9560
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 13084 9444 13136 9450
rect 13084 9386 13136 9392
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12636 9110 12664 9318
rect 12703 9276 13011 9285
rect 12703 9274 12709 9276
rect 12765 9274 12789 9276
rect 12845 9274 12869 9276
rect 12925 9274 12949 9276
rect 13005 9274 13011 9276
rect 12765 9222 12767 9274
rect 12947 9222 12949 9274
rect 12703 9220 12709 9222
rect 12765 9220 12789 9222
rect 12845 9220 12869 9222
rect 12925 9220 12949 9222
rect 13005 9220 13011 9222
rect 12703 9211 13011 9220
rect 12624 9104 12676 9110
rect 12624 9046 12676 9052
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12624 8968 12676 8974
rect 12624 8910 12676 8916
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8498 12572 8774
rect 12636 8566 12664 8910
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 7954 12572 8434
rect 12703 8188 13011 8197
rect 12703 8186 12709 8188
rect 12765 8186 12789 8188
rect 12845 8186 12869 8188
rect 12925 8186 12949 8188
rect 13005 8186 13011 8188
rect 12765 8134 12767 8186
rect 12947 8134 12949 8186
rect 12703 8132 12709 8134
rect 12765 8132 12789 8134
rect 12845 8132 12869 8134
rect 12925 8132 12949 8134
rect 13005 8132 13011 8134
rect 12703 8123 13011 8132
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12544 7546 12572 7890
rect 13096 7546 13124 9386
rect 13188 8838 13216 11290
rect 13280 10674 13308 13246
rect 13372 10674 13400 13670
rect 13464 13530 13492 15014
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13556 14618 13584 14894
rect 13544 14612 13596 14618
rect 13544 14554 13596 14560
rect 13452 13524 13504 13530
rect 13452 13466 13504 13472
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13544 12776 13596 12782
rect 13544 12718 13596 12724
rect 13464 12209 13492 12718
rect 13450 12200 13506 12209
rect 13450 12135 13506 12144
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13360 10668 13412 10674
rect 13360 10610 13412 10616
rect 13266 9752 13322 9761
rect 13322 9710 13400 9738
rect 13266 9687 13322 9696
rect 13266 9616 13322 9625
rect 13266 9551 13322 9560
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13280 8378 13308 9551
rect 13188 8350 13308 8378
rect 13188 7750 13216 8350
rect 13268 7880 13320 7886
rect 13268 7822 13320 7828
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 12703 7100 13011 7109
rect 12703 7098 12709 7100
rect 12765 7098 12789 7100
rect 12845 7098 12869 7100
rect 12925 7098 12949 7100
rect 13005 7098 13011 7100
rect 12765 7046 12767 7098
rect 12947 7046 12949 7098
rect 12703 7044 12709 7046
rect 12765 7044 12789 7046
rect 12845 7044 12869 7046
rect 12925 7044 12949 7046
rect 13005 7044 13011 7046
rect 12703 7035 13011 7044
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12530 6216 12586 6225
rect 12530 6151 12586 6160
rect 12544 5930 12572 6151
rect 12636 6118 12664 6598
rect 13188 6440 13216 7482
rect 13096 6412 13216 6440
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12703 6012 13011 6021
rect 12703 6010 12709 6012
rect 12765 6010 12789 6012
rect 12845 6010 12869 6012
rect 12925 6010 12949 6012
rect 13005 6010 13011 6012
rect 12765 5958 12767 6010
rect 12947 5958 12949 6010
rect 12703 5956 12709 5958
rect 12765 5956 12789 5958
rect 12845 5956 12869 5958
rect 12925 5956 12949 5958
rect 13005 5956 13011 5958
rect 12703 5947 13011 5956
rect 12544 5902 12664 5930
rect 12346 5743 12402 5752
rect 12440 5772 12492 5778
rect 12360 4554 12388 5743
rect 12440 5714 12492 5720
rect 12636 5692 12664 5902
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12808 5704 12860 5710
rect 12438 5672 12494 5681
rect 12636 5664 12808 5692
rect 12808 5646 12860 5652
rect 12438 5607 12440 5616
rect 12492 5607 12494 5616
rect 12440 5578 12492 5584
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12728 5166 12756 5510
rect 12716 5160 12768 5166
rect 12636 5120 12716 5148
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 4826 12572 4966
rect 12532 4820 12584 4826
rect 12532 4762 12584 4768
rect 12636 4622 12664 5120
rect 12716 5102 12768 5108
rect 12912 5030 12940 5850
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12703 4924 13011 4933
rect 12703 4922 12709 4924
rect 12765 4922 12789 4924
rect 12845 4922 12869 4924
rect 12925 4922 12949 4924
rect 13005 4922 13011 4924
rect 12765 4870 12767 4922
rect 12947 4870 12949 4922
rect 12703 4868 12709 4870
rect 12765 4868 12789 4870
rect 12845 4868 12869 4870
rect 12925 4868 12949 4870
rect 13005 4868 13011 4870
rect 12703 4859 13011 4868
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12348 4548 12400 4554
rect 12348 4490 12400 4496
rect 12532 4548 12584 4554
rect 12532 4490 12584 4496
rect 12268 4406 12388 4434
rect 12360 4214 12388 4406
rect 12544 4282 12572 4490
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12348 4208 12400 4214
rect 12348 4150 12400 4156
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 9345 3836 9653 3845
rect 9345 3834 9351 3836
rect 9407 3834 9431 3836
rect 9487 3834 9511 3836
rect 9567 3834 9591 3836
rect 9647 3834 9653 3836
rect 9407 3782 9409 3834
rect 9589 3782 9591 3834
rect 9345 3780 9351 3782
rect 9407 3780 9431 3782
rect 9487 3780 9511 3782
rect 9567 3780 9591 3782
rect 9647 3780 9653 3782
rect 9345 3771 9653 3780
rect 12703 3836 13011 3845
rect 12703 3834 12709 3836
rect 12765 3834 12789 3836
rect 12845 3834 12869 3836
rect 12925 3834 12949 3836
rect 13005 3834 13011 3836
rect 12765 3782 12767 3834
rect 12947 3782 12949 3834
rect 12703 3780 12709 3782
rect 12765 3780 12789 3782
rect 12845 3780 12869 3782
rect 12925 3780 12949 3782
rect 13005 3780 13011 3782
rect 12703 3771 13011 3780
rect 11024 3292 11332 3301
rect 11024 3290 11030 3292
rect 11086 3290 11110 3292
rect 11166 3290 11190 3292
rect 11246 3290 11270 3292
rect 11326 3290 11332 3292
rect 11086 3238 11088 3290
rect 11268 3238 11270 3290
rect 11024 3236 11030 3238
rect 11086 3236 11110 3238
rect 11166 3236 11190 3238
rect 11246 3236 11270 3238
rect 11326 3236 11332 3238
rect 11024 3227 11332 3236
rect 13096 2854 13124 6412
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13188 5370 13216 6258
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13280 4622 13308 7822
rect 13372 6848 13400 9710
rect 13464 9586 13492 12038
rect 13556 11898 13584 12718
rect 13648 12102 13676 16487
rect 13740 15484 13768 16612
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 15609 13860 16390
rect 13924 15706 13952 17070
rect 14016 16697 14044 17138
rect 14002 16688 14058 16697
rect 14002 16623 14058 16632
rect 13912 15700 13964 15706
rect 13912 15642 13964 15648
rect 13818 15600 13874 15609
rect 13818 15535 13874 15544
rect 13740 15456 14044 15484
rect 13820 15360 13872 15366
rect 13726 15328 13782 15337
rect 13820 15302 13872 15308
rect 13726 15263 13782 15272
rect 13740 13258 13768 15263
rect 13832 14482 13860 15302
rect 13910 15056 13966 15065
rect 13910 14991 13966 15000
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13924 14006 13952 14991
rect 13912 14000 13964 14006
rect 13912 13942 13964 13948
rect 14016 13852 14044 15456
rect 14108 15201 14136 19314
rect 14094 15192 14150 15201
rect 14094 15127 14150 15136
rect 14094 13968 14150 13977
rect 14094 13903 14150 13912
rect 13924 13824 14044 13852
rect 13728 13252 13780 13258
rect 13728 13194 13780 13200
rect 13726 12472 13782 12481
rect 13726 12407 13782 12416
rect 13740 12238 13768 12407
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13726 12064 13782 12073
rect 13726 11999 13782 12008
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13544 10600 13596 10606
rect 13544 10542 13596 10548
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13556 8634 13584 10542
rect 13634 9888 13690 9897
rect 13634 9823 13690 9832
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13648 8498 13676 9823
rect 13740 9625 13768 11999
rect 13820 9716 13872 9722
rect 13820 9658 13872 9664
rect 13726 9616 13782 9625
rect 13726 9551 13782 9560
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13740 8090 13768 9454
rect 13832 9178 13860 9658
rect 13820 9172 13872 9178
rect 13820 9114 13872 9120
rect 13924 9042 13952 13824
rect 14002 13424 14058 13433
rect 14002 13359 14058 13368
rect 14016 12986 14044 13359
rect 14004 12980 14056 12986
rect 14004 12922 14056 12928
rect 14108 12434 14136 13903
rect 14016 12406 14136 12434
rect 14016 11762 14044 12406
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 14004 10464 14056 10470
rect 14004 10406 14056 10412
rect 14094 10432 14150 10441
rect 14016 10169 14044 10406
rect 14094 10367 14150 10376
rect 14002 10160 14058 10169
rect 14108 10130 14136 10367
rect 14002 10095 14058 10104
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14200 9654 14228 20198
rect 14292 10810 14320 20318
rect 14382 19612 14690 19621
rect 14382 19610 14388 19612
rect 14444 19610 14468 19612
rect 14524 19610 14548 19612
rect 14604 19610 14628 19612
rect 14684 19610 14690 19612
rect 14444 19558 14446 19610
rect 14626 19558 14628 19610
rect 14382 19556 14388 19558
rect 14444 19556 14468 19558
rect 14524 19556 14548 19558
rect 14604 19556 14628 19558
rect 14684 19556 14690 19558
rect 14382 19547 14690 19556
rect 14370 19272 14426 19281
rect 14370 19207 14426 19216
rect 14384 18766 14412 19207
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14382 18524 14690 18533
rect 14382 18522 14388 18524
rect 14444 18522 14468 18524
rect 14524 18522 14548 18524
rect 14604 18522 14628 18524
rect 14684 18522 14690 18524
rect 14444 18470 14446 18522
rect 14626 18470 14628 18522
rect 14382 18468 14388 18470
rect 14444 18468 14468 18470
rect 14524 18468 14548 18470
rect 14604 18468 14628 18470
rect 14684 18468 14690 18470
rect 14382 18459 14690 18468
rect 14382 17436 14690 17445
rect 14382 17434 14388 17436
rect 14444 17434 14468 17436
rect 14524 17434 14548 17436
rect 14604 17434 14628 17436
rect 14684 17434 14690 17436
rect 14444 17382 14446 17434
rect 14626 17382 14628 17434
rect 14382 17380 14388 17382
rect 14444 17380 14468 17382
rect 14524 17380 14548 17382
rect 14604 17380 14628 17382
rect 14684 17380 14690 17382
rect 14382 17371 14690 17380
rect 14382 16348 14690 16357
rect 14382 16346 14388 16348
rect 14444 16346 14468 16348
rect 14524 16346 14548 16348
rect 14604 16346 14628 16348
rect 14684 16346 14690 16348
rect 14444 16294 14446 16346
rect 14626 16294 14628 16346
rect 14382 16292 14388 16294
rect 14444 16292 14468 16294
rect 14524 16292 14548 16294
rect 14604 16292 14628 16294
rect 14684 16292 14690 16294
rect 14382 16283 14690 16292
rect 14646 16144 14702 16153
rect 14646 16079 14702 16088
rect 14660 15502 14688 16079
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14382 15260 14690 15269
rect 14382 15258 14388 15260
rect 14444 15258 14468 15260
rect 14524 15258 14548 15260
rect 14604 15258 14628 15260
rect 14684 15258 14690 15260
rect 14444 15206 14446 15258
rect 14626 15206 14628 15258
rect 14382 15204 14388 15206
rect 14444 15204 14468 15206
rect 14524 15204 14548 15206
rect 14604 15204 14628 15206
rect 14684 15204 14690 15206
rect 14382 15195 14690 15204
rect 14372 14816 14424 14822
rect 14370 14784 14372 14793
rect 14424 14784 14426 14793
rect 14370 14719 14426 14728
rect 14382 14172 14690 14181
rect 14382 14170 14388 14172
rect 14444 14170 14468 14172
rect 14524 14170 14548 14172
rect 14604 14170 14628 14172
rect 14684 14170 14690 14172
rect 14444 14118 14446 14170
rect 14626 14118 14628 14170
rect 14382 14116 14388 14118
rect 14444 14116 14468 14118
rect 14524 14116 14548 14118
rect 14604 14116 14628 14118
rect 14684 14116 14690 14118
rect 14382 14107 14690 14116
rect 14370 13696 14426 13705
rect 14370 13631 14426 13640
rect 14384 13326 14412 13631
rect 14372 13320 14424 13326
rect 14372 13262 14424 13268
rect 14382 13084 14690 13093
rect 14382 13082 14388 13084
rect 14444 13082 14468 13084
rect 14524 13082 14548 13084
rect 14604 13082 14628 13084
rect 14684 13082 14690 13084
rect 14444 13030 14446 13082
rect 14626 13030 14628 13082
rect 14382 13028 14388 13030
rect 14444 13028 14468 13030
rect 14524 13028 14548 13030
rect 14604 13028 14628 13030
rect 14684 13028 14690 13030
rect 14382 13019 14690 13028
rect 14382 11996 14690 12005
rect 14382 11994 14388 11996
rect 14444 11994 14468 11996
rect 14524 11994 14548 11996
rect 14604 11994 14628 11996
rect 14684 11994 14690 11996
rect 14444 11942 14446 11994
rect 14626 11942 14628 11994
rect 14382 11940 14388 11942
rect 14444 11940 14468 11942
rect 14524 11940 14548 11942
rect 14604 11940 14628 11942
rect 14684 11940 14690 11942
rect 14382 11931 14690 11940
rect 14382 10908 14690 10917
rect 14382 10906 14388 10908
rect 14444 10906 14468 10908
rect 14524 10906 14548 10908
rect 14604 10906 14628 10908
rect 14684 10906 14690 10908
rect 14444 10854 14446 10906
rect 14626 10854 14628 10906
rect 14382 10852 14388 10854
rect 14444 10852 14468 10854
rect 14524 10852 14548 10854
rect 14604 10852 14628 10854
rect 14684 10852 14690 10854
rect 14382 10843 14690 10852
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14382 9820 14690 9829
rect 14382 9818 14388 9820
rect 14444 9818 14468 9820
rect 14524 9818 14548 9820
rect 14604 9818 14628 9820
rect 14684 9818 14690 9820
rect 14444 9766 14446 9818
rect 14626 9766 14628 9818
rect 14382 9764 14388 9766
rect 14444 9764 14468 9766
rect 14524 9764 14548 9766
rect 14604 9764 14628 9766
rect 14684 9764 14690 9766
rect 14382 9755 14690 9764
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14004 9376 14056 9382
rect 14002 9344 14004 9353
rect 14056 9344 14058 9353
rect 14002 9279 14058 9288
rect 14752 9194 14780 36094
rect 14292 9166 14780 9194
rect 13912 9036 13964 9042
rect 13912 8978 13964 8984
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 14200 8537 14228 8842
rect 14186 8528 14242 8537
rect 14186 8463 14242 8472
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13648 7410 13676 7754
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13740 7154 13768 7686
rect 14292 7546 14320 9166
rect 14844 9058 14872 36502
rect 15028 36009 15056 36722
rect 15014 36000 15070 36009
rect 15014 35935 15070 35944
rect 14924 34604 14976 34610
rect 14924 34546 14976 34552
rect 14936 30297 14964 34546
rect 15016 33312 15068 33318
rect 15016 33254 15068 33260
rect 14922 30288 14978 30297
rect 14922 30223 14978 30232
rect 14924 29844 14976 29850
rect 14924 29786 14976 29792
rect 14936 23089 14964 29786
rect 15028 29753 15056 33254
rect 15108 32428 15160 32434
rect 15108 32370 15160 32376
rect 15014 29744 15070 29753
rect 15014 29679 15070 29688
rect 15016 28620 15068 28626
rect 15016 28562 15068 28568
rect 15028 26217 15056 28562
rect 15014 26208 15070 26217
rect 15014 26143 15070 26152
rect 15016 24880 15068 24886
rect 15016 24822 15068 24828
rect 14922 23080 14978 23089
rect 14922 23015 14978 23024
rect 14922 22944 14978 22953
rect 14922 22879 14978 22888
rect 14936 22778 14964 22879
rect 14924 22772 14976 22778
rect 14924 22714 14976 22720
rect 14924 22568 14976 22574
rect 14924 22510 14976 22516
rect 14936 12434 14964 22510
rect 15028 21146 15056 24822
rect 15016 21140 15068 21146
rect 15016 21082 15068 21088
rect 15016 21004 15068 21010
rect 15016 20946 15068 20952
rect 15028 20777 15056 20946
rect 15014 20768 15070 20777
rect 15014 20703 15070 20712
rect 15014 18592 15070 18601
rect 15014 18527 15070 18536
rect 15028 18426 15056 18527
rect 15016 18420 15068 18426
rect 15016 18362 15068 18368
rect 15014 17232 15070 17241
rect 15014 17167 15070 17176
rect 15028 16833 15056 17167
rect 15014 16824 15070 16833
rect 15014 16759 15070 16768
rect 15014 16416 15070 16425
rect 15014 16351 15070 16360
rect 15028 16182 15056 16351
rect 15016 16176 15068 16182
rect 15016 16118 15068 16124
rect 15016 14340 15068 14346
rect 15016 14282 15068 14288
rect 15028 14249 15056 14282
rect 15014 14240 15070 14249
rect 15014 14175 15070 14184
rect 14936 12406 15056 12434
rect 14752 9030 14872 9058
rect 14382 8732 14690 8741
rect 14382 8730 14388 8732
rect 14444 8730 14468 8732
rect 14524 8730 14548 8732
rect 14604 8730 14628 8732
rect 14684 8730 14690 8732
rect 14444 8678 14446 8730
rect 14626 8678 14628 8730
rect 14382 8676 14388 8678
rect 14444 8676 14468 8678
rect 14524 8676 14548 8678
rect 14604 8676 14628 8678
rect 14684 8676 14690 8678
rect 14382 8667 14690 8676
rect 14382 7644 14690 7653
rect 14382 7642 14388 7644
rect 14444 7642 14468 7644
rect 14524 7642 14548 7644
rect 14604 7642 14628 7644
rect 14684 7642 14690 7644
rect 14444 7590 14446 7642
rect 14626 7590 14628 7642
rect 14382 7588 14388 7590
rect 14444 7588 14468 7590
rect 14524 7588 14548 7590
rect 14604 7588 14628 7590
rect 14684 7588 14690 7590
rect 14382 7579 14690 7588
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 13740 7126 13860 7154
rect 13372 6820 13492 6848
rect 13464 6730 13492 6820
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13452 6724 13504 6730
rect 13504 6684 13584 6712
rect 13452 6666 13504 6672
rect 13372 4826 13400 6666
rect 13450 6488 13506 6497
rect 13450 6423 13506 6432
rect 13464 6390 13492 6423
rect 13452 6384 13504 6390
rect 13452 6326 13504 6332
rect 13556 5828 13584 6684
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13648 5914 13676 6326
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 13464 5800 13584 5828
rect 13360 4820 13412 4826
rect 13360 4762 13412 4768
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13464 4146 13492 5800
rect 13740 5710 13768 6258
rect 13728 5704 13780 5710
rect 13634 5672 13690 5681
rect 13728 5646 13780 5652
rect 13634 5607 13690 5616
rect 13648 4146 13676 5607
rect 13726 5264 13782 5273
rect 13726 5199 13782 5208
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13740 3534 13768 5199
rect 13832 3942 13860 7126
rect 14382 6556 14690 6565
rect 14382 6554 14388 6556
rect 14444 6554 14468 6556
rect 14524 6554 14548 6556
rect 14604 6554 14628 6556
rect 14684 6554 14690 6556
rect 14444 6502 14446 6554
rect 14626 6502 14628 6554
rect 14382 6500 14388 6502
rect 14444 6500 14468 6502
rect 14524 6500 14548 6502
rect 14604 6500 14628 6502
rect 14684 6500 14690 6502
rect 14382 6491 14690 6500
rect 14382 5468 14690 5477
rect 14382 5466 14388 5468
rect 14444 5466 14468 5468
rect 14524 5466 14548 5468
rect 14604 5466 14628 5468
rect 14684 5466 14690 5468
rect 14444 5414 14446 5466
rect 14626 5414 14628 5466
rect 14382 5412 14388 5414
rect 14444 5412 14468 5414
rect 14524 5412 14548 5414
rect 14604 5412 14628 5414
rect 14684 5412 14690 5414
rect 14382 5403 14690 5412
rect 13910 4992 13966 5001
rect 13910 4927 13966 4936
rect 13924 4214 13952 4927
rect 14382 4380 14690 4389
rect 14382 4378 14388 4380
rect 14444 4378 14468 4380
rect 14524 4378 14548 4380
rect 14604 4378 14628 4380
rect 14684 4378 14690 4380
rect 14444 4326 14446 4378
rect 14626 4326 14628 4378
rect 14382 4324 14388 4326
rect 14444 4324 14468 4326
rect 14524 4324 14548 4326
rect 14604 4324 14628 4326
rect 14684 4324 14690 4326
rect 14382 4315 14690 4324
rect 13912 4208 13964 4214
rect 13912 4150 13964 4156
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 14382 3292 14690 3301
rect 14382 3290 14388 3292
rect 14444 3290 14468 3292
rect 14524 3290 14548 3292
rect 14604 3290 14628 3292
rect 14684 3290 14690 3292
rect 14444 3238 14446 3290
rect 14626 3238 14628 3290
rect 14382 3236 14388 3238
rect 14444 3236 14468 3238
rect 14524 3236 14548 3238
rect 14604 3236 14628 3238
rect 14684 3236 14690 3238
rect 14382 3227 14690 3236
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 9345 2748 9653 2757
rect 9345 2746 9351 2748
rect 9407 2746 9431 2748
rect 9487 2746 9511 2748
rect 9567 2746 9591 2748
rect 9647 2746 9653 2748
rect 9407 2694 9409 2746
rect 9589 2694 9591 2746
rect 9345 2692 9351 2694
rect 9407 2692 9431 2694
rect 9487 2692 9511 2694
rect 9567 2692 9591 2694
rect 9647 2692 9653 2694
rect 9345 2683 9653 2692
rect 12703 2748 13011 2757
rect 12703 2746 12709 2748
rect 12765 2746 12789 2748
rect 12845 2746 12869 2748
rect 12925 2746 12949 2748
rect 13005 2746 13011 2748
rect 12765 2694 12767 2746
rect 12947 2694 12949 2746
rect 12703 2692 12709 2694
rect 12765 2692 12789 2694
rect 12845 2692 12869 2694
rect 12925 2692 12949 2694
rect 13005 2692 13011 2694
rect 10874 2680 10930 2689
rect 12703 2683 13011 2692
rect 10874 2615 10930 2624
rect 9402 2544 9458 2553
rect 9402 2479 9458 2488
rect 9416 2106 9444 2479
rect 10888 2106 10916 2615
rect 11024 2204 11332 2213
rect 11024 2202 11030 2204
rect 11086 2202 11110 2204
rect 11166 2202 11190 2204
rect 11246 2202 11270 2204
rect 11326 2202 11332 2204
rect 11086 2150 11088 2202
rect 11268 2150 11270 2202
rect 11024 2148 11030 2150
rect 11086 2148 11110 2150
rect 11166 2148 11190 2150
rect 11246 2148 11270 2150
rect 11326 2148 11332 2150
rect 11024 2139 11332 2148
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 10140 2100 10192 2106
rect 10140 2042 10192 2048
rect 10876 2100 10928 2106
rect 13372 2088 13400 2790
rect 14382 2204 14690 2213
rect 14382 2202 14388 2204
rect 14444 2202 14468 2204
rect 14524 2202 14548 2204
rect 14604 2202 14628 2204
rect 14684 2202 14690 2204
rect 14444 2150 14446 2202
rect 14626 2150 14628 2202
rect 14382 2148 14388 2150
rect 14444 2148 14468 2150
rect 14524 2148 14548 2150
rect 14604 2148 14628 2150
rect 14684 2148 14690 2150
rect 14382 2139 14690 2148
rect 13452 2100 13504 2106
rect 13372 2060 13452 2088
rect 10876 2042 10928 2048
rect 13452 2042 13504 2048
rect 10152 2009 10180 2042
rect 10138 2000 10194 2009
rect 9220 1964 9272 1970
rect 9220 1906 9272 1912
rect 10048 1964 10100 1970
rect 10138 1935 10194 1944
rect 10784 1964 10836 1970
rect 10048 1906 10100 1912
rect 10784 1906 10836 1912
rect 11612 1964 11664 1970
rect 11612 1906 11664 1912
rect 12256 1964 12308 1970
rect 12256 1906 12308 1912
rect 13084 1964 13136 1970
rect 13084 1906 13136 1912
rect 13728 1964 13780 1970
rect 13728 1906 13780 1912
rect 14188 1964 14240 1970
rect 14188 1906 14240 1912
rect 9232 1562 9260 1906
rect 9345 1660 9653 1669
rect 9345 1658 9351 1660
rect 9407 1658 9431 1660
rect 9487 1658 9511 1660
rect 9567 1658 9591 1660
rect 9647 1658 9653 1660
rect 9407 1606 9409 1658
rect 9589 1606 9591 1658
rect 9345 1604 9351 1606
rect 9407 1604 9431 1606
rect 9487 1604 9511 1606
rect 9567 1604 9591 1606
rect 9647 1604 9653 1606
rect 9345 1595 9653 1604
rect 10060 1562 10088 1906
rect 10796 1562 10824 1906
rect 11624 1562 11652 1906
rect 12268 1562 12296 1906
rect 12703 1660 13011 1669
rect 12703 1658 12709 1660
rect 12765 1658 12789 1660
rect 12845 1658 12869 1660
rect 12925 1658 12949 1660
rect 13005 1658 13011 1660
rect 12765 1606 12767 1658
rect 12947 1606 12949 1658
rect 12703 1604 12709 1606
rect 12765 1604 12789 1606
rect 12845 1604 12869 1606
rect 12925 1604 12949 1606
rect 13005 1604 13011 1606
rect 12703 1595 13011 1604
rect 13096 1562 13124 1906
rect 13740 1562 13768 1906
rect 9220 1556 9272 1562
rect 9220 1498 9272 1504
rect 10048 1556 10100 1562
rect 10048 1498 10100 1504
rect 10784 1556 10836 1562
rect 10784 1498 10836 1504
rect 11612 1556 11664 1562
rect 11612 1498 11664 1504
rect 12256 1556 12308 1562
rect 12256 1498 12308 1504
rect 13084 1556 13136 1562
rect 13084 1498 13136 1504
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 9128 1488 9180 1494
rect 9128 1430 9180 1436
rect 2504 1352 2556 1358
rect 2504 1294 2556 1300
rect 2688 1352 2740 1358
rect 2688 1294 2740 1300
rect 3792 1352 3844 1358
rect 4620 1352 4672 1358
rect 3792 1294 3844 1300
rect 4618 1320 4620 1329
rect 5172 1352 5224 1358
rect 4672 1320 4674 1329
rect 2320 1284 2372 1290
rect 2320 1226 2372 1232
rect 2700 160 2728 1294
rect 478 -300 534 160
rect 1214 -300 1270 160
rect 1950 -300 2006 160
rect 2686 -300 2742 160
rect 3422 82 3478 160
rect 3804 82 3832 1294
rect 4160 1284 4212 1290
rect 5170 1320 5172 1329
rect 6184 1352 6236 1358
rect 5224 1320 5226 1329
rect 4618 1255 4674 1264
rect 5080 1284 5132 1290
rect 4160 1226 4212 1232
rect 6644 1352 6696 1358
rect 6184 1294 6236 1300
rect 6642 1320 6644 1329
rect 7104 1352 7156 1358
rect 6696 1320 6698 1329
rect 5170 1255 5226 1264
rect 5632 1284 5684 1290
rect 5080 1226 5132 1232
rect 5632 1226 5684 1232
rect 4172 160 4200 1226
rect 4308 1116 4616 1125
rect 4308 1114 4314 1116
rect 4370 1114 4394 1116
rect 4450 1114 4474 1116
rect 4530 1114 4554 1116
rect 4610 1114 4616 1116
rect 4370 1062 4372 1114
rect 4552 1062 4554 1114
rect 4308 1060 4314 1062
rect 4370 1060 4394 1062
rect 4450 1060 4474 1062
rect 4530 1060 4554 1062
rect 4610 1060 4616 1062
rect 4308 1051 4616 1060
rect 3422 54 3832 82
rect 3422 -300 3478 54
rect 4158 -300 4214 160
rect 4894 82 4950 160
rect 5092 82 5120 1226
rect 5644 160 5672 1226
rect 4894 54 5120 82
rect 4894 -300 4950 54
rect 5630 -300 5686 160
rect 6196 82 6224 1294
rect 7104 1294 7156 1300
rect 8116 1352 8168 1358
rect 8116 1294 8168 1300
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 9312 1352 9364 1358
rect 9312 1294 9364 1300
rect 10048 1352 10100 1358
rect 10048 1294 10100 1300
rect 10784 1352 10836 1358
rect 10784 1294 10836 1300
rect 11520 1352 11572 1358
rect 11520 1294 11572 1300
rect 12256 1352 12308 1358
rect 12256 1294 12308 1300
rect 13268 1352 13320 1358
rect 13268 1294 13320 1300
rect 13544 1352 13596 1358
rect 13596 1312 13768 1340
rect 13544 1294 13596 1300
rect 6642 1255 6698 1264
rect 7116 160 7144 1294
rect 7666 1116 7974 1125
rect 7666 1114 7672 1116
rect 7728 1114 7752 1116
rect 7808 1114 7832 1116
rect 7888 1114 7912 1116
rect 7968 1114 7974 1116
rect 7728 1062 7730 1114
rect 7910 1062 7912 1114
rect 7666 1060 7672 1062
rect 7728 1060 7752 1062
rect 7808 1060 7832 1062
rect 7888 1060 7912 1062
rect 7968 1060 7974 1062
rect 7666 1051 7974 1060
rect 7852 190 7972 218
rect 7852 160 7880 190
rect 6366 82 6422 160
rect 6196 54 6422 82
rect 6366 -300 6422 54
rect 7102 -300 7158 160
rect 7838 -300 7894 160
rect 7944 82 7972 190
rect 8128 82 8156 1294
rect 8588 160 8616 1294
rect 9324 160 9352 1294
rect 10060 160 10088 1294
rect 10796 160 10824 1294
rect 11024 1116 11332 1125
rect 11024 1114 11030 1116
rect 11086 1114 11110 1116
rect 11166 1114 11190 1116
rect 11246 1114 11270 1116
rect 11326 1114 11332 1116
rect 11086 1062 11088 1114
rect 11268 1062 11270 1114
rect 11024 1060 11030 1062
rect 11086 1060 11110 1062
rect 11166 1060 11190 1062
rect 11246 1060 11270 1062
rect 11326 1060 11332 1062
rect 11024 1051 11332 1060
rect 11532 160 11560 1294
rect 12268 160 12296 1294
rect 13004 190 13124 218
rect 13004 160 13032 190
rect 7944 54 8156 82
rect 8574 -300 8630 160
rect 9310 -300 9366 160
rect 10046 -300 10102 160
rect 10782 -300 10838 160
rect 11518 -300 11574 160
rect 12254 -300 12310 160
rect 12990 -300 13046 160
rect 13096 82 13124 190
rect 13280 82 13308 1294
rect 13740 160 13768 1312
rect 13818 1320 13874 1329
rect 13818 1255 13874 1264
rect 13832 1222 13860 1255
rect 13820 1216 13872 1222
rect 13820 1158 13872 1164
rect 13096 54 13308 82
rect 13726 -300 13782 160
rect 14200 82 14228 1906
rect 14752 1902 14780 9030
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8809 14872 8910
rect 14830 8800 14886 8809
rect 14830 8735 14886 8744
rect 14830 7712 14886 7721
rect 14830 7647 14886 7656
rect 14844 7478 14872 7647
rect 14832 7472 14884 7478
rect 14832 7414 14884 7420
rect 15028 6662 15056 12406
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15120 6458 15148 32370
rect 15200 32224 15252 32230
rect 15200 32166 15252 32172
rect 15304 32178 15332 41386
rect 15212 27305 15240 32166
rect 15304 32150 15516 32178
rect 15384 32020 15436 32026
rect 15384 31962 15436 31968
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15198 27296 15254 27305
rect 15198 27231 15254 27240
rect 15304 25650 15332 31758
rect 15396 28665 15424 31962
rect 15488 31396 15516 32150
rect 15580 31754 15608 42502
rect 15568 31748 15620 31754
rect 15568 31690 15620 31696
rect 15488 31368 15700 31396
rect 15568 31136 15620 31142
rect 15568 31078 15620 31084
rect 15476 30660 15528 30666
rect 15476 30602 15528 30608
rect 15382 28656 15438 28665
rect 15382 28591 15438 28600
rect 15382 27568 15438 27577
rect 15488 27554 15516 30602
rect 15438 27526 15516 27554
rect 15382 27503 15438 27512
rect 15304 25622 15424 25650
rect 15396 25378 15424 25622
rect 15304 25350 15424 25378
rect 15200 24812 15252 24818
rect 15200 24754 15252 24760
rect 15212 22982 15240 24754
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15304 22574 15332 25350
rect 15580 24936 15608 31078
rect 15488 24908 15608 24936
rect 15488 24698 15516 24908
rect 15568 24812 15620 24818
rect 15672 24800 15700 31368
rect 15620 24772 15700 24800
rect 15568 24754 15620 24760
rect 15488 24670 15608 24698
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15396 22094 15424 22578
rect 15304 22066 15424 22094
rect 15304 21978 15332 22066
rect 15212 21950 15332 21978
rect 15212 21457 15240 21950
rect 15384 21888 15436 21894
rect 15290 21856 15346 21865
rect 15384 21830 15436 21836
rect 15290 21791 15346 21800
rect 15198 21448 15254 21457
rect 15198 21383 15254 21392
rect 15200 21140 15252 21146
rect 15200 21082 15252 21088
rect 15212 15162 15240 21082
rect 15304 20806 15332 21791
rect 15292 20800 15344 20806
rect 15292 20742 15344 20748
rect 15290 18320 15346 18329
rect 15290 18255 15346 18264
rect 15304 16250 15332 18255
rect 15396 16561 15424 21830
rect 15488 21690 15516 24346
rect 15476 21684 15528 21690
rect 15476 21626 15528 21632
rect 15476 21480 15528 21486
rect 15476 21422 15528 21428
rect 15382 16552 15438 16561
rect 15382 16487 15438 16496
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15488 16182 15516 21422
rect 15580 18884 15608 24670
rect 15580 18856 15700 18884
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15580 17134 15608 18702
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15568 16176 15620 16182
rect 15672 16164 15700 18856
rect 15620 16136 15700 16164
rect 15568 16118 15620 16124
rect 15384 16040 15436 16046
rect 15290 16008 15346 16017
rect 15384 15982 15436 15988
rect 15290 15943 15346 15952
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15304 13530 15332 15943
rect 15396 14770 15424 15982
rect 15568 15972 15620 15978
rect 15568 15914 15620 15920
rect 15580 15858 15608 15914
rect 15580 15830 15700 15858
rect 15396 14742 15516 14770
rect 15382 14648 15438 14657
rect 15382 14583 15438 14592
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15290 9616 15346 9625
rect 15290 9551 15346 9560
rect 15108 6452 15160 6458
rect 15108 6394 15160 6400
rect 14830 5672 14886 5681
rect 14830 5607 14886 5616
rect 14740 1896 14792 1902
rect 14740 1838 14792 1844
rect 14844 1766 14872 5607
rect 15304 4214 15332 9551
rect 15292 4208 15344 4214
rect 15292 4150 15344 4156
rect 15396 4146 15424 14583
rect 15488 12986 15516 14742
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15672 9674 15700 15830
rect 15580 9646 15700 9674
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15580 1902 15608 9646
rect 15568 1896 15620 1902
rect 15568 1838 15620 1844
rect 14832 1760 14884 1766
rect 14832 1702 14884 1708
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 14382 1116 14690 1125
rect 14382 1114 14388 1116
rect 14444 1114 14468 1116
rect 14524 1114 14548 1116
rect 14604 1114 14628 1116
rect 14684 1114 14690 1116
rect 14444 1062 14446 1114
rect 14626 1062 14628 1114
rect 14382 1060 14388 1062
rect 14444 1060 14468 1062
rect 14524 1060 14548 1062
rect 14604 1060 14628 1062
rect 14684 1060 14690 1062
rect 14382 1051 14690 1060
rect 15212 160 15240 1294
rect 14462 82 14518 160
rect 14200 54 14518 82
rect 14462 -300 14518 54
rect 15198 -300 15254 160
<< via2 >>
rect 1398 41384 1454 41440
rect 754 40568 810 40624
rect 1490 39888 1546 39944
rect 754 38936 810 38992
rect 754 38120 810 38176
rect 754 37304 810 37360
rect 754 36488 810 36544
rect 1490 35808 1546 35864
rect 754 34856 810 34912
rect 1398 34448 1454 34504
rect 754 33224 810 33280
rect 4314 43546 4370 43548
rect 4394 43546 4450 43548
rect 4474 43546 4530 43548
rect 4554 43546 4610 43548
rect 4314 43494 4360 43546
rect 4360 43494 4370 43546
rect 4394 43494 4424 43546
rect 4424 43494 4436 43546
rect 4436 43494 4450 43546
rect 4474 43494 4488 43546
rect 4488 43494 4500 43546
rect 4500 43494 4530 43546
rect 4554 43494 4564 43546
rect 4564 43494 4610 43546
rect 4314 43492 4370 43494
rect 4394 43492 4450 43494
rect 4474 43492 4530 43494
rect 4554 43492 4610 43494
rect 7672 43546 7728 43548
rect 7752 43546 7808 43548
rect 7832 43546 7888 43548
rect 7912 43546 7968 43548
rect 7672 43494 7718 43546
rect 7718 43494 7728 43546
rect 7752 43494 7782 43546
rect 7782 43494 7794 43546
rect 7794 43494 7808 43546
rect 7832 43494 7846 43546
rect 7846 43494 7858 43546
rect 7858 43494 7888 43546
rect 7912 43494 7922 43546
rect 7922 43494 7968 43546
rect 7672 43492 7728 43494
rect 7752 43492 7808 43494
rect 7832 43492 7888 43494
rect 7912 43492 7968 43494
rect 11030 43546 11086 43548
rect 11110 43546 11166 43548
rect 11190 43546 11246 43548
rect 11270 43546 11326 43548
rect 11030 43494 11076 43546
rect 11076 43494 11086 43546
rect 11110 43494 11140 43546
rect 11140 43494 11152 43546
rect 11152 43494 11166 43546
rect 11190 43494 11204 43546
rect 11204 43494 11216 43546
rect 11216 43494 11246 43546
rect 11270 43494 11280 43546
rect 11280 43494 11326 43546
rect 11030 43492 11086 43494
rect 11110 43492 11166 43494
rect 11190 43492 11246 43494
rect 11270 43492 11326 43494
rect 2635 43002 2691 43004
rect 2715 43002 2771 43004
rect 2795 43002 2851 43004
rect 2875 43002 2931 43004
rect 2635 42950 2681 43002
rect 2681 42950 2691 43002
rect 2715 42950 2745 43002
rect 2745 42950 2757 43002
rect 2757 42950 2771 43002
rect 2795 42950 2809 43002
rect 2809 42950 2821 43002
rect 2821 42950 2851 43002
rect 2875 42950 2885 43002
rect 2885 42950 2931 43002
rect 2635 42948 2691 42950
rect 2715 42948 2771 42950
rect 2795 42948 2851 42950
rect 2875 42948 2931 42950
rect 754 32408 810 32464
rect 1398 31592 1454 31648
rect 754 30776 810 30832
rect 754 29960 810 30016
rect 754 29144 810 29200
rect 1766 29008 1822 29064
rect 1582 28464 1638 28520
rect 754 28328 810 28384
rect 1398 27512 1454 27568
rect 754 26696 810 26752
rect 1490 26152 1546 26208
rect 754 25064 810 25120
rect 754 24248 810 24304
rect 754 23432 810 23488
rect 754 22616 810 22672
rect 754 21800 810 21856
rect 754 20984 810 21040
rect 754 20168 810 20224
rect 754 19352 810 19408
rect 754 18536 810 18592
rect 754 16904 810 16960
rect 754 16088 810 16144
rect 754 15272 810 15328
rect 1490 17856 1546 17912
rect 846 14456 902 14512
rect 2635 41914 2691 41916
rect 2715 41914 2771 41916
rect 2795 41914 2851 41916
rect 2875 41914 2931 41916
rect 2635 41862 2681 41914
rect 2681 41862 2691 41914
rect 2715 41862 2745 41914
rect 2745 41862 2757 41914
rect 2757 41862 2771 41914
rect 2795 41862 2809 41914
rect 2809 41862 2821 41914
rect 2821 41862 2851 41914
rect 2875 41862 2885 41914
rect 2885 41862 2931 41914
rect 2635 41860 2691 41862
rect 2715 41860 2771 41862
rect 2795 41860 2851 41862
rect 2875 41860 2931 41862
rect 2635 40826 2691 40828
rect 2715 40826 2771 40828
rect 2795 40826 2851 40828
rect 2875 40826 2931 40828
rect 2635 40774 2681 40826
rect 2681 40774 2691 40826
rect 2715 40774 2745 40826
rect 2745 40774 2757 40826
rect 2757 40774 2771 40826
rect 2795 40774 2809 40826
rect 2809 40774 2821 40826
rect 2821 40774 2851 40826
rect 2875 40774 2885 40826
rect 2885 40774 2931 40826
rect 2635 40772 2691 40774
rect 2715 40772 2771 40774
rect 2795 40772 2851 40774
rect 2875 40772 2931 40774
rect 2635 39738 2691 39740
rect 2715 39738 2771 39740
rect 2795 39738 2851 39740
rect 2875 39738 2931 39740
rect 2635 39686 2681 39738
rect 2681 39686 2691 39738
rect 2715 39686 2745 39738
rect 2745 39686 2757 39738
rect 2757 39686 2771 39738
rect 2795 39686 2809 39738
rect 2809 39686 2821 39738
rect 2821 39686 2851 39738
rect 2875 39686 2885 39738
rect 2885 39686 2931 39738
rect 2635 39684 2691 39686
rect 2715 39684 2771 39686
rect 2795 39684 2851 39686
rect 2875 39684 2931 39686
rect 2635 38650 2691 38652
rect 2715 38650 2771 38652
rect 2795 38650 2851 38652
rect 2875 38650 2931 38652
rect 2635 38598 2681 38650
rect 2681 38598 2691 38650
rect 2715 38598 2745 38650
rect 2745 38598 2757 38650
rect 2757 38598 2771 38650
rect 2795 38598 2809 38650
rect 2809 38598 2821 38650
rect 2821 38598 2851 38650
rect 2875 38598 2885 38650
rect 2885 38598 2931 38650
rect 2635 38596 2691 38598
rect 2715 38596 2771 38598
rect 2795 38596 2851 38598
rect 2875 38596 2931 38598
rect 2635 37562 2691 37564
rect 2715 37562 2771 37564
rect 2795 37562 2851 37564
rect 2875 37562 2931 37564
rect 2635 37510 2681 37562
rect 2681 37510 2691 37562
rect 2715 37510 2745 37562
rect 2745 37510 2757 37562
rect 2757 37510 2771 37562
rect 2795 37510 2809 37562
rect 2809 37510 2821 37562
rect 2821 37510 2851 37562
rect 2875 37510 2885 37562
rect 2885 37510 2931 37562
rect 2635 37508 2691 37510
rect 2715 37508 2771 37510
rect 2795 37508 2851 37510
rect 2875 37508 2931 37510
rect 2635 36474 2691 36476
rect 2715 36474 2771 36476
rect 2795 36474 2851 36476
rect 2875 36474 2931 36476
rect 2635 36422 2681 36474
rect 2681 36422 2691 36474
rect 2715 36422 2745 36474
rect 2745 36422 2757 36474
rect 2757 36422 2771 36474
rect 2795 36422 2809 36474
rect 2809 36422 2821 36474
rect 2821 36422 2851 36474
rect 2875 36422 2885 36474
rect 2885 36422 2931 36474
rect 2635 36420 2691 36422
rect 2715 36420 2771 36422
rect 2795 36420 2851 36422
rect 2875 36420 2931 36422
rect 2635 35386 2691 35388
rect 2715 35386 2771 35388
rect 2795 35386 2851 35388
rect 2875 35386 2931 35388
rect 2635 35334 2681 35386
rect 2681 35334 2691 35386
rect 2715 35334 2745 35386
rect 2745 35334 2757 35386
rect 2757 35334 2771 35386
rect 2795 35334 2809 35386
rect 2809 35334 2821 35386
rect 2821 35334 2851 35386
rect 2875 35334 2885 35386
rect 2885 35334 2931 35386
rect 2635 35332 2691 35334
rect 2715 35332 2771 35334
rect 2795 35332 2851 35334
rect 2875 35332 2931 35334
rect 2635 34298 2691 34300
rect 2715 34298 2771 34300
rect 2795 34298 2851 34300
rect 2875 34298 2931 34300
rect 2635 34246 2681 34298
rect 2681 34246 2691 34298
rect 2715 34246 2745 34298
rect 2745 34246 2757 34298
rect 2757 34246 2771 34298
rect 2795 34246 2809 34298
rect 2809 34246 2821 34298
rect 2821 34246 2851 34298
rect 2875 34246 2885 34298
rect 2885 34246 2931 34298
rect 2635 34244 2691 34246
rect 2715 34244 2771 34246
rect 2795 34244 2851 34246
rect 2875 34244 2931 34246
rect 2635 33210 2691 33212
rect 2715 33210 2771 33212
rect 2795 33210 2851 33212
rect 2875 33210 2931 33212
rect 2635 33158 2681 33210
rect 2681 33158 2691 33210
rect 2715 33158 2745 33210
rect 2745 33158 2757 33210
rect 2757 33158 2771 33210
rect 2795 33158 2809 33210
rect 2809 33158 2821 33210
rect 2821 33158 2851 33210
rect 2875 33158 2885 33210
rect 2885 33158 2931 33210
rect 2635 33156 2691 33158
rect 2715 33156 2771 33158
rect 2795 33156 2851 33158
rect 2875 33156 2931 33158
rect 2635 32122 2691 32124
rect 2715 32122 2771 32124
rect 2795 32122 2851 32124
rect 2875 32122 2931 32124
rect 2635 32070 2681 32122
rect 2681 32070 2691 32122
rect 2715 32070 2745 32122
rect 2745 32070 2757 32122
rect 2757 32070 2771 32122
rect 2795 32070 2809 32122
rect 2809 32070 2821 32122
rect 2821 32070 2851 32122
rect 2875 32070 2885 32122
rect 2885 32070 2931 32122
rect 2635 32068 2691 32070
rect 2715 32068 2771 32070
rect 2795 32068 2851 32070
rect 2875 32068 2931 32070
rect 2635 31034 2691 31036
rect 2715 31034 2771 31036
rect 2795 31034 2851 31036
rect 2875 31034 2931 31036
rect 2635 30982 2681 31034
rect 2681 30982 2691 31034
rect 2715 30982 2745 31034
rect 2745 30982 2757 31034
rect 2757 30982 2771 31034
rect 2795 30982 2809 31034
rect 2809 30982 2821 31034
rect 2821 30982 2851 31034
rect 2875 30982 2885 31034
rect 2885 30982 2931 31034
rect 2635 30980 2691 30982
rect 2715 30980 2771 30982
rect 2795 30980 2851 30982
rect 2875 30980 2931 30982
rect 2635 29946 2691 29948
rect 2715 29946 2771 29948
rect 2795 29946 2851 29948
rect 2875 29946 2931 29948
rect 2635 29894 2681 29946
rect 2681 29894 2691 29946
rect 2715 29894 2745 29946
rect 2745 29894 2757 29946
rect 2757 29894 2771 29946
rect 2795 29894 2809 29946
rect 2809 29894 2821 29946
rect 2821 29894 2851 29946
rect 2875 29894 2885 29946
rect 2885 29894 2931 29946
rect 2635 29892 2691 29894
rect 2715 29892 2771 29894
rect 2795 29892 2851 29894
rect 2875 29892 2931 29894
rect 846 12824 902 12880
rect 2635 28858 2691 28860
rect 2715 28858 2771 28860
rect 2795 28858 2851 28860
rect 2875 28858 2931 28860
rect 2635 28806 2681 28858
rect 2681 28806 2691 28858
rect 2715 28806 2745 28858
rect 2745 28806 2757 28858
rect 2757 28806 2771 28858
rect 2795 28806 2809 28858
rect 2809 28806 2821 28858
rect 2821 28806 2851 28858
rect 2875 28806 2885 28858
rect 2885 28806 2931 28858
rect 2635 28804 2691 28806
rect 2715 28804 2771 28806
rect 2795 28804 2851 28806
rect 2875 28804 2931 28806
rect 2635 27770 2691 27772
rect 2715 27770 2771 27772
rect 2795 27770 2851 27772
rect 2875 27770 2931 27772
rect 2635 27718 2681 27770
rect 2681 27718 2691 27770
rect 2715 27718 2745 27770
rect 2745 27718 2757 27770
rect 2757 27718 2771 27770
rect 2795 27718 2809 27770
rect 2809 27718 2821 27770
rect 2821 27718 2851 27770
rect 2875 27718 2885 27770
rect 2885 27718 2931 27770
rect 2635 27716 2691 27718
rect 2715 27716 2771 27718
rect 2795 27716 2851 27718
rect 2875 27716 2931 27718
rect 2635 26682 2691 26684
rect 2715 26682 2771 26684
rect 2795 26682 2851 26684
rect 2875 26682 2931 26684
rect 2635 26630 2681 26682
rect 2681 26630 2691 26682
rect 2715 26630 2745 26682
rect 2745 26630 2757 26682
rect 2757 26630 2771 26682
rect 2795 26630 2809 26682
rect 2809 26630 2821 26682
rect 2821 26630 2851 26682
rect 2875 26630 2885 26682
rect 2885 26630 2931 26682
rect 2635 26628 2691 26630
rect 2715 26628 2771 26630
rect 2795 26628 2851 26630
rect 2875 26628 2931 26630
rect 2635 25594 2691 25596
rect 2715 25594 2771 25596
rect 2795 25594 2851 25596
rect 2875 25594 2931 25596
rect 2635 25542 2681 25594
rect 2681 25542 2691 25594
rect 2715 25542 2745 25594
rect 2745 25542 2757 25594
rect 2757 25542 2771 25594
rect 2795 25542 2809 25594
rect 2809 25542 2821 25594
rect 2821 25542 2851 25594
rect 2875 25542 2885 25594
rect 2885 25542 2931 25594
rect 2635 25540 2691 25542
rect 2715 25540 2771 25542
rect 2795 25540 2851 25542
rect 2875 25540 2931 25542
rect 2635 24506 2691 24508
rect 2715 24506 2771 24508
rect 2795 24506 2851 24508
rect 2875 24506 2931 24508
rect 2635 24454 2681 24506
rect 2681 24454 2691 24506
rect 2715 24454 2745 24506
rect 2745 24454 2757 24506
rect 2757 24454 2771 24506
rect 2795 24454 2809 24506
rect 2809 24454 2821 24506
rect 2821 24454 2851 24506
rect 2875 24454 2885 24506
rect 2885 24454 2931 24506
rect 2635 24452 2691 24454
rect 2715 24452 2771 24454
rect 2795 24452 2851 24454
rect 2875 24452 2931 24454
rect 2635 23418 2691 23420
rect 2715 23418 2771 23420
rect 2795 23418 2851 23420
rect 2875 23418 2931 23420
rect 2635 23366 2681 23418
rect 2681 23366 2691 23418
rect 2715 23366 2745 23418
rect 2745 23366 2757 23418
rect 2757 23366 2771 23418
rect 2795 23366 2809 23418
rect 2809 23366 2821 23418
rect 2821 23366 2851 23418
rect 2875 23366 2885 23418
rect 2885 23366 2931 23418
rect 2635 23364 2691 23366
rect 2715 23364 2771 23366
rect 2795 23364 2851 23366
rect 2875 23364 2931 23366
rect 2410 17040 2466 17096
rect 2635 22330 2691 22332
rect 2715 22330 2771 22332
rect 2795 22330 2851 22332
rect 2875 22330 2931 22332
rect 2635 22278 2681 22330
rect 2681 22278 2691 22330
rect 2715 22278 2745 22330
rect 2745 22278 2757 22330
rect 2757 22278 2771 22330
rect 2795 22278 2809 22330
rect 2809 22278 2821 22330
rect 2821 22278 2851 22330
rect 2875 22278 2885 22330
rect 2885 22278 2931 22330
rect 2635 22276 2691 22278
rect 2715 22276 2771 22278
rect 2795 22276 2851 22278
rect 2875 22276 2931 22278
rect 2635 21242 2691 21244
rect 2715 21242 2771 21244
rect 2795 21242 2851 21244
rect 2875 21242 2931 21244
rect 2635 21190 2681 21242
rect 2681 21190 2691 21242
rect 2715 21190 2745 21242
rect 2745 21190 2757 21242
rect 2757 21190 2771 21242
rect 2795 21190 2809 21242
rect 2809 21190 2821 21242
rect 2821 21190 2851 21242
rect 2875 21190 2885 21242
rect 2885 21190 2931 21242
rect 2635 21188 2691 21190
rect 2715 21188 2771 21190
rect 2795 21188 2851 21190
rect 2875 21188 2931 21190
rect 2635 20154 2691 20156
rect 2715 20154 2771 20156
rect 2795 20154 2851 20156
rect 2875 20154 2931 20156
rect 2635 20102 2681 20154
rect 2681 20102 2691 20154
rect 2715 20102 2745 20154
rect 2745 20102 2757 20154
rect 2757 20102 2771 20154
rect 2795 20102 2809 20154
rect 2809 20102 2821 20154
rect 2821 20102 2851 20154
rect 2875 20102 2885 20154
rect 2885 20102 2931 20154
rect 2635 20100 2691 20102
rect 2715 20100 2771 20102
rect 2795 20100 2851 20102
rect 2875 20100 2931 20102
rect 2635 19066 2691 19068
rect 2715 19066 2771 19068
rect 2795 19066 2851 19068
rect 2875 19066 2931 19068
rect 2635 19014 2681 19066
rect 2681 19014 2691 19066
rect 2715 19014 2745 19066
rect 2745 19014 2757 19066
rect 2757 19014 2771 19066
rect 2795 19014 2809 19066
rect 2809 19014 2821 19066
rect 2821 19014 2851 19066
rect 2875 19014 2885 19066
rect 2885 19014 2931 19066
rect 2635 19012 2691 19014
rect 2715 19012 2771 19014
rect 2795 19012 2851 19014
rect 2875 19012 2931 19014
rect 2635 17978 2691 17980
rect 2715 17978 2771 17980
rect 2795 17978 2851 17980
rect 2875 17978 2931 17980
rect 2635 17926 2681 17978
rect 2681 17926 2691 17978
rect 2715 17926 2745 17978
rect 2745 17926 2757 17978
rect 2757 17926 2771 17978
rect 2795 17926 2809 17978
rect 2809 17926 2821 17978
rect 2821 17926 2851 17978
rect 2875 17926 2885 17978
rect 2885 17926 2931 17978
rect 2635 17924 2691 17926
rect 2715 17924 2771 17926
rect 2795 17924 2851 17926
rect 2875 17924 2931 17926
rect 2635 16890 2691 16892
rect 2715 16890 2771 16892
rect 2795 16890 2851 16892
rect 2875 16890 2931 16892
rect 2635 16838 2681 16890
rect 2681 16838 2691 16890
rect 2715 16838 2745 16890
rect 2745 16838 2757 16890
rect 2757 16838 2771 16890
rect 2795 16838 2809 16890
rect 2809 16838 2821 16890
rect 2821 16838 2851 16890
rect 2875 16838 2885 16890
rect 2885 16838 2931 16890
rect 2635 16836 2691 16838
rect 2715 16836 2771 16838
rect 2795 16836 2851 16838
rect 2875 16836 2931 16838
rect 2635 15802 2691 15804
rect 2715 15802 2771 15804
rect 2795 15802 2851 15804
rect 2875 15802 2931 15804
rect 2635 15750 2681 15802
rect 2681 15750 2691 15802
rect 2715 15750 2745 15802
rect 2745 15750 2757 15802
rect 2757 15750 2771 15802
rect 2795 15750 2809 15802
rect 2809 15750 2821 15802
rect 2821 15750 2851 15802
rect 2875 15750 2885 15802
rect 2885 15750 2931 15802
rect 2635 15748 2691 15750
rect 2715 15748 2771 15750
rect 2795 15748 2851 15750
rect 2875 15748 2931 15750
rect 1582 13676 1584 13696
rect 1584 13676 1636 13696
rect 1636 13676 1638 13696
rect 1582 13640 1638 13676
rect 846 12044 848 12064
rect 848 12044 900 12064
rect 900 12044 902 12064
rect 846 12008 902 12044
rect 846 11192 902 11248
rect 846 10412 848 10432
rect 848 10412 900 10432
rect 900 10412 902 10432
rect 846 10376 902 10412
rect 2635 14714 2691 14716
rect 2715 14714 2771 14716
rect 2795 14714 2851 14716
rect 2875 14714 2931 14716
rect 2635 14662 2681 14714
rect 2681 14662 2691 14714
rect 2715 14662 2745 14714
rect 2745 14662 2757 14714
rect 2757 14662 2771 14714
rect 2795 14662 2809 14714
rect 2809 14662 2821 14714
rect 2821 14662 2851 14714
rect 2875 14662 2885 14714
rect 2885 14662 2931 14714
rect 2635 14660 2691 14662
rect 2715 14660 2771 14662
rect 2795 14660 2851 14662
rect 2875 14660 2931 14662
rect 2635 13626 2691 13628
rect 2715 13626 2771 13628
rect 2795 13626 2851 13628
rect 2875 13626 2931 13628
rect 2635 13574 2681 13626
rect 2681 13574 2691 13626
rect 2715 13574 2745 13626
rect 2745 13574 2757 13626
rect 2757 13574 2771 13626
rect 2795 13574 2809 13626
rect 2809 13574 2821 13626
rect 2821 13574 2851 13626
rect 2875 13574 2885 13626
rect 2885 13574 2931 13626
rect 2635 13572 2691 13574
rect 2715 13572 2771 13574
rect 2795 13572 2851 13574
rect 2875 13572 2931 13574
rect 2635 12538 2691 12540
rect 2715 12538 2771 12540
rect 2795 12538 2851 12540
rect 2875 12538 2931 12540
rect 2635 12486 2681 12538
rect 2681 12486 2691 12538
rect 2715 12486 2745 12538
rect 2745 12486 2757 12538
rect 2757 12486 2771 12538
rect 2795 12486 2809 12538
rect 2809 12486 2821 12538
rect 2821 12486 2851 12538
rect 2875 12486 2885 12538
rect 2885 12486 2931 12538
rect 2635 12484 2691 12486
rect 2715 12484 2771 12486
rect 2795 12484 2851 12486
rect 2875 12484 2931 12486
rect 2635 11450 2691 11452
rect 2715 11450 2771 11452
rect 2795 11450 2851 11452
rect 2875 11450 2931 11452
rect 2635 11398 2681 11450
rect 2681 11398 2691 11450
rect 2715 11398 2745 11450
rect 2745 11398 2757 11450
rect 2757 11398 2771 11450
rect 2795 11398 2809 11450
rect 2809 11398 2821 11450
rect 2821 11398 2851 11450
rect 2875 11398 2885 11450
rect 2885 11398 2931 11450
rect 2635 11396 2691 11398
rect 2715 11396 2771 11398
rect 2795 11396 2851 11398
rect 2875 11396 2931 11398
rect 1858 10648 1914 10704
rect 846 8780 848 8800
rect 848 8780 900 8800
rect 900 8780 902 8800
rect 846 8744 902 8780
rect 2635 10362 2691 10364
rect 2715 10362 2771 10364
rect 2795 10362 2851 10364
rect 2875 10362 2931 10364
rect 2635 10310 2681 10362
rect 2681 10310 2691 10362
rect 2715 10310 2745 10362
rect 2745 10310 2757 10362
rect 2757 10310 2771 10362
rect 2795 10310 2809 10362
rect 2809 10310 2821 10362
rect 2821 10310 2851 10362
rect 2875 10310 2885 10362
rect 2885 10310 2931 10362
rect 2635 10308 2691 10310
rect 2715 10308 2771 10310
rect 2795 10308 2851 10310
rect 2875 10308 2931 10310
rect 2778 9560 2834 9616
rect 2635 9274 2691 9276
rect 2715 9274 2771 9276
rect 2795 9274 2851 9276
rect 2875 9274 2931 9276
rect 2635 9222 2681 9274
rect 2681 9222 2691 9274
rect 2715 9222 2745 9274
rect 2745 9222 2757 9274
rect 2757 9222 2771 9274
rect 2795 9222 2809 9274
rect 2809 9222 2821 9274
rect 2821 9222 2851 9274
rect 2875 9222 2885 9274
rect 2885 9222 2931 9274
rect 2635 9220 2691 9222
rect 2715 9220 2771 9222
rect 2795 9220 2851 9222
rect 2875 9220 2931 9222
rect 1674 8200 1730 8256
rect 2635 8186 2691 8188
rect 2715 8186 2771 8188
rect 2795 8186 2851 8188
rect 2875 8186 2931 8188
rect 2635 8134 2681 8186
rect 2681 8134 2691 8186
rect 2715 8134 2745 8186
rect 2745 8134 2757 8186
rect 2757 8134 2771 8186
rect 2795 8134 2809 8186
rect 2809 8134 2821 8186
rect 2821 8134 2851 8186
rect 2875 8134 2885 8186
rect 2885 8134 2931 8186
rect 2635 8132 2691 8134
rect 2715 8132 2771 8134
rect 2795 8132 2851 8134
rect 2875 8132 2931 8134
rect 846 7148 848 7168
rect 848 7148 900 7168
rect 900 7148 902 7168
rect 846 7112 902 7148
rect 846 6296 902 6352
rect 2635 7098 2691 7100
rect 2715 7098 2771 7100
rect 2795 7098 2851 7100
rect 2875 7098 2931 7100
rect 2635 7046 2681 7098
rect 2681 7046 2691 7098
rect 2715 7046 2745 7098
rect 2745 7046 2757 7098
rect 2757 7046 2771 7098
rect 2795 7046 2809 7098
rect 2809 7046 2821 7098
rect 2821 7046 2851 7098
rect 2875 7046 2885 7098
rect 2885 7046 2931 7098
rect 2635 7044 2691 7046
rect 2715 7044 2771 7046
rect 2795 7044 2851 7046
rect 2875 7044 2931 7046
rect 1582 5516 1584 5536
rect 1584 5516 1636 5536
rect 1636 5516 1638 5536
rect 1582 5480 1638 5516
rect 846 4664 902 4720
rect 754 3848 810 3904
rect 2635 6010 2691 6012
rect 2715 6010 2771 6012
rect 2795 6010 2851 6012
rect 2875 6010 2931 6012
rect 2635 5958 2681 6010
rect 2681 5958 2691 6010
rect 2715 5958 2745 6010
rect 2745 5958 2757 6010
rect 2757 5958 2771 6010
rect 2795 5958 2809 6010
rect 2809 5958 2821 6010
rect 2821 5958 2851 6010
rect 2875 5958 2885 6010
rect 2885 5958 2931 6010
rect 2635 5956 2691 5958
rect 2715 5956 2771 5958
rect 2795 5956 2851 5958
rect 2875 5956 2931 5958
rect 2635 4922 2691 4924
rect 2715 4922 2771 4924
rect 2795 4922 2851 4924
rect 2875 4922 2931 4924
rect 2635 4870 2681 4922
rect 2681 4870 2691 4922
rect 2715 4870 2745 4922
rect 2745 4870 2757 4922
rect 2757 4870 2771 4922
rect 2795 4870 2809 4922
rect 2809 4870 2821 4922
rect 2821 4870 2851 4922
rect 2875 4870 2885 4922
rect 2885 4870 2931 4922
rect 2635 4868 2691 4870
rect 2715 4868 2771 4870
rect 2795 4868 2851 4870
rect 2875 4868 2931 4870
rect 4314 42458 4370 42460
rect 4394 42458 4450 42460
rect 4474 42458 4530 42460
rect 4554 42458 4610 42460
rect 4314 42406 4360 42458
rect 4360 42406 4370 42458
rect 4394 42406 4424 42458
rect 4424 42406 4436 42458
rect 4436 42406 4450 42458
rect 4474 42406 4488 42458
rect 4488 42406 4500 42458
rect 4500 42406 4530 42458
rect 4554 42406 4564 42458
rect 4564 42406 4610 42458
rect 4314 42404 4370 42406
rect 4394 42404 4450 42406
rect 4474 42404 4530 42406
rect 4554 42404 4610 42406
rect 3698 18672 3754 18728
rect 3606 18264 3662 18320
rect 4250 41520 4306 41576
rect 4894 41384 4950 41440
rect 4314 41370 4370 41372
rect 4394 41370 4450 41372
rect 4474 41370 4530 41372
rect 4554 41370 4610 41372
rect 4314 41318 4360 41370
rect 4360 41318 4370 41370
rect 4394 41318 4424 41370
rect 4424 41318 4436 41370
rect 4436 41318 4450 41370
rect 4474 41318 4488 41370
rect 4488 41318 4500 41370
rect 4500 41318 4530 41370
rect 4554 41318 4564 41370
rect 4564 41318 4610 41370
rect 4314 41316 4370 41318
rect 4394 41316 4450 41318
rect 4474 41316 4530 41318
rect 4554 41316 4610 41318
rect 4314 40282 4370 40284
rect 4394 40282 4450 40284
rect 4474 40282 4530 40284
rect 4554 40282 4610 40284
rect 4314 40230 4360 40282
rect 4360 40230 4370 40282
rect 4394 40230 4424 40282
rect 4424 40230 4436 40282
rect 4436 40230 4450 40282
rect 4474 40230 4488 40282
rect 4488 40230 4500 40282
rect 4500 40230 4530 40282
rect 4554 40230 4564 40282
rect 4564 40230 4610 40282
rect 4314 40228 4370 40230
rect 4394 40228 4450 40230
rect 4474 40228 4530 40230
rect 4554 40228 4610 40230
rect 4314 39194 4370 39196
rect 4394 39194 4450 39196
rect 4474 39194 4530 39196
rect 4554 39194 4610 39196
rect 4314 39142 4360 39194
rect 4360 39142 4370 39194
rect 4394 39142 4424 39194
rect 4424 39142 4436 39194
rect 4436 39142 4450 39194
rect 4474 39142 4488 39194
rect 4488 39142 4500 39194
rect 4500 39142 4530 39194
rect 4554 39142 4564 39194
rect 4564 39142 4610 39194
rect 4314 39140 4370 39142
rect 4394 39140 4450 39142
rect 4474 39140 4530 39142
rect 4554 39140 4610 39142
rect 4314 38106 4370 38108
rect 4394 38106 4450 38108
rect 4474 38106 4530 38108
rect 4554 38106 4610 38108
rect 4314 38054 4360 38106
rect 4360 38054 4370 38106
rect 4394 38054 4424 38106
rect 4424 38054 4436 38106
rect 4436 38054 4450 38106
rect 4474 38054 4488 38106
rect 4488 38054 4500 38106
rect 4500 38054 4530 38106
rect 4554 38054 4564 38106
rect 4564 38054 4610 38106
rect 4314 38052 4370 38054
rect 4394 38052 4450 38054
rect 4474 38052 4530 38054
rect 4554 38052 4610 38054
rect 4314 37018 4370 37020
rect 4394 37018 4450 37020
rect 4474 37018 4530 37020
rect 4554 37018 4610 37020
rect 4314 36966 4360 37018
rect 4360 36966 4370 37018
rect 4394 36966 4424 37018
rect 4424 36966 4436 37018
rect 4436 36966 4450 37018
rect 4474 36966 4488 37018
rect 4488 36966 4500 37018
rect 4500 36966 4530 37018
rect 4554 36966 4564 37018
rect 4564 36966 4610 37018
rect 4314 36964 4370 36966
rect 4394 36964 4450 36966
rect 4474 36964 4530 36966
rect 4554 36964 4610 36966
rect 4314 35930 4370 35932
rect 4394 35930 4450 35932
rect 4474 35930 4530 35932
rect 4554 35930 4610 35932
rect 4314 35878 4360 35930
rect 4360 35878 4370 35930
rect 4394 35878 4424 35930
rect 4424 35878 4436 35930
rect 4436 35878 4450 35930
rect 4474 35878 4488 35930
rect 4488 35878 4500 35930
rect 4500 35878 4530 35930
rect 4554 35878 4564 35930
rect 4564 35878 4610 35930
rect 4314 35876 4370 35878
rect 4394 35876 4450 35878
rect 4474 35876 4530 35878
rect 4554 35876 4610 35878
rect 4314 34842 4370 34844
rect 4394 34842 4450 34844
rect 4474 34842 4530 34844
rect 4554 34842 4610 34844
rect 4314 34790 4360 34842
rect 4360 34790 4370 34842
rect 4394 34790 4424 34842
rect 4424 34790 4436 34842
rect 4436 34790 4450 34842
rect 4474 34790 4488 34842
rect 4488 34790 4500 34842
rect 4500 34790 4530 34842
rect 4554 34790 4564 34842
rect 4564 34790 4610 34842
rect 4314 34788 4370 34790
rect 4394 34788 4450 34790
rect 4474 34788 4530 34790
rect 4554 34788 4610 34790
rect 4314 33754 4370 33756
rect 4394 33754 4450 33756
rect 4474 33754 4530 33756
rect 4554 33754 4610 33756
rect 4314 33702 4360 33754
rect 4360 33702 4370 33754
rect 4394 33702 4424 33754
rect 4424 33702 4436 33754
rect 4436 33702 4450 33754
rect 4474 33702 4488 33754
rect 4488 33702 4500 33754
rect 4500 33702 4530 33754
rect 4554 33702 4564 33754
rect 4564 33702 4610 33754
rect 4314 33700 4370 33702
rect 4394 33700 4450 33702
rect 4474 33700 4530 33702
rect 4554 33700 4610 33702
rect 4314 32666 4370 32668
rect 4394 32666 4450 32668
rect 4474 32666 4530 32668
rect 4554 32666 4610 32668
rect 4314 32614 4360 32666
rect 4360 32614 4370 32666
rect 4394 32614 4424 32666
rect 4424 32614 4436 32666
rect 4436 32614 4450 32666
rect 4474 32614 4488 32666
rect 4488 32614 4500 32666
rect 4500 32614 4530 32666
rect 4554 32614 4564 32666
rect 4564 32614 4610 32666
rect 4314 32612 4370 32614
rect 4394 32612 4450 32614
rect 4474 32612 4530 32614
rect 4554 32612 4610 32614
rect 4314 31578 4370 31580
rect 4394 31578 4450 31580
rect 4474 31578 4530 31580
rect 4554 31578 4610 31580
rect 4314 31526 4360 31578
rect 4360 31526 4370 31578
rect 4394 31526 4424 31578
rect 4424 31526 4436 31578
rect 4436 31526 4450 31578
rect 4474 31526 4488 31578
rect 4488 31526 4500 31578
rect 4500 31526 4530 31578
rect 4554 31526 4564 31578
rect 4564 31526 4610 31578
rect 4314 31524 4370 31526
rect 4394 31524 4450 31526
rect 4474 31524 4530 31526
rect 4554 31524 4610 31526
rect 4314 30490 4370 30492
rect 4394 30490 4450 30492
rect 4474 30490 4530 30492
rect 4554 30490 4610 30492
rect 4314 30438 4360 30490
rect 4360 30438 4370 30490
rect 4394 30438 4424 30490
rect 4424 30438 4436 30490
rect 4436 30438 4450 30490
rect 4474 30438 4488 30490
rect 4488 30438 4500 30490
rect 4500 30438 4530 30490
rect 4554 30438 4564 30490
rect 4564 30438 4610 30490
rect 4314 30436 4370 30438
rect 4394 30436 4450 30438
rect 4474 30436 4530 30438
rect 4554 30436 4610 30438
rect 4314 29402 4370 29404
rect 4394 29402 4450 29404
rect 4474 29402 4530 29404
rect 4554 29402 4610 29404
rect 4314 29350 4360 29402
rect 4360 29350 4370 29402
rect 4394 29350 4424 29402
rect 4424 29350 4436 29402
rect 4436 29350 4450 29402
rect 4474 29350 4488 29402
rect 4488 29350 4500 29402
rect 4500 29350 4530 29402
rect 4554 29350 4564 29402
rect 4564 29350 4610 29402
rect 4314 29348 4370 29350
rect 4394 29348 4450 29350
rect 4474 29348 4530 29350
rect 4554 29348 4610 29350
rect 4314 28314 4370 28316
rect 4394 28314 4450 28316
rect 4474 28314 4530 28316
rect 4554 28314 4610 28316
rect 4314 28262 4360 28314
rect 4360 28262 4370 28314
rect 4394 28262 4424 28314
rect 4424 28262 4436 28314
rect 4436 28262 4450 28314
rect 4474 28262 4488 28314
rect 4488 28262 4500 28314
rect 4500 28262 4530 28314
rect 4554 28262 4564 28314
rect 4564 28262 4610 28314
rect 4314 28260 4370 28262
rect 4394 28260 4450 28262
rect 4474 28260 4530 28262
rect 4554 28260 4610 28262
rect 4066 27920 4122 27976
rect 3974 17040 4030 17096
rect 4314 27226 4370 27228
rect 4394 27226 4450 27228
rect 4474 27226 4530 27228
rect 4554 27226 4610 27228
rect 4314 27174 4360 27226
rect 4360 27174 4370 27226
rect 4394 27174 4424 27226
rect 4424 27174 4436 27226
rect 4436 27174 4450 27226
rect 4474 27174 4488 27226
rect 4488 27174 4500 27226
rect 4500 27174 4530 27226
rect 4554 27174 4564 27226
rect 4564 27174 4610 27226
rect 4314 27172 4370 27174
rect 4394 27172 4450 27174
rect 4474 27172 4530 27174
rect 4554 27172 4610 27174
rect 4314 26138 4370 26140
rect 4394 26138 4450 26140
rect 4474 26138 4530 26140
rect 4554 26138 4610 26140
rect 4314 26086 4360 26138
rect 4360 26086 4370 26138
rect 4394 26086 4424 26138
rect 4424 26086 4436 26138
rect 4436 26086 4450 26138
rect 4474 26086 4488 26138
rect 4488 26086 4500 26138
rect 4500 26086 4530 26138
rect 4554 26086 4564 26138
rect 4564 26086 4610 26138
rect 4314 26084 4370 26086
rect 4394 26084 4450 26086
rect 4474 26084 4530 26086
rect 4554 26084 4610 26086
rect 4314 25050 4370 25052
rect 4394 25050 4450 25052
rect 4474 25050 4530 25052
rect 4554 25050 4610 25052
rect 4314 24998 4360 25050
rect 4360 24998 4370 25050
rect 4394 24998 4424 25050
rect 4424 24998 4436 25050
rect 4436 24998 4450 25050
rect 4474 24998 4488 25050
rect 4488 24998 4500 25050
rect 4500 24998 4530 25050
rect 4554 24998 4564 25050
rect 4564 24998 4610 25050
rect 4314 24996 4370 24998
rect 4394 24996 4450 24998
rect 4474 24996 4530 24998
rect 4554 24996 4610 24998
rect 5993 43002 6049 43004
rect 6073 43002 6129 43004
rect 6153 43002 6209 43004
rect 6233 43002 6289 43004
rect 5993 42950 6039 43002
rect 6039 42950 6049 43002
rect 6073 42950 6103 43002
rect 6103 42950 6115 43002
rect 6115 42950 6129 43002
rect 6153 42950 6167 43002
rect 6167 42950 6179 43002
rect 6179 42950 6209 43002
rect 6233 42950 6243 43002
rect 6243 42950 6289 43002
rect 5993 42948 6049 42950
rect 6073 42948 6129 42950
rect 6153 42948 6209 42950
rect 6233 42948 6289 42950
rect 9351 43002 9407 43004
rect 9431 43002 9487 43004
rect 9511 43002 9567 43004
rect 9591 43002 9647 43004
rect 9351 42950 9397 43002
rect 9397 42950 9407 43002
rect 9431 42950 9461 43002
rect 9461 42950 9473 43002
rect 9473 42950 9487 43002
rect 9511 42950 9525 43002
rect 9525 42950 9537 43002
rect 9537 42950 9567 43002
rect 9591 42950 9601 43002
rect 9601 42950 9647 43002
rect 9351 42948 9407 42950
rect 9431 42948 9487 42950
rect 9511 42948 9567 42950
rect 9591 42948 9647 42950
rect 12709 43002 12765 43004
rect 12789 43002 12845 43004
rect 12869 43002 12925 43004
rect 12949 43002 13005 43004
rect 12709 42950 12755 43002
rect 12755 42950 12765 43002
rect 12789 42950 12819 43002
rect 12819 42950 12831 43002
rect 12831 42950 12845 43002
rect 12869 42950 12883 43002
rect 12883 42950 12895 43002
rect 12895 42950 12925 43002
rect 12949 42950 12959 43002
rect 12959 42950 13005 43002
rect 12709 42948 12765 42950
rect 12789 42948 12845 42950
rect 12869 42948 12925 42950
rect 12949 42948 13005 42950
rect 10046 42744 10102 42800
rect 7930 42644 7932 42664
rect 7932 42644 7984 42664
rect 7984 42644 7986 42664
rect 4314 23962 4370 23964
rect 4394 23962 4450 23964
rect 4474 23962 4530 23964
rect 4554 23962 4610 23964
rect 4314 23910 4360 23962
rect 4360 23910 4370 23962
rect 4394 23910 4424 23962
rect 4424 23910 4436 23962
rect 4436 23910 4450 23962
rect 4474 23910 4488 23962
rect 4488 23910 4500 23962
rect 4500 23910 4530 23962
rect 4554 23910 4564 23962
rect 4564 23910 4610 23962
rect 4314 23908 4370 23910
rect 4394 23908 4450 23910
rect 4474 23908 4530 23910
rect 4554 23908 4610 23910
rect 4314 22874 4370 22876
rect 4394 22874 4450 22876
rect 4474 22874 4530 22876
rect 4554 22874 4610 22876
rect 4314 22822 4360 22874
rect 4360 22822 4370 22874
rect 4394 22822 4424 22874
rect 4424 22822 4436 22874
rect 4436 22822 4450 22874
rect 4474 22822 4488 22874
rect 4488 22822 4500 22874
rect 4500 22822 4530 22874
rect 4554 22822 4564 22874
rect 4564 22822 4610 22874
rect 4314 22820 4370 22822
rect 4394 22820 4450 22822
rect 4474 22820 4530 22822
rect 4554 22820 4610 22822
rect 4314 21786 4370 21788
rect 4394 21786 4450 21788
rect 4474 21786 4530 21788
rect 4554 21786 4610 21788
rect 4314 21734 4360 21786
rect 4360 21734 4370 21786
rect 4394 21734 4424 21786
rect 4424 21734 4436 21786
rect 4436 21734 4450 21786
rect 4474 21734 4488 21786
rect 4488 21734 4500 21786
rect 4500 21734 4530 21786
rect 4554 21734 4564 21786
rect 4564 21734 4610 21786
rect 4314 21732 4370 21734
rect 4394 21732 4450 21734
rect 4474 21732 4530 21734
rect 4554 21732 4610 21734
rect 4526 21564 4528 21584
rect 4528 21564 4580 21584
rect 4580 21564 4582 21584
rect 4526 21528 4582 21564
rect 4314 20698 4370 20700
rect 4394 20698 4450 20700
rect 4474 20698 4530 20700
rect 4554 20698 4610 20700
rect 4314 20646 4360 20698
rect 4360 20646 4370 20698
rect 4394 20646 4424 20698
rect 4424 20646 4436 20698
rect 4436 20646 4450 20698
rect 4474 20646 4488 20698
rect 4488 20646 4500 20698
rect 4500 20646 4530 20698
rect 4554 20646 4564 20698
rect 4564 20646 4610 20698
rect 4314 20644 4370 20646
rect 4394 20644 4450 20646
rect 4474 20644 4530 20646
rect 4554 20644 4610 20646
rect 4158 20440 4214 20496
rect 4314 19610 4370 19612
rect 4394 19610 4450 19612
rect 4474 19610 4530 19612
rect 4554 19610 4610 19612
rect 4314 19558 4360 19610
rect 4360 19558 4370 19610
rect 4394 19558 4424 19610
rect 4424 19558 4436 19610
rect 4436 19558 4450 19610
rect 4474 19558 4488 19610
rect 4488 19558 4500 19610
rect 4500 19558 4530 19610
rect 4554 19558 4564 19610
rect 4564 19558 4610 19610
rect 4314 19556 4370 19558
rect 4394 19556 4450 19558
rect 4474 19556 4530 19558
rect 4554 19556 4610 19558
rect 4314 18522 4370 18524
rect 4394 18522 4450 18524
rect 4474 18522 4530 18524
rect 4554 18522 4610 18524
rect 4314 18470 4360 18522
rect 4360 18470 4370 18522
rect 4394 18470 4424 18522
rect 4424 18470 4436 18522
rect 4436 18470 4450 18522
rect 4474 18470 4488 18522
rect 4488 18470 4500 18522
rect 4500 18470 4530 18522
rect 4554 18470 4564 18522
rect 4564 18470 4610 18522
rect 4314 18468 4370 18470
rect 4394 18468 4450 18470
rect 4474 18468 4530 18470
rect 4554 18468 4610 18470
rect 3882 10512 3938 10568
rect 2635 3834 2691 3836
rect 2715 3834 2771 3836
rect 2795 3834 2851 3836
rect 2875 3834 2931 3836
rect 2635 3782 2681 3834
rect 2681 3782 2691 3834
rect 2715 3782 2745 3834
rect 2745 3782 2757 3834
rect 2757 3782 2771 3834
rect 2795 3782 2809 3834
rect 2809 3782 2821 3834
rect 2821 3782 2851 3834
rect 2875 3782 2885 3834
rect 2885 3782 2931 3834
rect 2635 3780 2691 3782
rect 2715 3780 2771 3782
rect 2795 3780 2851 3782
rect 2875 3780 2931 3782
rect 2635 2746 2691 2748
rect 2715 2746 2771 2748
rect 2795 2746 2851 2748
rect 2875 2746 2931 2748
rect 2635 2694 2681 2746
rect 2681 2694 2691 2746
rect 2715 2694 2745 2746
rect 2745 2694 2757 2746
rect 2757 2694 2771 2746
rect 2795 2694 2809 2746
rect 2809 2694 2821 2746
rect 2821 2694 2851 2746
rect 2875 2694 2885 2746
rect 2885 2694 2931 2746
rect 2635 2692 2691 2694
rect 2715 2692 2771 2694
rect 2795 2692 2851 2694
rect 2875 2692 2931 2694
rect 4314 17434 4370 17436
rect 4394 17434 4450 17436
rect 4474 17434 4530 17436
rect 4554 17434 4610 17436
rect 4314 17382 4360 17434
rect 4360 17382 4370 17434
rect 4394 17382 4424 17434
rect 4424 17382 4436 17434
rect 4436 17382 4450 17434
rect 4474 17382 4488 17434
rect 4488 17382 4500 17434
rect 4500 17382 4530 17434
rect 4554 17382 4564 17434
rect 4564 17382 4610 17434
rect 4314 17380 4370 17382
rect 4394 17380 4450 17382
rect 4474 17380 4530 17382
rect 4554 17380 4610 17382
rect 4314 16346 4370 16348
rect 4394 16346 4450 16348
rect 4474 16346 4530 16348
rect 4554 16346 4610 16348
rect 4314 16294 4360 16346
rect 4360 16294 4370 16346
rect 4394 16294 4424 16346
rect 4424 16294 4436 16346
rect 4436 16294 4450 16346
rect 4474 16294 4488 16346
rect 4488 16294 4500 16346
rect 4500 16294 4530 16346
rect 4554 16294 4564 16346
rect 4564 16294 4610 16346
rect 4314 16292 4370 16294
rect 4394 16292 4450 16294
rect 4474 16292 4530 16294
rect 4554 16292 4610 16294
rect 4314 15258 4370 15260
rect 4394 15258 4450 15260
rect 4474 15258 4530 15260
rect 4554 15258 4610 15260
rect 4314 15206 4360 15258
rect 4360 15206 4370 15258
rect 4394 15206 4424 15258
rect 4424 15206 4436 15258
rect 4436 15206 4450 15258
rect 4474 15206 4488 15258
rect 4488 15206 4500 15258
rect 4500 15206 4530 15258
rect 4554 15206 4564 15258
rect 4564 15206 4610 15258
rect 4314 15204 4370 15206
rect 4394 15204 4450 15206
rect 4474 15204 4530 15206
rect 4554 15204 4610 15206
rect 4314 14170 4370 14172
rect 4394 14170 4450 14172
rect 4474 14170 4530 14172
rect 4554 14170 4610 14172
rect 4314 14118 4360 14170
rect 4360 14118 4370 14170
rect 4394 14118 4424 14170
rect 4424 14118 4436 14170
rect 4436 14118 4450 14170
rect 4474 14118 4488 14170
rect 4488 14118 4500 14170
rect 4500 14118 4530 14170
rect 4554 14118 4564 14170
rect 4564 14118 4610 14170
rect 4314 14116 4370 14118
rect 4394 14116 4450 14118
rect 4474 14116 4530 14118
rect 4554 14116 4610 14118
rect 4314 13082 4370 13084
rect 4394 13082 4450 13084
rect 4474 13082 4530 13084
rect 4554 13082 4610 13084
rect 4314 13030 4360 13082
rect 4360 13030 4370 13082
rect 4394 13030 4424 13082
rect 4424 13030 4436 13082
rect 4436 13030 4450 13082
rect 4474 13030 4488 13082
rect 4488 13030 4500 13082
rect 4500 13030 4530 13082
rect 4554 13030 4564 13082
rect 4564 13030 4610 13082
rect 4314 13028 4370 13030
rect 4394 13028 4450 13030
rect 4474 13028 4530 13030
rect 4554 13028 4610 13030
rect 4986 18808 5042 18864
rect 4314 11994 4370 11996
rect 4394 11994 4450 11996
rect 4474 11994 4530 11996
rect 4554 11994 4610 11996
rect 4314 11942 4360 11994
rect 4360 11942 4370 11994
rect 4394 11942 4424 11994
rect 4424 11942 4436 11994
rect 4436 11942 4450 11994
rect 4474 11942 4488 11994
rect 4488 11942 4500 11994
rect 4500 11942 4530 11994
rect 4554 11942 4564 11994
rect 4564 11942 4610 11994
rect 4314 11940 4370 11942
rect 4394 11940 4450 11942
rect 4474 11940 4530 11942
rect 4554 11940 4610 11942
rect 4314 10906 4370 10908
rect 4394 10906 4450 10908
rect 4474 10906 4530 10908
rect 4554 10906 4610 10908
rect 4314 10854 4360 10906
rect 4360 10854 4370 10906
rect 4394 10854 4424 10906
rect 4424 10854 4436 10906
rect 4436 10854 4450 10906
rect 4474 10854 4488 10906
rect 4488 10854 4500 10906
rect 4500 10854 4530 10906
rect 4554 10854 4564 10906
rect 4564 10854 4610 10906
rect 4314 10852 4370 10854
rect 4394 10852 4450 10854
rect 4474 10852 4530 10854
rect 4554 10852 4610 10854
rect 4314 9818 4370 9820
rect 4394 9818 4450 9820
rect 4474 9818 4530 9820
rect 4554 9818 4610 9820
rect 4314 9766 4360 9818
rect 4360 9766 4370 9818
rect 4394 9766 4424 9818
rect 4424 9766 4436 9818
rect 4436 9766 4450 9818
rect 4474 9766 4488 9818
rect 4488 9766 4500 9818
rect 4500 9766 4530 9818
rect 4554 9766 4564 9818
rect 4564 9766 4610 9818
rect 4314 9764 4370 9766
rect 4394 9764 4450 9766
rect 4474 9764 4530 9766
rect 4554 9764 4610 9766
rect 4314 8730 4370 8732
rect 4394 8730 4450 8732
rect 4474 8730 4530 8732
rect 4554 8730 4610 8732
rect 4314 8678 4360 8730
rect 4360 8678 4370 8730
rect 4394 8678 4424 8730
rect 4424 8678 4436 8730
rect 4436 8678 4450 8730
rect 4474 8678 4488 8730
rect 4488 8678 4500 8730
rect 4500 8678 4530 8730
rect 4554 8678 4564 8730
rect 4564 8678 4610 8730
rect 4314 8676 4370 8678
rect 4394 8676 4450 8678
rect 4474 8676 4530 8678
rect 4554 8676 4610 8678
rect 4314 7642 4370 7644
rect 4394 7642 4450 7644
rect 4474 7642 4530 7644
rect 4554 7642 4610 7644
rect 4314 7590 4360 7642
rect 4360 7590 4370 7642
rect 4394 7590 4424 7642
rect 4424 7590 4436 7642
rect 4436 7590 4450 7642
rect 4474 7590 4488 7642
rect 4488 7590 4500 7642
rect 4500 7590 4530 7642
rect 4554 7590 4564 7642
rect 4564 7590 4610 7642
rect 4314 7588 4370 7590
rect 4394 7588 4450 7590
rect 4474 7588 4530 7590
rect 4554 7588 4610 7590
rect 4314 6554 4370 6556
rect 4394 6554 4450 6556
rect 4474 6554 4530 6556
rect 4554 6554 4610 6556
rect 4314 6502 4360 6554
rect 4360 6502 4370 6554
rect 4394 6502 4424 6554
rect 4424 6502 4436 6554
rect 4436 6502 4450 6554
rect 4474 6502 4488 6554
rect 4488 6502 4500 6554
rect 4500 6502 4530 6554
rect 4554 6502 4564 6554
rect 4564 6502 4610 6554
rect 4314 6500 4370 6502
rect 4394 6500 4450 6502
rect 4474 6500 4530 6502
rect 4554 6500 4610 6502
rect 4314 5466 4370 5468
rect 4394 5466 4450 5468
rect 4474 5466 4530 5468
rect 4554 5466 4610 5468
rect 4314 5414 4360 5466
rect 4360 5414 4370 5466
rect 4394 5414 4424 5466
rect 4424 5414 4436 5466
rect 4436 5414 4450 5466
rect 4474 5414 4488 5466
rect 4488 5414 4500 5466
rect 4500 5414 4530 5466
rect 4554 5414 4564 5466
rect 4564 5414 4610 5466
rect 4314 5412 4370 5414
rect 4394 5412 4450 5414
rect 4474 5412 4530 5414
rect 4554 5412 4610 5414
rect 4314 4378 4370 4380
rect 4394 4378 4450 4380
rect 4474 4378 4530 4380
rect 4554 4378 4610 4380
rect 4314 4326 4360 4378
rect 4360 4326 4370 4378
rect 4394 4326 4424 4378
rect 4424 4326 4436 4378
rect 4436 4326 4450 4378
rect 4474 4326 4488 4378
rect 4488 4326 4500 4378
rect 4500 4326 4530 4378
rect 4554 4326 4564 4378
rect 4564 4326 4610 4378
rect 4314 4324 4370 4326
rect 4394 4324 4450 4326
rect 4474 4324 4530 4326
rect 4554 4324 4610 4326
rect 5446 20304 5502 20360
rect 5993 41914 6049 41916
rect 6073 41914 6129 41916
rect 6153 41914 6209 41916
rect 6233 41914 6289 41916
rect 5993 41862 6039 41914
rect 6039 41862 6049 41914
rect 6073 41862 6103 41914
rect 6103 41862 6115 41914
rect 6115 41862 6129 41914
rect 6153 41862 6167 41914
rect 6167 41862 6179 41914
rect 6179 41862 6209 41914
rect 6233 41862 6243 41914
rect 6243 41862 6289 41914
rect 5993 41860 6049 41862
rect 6073 41860 6129 41862
rect 6153 41860 6209 41862
rect 6233 41860 6289 41862
rect 7930 42608 7986 42644
rect 7672 42458 7728 42460
rect 7752 42458 7808 42460
rect 7832 42458 7888 42460
rect 7912 42458 7968 42460
rect 7672 42406 7718 42458
rect 7718 42406 7728 42458
rect 7752 42406 7782 42458
rect 7782 42406 7794 42458
rect 7794 42406 7808 42458
rect 7832 42406 7846 42458
rect 7846 42406 7858 42458
rect 7858 42406 7888 42458
rect 7912 42406 7922 42458
rect 7922 42406 7968 42458
rect 7672 42404 7728 42406
rect 7752 42404 7808 42406
rect 7832 42404 7888 42406
rect 7912 42404 7968 42406
rect 11030 42458 11086 42460
rect 11110 42458 11166 42460
rect 11190 42458 11246 42460
rect 11270 42458 11326 42460
rect 11030 42406 11076 42458
rect 11076 42406 11086 42458
rect 11110 42406 11140 42458
rect 11140 42406 11152 42458
rect 11152 42406 11166 42458
rect 11190 42406 11204 42458
rect 11204 42406 11216 42458
rect 11216 42406 11246 42458
rect 11270 42406 11280 42458
rect 11280 42406 11326 42458
rect 11030 42404 11086 42406
rect 11110 42404 11166 42406
rect 11190 42404 11246 42406
rect 11270 42404 11326 42406
rect 8666 42064 8722 42120
rect 9351 41914 9407 41916
rect 9431 41914 9487 41916
rect 9511 41914 9567 41916
rect 9591 41914 9647 41916
rect 9351 41862 9397 41914
rect 9397 41862 9407 41914
rect 9431 41862 9461 41914
rect 9461 41862 9473 41914
rect 9473 41862 9487 41914
rect 9511 41862 9525 41914
rect 9525 41862 9537 41914
rect 9537 41862 9567 41914
rect 9591 41862 9601 41914
rect 9601 41862 9647 41914
rect 9351 41860 9407 41862
rect 9431 41860 9487 41862
rect 9511 41860 9567 41862
rect 9591 41860 9647 41862
rect 12709 41914 12765 41916
rect 12789 41914 12845 41916
rect 12869 41914 12925 41916
rect 12949 41914 13005 41916
rect 12709 41862 12755 41914
rect 12755 41862 12765 41914
rect 12789 41862 12819 41914
rect 12819 41862 12831 41914
rect 12831 41862 12845 41914
rect 12869 41862 12883 41914
rect 12883 41862 12895 41914
rect 12895 41862 12925 41914
rect 12949 41862 12959 41914
rect 12959 41862 13005 41914
rect 12709 41860 12765 41862
rect 12789 41860 12845 41862
rect 12869 41860 12925 41862
rect 12949 41860 13005 41862
rect 14388 43546 14444 43548
rect 14468 43546 14524 43548
rect 14548 43546 14604 43548
rect 14628 43546 14684 43548
rect 14388 43494 14434 43546
rect 14434 43494 14444 43546
rect 14468 43494 14498 43546
rect 14498 43494 14510 43546
rect 14510 43494 14524 43546
rect 14548 43494 14562 43546
rect 14562 43494 14574 43546
rect 14574 43494 14604 43546
rect 14628 43494 14638 43546
rect 14638 43494 14684 43546
rect 14388 43492 14444 43494
rect 14468 43492 14524 43494
rect 14548 43492 14604 43494
rect 14628 43492 14684 43494
rect 7194 41656 7250 41712
rect 14388 42458 14444 42460
rect 14468 42458 14524 42460
rect 14548 42458 14604 42460
rect 14628 42458 14684 42460
rect 14388 42406 14434 42458
rect 14434 42406 14444 42458
rect 14468 42406 14498 42458
rect 14498 42406 14510 42458
rect 14510 42406 14524 42458
rect 14548 42406 14562 42458
rect 14562 42406 14574 42458
rect 14574 42406 14604 42458
rect 14628 42406 14638 42458
rect 14638 42406 14684 42458
rect 14388 42404 14444 42406
rect 14468 42404 14524 42406
rect 14548 42404 14604 42406
rect 14628 42404 14684 42406
rect 13818 41520 13874 41576
rect 6458 41384 6514 41440
rect 7672 41370 7728 41372
rect 7752 41370 7808 41372
rect 7832 41370 7888 41372
rect 7912 41370 7968 41372
rect 7672 41318 7718 41370
rect 7718 41318 7728 41370
rect 7752 41318 7782 41370
rect 7782 41318 7794 41370
rect 7794 41318 7808 41370
rect 7832 41318 7846 41370
rect 7846 41318 7858 41370
rect 7858 41318 7888 41370
rect 7912 41318 7922 41370
rect 7922 41318 7968 41370
rect 7672 41316 7728 41318
rect 7752 41316 7808 41318
rect 7832 41316 7888 41318
rect 7912 41316 7968 41318
rect 11030 41370 11086 41372
rect 11110 41370 11166 41372
rect 11190 41370 11246 41372
rect 11270 41370 11326 41372
rect 11030 41318 11076 41370
rect 11076 41318 11086 41370
rect 11110 41318 11140 41370
rect 11140 41318 11152 41370
rect 11152 41318 11166 41370
rect 11190 41318 11204 41370
rect 11204 41318 11216 41370
rect 11216 41318 11246 41370
rect 11270 41318 11280 41370
rect 11280 41318 11326 41370
rect 11030 41316 11086 41318
rect 11110 41316 11166 41318
rect 11190 41316 11246 41318
rect 11270 41316 11326 41318
rect 5993 40826 6049 40828
rect 6073 40826 6129 40828
rect 6153 40826 6209 40828
rect 6233 40826 6289 40828
rect 5993 40774 6039 40826
rect 6039 40774 6049 40826
rect 6073 40774 6103 40826
rect 6103 40774 6115 40826
rect 6115 40774 6129 40826
rect 6153 40774 6167 40826
rect 6167 40774 6179 40826
rect 6179 40774 6209 40826
rect 6233 40774 6243 40826
rect 6243 40774 6289 40826
rect 5993 40772 6049 40774
rect 6073 40772 6129 40774
rect 6153 40772 6209 40774
rect 6233 40772 6289 40774
rect 5993 39738 6049 39740
rect 6073 39738 6129 39740
rect 6153 39738 6209 39740
rect 6233 39738 6289 39740
rect 5993 39686 6039 39738
rect 6039 39686 6049 39738
rect 6073 39686 6103 39738
rect 6103 39686 6115 39738
rect 6115 39686 6129 39738
rect 6153 39686 6167 39738
rect 6167 39686 6179 39738
rect 6179 39686 6209 39738
rect 6233 39686 6243 39738
rect 6243 39686 6289 39738
rect 5993 39684 6049 39686
rect 6073 39684 6129 39686
rect 6153 39684 6209 39686
rect 6233 39684 6289 39686
rect 9351 40826 9407 40828
rect 9431 40826 9487 40828
rect 9511 40826 9567 40828
rect 9591 40826 9647 40828
rect 9351 40774 9397 40826
rect 9397 40774 9407 40826
rect 9431 40774 9461 40826
rect 9461 40774 9473 40826
rect 9473 40774 9487 40826
rect 9511 40774 9525 40826
rect 9525 40774 9537 40826
rect 9537 40774 9567 40826
rect 9591 40774 9601 40826
rect 9601 40774 9647 40826
rect 9351 40772 9407 40774
rect 9431 40772 9487 40774
rect 9511 40772 9567 40774
rect 9591 40772 9647 40774
rect 12709 40826 12765 40828
rect 12789 40826 12845 40828
rect 12869 40826 12925 40828
rect 12949 40826 13005 40828
rect 12709 40774 12755 40826
rect 12755 40774 12765 40826
rect 12789 40774 12819 40826
rect 12819 40774 12831 40826
rect 12831 40774 12845 40826
rect 12869 40774 12883 40826
rect 12883 40774 12895 40826
rect 12895 40774 12925 40826
rect 12949 40774 12959 40826
rect 12959 40774 13005 40826
rect 12709 40772 12765 40774
rect 12789 40772 12845 40774
rect 12869 40772 12925 40774
rect 12949 40772 13005 40774
rect 7672 40282 7728 40284
rect 7752 40282 7808 40284
rect 7832 40282 7888 40284
rect 7912 40282 7968 40284
rect 7672 40230 7718 40282
rect 7718 40230 7728 40282
rect 7752 40230 7782 40282
rect 7782 40230 7794 40282
rect 7794 40230 7808 40282
rect 7832 40230 7846 40282
rect 7846 40230 7858 40282
rect 7858 40230 7888 40282
rect 7912 40230 7922 40282
rect 7922 40230 7968 40282
rect 7672 40228 7728 40230
rect 7752 40228 7808 40230
rect 7832 40228 7888 40230
rect 7912 40228 7968 40230
rect 11030 40282 11086 40284
rect 11110 40282 11166 40284
rect 11190 40282 11246 40284
rect 11270 40282 11326 40284
rect 11030 40230 11076 40282
rect 11076 40230 11086 40282
rect 11110 40230 11140 40282
rect 11140 40230 11152 40282
rect 11152 40230 11166 40282
rect 11190 40230 11204 40282
rect 11204 40230 11216 40282
rect 11216 40230 11246 40282
rect 11270 40230 11280 40282
rect 11280 40230 11326 40282
rect 11030 40228 11086 40230
rect 11110 40228 11166 40230
rect 11190 40228 11246 40230
rect 11270 40228 11326 40230
rect 5993 38650 6049 38652
rect 6073 38650 6129 38652
rect 6153 38650 6209 38652
rect 6233 38650 6289 38652
rect 5993 38598 6039 38650
rect 6039 38598 6049 38650
rect 6073 38598 6103 38650
rect 6103 38598 6115 38650
rect 6115 38598 6129 38650
rect 6153 38598 6167 38650
rect 6167 38598 6179 38650
rect 6179 38598 6209 38650
rect 6233 38598 6243 38650
rect 6243 38598 6289 38650
rect 9351 39738 9407 39740
rect 9431 39738 9487 39740
rect 9511 39738 9567 39740
rect 9591 39738 9647 39740
rect 9351 39686 9397 39738
rect 9397 39686 9407 39738
rect 9431 39686 9461 39738
rect 9461 39686 9473 39738
rect 9473 39686 9487 39738
rect 9511 39686 9525 39738
rect 9525 39686 9537 39738
rect 9537 39686 9567 39738
rect 9591 39686 9601 39738
rect 9601 39686 9647 39738
rect 9351 39684 9407 39686
rect 9431 39684 9487 39686
rect 9511 39684 9567 39686
rect 9591 39684 9647 39686
rect 12709 39738 12765 39740
rect 12789 39738 12845 39740
rect 12869 39738 12925 39740
rect 12949 39738 13005 39740
rect 12709 39686 12755 39738
rect 12755 39686 12765 39738
rect 12789 39686 12819 39738
rect 12819 39686 12831 39738
rect 12831 39686 12845 39738
rect 12869 39686 12883 39738
rect 12883 39686 12895 39738
rect 12895 39686 12925 39738
rect 12949 39686 12959 39738
rect 12959 39686 13005 39738
rect 12709 39684 12765 39686
rect 12789 39684 12845 39686
rect 12869 39684 12925 39686
rect 12949 39684 13005 39686
rect 5993 38596 6049 38598
rect 6073 38596 6129 38598
rect 6153 38596 6209 38598
rect 6233 38596 6289 38598
rect 5993 37562 6049 37564
rect 6073 37562 6129 37564
rect 6153 37562 6209 37564
rect 6233 37562 6289 37564
rect 5993 37510 6039 37562
rect 6039 37510 6049 37562
rect 6073 37510 6103 37562
rect 6103 37510 6115 37562
rect 6115 37510 6129 37562
rect 6153 37510 6167 37562
rect 6167 37510 6179 37562
rect 6179 37510 6209 37562
rect 6233 37510 6243 37562
rect 6243 37510 6289 37562
rect 5993 37508 6049 37510
rect 6073 37508 6129 37510
rect 6153 37508 6209 37510
rect 6233 37508 6289 37510
rect 5993 36474 6049 36476
rect 6073 36474 6129 36476
rect 6153 36474 6209 36476
rect 6233 36474 6289 36476
rect 5993 36422 6039 36474
rect 6039 36422 6049 36474
rect 6073 36422 6103 36474
rect 6103 36422 6115 36474
rect 6115 36422 6129 36474
rect 6153 36422 6167 36474
rect 6167 36422 6179 36474
rect 6179 36422 6209 36474
rect 6233 36422 6243 36474
rect 6243 36422 6289 36474
rect 5993 36420 6049 36422
rect 6073 36420 6129 36422
rect 6153 36420 6209 36422
rect 6233 36420 6289 36422
rect 6458 35536 6514 35592
rect 5993 35386 6049 35388
rect 6073 35386 6129 35388
rect 6153 35386 6209 35388
rect 6233 35386 6289 35388
rect 5993 35334 6039 35386
rect 6039 35334 6049 35386
rect 6073 35334 6103 35386
rect 6103 35334 6115 35386
rect 6115 35334 6129 35386
rect 6153 35334 6167 35386
rect 6167 35334 6179 35386
rect 6179 35334 6209 35386
rect 6233 35334 6243 35386
rect 6243 35334 6289 35386
rect 5993 35332 6049 35334
rect 6073 35332 6129 35334
rect 6153 35332 6209 35334
rect 6233 35332 6289 35334
rect 5722 34604 5778 34640
rect 5722 34584 5724 34604
rect 5724 34584 5776 34604
rect 5776 34584 5778 34604
rect 5993 34298 6049 34300
rect 6073 34298 6129 34300
rect 6153 34298 6209 34300
rect 6233 34298 6289 34300
rect 5993 34246 6039 34298
rect 6039 34246 6049 34298
rect 6073 34246 6103 34298
rect 6103 34246 6115 34298
rect 6115 34246 6129 34298
rect 6153 34246 6167 34298
rect 6167 34246 6179 34298
rect 6179 34246 6209 34298
rect 6233 34246 6243 34298
rect 6243 34246 6289 34298
rect 5993 34244 6049 34246
rect 6073 34244 6129 34246
rect 6153 34244 6209 34246
rect 6233 34244 6289 34246
rect 5993 33210 6049 33212
rect 6073 33210 6129 33212
rect 6153 33210 6209 33212
rect 6233 33210 6289 33212
rect 5993 33158 6039 33210
rect 6039 33158 6049 33210
rect 6073 33158 6103 33210
rect 6103 33158 6115 33210
rect 6115 33158 6129 33210
rect 6153 33158 6167 33210
rect 6167 33158 6179 33210
rect 6179 33158 6209 33210
rect 6233 33158 6243 33210
rect 6243 33158 6289 33210
rect 5993 33156 6049 33158
rect 6073 33156 6129 33158
rect 6153 33156 6209 33158
rect 6233 33156 6289 33158
rect 5993 32122 6049 32124
rect 6073 32122 6129 32124
rect 6153 32122 6209 32124
rect 6233 32122 6289 32124
rect 5993 32070 6039 32122
rect 6039 32070 6049 32122
rect 6073 32070 6103 32122
rect 6103 32070 6115 32122
rect 6115 32070 6129 32122
rect 6153 32070 6167 32122
rect 6167 32070 6179 32122
rect 6179 32070 6209 32122
rect 6233 32070 6243 32122
rect 6243 32070 6289 32122
rect 5993 32068 6049 32070
rect 6073 32068 6129 32070
rect 6153 32068 6209 32070
rect 6233 32068 6289 32070
rect 7672 39194 7728 39196
rect 7752 39194 7808 39196
rect 7832 39194 7888 39196
rect 7912 39194 7968 39196
rect 7672 39142 7718 39194
rect 7718 39142 7728 39194
rect 7752 39142 7782 39194
rect 7782 39142 7794 39194
rect 7794 39142 7808 39194
rect 7832 39142 7846 39194
rect 7846 39142 7858 39194
rect 7858 39142 7888 39194
rect 7912 39142 7922 39194
rect 7922 39142 7968 39194
rect 7672 39140 7728 39142
rect 7752 39140 7808 39142
rect 7832 39140 7888 39142
rect 7912 39140 7968 39142
rect 11030 39194 11086 39196
rect 11110 39194 11166 39196
rect 11190 39194 11246 39196
rect 11270 39194 11326 39196
rect 11030 39142 11076 39194
rect 11076 39142 11086 39194
rect 11110 39142 11140 39194
rect 11140 39142 11152 39194
rect 11152 39142 11166 39194
rect 11190 39142 11204 39194
rect 11204 39142 11216 39194
rect 11216 39142 11246 39194
rect 11270 39142 11280 39194
rect 11280 39142 11326 39194
rect 11030 39140 11086 39142
rect 11110 39140 11166 39142
rect 11190 39140 11246 39142
rect 11270 39140 11326 39142
rect 9351 38650 9407 38652
rect 9431 38650 9487 38652
rect 9511 38650 9567 38652
rect 9591 38650 9647 38652
rect 9351 38598 9397 38650
rect 9397 38598 9407 38650
rect 9431 38598 9461 38650
rect 9461 38598 9473 38650
rect 9473 38598 9487 38650
rect 9511 38598 9525 38650
rect 9525 38598 9537 38650
rect 9537 38598 9567 38650
rect 9591 38598 9601 38650
rect 9601 38598 9647 38650
rect 9351 38596 9407 38598
rect 9431 38596 9487 38598
rect 9511 38596 9567 38598
rect 9591 38596 9647 38598
rect 7672 38106 7728 38108
rect 7752 38106 7808 38108
rect 7832 38106 7888 38108
rect 7912 38106 7968 38108
rect 7672 38054 7718 38106
rect 7718 38054 7728 38106
rect 7752 38054 7782 38106
rect 7782 38054 7794 38106
rect 7794 38054 7808 38106
rect 7832 38054 7846 38106
rect 7846 38054 7858 38106
rect 7858 38054 7888 38106
rect 7912 38054 7922 38106
rect 7922 38054 7968 38106
rect 7672 38052 7728 38054
rect 7752 38052 7808 38054
rect 7832 38052 7888 38054
rect 7912 38052 7968 38054
rect 11030 38106 11086 38108
rect 11110 38106 11166 38108
rect 11190 38106 11246 38108
rect 11270 38106 11326 38108
rect 11030 38054 11076 38106
rect 11076 38054 11086 38106
rect 11110 38054 11140 38106
rect 11140 38054 11152 38106
rect 11152 38054 11166 38106
rect 11190 38054 11204 38106
rect 11204 38054 11216 38106
rect 11216 38054 11246 38106
rect 11270 38054 11280 38106
rect 11280 38054 11326 38106
rect 11030 38052 11086 38054
rect 11110 38052 11166 38054
rect 11190 38052 11246 38054
rect 11270 38052 11326 38054
rect 9351 37562 9407 37564
rect 9431 37562 9487 37564
rect 9511 37562 9567 37564
rect 9591 37562 9647 37564
rect 9351 37510 9397 37562
rect 9397 37510 9407 37562
rect 9431 37510 9461 37562
rect 9461 37510 9473 37562
rect 9473 37510 9487 37562
rect 9511 37510 9525 37562
rect 9525 37510 9537 37562
rect 9537 37510 9567 37562
rect 9591 37510 9601 37562
rect 9601 37510 9647 37562
rect 9351 37508 9407 37510
rect 9431 37508 9487 37510
rect 9511 37508 9567 37510
rect 9591 37508 9647 37510
rect 10414 37304 10470 37360
rect 7672 37018 7728 37020
rect 7752 37018 7808 37020
rect 7832 37018 7888 37020
rect 7912 37018 7968 37020
rect 7672 36966 7718 37018
rect 7718 36966 7728 37018
rect 7752 36966 7782 37018
rect 7782 36966 7794 37018
rect 7794 36966 7808 37018
rect 7832 36966 7846 37018
rect 7846 36966 7858 37018
rect 7858 36966 7888 37018
rect 7912 36966 7922 37018
rect 7922 36966 7968 37018
rect 7672 36964 7728 36966
rect 7752 36964 7808 36966
rect 7832 36964 7888 36966
rect 7912 36964 7968 36966
rect 5993 31034 6049 31036
rect 6073 31034 6129 31036
rect 6153 31034 6209 31036
rect 6233 31034 6289 31036
rect 5993 30982 6039 31034
rect 6039 30982 6049 31034
rect 6073 30982 6103 31034
rect 6103 30982 6115 31034
rect 6115 30982 6129 31034
rect 6153 30982 6167 31034
rect 6167 30982 6179 31034
rect 6179 30982 6209 31034
rect 6233 30982 6243 31034
rect 6243 30982 6289 31034
rect 5993 30980 6049 30982
rect 6073 30980 6129 30982
rect 6153 30980 6209 30982
rect 6233 30980 6289 30982
rect 5993 29946 6049 29948
rect 6073 29946 6129 29948
rect 6153 29946 6209 29948
rect 6233 29946 6289 29948
rect 5993 29894 6039 29946
rect 6039 29894 6049 29946
rect 6073 29894 6103 29946
rect 6103 29894 6115 29946
rect 6115 29894 6129 29946
rect 6153 29894 6167 29946
rect 6167 29894 6179 29946
rect 6179 29894 6209 29946
rect 6233 29894 6243 29946
rect 6243 29894 6289 29946
rect 5993 29892 6049 29894
rect 6073 29892 6129 29894
rect 6153 29892 6209 29894
rect 6233 29892 6289 29894
rect 5993 28858 6049 28860
rect 6073 28858 6129 28860
rect 6153 28858 6209 28860
rect 6233 28858 6289 28860
rect 5993 28806 6039 28858
rect 6039 28806 6049 28858
rect 6073 28806 6103 28858
rect 6103 28806 6115 28858
rect 6115 28806 6129 28858
rect 6153 28806 6167 28858
rect 6167 28806 6179 28858
rect 6179 28806 6209 28858
rect 6233 28806 6243 28858
rect 6243 28806 6289 28858
rect 5993 28804 6049 28806
rect 6073 28804 6129 28806
rect 6153 28804 6209 28806
rect 6233 28804 6289 28806
rect 5993 27770 6049 27772
rect 6073 27770 6129 27772
rect 6153 27770 6209 27772
rect 6233 27770 6289 27772
rect 5993 27718 6039 27770
rect 6039 27718 6049 27770
rect 6073 27718 6103 27770
rect 6103 27718 6115 27770
rect 6115 27718 6129 27770
rect 6153 27718 6167 27770
rect 6167 27718 6179 27770
rect 6179 27718 6209 27770
rect 6233 27718 6243 27770
rect 6243 27718 6289 27770
rect 5993 27716 6049 27718
rect 6073 27716 6129 27718
rect 6153 27716 6209 27718
rect 6233 27716 6289 27718
rect 5993 26682 6049 26684
rect 6073 26682 6129 26684
rect 6153 26682 6209 26684
rect 6233 26682 6289 26684
rect 5993 26630 6039 26682
rect 6039 26630 6049 26682
rect 6073 26630 6103 26682
rect 6103 26630 6115 26682
rect 6115 26630 6129 26682
rect 6153 26630 6167 26682
rect 6167 26630 6179 26682
rect 6179 26630 6209 26682
rect 6233 26630 6243 26682
rect 6243 26630 6289 26682
rect 5993 26628 6049 26630
rect 6073 26628 6129 26630
rect 6153 26628 6209 26630
rect 6233 26628 6289 26630
rect 5993 25594 6049 25596
rect 6073 25594 6129 25596
rect 6153 25594 6209 25596
rect 6233 25594 6289 25596
rect 5993 25542 6039 25594
rect 6039 25542 6049 25594
rect 6073 25542 6103 25594
rect 6103 25542 6115 25594
rect 6115 25542 6129 25594
rect 6153 25542 6167 25594
rect 6167 25542 6179 25594
rect 6179 25542 6209 25594
rect 6233 25542 6243 25594
rect 6243 25542 6289 25594
rect 5993 25540 6049 25542
rect 6073 25540 6129 25542
rect 6153 25540 6209 25542
rect 6233 25540 6289 25542
rect 5993 24506 6049 24508
rect 6073 24506 6129 24508
rect 6153 24506 6209 24508
rect 6233 24506 6289 24508
rect 5993 24454 6039 24506
rect 6039 24454 6049 24506
rect 6073 24454 6103 24506
rect 6103 24454 6115 24506
rect 6115 24454 6129 24506
rect 6153 24454 6167 24506
rect 6167 24454 6179 24506
rect 6179 24454 6209 24506
rect 6233 24454 6243 24506
rect 6243 24454 6289 24506
rect 5993 24452 6049 24454
rect 6073 24452 6129 24454
rect 6153 24452 6209 24454
rect 6233 24452 6289 24454
rect 5993 23418 6049 23420
rect 6073 23418 6129 23420
rect 6153 23418 6209 23420
rect 6233 23418 6289 23420
rect 5993 23366 6039 23418
rect 6039 23366 6049 23418
rect 6073 23366 6103 23418
rect 6103 23366 6115 23418
rect 6115 23366 6129 23418
rect 6153 23366 6167 23418
rect 6167 23366 6179 23418
rect 6179 23366 6209 23418
rect 6233 23366 6243 23418
rect 6243 23366 6289 23418
rect 5993 23364 6049 23366
rect 6073 23364 6129 23366
rect 6153 23364 6209 23366
rect 6233 23364 6289 23366
rect 5993 22330 6049 22332
rect 6073 22330 6129 22332
rect 6153 22330 6209 22332
rect 6233 22330 6289 22332
rect 5993 22278 6039 22330
rect 6039 22278 6049 22330
rect 6073 22278 6103 22330
rect 6103 22278 6115 22330
rect 6115 22278 6129 22330
rect 6153 22278 6167 22330
rect 6167 22278 6179 22330
rect 6179 22278 6209 22330
rect 6233 22278 6243 22330
rect 6243 22278 6289 22330
rect 5993 22276 6049 22278
rect 6073 22276 6129 22278
rect 6153 22276 6209 22278
rect 6233 22276 6289 22278
rect 5993 21242 6049 21244
rect 6073 21242 6129 21244
rect 6153 21242 6209 21244
rect 6233 21242 6289 21244
rect 5993 21190 6039 21242
rect 6039 21190 6049 21242
rect 6073 21190 6103 21242
rect 6103 21190 6115 21242
rect 6115 21190 6129 21242
rect 6153 21190 6167 21242
rect 6167 21190 6179 21242
rect 6179 21190 6209 21242
rect 6233 21190 6243 21242
rect 6243 21190 6289 21242
rect 5993 21188 6049 21190
rect 6073 21188 6129 21190
rect 6153 21188 6209 21190
rect 6233 21188 6289 21190
rect 5993 20154 6049 20156
rect 6073 20154 6129 20156
rect 6153 20154 6209 20156
rect 6233 20154 6289 20156
rect 5993 20102 6039 20154
rect 6039 20102 6049 20154
rect 6073 20102 6103 20154
rect 6103 20102 6115 20154
rect 6115 20102 6129 20154
rect 6153 20102 6167 20154
rect 6167 20102 6179 20154
rect 6179 20102 6209 20154
rect 6233 20102 6243 20154
rect 6243 20102 6289 20154
rect 5993 20100 6049 20102
rect 6073 20100 6129 20102
rect 6153 20100 6209 20102
rect 6233 20100 6289 20102
rect 5993 19066 6049 19068
rect 6073 19066 6129 19068
rect 6153 19066 6209 19068
rect 6233 19066 6289 19068
rect 5993 19014 6039 19066
rect 6039 19014 6049 19066
rect 6073 19014 6103 19066
rect 6103 19014 6115 19066
rect 6115 19014 6129 19066
rect 6153 19014 6167 19066
rect 6167 19014 6179 19066
rect 6179 19014 6209 19066
rect 6233 19014 6243 19066
rect 6243 19014 6289 19066
rect 5993 19012 6049 19014
rect 6073 19012 6129 19014
rect 6153 19012 6209 19014
rect 6233 19012 6289 19014
rect 5993 17978 6049 17980
rect 6073 17978 6129 17980
rect 6153 17978 6209 17980
rect 6233 17978 6289 17980
rect 5993 17926 6039 17978
rect 6039 17926 6049 17978
rect 6073 17926 6103 17978
rect 6103 17926 6115 17978
rect 6115 17926 6129 17978
rect 6153 17926 6167 17978
rect 6167 17926 6179 17978
rect 6179 17926 6209 17978
rect 6233 17926 6243 17978
rect 6243 17926 6289 17978
rect 5993 17924 6049 17926
rect 6073 17924 6129 17926
rect 6153 17924 6209 17926
rect 6233 17924 6289 17926
rect 5993 16890 6049 16892
rect 6073 16890 6129 16892
rect 6153 16890 6209 16892
rect 6233 16890 6289 16892
rect 5993 16838 6039 16890
rect 6039 16838 6049 16890
rect 6073 16838 6103 16890
rect 6103 16838 6115 16890
rect 6115 16838 6129 16890
rect 6153 16838 6167 16890
rect 6167 16838 6179 16890
rect 6179 16838 6209 16890
rect 6233 16838 6243 16890
rect 6243 16838 6289 16890
rect 5993 16836 6049 16838
rect 6073 16836 6129 16838
rect 6153 16836 6209 16838
rect 6233 16836 6289 16838
rect 5993 15802 6049 15804
rect 6073 15802 6129 15804
rect 6153 15802 6209 15804
rect 6233 15802 6289 15804
rect 5993 15750 6039 15802
rect 6039 15750 6049 15802
rect 6073 15750 6103 15802
rect 6103 15750 6115 15802
rect 6115 15750 6129 15802
rect 6153 15750 6167 15802
rect 6167 15750 6179 15802
rect 6179 15750 6209 15802
rect 6233 15750 6243 15802
rect 6243 15750 6289 15802
rect 5993 15748 6049 15750
rect 6073 15748 6129 15750
rect 6153 15748 6209 15750
rect 6233 15748 6289 15750
rect 5993 14714 6049 14716
rect 6073 14714 6129 14716
rect 6153 14714 6209 14716
rect 6233 14714 6289 14716
rect 5993 14662 6039 14714
rect 6039 14662 6049 14714
rect 6073 14662 6103 14714
rect 6103 14662 6115 14714
rect 6115 14662 6129 14714
rect 6153 14662 6167 14714
rect 6167 14662 6179 14714
rect 6179 14662 6209 14714
rect 6233 14662 6243 14714
rect 6243 14662 6289 14714
rect 5993 14660 6049 14662
rect 6073 14660 6129 14662
rect 6153 14660 6209 14662
rect 6233 14660 6289 14662
rect 5993 13626 6049 13628
rect 6073 13626 6129 13628
rect 6153 13626 6209 13628
rect 6233 13626 6289 13628
rect 5993 13574 6039 13626
rect 6039 13574 6049 13626
rect 6073 13574 6103 13626
rect 6103 13574 6115 13626
rect 6115 13574 6129 13626
rect 6153 13574 6167 13626
rect 6167 13574 6179 13626
rect 6179 13574 6209 13626
rect 6233 13574 6243 13626
rect 6243 13574 6289 13626
rect 5993 13572 6049 13574
rect 6073 13572 6129 13574
rect 6153 13572 6209 13574
rect 6233 13572 6289 13574
rect 6918 29008 6974 29064
rect 6826 28464 6882 28520
rect 5993 12538 6049 12540
rect 6073 12538 6129 12540
rect 6153 12538 6209 12540
rect 6233 12538 6289 12540
rect 5993 12486 6039 12538
rect 6039 12486 6049 12538
rect 6073 12486 6103 12538
rect 6103 12486 6115 12538
rect 6115 12486 6129 12538
rect 6153 12486 6167 12538
rect 6167 12486 6179 12538
rect 6179 12486 6209 12538
rect 6233 12486 6243 12538
rect 6243 12486 6289 12538
rect 5993 12484 6049 12486
rect 6073 12484 6129 12486
rect 6153 12484 6209 12486
rect 6233 12484 6289 12486
rect 7672 35930 7728 35932
rect 7752 35930 7808 35932
rect 7832 35930 7888 35932
rect 7912 35930 7968 35932
rect 7672 35878 7718 35930
rect 7718 35878 7728 35930
rect 7752 35878 7782 35930
rect 7782 35878 7794 35930
rect 7794 35878 7808 35930
rect 7832 35878 7846 35930
rect 7846 35878 7858 35930
rect 7858 35878 7888 35930
rect 7912 35878 7922 35930
rect 7922 35878 7968 35930
rect 7672 35876 7728 35878
rect 7752 35876 7808 35878
rect 7832 35876 7888 35878
rect 7912 35876 7968 35878
rect 7672 34842 7728 34844
rect 7752 34842 7808 34844
rect 7832 34842 7888 34844
rect 7912 34842 7968 34844
rect 7672 34790 7718 34842
rect 7718 34790 7728 34842
rect 7752 34790 7782 34842
rect 7782 34790 7794 34842
rect 7794 34790 7808 34842
rect 7832 34790 7846 34842
rect 7846 34790 7858 34842
rect 7858 34790 7888 34842
rect 7912 34790 7922 34842
rect 7922 34790 7968 34842
rect 7672 34788 7728 34790
rect 7752 34788 7808 34790
rect 7832 34788 7888 34790
rect 7912 34788 7968 34790
rect 7672 33754 7728 33756
rect 7752 33754 7808 33756
rect 7832 33754 7888 33756
rect 7912 33754 7968 33756
rect 7672 33702 7718 33754
rect 7718 33702 7728 33754
rect 7752 33702 7782 33754
rect 7782 33702 7794 33754
rect 7794 33702 7808 33754
rect 7832 33702 7846 33754
rect 7846 33702 7858 33754
rect 7858 33702 7888 33754
rect 7912 33702 7922 33754
rect 7922 33702 7968 33754
rect 7672 33700 7728 33702
rect 7752 33700 7808 33702
rect 7832 33700 7888 33702
rect 7912 33700 7968 33702
rect 7672 32666 7728 32668
rect 7752 32666 7808 32668
rect 7832 32666 7888 32668
rect 7912 32666 7968 32668
rect 7672 32614 7718 32666
rect 7718 32614 7728 32666
rect 7752 32614 7782 32666
rect 7782 32614 7794 32666
rect 7794 32614 7808 32666
rect 7832 32614 7846 32666
rect 7846 32614 7858 32666
rect 7858 32614 7888 32666
rect 7912 32614 7922 32666
rect 7922 32614 7968 32666
rect 7672 32612 7728 32614
rect 7752 32612 7808 32614
rect 7832 32612 7888 32614
rect 7912 32612 7968 32614
rect 7672 31578 7728 31580
rect 7752 31578 7808 31580
rect 7832 31578 7888 31580
rect 7912 31578 7968 31580
rect 7672 31526 7718 31578
rect 7718 31526 7728 31578
rect 7752 31526 7782 31578
rect 7782 31526 7794 31578
rect 7794 31526 7808 31578
rect 7832 31526 7846 31578
rect 7846 31526 7858 31578
rect 7858 31526 7888 31578
rect 7912 31526 7922 31578
rect 7922 31526 7968 31578
rect 7672 31524 7728 31526
rect 7752 31524 7808 31526
rect 7832 31524 7888 31526
rect 7912 31524 7968 31526
rect 7194 28464 7250 28520
rect 7672 30490 7728 30492
rect 7752 30490 7808 30492
rect 7832 30490 7888 30492
rect 7912 30490 7968 30492
rect 7672 30438 7718 30490
rect 7718 30438 7728 30490
rect 7752 30438 7782 30490
rect 7782 30438 7794 30490
rect 7794 30438 7808 30490
rect 7832 30438 7846 30490
rect 7846 30438 7858 30490
rect 7858 30438 7888 30490
rect 7912 30438 7922 30490
rect 7922 30438 7968 30490
rect 7672 30436 7728 30438
rect 7752 30436 7808 30438
rect 7832 30436 7888 30438
rect 7912 30436 7968 30438
rect 7672 29402 7728 29404
rect 7752 29402 7808 29404
rect 7832 29402 7888 29404
rect 7912 29402 7968 29404
rect 7672 29350 7718 29402
rect 7718 29350 7728 29402
rect 7752 29350 7782 29402
rect 7782 29350 7794 29402
rect 7794 29350 7808 29402
rect 7832 29350 7846 29402
rect 7846 29350 7858 29402
rect 7858 29350 7888 29402
rect 7912 29350 7922 29402
rect 7922 29350 7968 29402
rect 7672 29348 7728 29350
rect 7752 29348 7808 29350
rect 7832 29348 7888 29350
rect 7912 29348 7968 29350
rect 7672 28314 7728 28316
rect 7752 28314 7808 28316
rect 7832 28314 7888 28316
rect 7912 28314 7968 28316
rect 7672 28262 7718 28314
rect 7718 28262 7728 28314
rect 7752 28262 7782 28314
rect 7782 28262 7794 28314
rect 7794 28262 7808 28314
rect 7832 28262 7846 28314
rect 7846 28262 7858 28314
rect 7858 28262 7888 28314
rect 7912 28262 7922 28314
rect 7922 28262 7968 28314
rect 7672 28260 7728 28262
rect 7752 28260 7808 28262
rect 7832 28260 7888 28262
rect 7912 28260 7968 28262
rect 7930 27784 7986 27840
rect 7672 27226 7728 27228
rect 7752 27226 7808 27228
rect 7832 27226 7888 27228
rect 7912 27226 7968 27228
rect 7672 27174 7718 27226
rect 7718 27174 7728 27226
rect 7752 27174 7782 27226
rect 7782 27174 7794 27226
rect 7794 27174 7808 27226
rect 7832 27174 7846 27226
rect 7846 27174 7858 27226
rect 7858 27174 7888 27226
rect 7912 27174 7922 27226
rect 7922 27174 7968 27226
rect 7672 27172 7728 27174
rect 7752 27172 7808 27174
rect 7832 27172 7888 27174
rect 7912 27172 7968 27174
rect 7286 26324 7288 26344
rect 7288 26324 7340 26344
rect 7340 26324 7342 26344
rect 7286 26288 7342 26324
rect 6918 20712 6974 20768
rect 6918 20440 6974 20496
rect 7010 19896 7066 19952
rect 7010 19216 7066 19272
rect 6826 19116 6828 19136
rect 6828 19116 6880 19136
rect 6880 19116 6882 19136
rect 6826 19080 6882 19116
rect 6918 17604 6974 17640
rect 6918 17584 6920 17604
rect 6920 17584 6972 17604
rect 6972 17584 6974 17604
rect 7672 26138 7728 26140
rect 7752 26138 7808 26140
rect 7832 26138 7888 26140
rect 7912 26138 7968 26140
rect 7672 26086 7718 26138
rect 7718 26086 7728 26138
rect 7752 26086 7782 26138
rect 7782 26086 7794 26138
rect 7794 26086 7808 26138
rect 7832 26086 7846 26138
rect 7846 26086 7858 26138
rect 7858 26086 7888 26138
rect 7912 26086 7922 26138
rect 7922 26086 7968 26138
rect 7672 26084 7728 26086
rect 7752 26084 7808 26086
rect 7832 26084 7888 26086
rect 7912 26084 7968 26086
rect 7672 25050 7728 25052
rect 7752 25050 7808 25052
rect 7832 25050 7888 25052
rect 7912 25050 7968 25052
rect 7672 24998 7718 25050
rect 7718 24998 7728 25050
rect 7752 24998 7782 25050
rect 7782 24998 7794 25050
rect 7794 24998 7808 25050
rect 7832 24998 7846 25050
rect 7846 24998 7858 25050
rect 7858 24998 7888 25050
rect 7912 24998 7922 25050
rect 7922 24998 7968 25050
rect 7672 24996 7728 24998
rect 7752 24996 7808 24998
rect 7832 24996 7888 24998
rect 7912 24996 7968 24998
rect 7672 23962 7728 23964
rect 7752 23962 7808 23964
rect 7832 23962 7888 23964
rect 7912 23962 7968 23964
rect 7672 23910 7718 23962
rect 7718 23910 7728 23962
rect 7752 23910 7782 23962
rect 7782 23910 7794 23962
rect 7794 23910 7808 23962
rect 7832 23910 7846 23962
rect 7846 23910 7858 23962
rect 7858 23910 7888 23962
rect 7912 23910 7922 23962
rect 7922 23910 7968 23962
rect 7672 23908 7728 23910
rect 7752 23908 7808 23910
rect 7832 23908 7888 23910
rect 7912 23908 7968 23910
rect 7562 23568 7618 23624
rect 7378 21800 7434 21856
rect 5993 11450 6049 11452
rect 6073 11450 6129 11452
rect 6153 11450 6209 11452
rect 6233 11450 6289 11452
rect 5993 11398 6039 11450
rect 6039 11398 6049 11450
rect 6073 11398 6103 11450
rect 6103 11398 6115 11450
rect 6115 11398 6129 11450
rect 6153 11398 6167 11450
rect 6167 11398 6179 11450
rect 6179 11398 6209 11450
rect 6233 11398 6243 11450
rect 6243 11398 6289 11450
rect 5993 11396 6049 11398
rect 6073 11396 6129 11398
rect 6153 11396 6209 11398
rect 6233 11396 6289 11398
rect 9351 36474 9407 36476
rect 9431 36474 9487 36476
rect 9511 36474 9567 36476
rect 9591 36474 9647 36476
rect 9351 36422 9397 36474
rect 9397 36422 9407 36474
rect 9431 36422 9461 36474
rect 9461 36422 9473 36474
rect 9473 36422 9487 36474
rect 9511 36422 9525 36474
rect 9525 36422 9537 36474
rect 9537 36422 9567 36474
rect 9591 36422 9601 36474
rect 9601 36422 9647 36474
rect 9351 36420 9407 36422
rect 9431 36420 9487 36422
rect 9511 36420 9567 36422
rect 9591 36420 9647 36422
rect 9351 35386 9407 35388
rect 9431 35386 9487 35388
rect 9511 35386 9567 35388
rect 9591 35386 9647 35388
rect 9351 35334 9397 35386
rect 9397 35334 9407 35386
rect 9431 35334 9461 35386
rect 9461 35334 9473 35386
rect 9473 35334 9487 35386
rect 9511 35334 9525 35386
rect 9525 35334 9537 35386
rect 9537 35334 9567 35386
rect 9591 35334 9601 35386
rect 9601 35334 9647 35386
rect 9351 35332 9407 35334
rect 9431 35332 9487 35334
rect 9511 35332 9567 35334
rect 9591 35332 9647 35334
rect 9351 34298 9407 34300
rect 9431 34298 9487 34300
rect 9511 34298 9567 34300
rect 9591 34298 9647 34300
rect 9351 34246 9397 34298
rect 9397 34246 9407 34298
rect 9431 34246 9461 34298
rect 9461 34246 9473 34298
rect 9473 34246 9487 34298
rect 9511 34246 9525 34298
rect 9525 34246 9537 34298
rect 9537 34246 9567 34298
rect 9591 34246 9601 34298
rect 9601 34246 9647 34298
rect 9351 34244 9407 34246
rect 9431 34244 9487 34246
rect 9511 34244 9567 34246
rect 9591 34244 9647 34246
rect 11794 37304 11850 37360
rect 11702 37168 11758 37224
rect 11030 37018 11086 37020
rect 11110 37018 11166 37020
rect 11190 37018 11246 37020
rect 11270 37018 11326 37020
rect 11030 36966 11076 37018
rect 11076 36966 11086 37018
rect 11110 36966 11140 37018
rect 11140 36966 11152 37018
rect 11152 36966 11166 37018
rect 11190 36966 11204 37018
rect 11204 36966 11216 37018
rect 11216 36966 11246 37018
rect 11270 36966 11280 37018
rect 11280 36966 11326 37018
rect 11030 36964 11086 36966
rect 11110 36964 11166 36966
rect 11190 36964 11246 36966
rect 11270 36964 11326 36966
rect 11426 36896 11482 36952
rect 9351 33210 9407 33212
rect 9431 33210 9487 33212
rect 9511 33210 9567 33212
rect 9591 33210 9647 33212
rect 9351 33158 9397 33210
rect 9397 33158 9407 33210
rect 9431 33158 9461 33210
rect 9461 33158 9473 33210
rect 9473 33158 9487 33210
rect 9511 33158 9525 33210
rect 9525 33158 9537 33210
rect 9537 33158 9567 33210
rect 9591 33158 9601 33210
rect 9601 33158 9647 33210
rect 9351 33156 9407 33158
rect 9431 33156 9487 33158
rect 9511 33156 9567 33158
rect 9591 33156 9647 33158
rect 8390 28056 8446 28112
rect 7672 22874 7728 22876
rect 7752 22874 7808 22876
rect 7832 22874 7888 22876
rect 7912 22874 7968 22876
rect 7672 22822 7718 22874
rect 7718 22822 7728 22874
rect 7752 22822 7782 22874
rect 7782 22822 7794 22874
rect 7794 22822 7808 22874
rect 7832 22822 7846 22874
rect 7846 22822 7858 22874
rect 7858 22822 7888 22874
rect 7912 22822 7922 22874
rect 7922 22822 7968 22874
rect 7672 22820 7728 22822
rect 7752 22820 7808 22822
rect 7832 22820 7888 22822
rect 7912 22820 7968 22822
rect 7470 19236 7526 19272
rect 7470 19216 7472 19236
rect 7472 19216 7524 19236
rect 7524 19216 7526 19236
rect 7672 21786 7728 21788
rect 7752 21786 7808 21788
rect 7832 21786 7888 21788
rect 7912 21786 7968 21788
rect 7672 21734 7718 21786
rect 7718 21734 7728 21786
rect 7752 21734 7782 21786
rect 7782 21734 7794 21786
rect 7794 21734 7808 21786
rect 7832 21734 7846 21786
rect 7846 21734 7858 21786
rect 7858 21734 7888 21786
rect 7912 21734 7922 21786
rect 7922 21734 7968 21786
rect 7672 21732 7728 21734
rect 7752 21732 7808 21734
rect 7832 21732 7888 21734
rect 7912 21732 7968 21734
rect 7672 20698 7728 20700
rect 7752 20698 7808 20700
rect 7832 20698 7888 20700
rect 7912 20698 7968 20700
rect 7672 20646 7718 20698
rect 7718 20646 7728 20698
rect 7752 20646 7782 20698
rect 7782 20646 7794 20698
rect 7794 20646 7808 20698
rect 7832 20646 7846 20698
rect 7846 20646 7858 20698
rect 7858 20646 7888 20698
rect 7912 20646 7922 20698
rect 7922 20646 7968 20698
rect 7672 20644 7728 20646
rect 7752 20644 7808 20646
rect 7832 20644 7888 20646
rect 7912 20644 7968 20646
rect 7930 20460 7986 20496
rect 7930 20440 7932 20460
rect 7932 20440 7984 20460
rect 7984 20440 7986 20460
rect 7672 19610 7728 19612
rect 7752 19610 7808 19612
rect 7832 19610 7888 19612
rect 7912 19610 7968 19612
rect 7672 19558 7718 19610
rect 7718 19558 7728 19610
rect 7752 19558 7782 19610
rect 7782 19558 7794 19610
rect 7794 19558 7808 19610
rect 7832 19558 7846 19610
rect 7846 19558 7858 19610
rect 7858 19558 7888 19610
rect 7912 19558 7922 19610
rect 7922 19558 7968 19610
rect 7672 19556 7728 19558
rect 7752 19556 7808 19558
rect 7832 19556 7888 19558
rect 7912 19556 7968 19558
rect 7562 18672 7618 18728
rect 7672 18522 7728 18524
rect 7752 18522 7808 18524
rect 7832 18522 7888 18524
rect 7912 18522 7968 18524
rect 7672 18470 7718 18522
rect 7718 18470 7728 18522
rect 7752 18470 7782 18522
rect 7782 18470 7794 18522
rect 7794 18470 7808 18522
rect 7832 18470 7846 18522
rect 7846 18470 7858 18522
rect 7858 18470 7888 18522
rect 7912 18470 7922 18522
rect 7922 18470 7968 18522
rect 7672 18468 7728 18470
rect 7752 18468 7808 18470
rect 7832 18468 7888 18470
rect 7912 18468 7968 18470
rect 8022 17992 8078 18048
rect 7672 17434 7728 17436
rect 7752 17434 7808 17436
rect 7832 17434 7888 17436
rect 7912 17434 7968 17436
rect 7672 17382 7718 17434
rect 7718 17382 7728 17434
rect 7752 17382 7782 17434
rect 7782 17382 7794 17434
rect 7794 17382 7808 17434
rect 7832 17382 7846 17434
rect 7846 17382 7858 17434
rect 7858 17382 7888 17434
rect 7912 17382 7922 17434
rect 7922 17382 7968 17434
rect 7672 17380 7728 17382
rect 7752 17380 7808 17382
rect 7832 17380 7888 17382
rect 7912 17380 7968 17382
rect 7672 16346 7728 16348
rect 7752 16346 7808 16348
rect 7832 16346 7888 16348
rect 7912 16346 7968 16348
rect 7672 16294 7718 16346
rect 7718 16294 7728 16346
rect 7752 16294 7782 16346
rect 7782 16294 7794 16346
rect 7794 16294 7808 16346
rect 7832 16294 7846 16346
rect 7846 16294 7858 16346
rect 7858 16294 7888 16346
rect 7912 16294 7922 16346
rect 7922 16294 7968 16346
rect 7672 16292 7728 16294
rect 7752 16292 7808 16294
rect 7832 16292 7888 16294
rect 7912 16292 7968 16294
rect 7562 15816 7618 15872
rect 7672 15258 7728 15260
rect 7752 15258 7808 15260
rect 7832 15258 7888 15260
rect 7912 15258 7968 15260
rect 7672 15206 7718 15258
rect 7718 15206 7728 15258
rect 7752 15206 7782 15258
rect 7782 15206 7794 15258
rect 7794 15206 7808 15258
rect 7832 15206 7846 15258
rect 7846 15206 7858 15258
rect 7858 15206 7888 15258
rect 7912 15206 7922 15258
rect 7922 15206 7968 15258
rect 7672 15204 7728 15206
rect 7752 15204 7808 15206
rect 7832 15204 7888 15206
rect 7912 15204 7968 15206
rect 9351 32122 9407 32124
rect 9431 32122 9487 32124
rect 9511 32122 9567 32124
rect 9591 32122 9647 32124
rect 9351 32070 9397 32122
rect 9397 32070 9407 32122
rect 9431 32070 9461 32122
rect 9461 32070 9473 32122
rect 9473 32070 9487 32122
rect 9511 32070 9525 32122
rect 9525 32070 9537 32122
rect 9537 32070 9567 32122
rect 9591 32070 9601 32122
rect 9601 32070 9647 32122
rect 9351 32068 9407 32070
rect 9431 32068 9487 32070
rect 9511 32068 9567 32070
rect 9591 32068 9647 32070
rect 8666 23568 8722 23624
rect 8574 21528 8630 21584
rect 8298 19352 8354 19408
rect 8206 18672 8262 18728
rect 7672 14170 7728 14172
rect 7752 14170 7808 14172
rect 7832 14170 7888 14172
rect 7912 14170 7968 14172
rect 7672 14118 7718 14170
rect 7718 14118 7728 14170
rect 7752 14118 7782 14170
rect 7782 14118 7794 14170
rect 7794 14118 7808 14170
rect 7832 14118 7846 14170
rect 7846 14118 7858 14170
rect 7858 14118 7888 14170
rect 7912 14118 7922 14170
rect 7922 14118 7968 14170
rect 7672 14116 7728 14118
rect 7752 14116 7808 14118
rect 7832 14116 7888 14118
rect 7912 14116 7968 14118
rect 7654 13912 7710 13968
rect 7562 13640 7618 13696
rect 7672 13082 7728 13084
rect 7752 13082 7808 13084
rect 7832 13082 7888 13084
rect 7912 13082 7968 13084
rect 7672 13030 7718 13082
rect 7718 13030 7728 13082
rect 7752 13030 7782 13082
rect 7782 13030 7794 13082
rect 7794 13030 7808 13082
rect 7832 13030 7846 13082
rect 7846 13030 7858 13082
rect 7858 13030 7888 13082
rect 7912 13030 7922 13082
rect 7922 13030 7968 13082
rect 7672 13028 7728 13030
rect 7752 13028 7808 13030
rect 7832 13028 7888 13030
rect 7912 13028 7968 13030
rect 5993 10362 6049 10364
rect 6073 10362 6129 10364
rect 6153 10362 6209 10364
rect 6233 10362 6289 10364
rect 5993 10310 6039 10362
rect 6039 10310 6049 10362
rect 6073 10310 6103 10362
rect 6103 10310 6115 10362
rect 6115 10310 6129 10362
rect 6153 10310 6167 10362
rect 6167 10310 6179 10362
rect 6179 10310 6209 10362
rect 6233 10310 6243 10362
rect 6243 10310 6289 10362
rect 5993 10308 6049 10310
rect 6073 10308 6129 10310
rect 6153 10308 6209 10310
rect 6233 10308 6289 10310
rect 5993 9274 6049 9276
rect 6073 9274 6129 9276
rect 6153 9274 6209 9276
rect 6233 9274 6289 9276
rect 5993 9222 6039 9274
rect 6039 9222 6049 9274
rect 6073 9222 6103 9274
rect 6103 9222 6115 9274
rect 6115 9222 6129 9274
rect 6153 9222 6167 9274
rect 6167 9222 6179 9274
rect 6179 9222 6209 9274
rect 6233 9222 6243 9274
rect 6243 9222 6289 9274
rect 5993 9220 6049 9222
rect 6073 9220 6129 9222
rect 6153 9220 6209 9222
rect 6233 9220 6289 9222
rect 5906 8508 5908 8528
rect 5908 8508 5960 8528
rect 5960 8508 5962 8528
rect 5906 8472 5962 8508
rect 5993 8186 6049 8188
rect 6073 8186 6129 8188
rect 6153 8186 6209 8188
rect 6233 8186 6289 8188
rect 5993 8134 6039 8186
rect 6039 8134 6049 8186
rect 6073 8134 6103 8186
rect 6103 8134 6115 8186
rect 6115 8134 6129 8186
rect 6153 8134 6167 8186
rect 6167 8134 6179 8186
rect 6179 8134 6209 8186
rect 6233 8134 6243 8186
rect 6243 8134 6289 8186
rect 5993 8132 6049 8134
rect 6073 8132 6129 8134
rect 6153 8132 6209 8134
rect 6233 8132 6289 8134
rect 5170 7248 5226 7304
rect 5993 7098 6049 7100
rect 6073 7098 6129 7100
rect 6153 7098 6209 7100
rect 6233 7098 6289 7100
rect 5993 7046 6039 7098
rect 6039 7046 6049 7098
rect 6073 7046 6103 7098
rect 6103 7046 6115 7098
rect 6115 7046 6129 7098
rect 6153 7046 6167 7098
rect 6167 7046 6179 7098
rect 6179 7046 6209 7098
rect 6233 7046 6243 7098
rect 6243 7046 6289 7098
rect 5993 7044 6049 7046
rect 6073 7044 6129 7046
rect 6153 7044 6209 7046
rect 6233 7044 6289 7046
rect 5993 6010 6049 6012
rect 6073 6010 6129 6012
rect 6153 6010 6209 6012
rect 6233 6010 6289 6012
rect 5993 5958 6039 6010
rect 6039 5958 6049 6010
rect 6073 5958 6103 6010
rect 6103 5958 6115 6010
rect 6115 5958 6129 6010
rect 6153 5958 6167 6010
rect 6167 5958 6179 6010
rect 6179 5958 6209 6010
rect 6233 5958 6243 6010
rect 6243 5958 6289 6010
rect 5993 5956 6049 5958
rect 6073 5956 6129 5958
rect 6153 5956 6209 5958
rect 6233 5956 6289 5958
rect 7672 11994 7728 11996
rect 7752 11994 7808 11996
rect 7832 11994 7888 11996
rect 7912 11994 7968 11996
rect 7672 11942 7718 11994
rect 7718 11942 7728 11994
rect 7752 11942 7782 11994
rect 7782 11942 7794 11994
rect 7794 11942 7808 11994
rect 7832 11942 7846 11994
rect 7846 11942 7858 11994
rect 7858 11942 7888 11994
rect 7912 11942 7922 11994
rect 7922 11942 7968 11994
rect 7672 11940 7728 11942
rect 7752 11940 7808 11942
rect 7832 11940 7888 11942
rect 7912 11940 7968 11942
rect 9351 31034 9407 31036
rect 9431 31034 9487 31036
rect 9511 31034 9567 31036
rect 9591 31034 9647 31036
rect 9351 30982 9397 31034
rect 9397 30982 9407 31034
rect 9431 30982 9461 31034
rect 9461 30982 9473 31034
rect 9473 30982 9487 31034
rect 9511 30982 9525 31034
rect 9525 30982 9537 31034
rect 9537 30982 9567 31034
rect 9591 30982 9601 31034
rect 9601 30982 9647 31034
rect 9351 30980 9407 30982
rect 9431 30980 9487 30982
rect 9511 30980 9567 30982
rect 9591 30980 9647 30982
rect 9862 33940 9864 33960
rect 9864 33940 9916 33960
rect 9916 33940 9918 33960
rect 9862 33904 9918 33940
rect 8942 28056 8998 28112
rect 8942 27820 8944 27840
rect 8944 27820 8996 27840
rect 8996 27820 8998 27840
rect 8942 27784 8998 27820
rect 9126 29008 9182 29064
rect 9351 29946 9407 29948
rect 9431 29946 9487 29948
rect 9511 29946 9567 29948
rect 9591 29946 9647 29948
rect 9351 29894 9397 29946
rect 9397 29894 9407 29946
rect 9431 29894 9461 29946
rect 9461 29894 9473 29946
rect 9473 29894 9487 29946
rect 9511 29894 9525 29946
rect 9525 29894 9537 29946
rect 9537 29894 9567 29946
rect 9591 29894 9601 29946
rect 9601 29894 9647 29946
rect 9351 29892 9407 29894
rect 9431 29892 9487 29894
rect 9511 29892 9567 29894
rect 9591 29892 9647 29894
rect 9034 27648 9090 27704
rect 9351 28858 9407 28860
rect 9431 28858 9487 28860
rect 9511 28858 9567 28860
rect 9591 28858 9647 28860
rect 9351 28806 9397 28858
rect 9397 28806 9407 28858
rect 9431 28806 9461 28858
rect 9461 28806 9473 28858
rect 9473 28806 9487 28858
rect 9511 28806 9525 28858
rect 9525 28806 9537 28858
rect 9537 28806 9567 28858
rect 9591 28806 9601 28858
rect 9601 28806 9647 28858
rect 9351 28804 9407 28806
rect 9431 28804 9487 28806
rect 9511 28804 9567 28806
rect 9591 28804 9647 28806
rect 9034 22480 9090 22536
rect 9678 27920 9734 27976
rect 9351 27770 9407 27772
rect 9431 27770 9487 27772
rect 9511 27770 9567 27772
rect 9591 27770 9647 27772
rect 9351 27718 9397 27770
rect 9397 27718 9407 27770
rect 9431 27718 9461 27770
rect 9461 27718 9473 27770
rect 9473 27718 9487 27770
rect 9511 27718 9525 27770
rect 9525 27718 9537 27770
rect 9537 27718 9567 27770
rect 9591 27718 9601 27770
rect 9601 27718 9647 27770
rect 9351 27716 9407 27718
rect 9431 27716 9487 27718
rect 9511 27716 9567 27718
rect 9591 27716 9647 27718
rect 9351 26682 9407 26684
rect 9431 26682 9487 26684
rect 9511 26682 9567 26684
rect 9591 26682 9647 26684
rect 9351 26630 9397 26682
rect 9397 26630 9407 26682
rect 9431 26630 9461 26682
rect 9461 26630 9473 26682
rect 9473 26630 9487 26682
rect 9511 26630 9525 26682
rect 9525 26630 9537 26682
rect 9537 26630 9567 26682
rect 9591 26630 9601 26682
rect 9601 26630 9647 26682
rect 9351 26628 9407 26630
rect 9431 26628 9487 26630
rect 9511 26628 9567 26630
rect 9591 26628 9647 26630
rect 9351 25594 9407 25596
rect 9431 25594 9487 25596
rect 9511 25594 9567 25596
rect 9591 25594 9647 25596
rect 9351 25542 9397 25594
rect 9397 25542 9407 25594
rect 9431 25542 9461 25594
rect 9461 25542 9473 25594
rect 9473 25542 9487 25594
rect 9511 25542 9525 25594
rect 9525 25542 9537 25594
rect 9537 25542 9567 25594
rect 9591 25542 9601 25594
rect 9601 25542 9647 25594
rect 9351 25540 9407 25542
rect 9431 25540 9487 25542
rect 9511 25540 9567 25542
rect 9591 25540 9647 25542
rect 9678 25200 9734 25256
rect 9351 24506 9407 24508
rect 9431 24506 9487 24508
rect 9511 24506 9567 24508
rect 9591 24506 9647 24508
rect 9351 24454 9397 24506
rect 9397 24454 9407 24506
rect 9431 24454 9461 24506
rect 9461 24454 9473 24506
rect 9473 24454 9487 24506
rect 9511 24454 9525 24506
rect 9525 24454 9537 24506
rect 9537 24454 9567 24506
rect 9591 24454 9601 24506
rect 9601 24454 9647 24506
rect 9351 24452 9407 24454
rect 9431 24452 9487 24454
rect 9511 24452 9567 24454
rect 9591 24452 9647 24454
rect 9678 23604 9680 23624
rect 9680 23604 9732 23624
rect 9732 23604 9734 23624
rect 9678 23568 9734 23604
rect 9351 23418 9407 23420
rect 9431 23418 9487 23420
rect 9511 23418 9567 23420
rect 9591 23418 9647 23420
rect 9351 23366 9397 23418
rect 9397 23366 9407 23418
rect 9431 23366 9461 23418
rect 9461 23366 9473 23418
rect 9473 23366 9487 23418
rect 9511 23366 9525 23418
rect 9525 23366 9537 23418
rect 9537 23366 9567 23418
rect 9591 23366 9601 23418
rect 9601 23366 9647 23418
rect 9351 23364 9407 23366
rect 9431 23364 9487 23366
rect 9511 23364 9567 23366
rect 9591 23364 9647 23366
rect 9351 22330 9407 22332
rect 9431 22330 9487 22332
rect 9511 22330 9567 22332
rect 9591 22330 9647 22332
rect 9351 22278 9397 22330
rect 9397 22278 9407 22330
rect 9431 22278 9461 22330
rect 9461 22278 9473 22330
rect 9473 22278 9487 22330
rect 9511 22278 9525 22330
rect 9525 22278 9537 22330
rect 9537 22278 9567 22330
rect 9591 22278 9601 22330
rect 9601 22278 9647 22330
rect 9351 22276 9407 22278
rect 9431 22276 9487 22278
rect 9511 22276 9567 22278
rect 9591 22276 9647 22278
rect 9402 21936 9458 21992
rect 8942 19916 8998 19952
rect 8942 19896 8944 19916
rect 8944 19896 8996 19916
rect 8996 19896 8998 19916
rect 8482 17992 8538 18048
rect 8850 19116 8852 19136
rect 8852 19116 8904 19136
rect 8904 19116 8906 19136
rect 8850 19080 8906 19116
rect 8758 18128 8814 18184
rect 7470 11056 7526 11112
rect 7102 7928 7158 7984
rect 7194 7792 7250 7848
rect 7286 7384 7342 7440
rect 5993 4922 6049 4924
rect 6073 4922 6129 4924
rect 6153 4922 6209 4924
rect 6233 4922 6289 4924
rect 5993 4870 6039 4922
rect 6039 4870 6049 4922
rect 6073 4870 6103 4922
rect 6103 4870 6115 4922
rect 6115 4870 6129 4922
rect 6153 4870 6167 4922
rect 6167 4870 6179 4922
rect 6179 4870 6209 4922
rect 6233 4870 6243 4922
rect 6243 4870 6289 4922
rect 5993 4868 6049 4870
rect 6073 4868 6129 4870
rect 6153 4868 6209 4870
rect 6233 4868 6289 4870
rect 5993 3834 6049 3836
rect 6073 3834 6129 3836
rect 6153 3834 6209 3836
rect 6233 3834 6289 3836
rect 5993 3782 6039 3834
rect 6039 3782 6049 3834
rect 6073 3782 6103 3834
rect 6103 3782 6115 3834
rect 6115 3782 6129 3834
rect 6153 3782 6167 3834
rect 6167 3782 6179 3834
rect 6179 3782 6209 3834
rect 6233 3782 6243 3834
rect 6243 3782 6289 3834
rect 5993 3780 6049 3782
rect 6073 3780 6129 3782
rect 6153 3780 6209 3782
rect 6233 3780 6289 3782
rect 4314 3290 4370 3292
rect 4394 3290 4450 3292
rect 4474 3290 4530 3292
rect 4554 3290 4610 3292
rect 4314 3238 4360 3290
rect 4360 3238 4370 3290
rect 4394 3238 4424 3290
rect 4424 3238 4436 3290
rect 4436 3238 4450 3290
rect 4474 3238 4488 3290
rect 4488 3238 4500 3290
rect 4500 3238 4530 3290
rect 4554 3238 4564 3290
rect 4564 3238 4610 3290
rect 4314 3236 4370 3238
rect 4394 3236 4450 3238
rect 4474 3236 4530 3238
rect 4554 3236 4610 3238
rect 5993 2746 6049 2748
rect 6073 2746 6129 2748
rect 6153 2746 6209 2748
rect 6233 2746 6289 2748
rect 5993 2694 6039 2746
rect 6039 2694 6049 2746
rect 6073 2694 6103 2746
rect 6103 2694 6115 2746
rect 6115 2694 6129 2746
rect 6153 2694 6167 2746
rect 6167 2694 6179 2746
rect 6179 2694 6209 2746
rect 6233 2694 6243 2746
rect 6243 2694 6289 2746
rect 5993 2692 6049 2694
rect 6073 2692 6129 2694
rect 6153 2692 6209 2694
rect 6233 2692 6289 2694
rect 6642 2624 6698 2680
rect 4314 2202 4370 2204
rect 4394 2202 4450 2204
rect 4474 2202 4530 2204
rect 4554 2202 4610 2204
rect 4314 2150 4360 2202
rect 4360 2150 4370 2202
rect 4394 2150 4424 2202
rect 4424 2150 4436 2202
rect 4436 2150 4450 2202
rect 4474 2150 4488 2202
rect 4488 2150 4500 2202
rect 4500 2150 4530 2202
rect 4554 2150 4564 2202
rect 4564 2150 4610 2202
rect 4314 2148 4370 2150
rect 4394 2148 4450 2150
rect 4474 2148 4530 2150
rect 4554 2148 4610 2150
rect 7194 2488 7250 2544
rect 7672 10906 7728 10908
rect 7752 10906 7808 10908
rect 7832 10906 7888 10908
rect 7912 10906 7968 10908
rect 7672 10854 7718 10906
rect 7718 10854 7728 10906
rect 7752 10854 7782 10906
rect 7782 10854 7794 10906
rect 7794 10854 7808 10906
rect 7832 10854 7846 10906
rect 7846 10854 7858 10906
rect 7858 10854 7888 10906
rect 7912 10854 7922 10906
rect 7922 10854 7968 10906
rect 7672 10852 7728 10854
rect 7752 10852 7808 10854
rect 7832 10852 7888 10854
rect 7912 10852 7968 10854
rect 7672 9818 7728 9820
rect 7752 9818 7808 9820
rect 7832 9818 7888 9820
rect 7912 9818 7968 9820
rect 7672 9766 7718 9818
rect 7718 9766 7728 9818
rect 7752 9766 7782 9818
rect 7782 9766 7794 9818
rect 7794 9766 7808 9818
rect 7832 9766 7846 9818
rect 7846 9766 7858 9818
rect 7858 9766 7888 9818
rect 7912 9766 7922 9818
rect 7922 9766 7968 9818
rect 7672 9764 7728 9766
rect 7752 9764 7808 9766
rect 7832 9764 7888 9766
rect 7912 9764 7968 9766
rect 7672 8730 7728 8732
rect 7752 8730 7808 8732
rect 7832 8730 7888 8732
rect 7912 8730 7968 8732
rect 7672 8678 7718 8730
rect 7718 8678 7728 8730
rect 7752 8678 7782 8730
rect 7782 8678 7794 8730
rect 7794 8678 7808 8730
rect 7832 8678 7846 8730
rect 7846 8678 7858 8730
rect 7858 8678 7888 8730
rect 7912 8678 7922 8730
rect 7922 8678 7968 8730
rect 7672 8676 7728 8678
rect 7752 8676 7808 8678
rect 7832 8676 7888 8678
rect 7912 8676 7968 8678
rect 8206 10648 8262 10704
rect 8574 13232 8630 13288
rect 8482 8744 8538 8800
rect 8022 8064 8078 8120
rect 7654 7792 7710 7848
rect 7672 7642 7728 7644
rect 7752 7642 7808 7644
rect 7832 7642 7888 7644
rect 7912 7642 7968 7644
rect 7672 7590 7718 7642
rect 7718 7590 7728 7642
rect 7752 7590 7782 7642
rect 7782 7590 7794 7642
rect 7794 7590 7808 7642
rect 7832 7590 7846 7642
rect 7846 7590 7858 7642
rect 7858 7590 7888 7642
rect 7912 7590 7922 7642
rect 7922 7590 7968 7642
rect 7672 7588 7728 7590
rect 7752 7588 7808 7590
rect 7832 7588 7888 7590
rect 7912 7588 7968 7590
rect 8114 7520 8170 7576
rect 7672 6554 7728 6556
rect 7752 6554 7808 6556
rect 7832 6554 7888 6556
rect 7912 6554 7968 6556
rect 7672 6502 7718 6554
rect 7718 6502 7728 6554
rect 7752 6502 7782 6554
rect 7782 6502 7794 6554
rect 7794 6502 7808 6554
rect 7832 6502 7846 6554
rect 7846 6502 7858 6554
rect 7858 6502 7888 6554
rect 7912 6502 7922 6554
rect 7922 6502 7968 6554
rect 7672 6500 7728 6502
rect 7752 6500 7808 6502
rect 7832 6500 7888 6502
rect 7912 6500 7968 6502
rect 8206 6160 8262 6216
rect 8298 5652 8300 5672
rect 8300 5652 8352 5672
rect 8352 5652 8354 5672
rect 8298 5616 8354 5652
rect 7672 5466 7728 5468
rect 7752 5466 7808 5468
rect 7832 5466 7888 5468
rect 7912 5466 7968 5468
rect 7672 5414 7718 5466
rect 7718 5414 7728 5466
rect 7752 5414 7782 5466
rect 7782 5414 7794 5466
rect 7794 5414 7808 5466
rect 7832 5414 7846 5466
rect 7846 5414 7858 5466
rect 7858 5414 7888 5466
rect 7912 5414 7922 5466
rect 7922 5414 7968 5466
rect 7672 5412 7728 5414
rect 7752 5412 7808 5414
rect 7832 5412 7888 5414
rect 7912 5412 7968 5414
rect 7672 4378 7728 4380
rect 7752 4378 7808 4380
rect 7832 4378 7888 4380
rect 7912 4378 7968 4380
rect 7672 4326 7718 4378
rect 7718 4326 7728 4378
rect 7752 4326 7782 4378
rect 7782 4326 7794 4378
rect 7794 4326 7808 4378
rect 7832 4326 7846 4378
rect 7846 4326 7858 4378
rect 7858 4326 7888 4378
rect 7912 4326 7922 4378
rect 7922 4326 7968 4378
rect 7672 4324 7728 4326
rect 7752 4324 7808 4326
rect 7832 4324 7888 4326
rect 7912 4324 7968 4326
rect 9351 21242 9407 21244
rect 9431 21242 9487 21244
rect 9511 21242 9567 21244
rect 9591 21242 9647 21244
rect 9351 21190 9397 21242
rect 9397 21190 9407 21242
rect 9431 21190 9461 21242
rect 9461 21190 9473 21242
rect 9473 21190 9487 21242
rect 9511 21190 9525 21242
rect 9525 21190 9537 21242
rect 9537 21190 9567 21242
rect 9591 21190 9601 21242
rect 9601 21190 9647 21242
rect 9351 21188 9407 21190
rect 9431 21188 9487 21190
rect 9511 21188 9567 21190
rect 9591 21188 9647 21190
rect 11030 35930 11086 35932
rect 11110 35930 11166 35932
rect 11190 35930 11246 35932
rect 11270 35930 11326 35932
rect 11030 35878 11076 35930
rect 11076 35878 11086 35930
rect 11110 35878 11140 35930
rect 11140 35878 11152 35930
rect 11152 35878 11166 35930
rect 11190 35878 11204 35930
rect 11204 35878 11216 35930
rect 11216 35878 11246 35930
rect 11270 35878 11280 35930
rect 11280 35878 11326 35930
rect 11030 35876 11086 35878
rect 11110 35876 11166 35878
rect 11190 35876 11246 35878
rect 11270 35876 11326 35878
rect 12709 38650 12765 38652
rect 12789 38650 12845 38652
rect 12869 38650 12925 38652
rect 12949 38650 13005 38652
rect 12709 38598 12755 38650
rect 12755 38598 12765 38650
rect 12789 38598 12819 38650
rect 12819 38598 12831 38650
rect 12831 38598 12845 38650
rect 12869 38598 12883 38650
rect 12883 38598 12895 38650
rect 12895 38598 12925 38650
rect 12949 38598 12959 38650
rect 12959 38598 13005 38650
rect 12709 38596 12765 38598
rect 12789 38596 12845 38598
rect 12869 38596 12925 38598
rect 12949 38596 13005 38598
rect 13910 38700 13912 38720
rect 13912 38700 13964 38720
rect 13964 38700 13966 38720
rect 13910 38664 13966 38700
rect 13358 38392 13414 38448
rect 12709 37562 12765 37564
rect 12789 37562 12845 37564
rect 12869 37562 12925 37564
rect 12949 37562 13005 37564
rect 12709 37510 12755 37562
rect 12755 37510 12765 37562
rect 12789 37510 12819 37562
rect 12819 37510 12831 37562
rect 12831 37510 12845 37562
rect 12869 37510 12883 37562
rect 12883 37510 12895 37562
rect 12895 37510 12925 37562
rect 12949 37510 12959 37562
rect 12959 37510 13005 37562
rect 12709 37508 12765 37510
rect 12789 37508 12845 37510
rect 12869 37508 12925 37510
rect 12949 37508 13005 37510
rect 12346 37168 12402 37224
rect 11030 34842 11086 34844
rect 11110 34842 11166 34844
rect 11190 34842 11246 34844
rect 11270 34842 11326 34844
rect 11030 34790 11076 34842
rect 11076 34790 11086 34842
rect 11110 34790 11140 34842
rect 11140 34790 11152 34842
rect 11152 34790 11166 34842
rect 11190 34790 11204 34842
rect 11204 34790 11216 34842
rect 11216 34790 11246 34842
rect 11270 34790 11280 34842
rect 11280 34790 11326 34842
rect 11030 34788 11086 34790
rect 11110 34788 11166 34790
rect 11190 34788 11246 34790
rect 11270 34788 11326 34790
rect 11334 34040 11390 34096
rect 11030 33754 11086 33756
rect 11110 33754 11166 33756
rect 11190 33754 11246 33756
rect 11270 33754 11326 33756
rect 11030 33702 11076 33754
rect 11076 33702 11086 33754
rect 11110 33702 11140 33754
rect 11140 33702 11152 33754
rect 11152 33702 11166 33754
rect 11190 33702 11204 33754
rect 11204 33702 11216 33754
rect 11216 33702 11246 33754
rect 11270 33702 11280 33754
rect 11280 33702 11326 33754
rect 11030 33700 11086 33702
rect 11110 33700 11166 33702
rect 11190 33700 11246 33702
rect 11270 33700 11326 33702
rect 10322 30776 10378 30832
rect 10046 28056 10102 28112
rect 9862 26424 9918 26480
rect 10046 25880 10102 25936
rect 10046 24148 10048 24168
rect 10048 24148 10100 24168
rect 10100 24148 10102 24168
rect 10046 24112 10102 24148
rect 9770 22480 9826 22536
rect 9678 20848 9734 20904
rect 9351 20154 9407 20156
rect 9431 20154 9487 20156
rect 9511 20154 9567 20156
rect 9591 20154 9647 20156
rect 9351 20102 9397 20154
rect 9397 20102 9407 20154
rect 9431 20102 9461 20154
rect 9461 20102 9473 20154
rect 9473 20102 9487 20154
rect 9511 20102 9525 20154
rect 9525 20102 9537 20154
rect 9537 20102 9567 20154
rect 9591 20102 9601 20154
rect 9601 20102 9647 20154
rect 9351 20100 9407 20102
rect 9431 20100 9487 20102
rect 9511 20100 9567 20102
rect 9591 20100 9647 20102
rect 9402 19216 9458 19272
rect 9351 19066 9407 19068
rect 9431 19066 9487 19068
rect 9511 19066 9567 19068
rect 9591 19066 9647 19068
rect 9351 19014 9397 19066
rect 9397 19014 9407 19066
rect 9431 19014 9461 19066
rect 9461 19014 9473 19066
rect 9473 19014 9487 19066
rect 9511 19014 9525 19066
rect 9525 19014 9537 19066
rect 9537 19014 9567 19066
rect 9591 19014 9601 19066
rect 9601 19014 9647 19066
rect 9351 19012 9407 19014
rect 9431 19012 9487 19014
rect 9511 19012 9567 19014
rect 9591 19012 9647 19014
rect 10230 23568 10286 23624
rect 10966 32852 10968 32872
rect 10968 32852 11020 32872
rect 11020 32852 11022 32872
rect 10966 32816 11022 32852
rect 11242 32816 11298 32872
rect 11030 32666 11086 32668
rect 11110 32666 11166 32668
rect 11190 32666 11246 32668
rect 11270 32666 11326 32668
rect 11030 32614 11076 32666
rect 11076 32614 11086 32666
rect 11110 32614 11140 32666
rect 11140 32614 11152 32666
rect 11152 32614 11166 32666
rect 11190 32614 11204 32666
rect 11204 32614 11216 32666
rect 11216 32614 11246 32666
rect 11270 32614 11280 32666
rect 11280 32614 11326 32666
rect 11030 32612 11086 32614
rect 11110 32612 11166 32614
rect 11190 32612 11246 32614
rect 11270 32612 11326 32614
rect 11030 31578 11086 31580
rect 11110 31578 11166 31580
rect 11190 31578 11246 31580
rect 11270 31578 11326 31580
rect 11030 31526 11076 31578
rect 11076 31526 11086 31578
rect 11110 31526 11140 31578
rect 11140 31526 11152 31578
rect 11152 31526 11166 31578
rect 11190 31526 11204 31578
rect 11204 31526 11216 31578
rect 11216 31526 11246 31578
rect 11270 31526 11280 31578
rect 11280 31526 11326 31578
rect 11030 31524 11086 31526
rect 11110 31524 11166 31526
rect 11190 31524 11246 31526
rect 11270 31524 11326 31526
rect 11030 30490 11086 30492
rect 11110 30490 11166 30492
rect 11190 30490 11246 30492
rect 11270 30490 11326 30492
rect 11030 30438 11076 30490
rect 11076 30438 11086 30490
rect 11110 30438 11140 30490
rect 11140 30438 11152 30490
rect 11152 30438 11166 30490
rect 11190 30438 11204 30490
rect 11204 30438 11216 30490
rect 11216 30438 11246 30490
rect 11270 30438 11280 30490
rect 11280 30438 11326 30490
rect 11030 30436 11086 30438
rect 11110 30436 11166 30438
rect 11190 30436 11246 30438
rect 11270 30436 11326 30438
rect 11030 29402 11086 29404
rect 11110 29402 11166 29404
rect 11190 29402 11246 29404
rect 11270 29402 11326 29404
rect 11030 29350 11076 29402
rect 11076 29350 11086 29402
rect 11110 29350 11140 29402
rect 11140 29350 11152 29402
rect 11152 29350 11166 29402
rect 11190 29350 11204 29402
rect 11204 29350 11216 29402
rect 11216 29350 11246 29402
rect 11270 29350 11280 29402
rect 11280 29350 11326 29402
rect 11030 29348 11086 29350
rect 11110 29348 11166 29350
rect 11190 29348 11246 29350
rect 11270 29348 11326 29350
rect 10690 28464 10746 28520
rect 11058 29164 11114 29200
rect 11058 29144 11060 29164
rect 11060 29144 11112 29164
rect 11112 29144 11114 29164
rect 11426 28600 11482 28656
rect 10690 27512 10746 27568
rect 10046 21292 10048 21312
rect 10048 21292 10100 21312
rect 10100 21292 10102 21312
rect 10046 21256 10102 21292
rect 9770 19352 9826 19408
rect 9862 18264 9918 18320
rect 9351 17978 9407 17980
rect 9431 17978 9487 17980
rect 9511 17978 9567 17980
rect 9591 17978 9647 17980
rect 9351 17926 9397 17978
rect 9397 17926 9407 17978
rect 9431 17926 9461 17978
rect 9461 17926 9473 17978
rect 9473 17926 9487 17978
rect 9511 17926 9525 17978
rect 9525 17926 9537 17978
rect 9537 17926 9567 17978
rect 9591 17926 9601 17978
rect 9601 17926 9647 17978
rect 9351 17924 9407 17926
rect 9431 17924 9487 17926
rect 9511 17924 9567 17926
rect 9591 17924 9647 17926
rect 9862 18128 9918 18184
rect 9770 17856 9826 17912
rect 9351 16890 9407 16892
rect 9431 16890 9487 16892
rect 9511 16890 9567 16892
rect 9591 16890 9647 16892
rect 9351 16838 9397 16890
rect 9397 16838 9407 16890
rect 9431 16838 9461 16890
rect 9461 16838 9473 16890
rect 9473 16838 9487 16890
rect 9511 16838 9525 16890
rect 9525 16838 9537 16890
rect 9537 16838 9567 16890
rect 9591 16838 9601 16890
rect 9601 16838 9647 16890
rect 9351 16836 9407 16838
rect 9431 16836 9487 16838
rect 9511 16836 9567 16838
rect 9591 16836 9647 16838
rect 9034 13232 9090 13288
rect 8850 11192 8906 11248
rect 9034 10920 9090 10976
rect 9678 16496 9734 16552
rect 9351 15802 9407 15804
rect 9431 15802 9487 15804
rect 9511 15802 9567 15804
rect 9591 15802 9647 15804
rect 9351 15750 9397 15802
rect 9397 15750 9407 15802
rect 9431 15750 9461 15802
rect 9461 15750 9473 15802
rect 9473 15750 9487 15802
rect 9511 15750 9525 15802
rect 9525 15750 9537 15802
rect 9537 15750 9567 15802
rect 9591 15750 9601 15802
rect 9601 15750 9647 15802
rect 9351 15748 9407 15750
rect 9431 15748 9487 15750
rect 9511 15748 9567 15750
rect 9591 15748 9647 15750
rect 9678 15544 9734 15600
rect 9862 15000 9918 15056
rect 9351 14714 9407 14716
rect 9431 14714 9487 14716
rect 9511 14714 9567 14716
rect 9591 14714 9647 14716
rect 9351 14662 9397 14714
rect 9397 14662 9407 14714
rect 9431 14662 9461 14714
rect 9461 14662 9473 14714
rect 9473 14662 9487 14714
rect 9511 14662 9525 14714
rect 9525 14662 9537 14714
rect 9537 14662 9567 14714
rect 9591 14662 9601 14714
rect 9601 14662 9647 14714
rect 9351 14660 9407 14662
rect 9431 14660 9487 14662
rect 9511 14660 9567 14662
rect 9591 14660 9647 14662
rect 9770 14728 9826 14784
rect 9678 14184 9734 14240
rect 9351 13626 9407 13628
rect 9431 13626 9487 13628
rect 9511 13626 9567 13628
rect 9591 13626 9647 13628
rect 9351 13574 9397 13626
rect 9397 13574 9407 13626
rect 9431 13574 9461 13626
rect 9461 13574 9473 13626
rect 9473 13574 9487 13626
rect 9511 13574 9525 13626
rect 9525 13574 9537 13626
rect 9537 13574 9567 13626
rect 9591 13574 9601 13626
rect 9601 13574 9647 13626
rect 9351 13572 9407 13574
rect 9431 13572 9487 13574
rect 9511 13572 9567 13574
rect 9591 13572 9647 13574
rect 9402 13368 9458 13424
rect 9351 12538 9407 12540
rect 9431 12538 9487 12540
rect 9511 12538 9567 12540
rect 9591 12538 9647 12540
rect 9351 12486 9397 12538
rect 9397 12486 9407 12538
rect 9431 12486 9461 12538
rect 9461 12486 9473 12538
rect 9473 12486 9487 12538
rect 9511 12486 9525 12538
rect 9525 12486 9537 12538
rect 9537 12486 9567 12538
rect 9591 12486 9601 12538
rect 9601 12486 9647 12538
rect 9351 12484 9407 12486
rect 9431 12484 9487 12486
rect 9511 12484 9567 12486
rect 9591 12484 9647 12486
rect 9402 12280 9458 12336
rect 9351 11450 9407 11452
rect 9431 11450 9487 11452
rect 9511 11450 9567 11452
rect 9591 11450 9647 11452
rect 9351 11398 9397 11450
rect 9397 11398 9407 11450
rect 9431 11398 9461 11450
rect 9461 11398 9473 11450
rect 9473 11398 9487 11450
rect 9511 11398 9525 11450
rect 9525 11398 9537 11450
rect 9537 11398 9567 11450
rect 9591 11398 9601 11450
rect 9601 11398 9647 11450
rect 9351 11396 9407 11398
rect 9431 11396 9487 11398
rect 9511 11396 9567 11398
rect 9591 11396 9647 11398
rect 9402 10512 9458 10568
rect 9351 10362 9407 10364
rect 9431 10362 9487 10364
rect 9511 10362 9567 10364
rect 9591 10362 9647 10364
rect 9351 10310 9397 10362
rect 9397 10310 9407 10362
rect 9431 10310 9461 10362
rect 9461 10310 9473 10362
rect 9473 10310 9487 10362
rect 9511 10310 9525 10362
rect 9525 10310 9537 10362
rect 9537 10310 9567 10362
rect 9591 10310 9601 10362
rect 9601 10310 9647 10362
rect 9351 10308 9407 10310
rect 9431 10308 9487 10310
rect 9511 10308 9567 10310
rect 9591 10308 9647 10310
rect 9586 9424 9642 9480
rect 9351 9274 9407 9276
rect 9431 9274 9487 9276
rect 9511 9274 9567 9276
rect 9591 9274 9647 9276
rect 9351 9222 9397 9274
rect 9397 9222 9407 9274
rect 9431 9222 9461 9274
rect 9461 9222 9473 9274
rect 9473 9222 9487 9274
rect 9511 9222 9525 9274
rect 9525 9222 9537 9274
rect 9537 9222 9567 9274
rect 9591 9222 9601 9274
rect 9601 9222 9647 9274
rect 9351 9220 9407 9222
rect 9431 9220 9487 9222
rect 9511 9220 9567 9222
rect 9591 9220 9647 9222
rect 9351 8186 9407 8188
rect 9431 8186 9487 8188
rect 9511 8186 9567 8188
rect 9591 8186 9647 8188
rect 9351 8134 9397 8186
rect 9397 8134 9407 8186
rect 9431 8134 9461 8186
rect 9461 8134 9473 8186
rect 9473 8134 9487 8186
rect 9511 8134 9525 8186
rect 9525 8134 9537 8186
rect 9537 8134 9567 8186
rect 9591 8134 9601 8186
rect 9601 8134 9647 8186
rect 9351 8132 9407 8134
rect 9431 8132 9487 8134
rect 9511 8132 9567 8134
rect 9591 8132 9647 8134
rect 7672 3290 7728 3292
rect 7752 3290 7808 3292
rect 7832 3290 7888 3292
rect 7912 3290 7968 3292
rect 7672 3238 7718 3290
rect 7718 3238 7728 3290
rect 7752 3238 7782 3290
rect 7782 3238 7794 3290
rect 7794 3238 7808 3290
rect 7832 3238 7846 3290
rect 7846 3238 7858 3290
rect 7858 3238 7888 3290
rect 7912 3238 7922 3290
rect 7922 3238 7968 3290
rect 7672 3236 7728 3238
rect 7752 3236 7808 3238
rect 7832 3236 7888 3238
rect 7912 3236 7968 3238
rect 8666 2352 8722 2408
rect 7672 2202 7728 2204
rect 7752 2202 7808 2204
rect 7832 2202 7888 2204
rect 7912 2202 7968 2204
rect 7672 2150 7718 2202
rect 7718 2150 7728 2202
rect 7752 2150 7782 2202
rect 7782 2150 7794 2202
rect 7794 2150 7808 2202
rect 7832 2150 7846 2202
rect 7846 2150 7858 2202
rect 7858 2150 7888 2202
rect 7912 2150 7922 2202
rect 7922 2150 7968 2202
rect 7672 2148 7728 2150
rect 7752 2148 7808 2150
rect 7832 2148 7888 2150
rect 7912 2148 7968 2150
rect 2635 1658 2691 1660
rect 2715 1658 2771 1660
rect 2795 1658 2851 1660
rect 2875 1658 2931 1660
rect 2635 1606 2681 1658
rect 2681 1606 2691 1658
rect 2715 1606 2745 1658
rect 2745 1606 2757 1658
rect 2757 1606 2771 1658
rect 2795 1606 2809 1658
rect 2809 1606 2821 1658
rect 2821 1606 2851 1658
rect 2875 1606 2885 1658
rect 2885 1606 2931 1658
rect 2635 1604 2691 1606
rect 2715 1604 2771 1606
rect 2795 1604 2851 1606
rect 2875 1604 2931 1606
rect 5993 1658 6049 1660
rect 6073 1658 6129 1660
rect 6153 1658 6209 1660
rect 6233 1658 6289 1660
rect 5993 1606 6039 1658
rect 6039 1606 6049 1658
rect 6073 1606 6103 1658
rect 6103 1606 6115 1658
rect 6115 1606 6129 1658
rect 6153 1606 6167 1658
rect 6167 1606 6179 1658
rect 6179 1606 6209 1658
rect 6233 1606 6243 1658
rect 6243 1606 6289 1658
rect 5993 1604 6049 1606
rect 6073 1604 6129 1606
rect 6153 1604 6209 1606
rect 6233 1604 6289 1606
rect 9862 8608 9918 8664
rect 9862 7928 9918 7984
rect 9678 7792 9734 7848
rect 9494 7656 9550 7712
rect 9310 7520 9366 7576
rect 9494 7384 9550 7440
rect 9632 7418 9688 7474
rect 9770 7384 9826 7440
rect 9678 7284 9680 7304
rect 9680 7284 9732 7304
rect 9732 7284 9734 7304
rect 9678 7248 9734 7284
rect 9351 7098 9407 7100
rect 9431 7098 9487 7100
rect 9511 7098 9567 7100
rect 9591 7098 9647 7100
rect 9351 7046 9397 7098
rect 9397 7046 9407 7098
rect 9431 7046 9461 7098
rect 9461 7046 9473 7098
rect 9473 7046 9487 7098
rect 9511 7046 9525 7098
rect 9525 7046 9537 7098
rect 9537 7046 9567 7098
rect 9591 7046 9601 7098
rect 9601 7046 9647 7098
rect 9351 7044 9407 7046
rect 9431 7044 9487 7046
rect 9511 7044 9567 7046
rect 9591 7044 9647 7046
rect 9310 6840 9366 6896
rect 9770 6976 9826 7032
rect 10598 22480 10654 22536
rect 11030 28314 11086 28316
rect 11110 28314 11166 28316
rect 11190 28314 11246 28316
rect 11270 28314 11326 28316
rect 11030 28262 11076 28314
rect 11076 28262 11086 28314
rect 11110 28262 11140 28314
rect 11140 28262 11152 28314
rect 11152 28262 11166 28314
rect 11190 28262 11204 28314
rect 11204 28262 11216 28314
rect 11216 28262 11246 28314
rect 11270 28262 11280 28314
rect 11280 28262 11326 28314
rect 11030 28260 11086 28262
rect 11110 28260 11166 28262
rect 11190 28260 11246 28262
rect 11270 28260 11326 28262
rect 11030 27226 11086 27228
rect 11110 27226 11166 27228
rect 11190 27226 11246 27228
rect 11270 27226 11326 27228
rect 11030 27174 11076 27226
rect 11076 27174 11086 27226
rect 11110 27174 11140 27226
rect 11140 27174 11152 27226
rect 11152 27174 11166 27226
rect 11190 27174 11204 27226
rect 11204 27174 11216 27226
rect 11216 27174 11246 27226
rect 11270 27174 11280 27226
rect 11280 27174 11326 27226
rect 11030 27172 11086 27174
rect 11110 27172 11166 27174
rect 11190 27172 11246 27174
rect 11270 27172 11326 27174
rect 11030 26138 11086 26140
rect 11110 26138 11166 26140
rect 11190 26138 11246 26140
rect 11270 26138 11326 26140
rect 11030 26086 11076 26138
rect 11076 26086 11086 26138
rect 11110 26086 11140 26138
rect 11140 26086 11152 26138
rect 11152 26086 11166 26138
rect 11190 26086 11204 26138
rect 11204 26086 11216 26138
rect 11216 26086 11246 26138
rect 11270 26086 11280 26138
rect 11280 26086 11326 26138
rect 11030 26084 11086 26086
rect 11110 26084 11166 26086
rect 11190 26084 11246 26086
rect 11270 26084 11326 26086
rect 11426 25336 11482 25392
rect 10966 25200 11022 25256
rect 11030 25050 11086 25052
rect 11110 25050 11166 25052
rect 11190 25050 11246 25052
rect 11270 25050 11326 25052
rect 11030 24998 11076 25050
rect 11076 24998 11086 25050
rect 11110 24998 11140 25050
rect 11140 24998 11152 25050
rect 11152 24998 11166 25050
rect 11190 24998 11204 25050
rect 11204 24998 11216 25050
rect 11216 24998 11246 25050
rect 11270 24998 11280 25050
rect 11280 24998 11326 25050
rect 11030 24996 11086 24998
rect 11110 24996 11166 24998
rect 11190 24996 11246 24998
rect 11270 24996 11326 24998
rect 11426 24112 11482 24168
rect 11030 23962 11086 23964
rect 11110 23962 11166 23964
rect 11190 23962 11246 23964
rect 11270 23962 11326 23964
rect 11030 23910 11076 23962
rect 11076 23910 11086 23962
rect 11110 23910 11140 23962
rect 11140 23910 11152 23962
rect 11152 23910 11166 23962
rect 11190 23910 11204 23962
rect 11204 23910 11216 23962
rect 11216 23910 11246 23962
rect 11270 23910 11280 23962
rect 11280 23910 11326 23962
rect 11030 23908 11086 23910
rect 11110 23908 11166 23910
rect 11190 23908 11246 23910
rect 11270 23908 11326 23910
rect 11030 22874 11086 22876
rect 11110 22874 11166 22876
rect 11190 22874 11246 22876
rect 11270 22874 11326 22876
rect 11030 22822 11076 22874
rect 11076 22822 11086 22874
rect 11110 22822 11140 22874
rect 11140 22822 11152 22874
rect 11152 22822 11166 22874
rect 11190 22822 11204 22874
rect 11204 22822 11216 22874
rect 11216 22822 11246 22874
rect 11270 22822 11280 22874
rect 11280 22822 11326 22874
rect 11030 22820 11086 22822
rect 11110 22820 11166 22822
rect 11190 22820 11246 22822
rect 11270 22820 11326 22822
rect 11030 21786 11086 21788
rect 11110 21786 11166 21788
rect 11190 21786 11246 21788
rect 11270 21786 11326 21788
rect 11030 21734 11076 21786
rect 11076 21734 11086 21786
rect 11110 21734 11140 21786
rect 11140 21734 11152 21786
rect 11152 21734 11166 21786
rect 11190 21734 11204 21786
rect 11204 21734 11216 21786
rect 11216 21734 11246 21786
rect 11270 21734 11280 21786
rect 11280 21734 11326 21786
rect 11030 21732 11086 21734
rect 11110 21732 11166 21734
rect 11190 21732 11246 21734
rect 11270 21732 11326 21734
rect 11030 20698 11086 20700
rect 11110 20698 11166 20700
rect 11190 20698 11246 20700
rect 11270 20698 11326 20700
rect 11030 20646 11076 20698
rect 11076 20646 11086 20698
rect 11110 20646 11140 20698
rect 11140 20646 11152 20698
rect 11152 20646 11166 20698
rect 11190 20646 11204 20698
rect 11204 20646 11216 20698
rect 11216 20646 11246 20698
rect 11270 20646 11280 20698
rect 11280 20646 11326 20698
rect 11030 20644 11086 20646
rect 11110 20644 11166 20646
rect 11190 20644 11246 20646
rect 11270 20644 11326 20646
rect 10506 17720 10562 17776
rect 11030 19610 11086 19612
rect 11110 19610 11166 19612
rect 11190 19610 11246 19612
rect 11270 19610 11326 19612
rect 11030 19558 11076 19610
rect 11076 19558 11086 19610
rect 11110 19558 11140 19610
rect 11140 19558 11152 19610
rect 11152 19558 11166 19610
rect 11190 19558 11204 19610
rect 11204 19558 11216 19610
rect 11216 19558 11246 19610
rect 11270 19558 11280 19610
rect 11280 19558 11326 19610
rect 11030 19556 11086 19558
rect 11110 19556 11166 19558
rect 11190 19556 11246 19558
rect 11270 19556 11326 19558
rect 11242 19352 11298 19408
rect 10690 18808 10746 18864
rect 11030 18522 11086 18524
rect 11110 18522 11166 18524
rect 11190 18522 11246 18524
rect 11270 18522 11326 18524
rect 11030 18470 11076 18522
rect 11076 18470 11086 18522
rect 11110 18470 11140 18522
rect 11140 18470 11152 18522
rect 11152 18470 11166 18522
rect 11190 18470 11204 18522
rect 11204 18470 11216 18522
rect 11216 18470 11246 18522
rect 11270 18470 11280 18522
rect 11280 18470 11326 18522
rect 11030 18468 11086 18470
rect 11110 18468 11166 18470
rect 11190 18468 11246 18470
rect 11270 18468 11326 18470
rect 10322 14728 10378 14784
rect 10322 14592 10378 14648
rect 10230 12280 10286 12336
rect 10598 14456 10654 14512
rect 10322 11056 10378 11112
rect 12070 33904 12126 33960
rect 12714 36896 12770 36952
rect 13358 37032 13414 37088
rect 13726 36760 13782 36816
rect 12709 36474 12765 36476
rect 12789 36474 12845 36476
rect 12869 36474 12925 36476
rect 12949 36474 13005 36476
rect 12709 36422 12755 36474
rect 12755 36422 12765 36474
rect 12789 36422 12819 36474
rect 12819 36422 12831 36474
rect 12831 36422 12845 36474
rect 12869 36422 12883 36474
rect 12883 36422 12895 36474
rect 12895 36422 12925 36474
rect 12949 36422 12959 36474
rect 12959 36422 13005 36474
rect 12709 36420 12765 36422
rect 12789 36420 12845 36422
rect 12869 36420 12925 36422
rect 12949 36420 13005 36422
rect 12622 35672 12678 35728
rect 12714 35536 12770 35592
rect 13174 35400 13230 35456
rect 12709 35386 12765 35388
rect 12789 35386 12845 35388
rect 12869 35386 12925 35388
rect 12949 35386 13005 35388
rect 12709 35334 12755 35386
rect 12755 35334 12765 35386
rect 12789 35334 12819 35386
rect 12819 35334 12831 35386
rect 12831 35334 12845 35386
rect 12869 35334 12883 35386
rect 12883 35334 12895 35386
rect 12895 35334 12925 35386
rect 12949 35334 12959 35386
rect 12959 35334 13005 35386
rect 12709 35332 12765 35334
rect 12789 35332 12845 35334
rect 12869 35332 12925 35334
rect 12949 35332 13005 35334
rect 13082 34584 13138 34640
rect 12709 34298 12765 34300
rect 12789 34298 12845 34300
rect 12869 34298 12925 34300
rect 12949 34298 13005 34300
rect 12709 34246 12755 34298
rect 12755 34246 12765 34298
rect 12789 34246 12819 34298
rect 12819 34246 12831 34298
rect 12831 34246 12845 34298
rect 12869 34246 12883 34298
rect 12883 34246 12895 34298
rect 12895 34246 12925 34298
rect 12949 34246 12959 34298
rect 12959 34246 13005 34298
rect 12709 34244 12765 34246
rect 12789 34244 12845 34246
rect 12869 34244 12925 34246
rect 12949 34244 13005 34246
rect 11794 30912 11850 30968
rect 11794 30676 11796 30696
rect 11796 30676 11848 30696
rect 11848 30676 11850 30696
rect 11794 30640 11850 30676
rect 11886 30368 11942 30424
rect 11610 29144 11666 29200
rect 12346 32952 12402 33008
rect 12254 32272 12310 32328
rect 12709 33210 12765 33212
rect 12789 33210 12845 33212
rect 12869 33210 12925 33212
rect 12949 33210 13005 33212
rect 12709 33158 12755 33210
rect 12755 33158 12765 33210
rect 12789 33158 12819 33210
rect 12819 33158 12831 33210
rect 12831 33158 12845 33210
rect 12869 33158 12883 33210
rect 12883 33158 12895 33210
rect 12895 33158 12925 33210
rect 12949 33158 12959 33210
rect 12959 33158 13005 33210
rect 12709 33156 12765 33158
rect 12789 33156 12845 33158
rect 12869 33156 12925 33158
rect 12949 33156 13005 33158
rect 13634 36488 13690 36544
rect 14388 41370 14444 41372
rect 14468 41370 14524 41372
rect 14548 41370 14604 41372
rect 14628 41370 14684 41372
rect 14388 41318 14434 41370
rect 14434 41318 14444 41370
rect 14468 41318 14498 41370
rect 14498 41318 14510 41370
rect 14510 41318 14524 41370
rect 14548 41318 14562 41370
rect 14562 41318 14574 41370
rect 14574 41318 14604 41370
rect 14628 41318 14638 41370
rect 14638 41318 14684 41370
rect 14388 41316 14444 41318
rect 14468 41316 14524 41318
rect 14548 41316 14604 41318
rect 14628 41316 14684 41318
rect 14388 40282 14444 40284
rect 14468 40282 14524 40284
rect 14548 40282 14604 40284
rect 14628 40282 14684 40284
rect 14388 40230 14434 40282
rect 14434 40230 14444 40282
rect 14468 40230 14498 40282
rect 14498 40230 14510 40282
rect 14510 40230 14524 40282
rect 14548 40230 14562 40282
rect 14562 40230 14574 40282
rect 14574 40230 14604 40282
rect 14628 40230 14638 40282
rect 14638 40230 14684 40282
rect 14388 40228 14444 40230
rect 14468 40228 14524 40230
rect 14548 40228 14604 40230
rect 14628 40228 14684 40230
rect 14094 39480 14150 39536
rect 14388 39194 14444 39196
rect 14468 39194 14524 39196
rect 14548 39194 14604 39196
rect 14628 39194 14684 39196
rect 14388 39142 14434 39194
rect 14434 39142 14444 39194
rect 14468 39142 14498 39194
rect 14498 39142 14510 39194
rect 14510 39142 14524 39194
rect 14548 39142 14562 39194
rect 14562 39142 14574 39194
rect 14574 39142 14604 39194
rect 14628 39142 14638 39194
rect 14638 39142 14684 39194
rect 14388 39140 14444 39142
rect 14468 39140 14524 39142
rect 14548 39140 14604 39142
rect 14628 39140 14684 39142
rect 14278 38936 14334 38992
rect 14388 38106 14444 38108
rect 14468 38106 14524 38108
rect 14548 38106 14604 38108
rect 14628 38106 14684 38108
rect 14388 38054 14434 38106
rect 14434 38054 14444 38106
rect 14468 38054 14498 38106
rect 14498 38054 14510 38106
rect 14510 38054 14524 38106
rect 14548 38054 14562 38106
rect 14562 38054 14574 38106
rect 14574 38054 14604 38106
rect 14628 38054 14638 38106
rect 14638 38054 14684 38106
rect 14388 38052 14444 38054
rect 14468 38052 14524 38054
rect 14548 38052 14604 38054
rect 14628 38052 14684 38054
rect 14278 37848 14334 37904
rect 14370 37576 14426 37632
rect 14186 37304 14242 37360
rect 14388 37018 14444 37020
rect 14468 37018 14524 37020
rect 14548 37018 14604 37020
rect 14628 37018 14684 37020
rect 14388 36966 14434 37018
rect 14434 36966 14444 37018
rect 14468 36966 14498 37018
rect 14498 36966 14510 37018
rect 14510 36966 14524 37018
rect 14548 36966 14562 37018
rect 14562 36966 14574 37018
rect 14574 36966 14604 37018
rect 14628 36966 14638 37018
rect 14638 36966 14684 37018
rect 14388 36964 14444 36966
rect 14468 36964 14524 36966
rect 14548 36964 14604 36966
rect 14628 36964 14684 36966
rect 14830 39208 14886 39264
rect 14830 38120 14886 38176
rect 14186 36216 14242 36272
rect 14388 35930 14444 35932
rect 14468 35930 14524 35932
rect 14548 35930 14604 35932
rect 14628 35930 14684 35932
rect 14388 35878 14434 35930
rect 14434 35878 14444 35930
rect 14468 35878 14498 35930
rect 14498 35878 14510 35930
rect 14510 35878 14524 35930
rect 14548 35878 14562 35930
rect 14562 35878 14574 35930
rect 14574 35878 14604 35930
rect 14628 35878 14638 35930
rect 14638 35878 14684 35930
rect 14388 35876 14444 35878
rect 14468 35876 14524 35878
rect 14548 35876 14604 35878
rect 14628 35876 14684 35878
rect 13726 34992 13782 35048
rect 13542 34584 13598 34640
rect 13266 34176 13322 34232
rect 12898 32408 12954 32464
rect 13450 34312 13506 34368
rect 13358 33088 13414 33144
rect 14002 35128 14058 35184
rect 13726 34176 13782 34232
rect 13726 33904 13782 33960
rect 13634 33496 13690 33552
rect 13450 32816 13506 32872
rect 12709 32122 12765 32124
rect 12789 32122 12845 32124
rect 12869 32122 12925 32124
rect 12949 32122 13005 32124
rect 12709 32070 12755 32122
rect 12755 32070 12765 32122
rect 12789 32070 12819 32122
rect 12819 32070 12831 32122
rect 12831 32070 12845 32122
rect 12869 32070 12883 32122
rect 12883 32070 12895 32122
rect 12895 32070 12925 32122
rect 12949 32070 12959 32122
rect 12959 32070 13005 32122
rect 12709 32068 12765 32070
rect 12789 32068 12845 32070
rect 12869 32068 12925 32070
rect 12949 32068 13005 32070
rect 12530 30912 12586 30968
rect 12254 30776 12310 30832
rect 11978 28736 12034 28792
rect 11610 26832 11666 26888
rect 11610 26696 11666 26752
rect 11978 27784 12034 27840
rect 11886 27412 11888 27432
rect 11888 27412 11940 27432
rect 11940 27412 11942 27432
rect 11886 27376 11942 27412
rect 11610 23160 11666 23216
rect 11610 23024 11666 23080
rect 11886 25336 11942 25392
rect 11610 20304 11666 20360
rect 12070 26968 12126 27024
rect 12254 28908 12256 28928
rect 12256 28908 12308 28928
rect 12308 28908 12310 28928
rect 12254 28872 12310 28908
rect 12254 28756 12310 28792
rect 12254 28736 12256 28756
rect 12256 28736 12308 28756
rect 12308 28736 12310 28756
rect 12346 28056 12402 28112
rect 12346 27648 12402 27704
rect 12990 31184 13046 31240
rect 12709 31034 12765 31036
rect 12789 31034 12845 31036
rect 12869 31034 12925 31036
rect 12949 31034 13005 31036
rect 12709 30982 12755 31034
rect 12755 30982 12765 31034
rect 12789 30982 12819 31034
rect 12819 30982 12831 31034
rect 12831 30982 12845 31034
rect 12869 30982 12883 31034
rect 12883 30982 12895 31034
rect 12895 30982 12925 31034
rect 12949 30982 12959 31034
rect 12959 30982 13005 31034
rect 12709 30980 12765 30982
rect 12789 30980 12845 30982
rect 12869 30980 12925 30982
rect 12949 30980 13005 30982
rect 13450 31864 13506 31920
rect 13634 31864 13690 31920
rect 13266 31320 13322 31376
rect 12530 29552 12586 29608
rect 12709 29946 12765 29948
rect 12789 29946 12845 29948
rect 12869 29946 12925 29948
rect 12949 29946 13005 29948
rect 12709 29894 12755 29946
rect 12755 29894 12765 29946
rect 12789 29894 12819 29946
rect 12819 29894 12831 29946
rect 12831 29894 12845 29946
rect 12869 29894 12883 29946
rect 12883 29894 12895 29946
rect 12895 29894 12925 29946
rect 12949 29894 12959 29946
rect 12959 29894 13005 29946
rect 12709 29892 12765 29894
rect 12789 29892 12845 29894
rect 12869 29892 12925 29894
rect 12949 29892 13005 29894
rect 12709 28858 12765 28860
rect 12789 28858 12845 28860
rect 12869 28858 12925 28860
rect 12949 28858 13005 28860
rect 12709 28806 12755 28858
rect 12755 28806 12765 28858
rect 12789 28806 12819 28858
rect 12819 28806 12831 28858
rect 12831 28806 12845 28858
rect 12869 28806 12883 28858
rect 12883 28806 12895 28858
rect 12895 28806 12925 28858
rect 12949 28806 12959 28858
rect 12959 28806 13005 28858
rect 12709 28804 12765 28806
rect 12789 28804 12845 28806
rect 12869 28804 12925 28806
rect 12949 28804 13005 28806
rect 12530 28736 12586 28792
rect 12714 28500 12716 28520
rect 12716 28500 12768 28520
rect 12768 28500 12770 28520
rect 12714 28464 12770 28500
rect 12530 27376 12586 27432
rect 12709 27770 12765 27772
rect 12789 27770 12845 27772
rect 12869 27770 12925 27772
rect 12949 27770 13005 27772
rect 12709 27718 12755 27770
rect 12755 27718 12765 27770
rect 12789 27718 12819 27770
rect 12819 27718 12831 27770
rect 12831 27718 12845 27770
rect 12869 27718 12883 27770
rect 12883 27718 12895 27770
rect 12895 27718 12925 27770
rect 12949 27718 12959 27770
rect 12959 27718 13005 27770
rect 12709 27716 12765 27718
rect 12789 27716 12845 27718
rect 12869 27716 12925 27718
rect 12949 27716 13005 27718
rect 12709 26682 12765 26684
rect 12789 26682 12845 26684
rect 12869 26682 12925 26684
rect 12949 26682 13005 26684
rect 12709 26630 12755 26682
rect 12755 26630 12765 26682
rect 12789 26630 12819 26682
rect 12819 26630 12831 26682
rect 12831 26630 12845 26682
rect 12869 26630 12883 26682
rect 12883 26630 12895 26682
rect 12895 26630 12925 26682
rect 12949 26630 12959 26682
rect 12959 26630 13005 26682
rect 12709 26628 12765 26630
rect 12789 26628 12845 26630
rect 12869 26628 12925 26630
rect 12949 26628 13005 26630
rect 12438 25900 12494 25936
rect 12438 25880 12440 25900
rect 12440 25880 12492 25900
rect 12492 25880 12494 25900
rect 12254 23568 12310 23624
rect 12898 26424 12954 26480
rect 12709 25594 12765 25596
rect 12789 25594 12845 25596
rect 12869 25594 12925 25596
rect 12949 25594 13005 25596
rect 12709 25542 12755 25594
rect 12755 25542 12765 25594
rect 12789 25542 12819 25594
rect 12819 25542 12831 25594
rect 12831 25542 12845 25594
rect 12869 25542 12883 25594
rect 12883 25542 12895 25594
rect 12895 25542 12925 25594
rect 12949 25542 12959 25594
rect 12959 25542 13005 25594
rect 12709 25540 12765 25542
rect 12789 25540 12845 25542
rect 12869 25540 12925 25542
rect 12949 25540 13005 25542
rect 12806 24928 12862 24984
rect 12709 24506 12765 24508
rect 12789 24506 12845 24508
rect 12869 24506 12925 24508
rect 12949 24506 13005 24508
rect 12709 24454 12755 24506
rect 12755 24454 12765 24506
rect 12789 24454 12819 24506
rect 12819 24454 12831 24506
rect 12831 24454 12845 24506
rect 12869 24454 12883 24506
rect 12883 24454 12895 24506
rect 12895 24454 12925 24506
rect 12949 24454 12959 24506
rect 12959 24454 13005 24506
rect 12709 24452 12765 24454
rect 12789 24452 12845 24454
rect 12869 24452 12925 24454
rect 12949 24452 13005 24454
rect 12709 23418 12765 23420
rect 12789 23418 12845 23420
rect 12869 23418 12925 23420
rect 12949 23418 13005 23420
rect 12709 23366 12755 23418
rect 12755 23366 12765 23418
rect 12789 23366 12819 23418
rect 12819 23366 12831 23418
rect 12831 23366 12845 23418
rect 12869 23366 12883 23418
rect 12883 23366 12895 23418
rect 12895 23366 12925 23418
rect 12949 23366 12959 23418
rect 12959 23366 13005 23418
rect 12709 23364 12765 23366
rect 12789 23364 12845 23366
rect 12869 23364 12925 23366
rect 12949 23364 13005 23366
rect 14388 34842 14444 34844
rect 14468 34842 14524 34844
rect 14548 34842 14604 34844
rect 14628 34842 14684 34844
rect 14388 34790 14434 34842
rect 14434 34790 14444 34842
rect 14468 34790 14498 34842
rect 14498 34790 14510 34842
rect 14510 34790 14524 34842
rect 14548 34790 14562 34842
rect 14562 34790 14574 34842
rect 14574 34790 14604 34842
rect 14628 34790 14638 34842
rect 14638 34790 14684 34842
rect 14388 34788 14444 34790
rect 14468 34788 14524 34790
rect 14548 34788 14604 34790
rect 14628 34788 14684 34790
rect 14388 33754 14444 33756
rect 14468 33754 14524 33756
rect 14548 33754 14604 33756
rect 14628 33754 14684 33756
rect 14388 33702 14434 33754
rect 14434 33702 14444 33754
rect 14468 33702 14498 33754
rect 14498 33702 14510 33754
rect 14510 33702 14524 33754
rect 14548 33702 14562 33754
rect 14562 33702 14574 33754
rect 14574 33702 14604 33754
rect 14628 33702 14638 33754
rect 14638 33702 14684 33754
rect 14388 33700 14444 33702
rect 14468 33700 14524 33702
rect 14548 33700 14604 33702
rect 14628 33700 14684 33702
rect 14094 33224 14150 33280
rect 13910 32952 13966 33008
rect 13450 28464 13506 28520
rect 14186 32000 14242 32056
rect 13450 27648 13506 27704
rect 13726 25880 13782 25936
rect 13910 27512 13966 27568
rect 14388 32666 14444 32668
rect 14468 32666 14524 32668
rect 14548 32666 14604 32668
rect 14628 32666 14684 32668
rect 14388 32614 14434 32666
rect 14434 32614 14444 32666
rect 14468 32614 14498 32666
rect 14498 32614 14510 32666
rect 14510 32614 14524 32666
rect 14548 32614 14562 32666
rect 14562 32614 14574 32666
rect 14574 32614 14604 32666
rect 14628 32614 14638 32666
rect 14638 32614 14684 32666
rect 14388 32612 14444 32614
rect 14468 32612 14524 32614
rect 14548 32612 14604 32614
rect 14628 32612 14684 32614
rect 14094 30232 14150 30288
rect 14388 31578 14444 31580
rect 14468 31578 14524 31580
rect 14548 31578 14604 31580
rect 14628 31578 14684 31580
rect 14388 31526 14434 31578
rect 14434 31526 14444 31578
rect 14468 31526 14498 31578
rect 14498 31526 14510 31578
rect 14510 31526 14524 31578
rect 14548 31526 14562 31578
rect 14562 31526 14574 31578
rect 14574 31526 14604 31578
rect 14628 31526 14638 31578
rect 14638 31526 14684 31578
rect 14388 31524 14444 31526
rect 14468 31524 14524 31526
rect 14548 31524 14604 31526
rect 14628 31524 14684 31526
rect 14388 30490 14444 30492
rect 14468 30490 14524 30492
rect 14548 30490 14604 30492
rect 14628 30490 14684 30492
rect 14388 30438 14434 30490
rect 14434 30438 14444 30490
rect 14468 30438 14498 30490
rect 14498 30438 14510 30490
rect 14510 30438 14524 30490
rect 14548 30438 14562 30490
rect 14562 30438 14574 30490
rect 14574 30438 14604 30490
rect 14628 30438 14638 30490
rect 14638 30438 14684 30490
rect 14388 30436 14444 30438
rect 14468 30436 14524 30438
rect 14548 30436 14604 30438
rect 14628 30436 14684 30438
rect 14388 29402 14444 29404
rect 14468 29402 14524 29404
rect 14548 29402 14604 29404
rect 14628 29402 14684 29404
rect 14388 29350 14434 29402
rect 14434 29350 14444 29402
rect 14468 29350 14498 29402
rect 14498 29350 14510 29402
rect 14510 29350 14524 29402
rect 14548 29350 14562 29402
rect 14562 29350 14574 29402
rect 14574 29350 14604 29402
rect 14628 29350 14638 29402
rect 14638 29350 14684 29402
rect 14388 29348 14444 29350
rect 14468 29348 14524 29350
rect 14548 29348 14604 29350
rect 14628 29348 14684 29350
rect 14388 28314 14444 28316
rect 14468 28314 14524 28316
rect 14548 28314 14604 28316
rect 14628 28314 14684 28316
rect 14388 28262 14434 28314
rect 14434 28262 14444 28314
rect 14468 28262 14498 28314
rect 14498 28262 14510 28314
rect 14510 28262 14524 28314
rect 14548 28262 14562 28314
rect 14562 28262 14574 28314
rect 14574 28262 14604 28314
rect 14628 28262 14638 28314
rect 14638 28262 14684 28314
rect 14388 28260 14444 28262
rect 14468 28260 14524 28262
rect 14548 28260 14604 28262
rect 14628 28260 14684 28262
rect 14278 28056 14334 28112
rect 14388 27226 14444 27228
rect 14468 27226 14524 27228
rect 14548 27226 14604 27228
rect 14628 27226 14684 27228
rect 14388 27174 14434 27226
rect 14434 27174 14444 27226
rect 14468 27174 14498 27226
rect 14498 27174 14510 27226
rect 14510 27174 14524 27226
rect 14548 27174 14562 27226
rect 14562 27174 14574 27226
rect 14574 27174 14604 27226
rect 14628 27174 14638 27226
rect 14638 27174 14684 27226
rect 14388 27172 14444 27174
rect 14468 27172 14524 27174
rect 14548 27172 14604 27174
rect 14628 27172 14684 27174
rect 13818 25608 13874 25664
rect 13450 24520 13506 24576
rect 13174 23160 13230 23216
rect 12709 22330 12765 22332
rect 12789 22330 12845 22332
rect 12869 22330 12925 22332
rect 12949 22330 13005 22332
rect 12709 22278 12755 22330
rect 12755 22278 12765 22330
rect 12789 22278 12819 22330
rect 12819 22278 12831 22330
rect 12831 22278 12845 22330
rect 12869 22278 12883 22330
rect 12883 22278 12895 22330
rect 12895 22278 12925 22330
rect 12949 22278 12959 22330
rect 12959 22278 13005 22330
rect 12709 22276 12765 22278
rect 12789 22276 12845 22278
rect 12869 22276 12925 22278
rect 12949 22276 13005 22278
rect 12254 21256 12310 21312
rect 12162 20576 12218 20632
rect 10874 17620 10876 17640
rect 10876 17620 10928 17640
rect 10928 17620 10930 17640
rect 10874 17584 10930 17620
rect 10782 17312 10838 17368
rect 11030 17434 11086 17436
rect 11110 17434 11166 17436
rect 11190 17434 11246 17436
rect 11270 17434 11326 17436
rect 11030 17382 11076 17434
rect 11076 17382 11086 17434
rect 11110 17382 11140 17434
rect 11140 17382 11152 17434
rect 11152 17382 11166 17434
rect 11190 17382 11204 17434
rect 11204 17382 11216 17434
rect 11216 17382 11246 17434
rect 11270 17382 11280 17434
rect 11280 17382 11326 17434
rect 11030 17380 11086 17382
rect 11110 17380 11166 17382
rect 11190 17380 11246 17382
rect 11270 17380 11326 17382
rect 11150 17040 11206 17096
rect 11150 16632 11206 16688
rect 11030 16346 11086 16348
rect 11110 16346 11166 16348
rect 11190 16346 11246 16348
rect 11270 16346 11326 16348
rect 11030 16294 11076 16346
rect 11076 16294 11086 16346
rect 11110 16294 11140 16346
rect 11140 16294 11152 16346
rect 11152 16294 11166 16346
rect 11190 16294 11204 16346
rect 11204 16294 11216 16346
rect 11216 16294 11246 16346
rect 11270 16294 11280 16346
rect 11280 16294 11326 16346
rect 11030 16292 11086 16294
rect 11110 16292 11166 16294
rect 11190 16292 11246 16294
rect 11270 16292 11326 16294
rect 11058 15564 11114 15600
rect 11058 15544 11060 15564
rect 11060 15544 11112 15564
rect 11112 15544 11114 15564
rect 11030 15258 11086 15260
rect 11110 15258 11166 15260
rect 11190 15258 11246 15260
rect 11270 15258 11326 15260
rect 11030 15206 11076 15258
rect 11076 15206 11086 15258
rect 11110 15206 11140 15258
rect 11140 15206 11152 15258
rect 11152 15206 11166 15258
rect 11190 15206 11204 15258
rect 11204 15206 11216 15258
rect 11216 15206 11246 15258
rect 11270 15206 11280 15258
rect 11280 15206 11326 15258
rect 11030 15204 11086 15206
rect 11110 15204 11166 15206
rect 11190 15204 11246 15206
rect 11270 15204 11326 15206
rect 10782 14864 10838 14920
rect 11058 14592 11114 14648
rect 11150 14456 11206 14512
rect 12162 19760 12218 19816
rect 12709 21242 12765 21244
rect 12789 21242 12845 21244
rect 12869 21242 12925 21244
rect 12949 21242 13005 21244
rect 12709 21190 12755 21242
rect 12755 21190 12765 21242
rect 12789 21190 12819 21242
rect 12819 21190 12831 21242
rect 12831 21190 12845 21242
rect 12869 21190 12883 21242
rect 12883 21190 12895 21242
rect 12895 21190 12925 21242
rect 12949 21190 12959 21242
rect 12959 21190 13005 21242
rect 12709 21188 12765 21190
rect 12789 21188 12845 21190
rect 12869 21188 12925 21190
rect 12949 21188 13005 21190
rect 12070 18808 12126 18864
rect 11702 17620 11704 17640
rect 11704 17620 11756 17640
rect 11756 17620 11758 17640
rect 11702 17584 11758 17620
rect 11702 17176 11758 17232
rect 11610 16396 11612 16416
rect 11612 16396 11664 16416
rect 11664 16396 11666 16416
rect 11610 16360 11666 16396
rect 11030 14170 11086 14172
rect 11110 14170 11166 14172
rect 11190 14170 11246 14172
rect 11270 14170 11326 14172
rect 11030 14118 11076 14170
rect 11076 14118 11086 14170
rect 11110 14118 11140 14170
rect 11140 14118 11152 14170
rect 11152 14118 11166 14170
rect 11190 14118 11204 14170
rect 11204 14118 11216 14170
rect 11216 14118 11246 14170
rect 11270 14118 11280 14170
rect 11280 14118 11326 14170
rect 11030 14116 11086 14118
rect 11110 14116 11166 14118
rect 11190 14116 11246 14118
rect 11270 14116 11326 14118
rect 11334 13912 11390 13968
rect 11886 17176 11942 17232
rect 12070 17584 12126 17640
rect 12714 20576 12770 20632
rect 12709 20154 12765 20156
rect 12789 20154 12845 20156
rect 12869 20154 12925 20156
rect 12949 20154 13005 20156
rect 12709 20102 12755 20154
rect 12755 20102 12765 20154
rect 12789 20102 12819 20154
rect 12819 20102 12831 20154
rect 12831 20102 12845 20154
rect 12869 20102 12883 20154
rect 12883 20102 12895 20154
rect 12895 20102 12925 20154
rect 12949 20102 12959 20154
rect 12959 20102 13005 20154
rect 12709 20100 12765 20102
rect 12789 20100 12845 20102
rect 12869 20100 12925 20102
rect 12949 20100 13005 20102
rect 12622 19916 12678 19952
rect 12622 19896 12624 19916
rect 12624 19896 12676 19916
rect 12676 19896 12678 19916
rect 13358 21428 13360 21448
rect 13360 21428 13412 21448
rect 13412 21428 13414 21448
rect 13358 21392 13414 21428
rect 13266 20984 13322 21040
rect 12709 19066 12765 19068
rect 12789 19066 12845 19068
rect 12869 19066 12925 19068
rect 12949 19066 13005 19068
rect 12709 19014 12755 19066
rect 12755 19014 12765 19066
rect 12789 19014 12819 19066
rect 12819 19014 12831 19066
rect 12831 19014 12845 19066
rect 12869 19014 12883 19066
rect 12883 19014 12895 19066
rect 12895 19014 12925 19066
rect 12949 19014 12959 19066
rect 12959 19014 13005 19066
rect 12709 19012 12765 19014
rect 12789 19012 12845 19014
rect 12869 19012 12925 19014
rect 12949 19012 13005 19014
rect 12346 18284 12402 18320
rect 12346 18264 12348 18284
rect 12348 18264 12400 18284
rect 12400 18264 12402 18284
rect 12346 18128 12402 18184
rect 11702 15408 11758 15464
rect 11702 14184 11758 14240
rect 12070 15564 12126 15600
rect 12070 15544 12072 15564
rect 12072 15544 12124 15564
rect 12124 15544 12126 15564
rect 12162 15136 12218 15192
rect 11886 14592 11942 14648
rect 11978 14456 12034 14512
rect 11242 13268 11244 13288
rect 11244 13268 11296 13288
rect 11296 13268 11298 13288
rect 11242 13232 11298 13268
rect 11030 13082 11086 13084
rect 11110 13082 11166 13084
rect 11190 13082 11246 13084
rect 11270 13082 11326 13084
rect 11030 13030 11076 13082
rect 11076 13030 11086 13082
rect 11110 13030 11140 13082
rect 11140 13030 11152 13082
rect 11152 13030 11166 13082
rect 11190 13030 11204 13082
rect 11204 13030 11216 13082
rect 11216 13030 11246 13082
rect 11270 13030 11280 13082
rect 11280 13030 11326 13082
rect 11030 13028 11086 13030
rect 11110 13028 11166 13030
rect 11190 13028 11246 13030
rect 11270 13028 11326 13030
rect 11334 12588 11336 12608
rect 11336 12588 11388 12608
rect 11388 12588 11390 12608
rect 11334 12552 11390 12588
rect 11030 11994 11086 11996
rect 11110 11994 11166 11996
rect 11190 11994 11246 11996
rect 11270 11994 11326 11996
rect 11030 11942 11076 11994
rect 11076 11942 11086 11994
rect 11110 11942 11140 11994
rect 11140 11942 11152 11994
rect 11152 11942 11166 11994
rect 11190 11942 11204 11994
rect 11204 11942 11216 11994
rect 11216 11942 11246 11994
rect 11270 11942 11280 11994
rect 11280 11942 11326 11994
rect 11030 11940 11086 11942
rect 11110 11940 11166 11942
rect 11190 11940 11246 11942
rect 11270 11940 11326 11942
rect 11610 12008 11666 12064
rect 12162 12280 12218 12336
rect 12070 11772 12072 11792
rect 12072 11772 12124 11792
rect 12124 11772 12126 11792
rect 12070 11736 12126 11772
rect 12070 11600 12126 11656
rect 11886 11464 11942 11520
rect 11794 11192 11850 11248
rect 10138 10004 10140 10024
rect 10140 10004 10192 10024
rect 10192 10004 10194 10024
rect 10138 9968 10194 10004
rect 10414 9968 10470 10024
rect 10138 9288 10194 9344
rect 9770 6704 9826 6760
rect 10506 9288 10562 9344
rect 11030 10906 11086 10908
rect 11110 10906 11166 10908
rect 11190 10906 11246 10908
rect 11270 10906 11326 10908
rect 11030 10854 11076 10906
rect 11076 10854 11086 10906
rect 11110 10854 11140 10906
rect 11140 10854 11152 10906
rect 11152 10854 11166 10906
rect 11190 10854 11204 10906
rect 11204 10854 11216 10906
rect 11216 10854 11246 10906
rect 11270 10854 11280 10906
rect 11280 10854 11326 10906
rect 11030 10852 11086 10854
rect 11110 10852 11166 10854
rect 11190 10852 11246 10854
rect 11270 10852 11326 10854
rect 11030 9818 11086 9820
rect 11110 9818 11166 9820
rect 11190 9818 11246 9820
rect 11270 9818 11326 9820
rect 11030 9766 11076 9818
rect 11076 9766 11086 9818
rect 11110 9766 11140 9818
rect 11140 9766 11152 9818
rect 11152 9766 11166 9818
rect 11190 9766 11204 9818
rect 11204 9766 11216 9818
rect 11216 9766 11246 9818
rect 11270 9766 11280 9818
rect 11280 9766 11326 9818
rect 11030 9764 11086 9766
rect 11110 9764 11166 9766
rect 11190 9764 11246 9766
rect 11270 9764 11326 9766
rect 11242 9016 11298 9072
rect 11426 9288 11482 9344
rect 11610 10124 11666 10160
rect 11610 10104 11612 10124
rect 11612 10104 11664 10124
rect 11664 10104 11666 10124
rect 11610 9424 11666 9480
rect 11030 8730 11086 8732
rect 11110 8730 11166 8732
rect 11190 8730 11246 8732
rect 11270 8730 11326 8732
rect 11030 8678 11076 8730
rect 11076 8678 11086 8730
rect 11110 8678 11140 8730
rect 11140 8678 11152 8730
rect 11152 8678 11166 8730
rect 11190 8678 11204 8730
rect 11204 8678 11216 8730
rect 11216 8678 11246 8730
rect 11270 8678 11280 8730
rect 11280 8678 11326 8730
rect 11030 8676 11086 8678
rect 11110 8676 11166 8678
rect 11190 8676 11246 8678
rect 11270 8676 11326 8678
rect 11334 8472 11390 8528
rect 10782 7692 10784 7712
rect 10784 7692 10836 7712
rect 10836 7692 10838 7712
rect 10782 7656 10838 7692
rect 10782 7384 10838 7440
rect 10322 6316 10378 6352
rect 10322 6296 10324 6316
rect 10324 6296 10376 6316
rect 10376 6296 10378 6316
rect 9351 6010 9407 6012
rect 9431 6010 9487 6012
rect 9511 6010 9567 6012
rect 9591 6010 9647 6012
rect 9351 5958 9397 6010
rect 9397 5958 9407 6010
rect 9431 5958 9461 6010
rect 9461 5958 9473 6010
rect 9473 5958 9487 6010
rect 9511 5958 9525 6010
rect 9525 5958 9537 6010
rect 9537 5958 9567 6010
rect 9591 5958 9601 6010
rect 9601 5958 9647 6010
rect 9351 5956 9407 5958
rect 9431 5956 9487 5958
rect 9511 5956 9567 5958
rect 9591 5956 9647 5958
rect 9351 4922 9407 4924
rect 9431 4922 9487 4924
rect 9511 4922 9567 4924
rect 9591 4922 9647 4924
rect 9351 4870 9397 4922
rect 9397 4870 9407 4922
rect 9431 4870 9461 4922
rect 9461 4870 9473 4922
rect 9473 4870 9487 4922
rect 9511 4870 9525 4922
rect 9525 4870 9537 4922
rect 9537 4870 9567 4922
rect 9591 4870 9601 4922
rect 9601 4870 9647 4922
rect 9351 4868 9407 4870
rect 9431 4868 9487 4870
rect 9511 4868 9567 4870
rect 9591 4868 9647 4870
rect 11242 7928 11298 7984
rect 11150 7792 11206 7848
rect 11030 7642 11086 7644
rect 11110 7642 11166 7644
rect 11190 7642 11246 7644
rect 11270 7642 11326 7644
rect 11030 7590 11076 7642
rect 11076 7590 11086 7642
rect 11110 7590 11140 7642
rect 11140 7590 11152 7642
rect 11152 7590 11166 7642
rect 11190 7590 11204 7642
rect 11204 7590 11216 7642
rect 11216 7590 11246 7642
rect 11270 7590 11280 7642
rect 11280 7590 11326 7642
rect 11030 7588 11086 7590
rect 11110 7588 11166 7590
rect 11190 7588 11246 7590
rect 11270 7588 11326 7590
rect 11030 6554 11086 6556
rect 11110 6554 11166 6556
rect 11190 6554 11246 6556
rect 11270 6554 11326 6556
rect 11030 6502 11076 6554
rect 11076 6502 11086 6554
rect 11110 6502 11140 6554
rect 11140 6502 11152 6554
rect 11152 6502 11166 6554
rect 11190 6502 11204 6554
rect 11204 6502 11216 6554
rect 11216 6502 11246 6554
rect 11270 6502 11280 6554
rect 11280 6502 11326 6554
rect 11030 6500 11086 6502
rect 11110 6500 11166 6502
rect 11190 6500 11246 6502
rect 11270 6500 11326 6502
rect 11978 10920 12034 10976
rect 11886 10668 11942 10704
rect 11886 10648 11888 10668
rect 11888 10648 11940 10668
rect 11940 10648 11942 10668
rect 12709 17978 12765 17980
rect 12789 17978 12845 17980
rect 12869 17978 12925 17980
rect 12949 17978 13005 17980
rect 12709 17926 12755 17978
rect 12755 17926 12765 17978
rect 12789 17926 12819 17978
rect 12819 17926 12831 17978
rect 12831 17926 12845 17978
rect 12869 17926 12883 17978
rect 12883 17926 12895 17978
rect 12895 17926 12925 17978
rect 12949 17926 12959 17978
rect 12959 17926 13005 17978
rect 12709 17924 12765 17926
rect 12789 17924 12845 17926
rect 12869 17924 12925 17926
rect 12949 17924 13005 17926
rect 12530 15020 12586 15056
rect 12530 15000 12532 15020
rect 12532 15000 12584 15020
rect 12584 15000 12586 15020
rect 12438 14592 12494 14648
rect 12438 13948 12440 13968
rect 12440 13948 12492 13968
rect 12492 13948 12494 13968
rect 12438 13912 12494 13948
rect 12346 12824 12402 12880
rect 12990 17448 13046 17504
rect 12709 16890 12765 16892
rect 12789 16890 12845 16892
rect 12869 16890 12925 16892
rect 12949 16890 13005 16892
rect 12709 16838 12755 16890
rect 12755 16838 12765 16890
rect 12789 16838 12819 16890
rect 12819 16838 12831 16890
rect 12831 16838 12845 16890
rect 12869 16838 12883 16890
rect 12883 16838 12895 16890
rect 12895 16838 12925 16890
rect 12949 16838 12959 16890
rect 12959 16838 13005 16890
rect 12709 16836 12765 16838
rect 12789 16836 12845 16838
rect 12869 16836 12925 16838
rect 12949 16836 13005 16838
rect 13082 15816 13138 15872
rect 12709 15802 12765 15804
rect 12789 15802 12845 15804
rect 12869 15802 12925 15804
rect 12949 15802 13005 15804
rect 12709 15750 12755 15802
rect 12755 15750 12765 15802
rect 12789 15750 12819 15802
rect 12819 15750 12831 15802
rect 12831 15750 12845 15802
rect 12869 15750 12883 15802
rect 12883 15750 12895 15802
rect 12895 15750 12925 15802
rect 12949 15750 12959 15802
rect 12959 15750 13005 15802
rect 12709 15748 12765 15750
rect 12789 15748 12845 15750
rect 12869 15748 12925 15750
rect 12949 15748 13005 15750
rect 12709 14714 12765 14716
rect 12789 14714 12845 14716
rect 12869 14714 12925 14716
rect 12949 14714 13005 14716
rect 12709 14662 12755 14714
rect 12755 14662 12765 14714
rect 12789 14662 12819 14714
rect 12819 14662 12831 14714
rect 12831 14662 12845 14714
rect 12869 14662 12883 14714
rect 12883 14662 12895 14714
rect 12895 14662 12925 14714
rect 12949 14662 12959 14714
rect 12959 14662 13005 14714
rect 12709 14660 12765 14662
rect 12789 14660 12845 14662
rect 12869 14660 12925 14662
rect 12949 14660 13005 14662
rect 12990 14456 13046 14512
rect 12709 13626 12765 13628
rect 12789 13626 12845 13628
rect 12869 13626 12925 13628
rect 12949 13626 13005 13628
rect 12709 13574 12755 13626
rect 12755 13574 12765 13626
rect 12789 13574 12819 13626
rect 12819 13574 12831 13626
rect 12831 13574 12845 13626
rect 12869 13574 12883 13626
rect 12883 13574 12895 13626
rect 12895 13574 12925 13626
rect 12949 13574 12959 13626
rect 12959 13574 13005 13626
rect 12709 13572 12765 13574
rect 12789 13572 12845 13574
rect 12869 13572 12925 13574
rect 12949 13572 13005 13574
rect 13818 23432 13874 23488
rect 13726 23160 13782 23216
rect 13726 22208 13782 22264
rect 13818 22072 13874 22128
rect 14002 26424 14058 26480
rect 14388 26138 14444 26140
rect 14468 26138 14524 26140
rect 14548 26138 14604 26140
rect 14628 26138 14684 26140
rect 14388 26086 14434 26138
rect 14434 26086 14444 26138
rect 14468 26086 14498 26138
rect 14498 26086 14510 26138
rect 14510 26086 14524 26138
rect 14548 26086 14562 26138
rect 14562 26086 14574 26138
rect 14574 26086 14604 26138
rect 14628 26086 14638 26138
rect 14638 26086 14684 26138
rect 14388 26084 14444 26086
rect 14468 26084 14524 26086
rect 14548 26084 14604 26086
rect 14628 26084 14684 26086
rect 14186 25200 14242 25256
rect 14388 25050 14444 25052
rect 14468 25050 14524 25052
rect 14548 25050 14604 25052
rect 14628 25050 14684 25052
rect 14388 24998 14434 25050
rect 14434 24998 14444 25050
rect 14468 24998 14498 25050
rect 14498 24998 14510 25050
rect 14510 24998 14524 25050
rect 14548 24998 14562 25050
rect 14562 24998 14574 25050
rect 14574 24998 14604 25050
rect 14628 24998 14638 25050
rect 14638 24998 14684 25050
rect 14388 24996 14444 24998
rect 14468 24996 14524 24998
rect 14548 24996 14604 24998
rect 14628 24996 14684 24998
rect 14002 24792 14058 24848
rect 14002 24248 14058 24304
rect 14388 23962 14444 23964
rect 14468 23962 14524 23964
rect 14548 23962 14604 23964
rect 14628 23962 14684 23964
rect 14388 23910 14434 23962
rect 14434 23910 14444 23962
rect 14468 23910 14498 23962
rect 14498 23910 14510 23962
rect 14510 23910 14524 23962
rect 14548 23910 14562 23962
rect 14562 23910 14574 23962
rect 14574 23910 14604 23962
rect 14628 23910 14638 23962
rect 14638 23910 14684 23962
rect 14388 23908 14444 23910
rect 14468 23908 14524 23910
rect 14548 23908 14604 23910
rect 14628 23908 14684 23910
rect 14278 23704 14334 23760
rect 13910 21936 13966 21992
rect 13726 21528 13782 21584
rect 13818 20712 13874 20768
rect 13450 18400 13506 18456
rect 13450 18284 13506 18320
rect 13450 18264 13452 18284
rect 13452 18264 13504 18284
rect 13504 18264 13506 18284
rect 13542 17312 13598 17368
rect 14002 21256 14058 21312
rect 14094 20984 14150 21040
rect 14388 22874 14444 22876
rect 14468 22874 14524 22876
rect 14548 22874 14604 22876
rect 14628 22874 14684 22876
rect 14388 22822 14434 22874
rect 14434 22822 14444 22874
rect 14468 22822 14498 22874
rect 14498 22822 14510 22874
rect 14510 22822 14524 22874
rect 14548 22822 14562 22874
rect 14562 22822 14574 22874
rect 14574 22822 14604 22874
rect 14628 22822 14638 22874
rect 14638 22822 14684 22874
rect 14388 22820 14444 22822
rect 14468 22820 14524 22822
rect 14548 22820 14604 22822
rect 14628 22820 14684 22822
rect 14278 22616 14334 22672
rect 14388 21786 14444 21788
rect 14468 21786 14524 21788
rect 14548 21786 14604 21788
rect 14628 21786 14684 21788
rect 14388 21734 14434 21786
rect 14434 21734 14444 21786
rect 14468 21734 14498 21786
rect 14498 21734 14510 21786
rect 14510 21734 14524 21786
rect 14548 21734 14562 21786
rect 14562 21734 14574 21786
rect 14574 21734 14604 21786
rect 14628 21734 14638 21786
rect 14638 21734 14684 21786
rect 14388 21732 14444 21734
rect 14468 21732 14524 21734
rect 14548 21732 14604 21734
rect 14628 21732 14684 21734
rect 14388 20698 14444 20700
rect 14468 20698 14524 20700
rect 14548 20698 14604 20700
rect 14628 20698 14684 20700
rect 14388 20646 14434 20698
rect 14434 20646 14444 20698
rect 14468 20646 14498 20698
rect 14498 20646 14510 20698
rect 14510 20646 14524 20698
rect 14548 20646 14562 20698
rect 14562 20646 14574 20698
rect 14574 20646 14604 20698
rect 14628 20646 14638 20698
rect 14638 20646 14684 20698
rect 14388 20644 14444 20646
rect 14468 20644 14524 20646
rect 14548 20644 14604 20646
rect 14628 20644 14684 20646
rect 14094 20168 14150 20224
rect 14002 19080 14058 19136
rect 13634 16496 13690 16552
rect 13082 13232 13138 13288
rect 12438 12416 12494 12472
rect 12714 12688 12770 12744
rect 12530 11464 12586 11520
rect 11702 7384 11758 7440
rect 12070 7248 12126 7304
rect 11702 6704 11758 6760
rect 11030 5466 11086 5468
rect 11110 5466 11166 5468
rect 11190 5466 11246 5468
rect 11270 5466 11326 5468
rect 11030 5414 11076 5466
rect 11076 5414 11086 5466
rect 11110 5414 11140 5466
rect 11140 5414 11152 5466
rect 11152 5414 11166 5466
rect 11190 5414 11204 5466
rect 11204 5414 11216 5466
rect 11216 5414 11246 5466
rect 11270 5414 11280 5466
rect 11280 5414 11326 5466
rect 11030 5412 11086 5414
rect 11110 5412 11166 5414
rect 11190 5412 11246 5414
rect 11270 5412 11326 5414
rect 11030 4378 11086 4380
rect 11110 4378 11166 4380
rect 11190 4378 11246 4380
rect 11270 4378 11326 4380
rect 11030 4326 11076 4378
rect 11076 4326 11086 4378
rect 11110 4326 11140 4378
rect 11140 4326 11152 4378
rect 11152 4326 11166 4378
rect 11190 4326 11204 4378
rect 11204 4326 11216 4378
rect 11216 4326 11246 4378
rect 11270 4326 11280 4378
rect 11280 4326 11326 4378
rect 11030 4324 11086 4326
rect 11110 4324 11166 4326
rect 11190 4324 11246 4326
rect 11270 4324 11326 4326
rect 12346 10648 12402 10704
rect 12346 10512 12402 10568
rect 12438 10104 12494 10160
rect 12438 9560 12494 9616
rect 12254 6296 12310 6352
rect 11978 5072 12034 5128
rect 12346 5752 12402 5808
rect 12709 12538 12765 12540
rect 12789 12538 12845 12540
rect 12869 12538 12925 12540
rect 12949 12538 13005 12540
rect 12709 12486 12755 12538
rect 12755 12486 12765 12538
rect 12789 12486 12819 12538
rect 12819 12486 12831 12538
rect 12831 12486 12845 12538
rect 12869 12486 12883 12538
rect 12883 12486 12895 12538
rect 12895 12486 12925 12538
rect 12949 12486 12959 12538
rect 12959 12486 13005 12538
rect 12709 12484 12765 12486
rect 12789 12484 12845 12486
rect 12869 12484 12925 12486
rect 12949 12484 13005 12486
rect 12709 11450 12765 11452
rect 12789 11450 12845 11452
rect 12869 11450 12925 11452
rect 12949 11450 13005 11452
rect 12709 11398 12755 11450
rect 12755 11398 12765 11450
rect 12789 11398 12819 11450
rect 12819 11398 12831 11450
rect 12831 11398 12845 11450
rect 12869 11398 12883 11450
rect 12883 11398 12895 11450
rect 12895 11398 12925 11450
rect 12949 11398 12959 11450
rect 12959 11398 13005 11450
rect 12709 11396 12765 11398
rect 12789 11396 12845 11398
rect 12869 11396 12925 11398
rect 12949 11396 13005 11398
rect 12714 11092 12716 11112
rect 12716 11092 12768 11112
rect 12768 11092 12770 11112
rect 12714 11056 12770 11092
rect 12709 10362 12765 10364
rect 12789 10362 12845 10364
rect 12869 10362 12925 10364
rect 12949 10362 13005 10364
rect 12709 10310 12755 10362
rect 12755 10310 12765 10362
rect 12789 10310 12819 10362
rect 12819 10310 12831 10362
rect 12831 10310 12845 10362
rect 12869 10310 12883 10362
rect 12883 10310 12895 10362
rect 12895 10310 12925 10362
rect 12949 10310 12959 10362
rect 12959 10310 13005 10362
rect 12709 10308 12765 10310
rect 12789 10308 12845 10310
rect 12869 10308 12925 10310
rect 12949 10308 13005 10310
rect 13082 9560 13138 9616
rect 12709 9274 12765 9276
rect 12789 9274 12845 9276
rect 12869 9274 12925 9276
rect 12949 9274 13005 9276
rect 12709 9222 12755 9274
rect 12755 9222 12765 9274
rect 12789 9222 12819 9274
rect 12819 9222 12831 9274
rect 12831 9222 12845 9274
rect 12869 9222 12883 9274
rect 12883 9222 12895 9274
rect 12895 9222 12925 9274
rect 12949 9222 12959 9274
rect 12959 9222 13005 9274
rect 12709 9220 12765 9222
rect 12789 9220 12845 9222
rect 12869 9220 12925 9222
rect 12949 9220 13005 9222
rect 12709 8186 12765 8188
rect 12789 8186 12845 8188
rect 12869 8186 12925 8188
rect 12949 8186 13005 8188
rect 12709 8134 12755 8186
rect 12755 8134 12765 8186
rect 12789 8134 12819 8186
rect 12819 8134 12831 8186
rect 12831 8134 12845 8186
rect 12869 8134 12883 8186
rect 12883 8134 12895 8186
rect 12895 8134 12925 8186
rect 12949 8134 12959 8186
rect 12959 8134 13005 8186
rect 12709 8132 12765 8134
rect 12789 8132 12845 8134
rect 12869 8132 12925 8134
rect 12949 8132 13005 8134
rect 13450 12144 13506 12200
rect 13266 9696 13322 9752
rect 13266 9560 13322 9616
rect 12709 7098 12765 7100
rect 12789 7098 12845 7100
rect 12869 7098 12925 7100
rect 12949 7098 13005 7100
rect 12709 7046 12755 7098
rect 12755 7046 12765 7098
rect 12789 7046 12819 7098
rect 12819 7046 12831 7098
rect 12831 7046 12845 7098
rect 12869 7046 12883 7098
rect 12883 7046 12895 7098
rect 12895 7046 12925 7098
rect 12949 7046 12959 7098
rect 12959 7046 13005 7098
rect 12709 7044 12765 7046
rect 12789 7044 12845 7046
rect 12869 7044 12925 7046
rect 12949 7044 13005 7046
rect 12530 6160 12586 6216
rect 12709 6010 12765 6012
rect 12789 6010 12845 6012
rect 12869 6010 12925 6012
rect 12949 6010 13005 6012
rect 12709 5958 12755 6010
rect 12755 5958 12765 6010
rect 12789 5958 12819 6010
rect 12819 5958 12831 6010
rect 12831 5958 12845 6010
rect 12869 5958 12883 6010
rect 12883 5958 12895 6010
rect 12895 5958 12925 6010
rect 12949 5958 12959 6010
rect 12959 5958 13005 6010
rect 12709 5956 12765 5958
rect 12789 5956 12845 5958
rect 12869 5956 12925 5958
rect 12949 5956 13005 5958
rect 12438 5636 12494 5672
rect 12438 5616 12440 5636
rect 12440 5616 12492 5636
rect 12492 5616 12494 5636
rect 12709 4922 12765 4924
rect 12789 4922 12845 4924
rect 12869 4922 12925 4924
rect 12949 4922 13005 4924
rect 12709 4870 12755 4922
rect 12755 4870 12765 4922
rect 12789 4870 12819 4922
rect 12819 4870 12831 4922
rect 12831 4870 12845 4922
rect 12869 4870 12883 4922
rect 12883 4870 12895 4922
rect 12895 4870 12925 4922
rect 12949 4870 12959 4922
rect 12959 4870 13005 4922
rect 12709 4868 12765 4870
rect 12789 4868 12845 4870
rect 12869 4868 12925 4870
rect 12949 4868 13005 4870
rect 9351 3834 9407 3836
rect 9431 3834 9487 3836
rect 9511 3834 9567 3836
rect 9591 3834 9647 3836
rect 9351 3782 9397 3834
rect 9397 3782 9407 3834
rect 9431 3782 9461 3834
rect 9461 3782 9473 3834
rect 9473 3782 9487 3834
rect 9511 3782 9525 3834
rect 9525 3782 9537 3834
rect 9537 3782 9567 3834
rect 9591 3782 9601 3834
rect 9601 3782 9647 3834
rect 9351 3780 9407 3782
rect 9431 3780 9487 3782
rect 9511 3780 9567 3782
rect 9591 3780 9647 3782
rect 12709 3834 12765 3836
rect 12789 3834 12845 3836
rect 12869 3834 12925 3836
rect 12949 3834 13005 3836
rect 12709 3782 12755 3834
rect 12755 3782 12765 3834
rect 12789 3782 12819 3834
rect 12819 3782 12831 3834
rect 12831 3782 12845 3834
rect 12869 3782 12883 3834
rect 12883 3782 12895 3834
rect 12895 3782 12925 3834
rect 12949 3782 12959 3834
rect 12959 3782 13005 3834
rect 12709 3780 12765 3782
rect 12789 3780 12845 3782
rect 12869 3780 12925 3782
rect 12949 3780 13005 3782
rect 11030 3290 11086 3292
rect 11110 3290 11166 3292
rect 11190 3290 11246 3292
rect 11270 3290 11326 3292
rect 11030 3238 11076 3290
rect 11076 3238 11086 3290
rect 11110 3238 11140 3290
rect 11140 3238 11152 3290
rect 11152 3238 11166 3290
rect 11190 3238 11204 3290
rect 11204 3238 11216 3290
rect 11216 3238 11246 3290
rect 11270 3238 11280 3290
rect 11280 3238 11326 3290
rect 11030 3236 11086 3238
rect 11110 3236 11166 3238
rect 11190 3236 11246 3238
rect 11270 3236 11326 3238
rect 14002 16632 14058 16688
rect 13818 15544 13874 15600
rect 13726 15272 13782 15328
rect 13910 15000 13966 15056
rect 14094 15136 14150 15192
rect 14094 13912 14150 13968
rect 13726 12416 13782 12472
rect 13726 12008 13782 12064
rect 13634 9832 13690 9888
rect 13726 9560 13782 9616
rect 14002 13368 14058 13424
rect 14094 10376 14150 10432
rect 14002 10104 14058 10160
rect 14388 19610 14444 19612
rect 14468 19610 14524 19612
rect 14548 19610 14604 19612
rect 14628 19610 14684 19612
rect 14388 19558 14434 19610
rect 14434 19558 14444 19610
rect 14468 19558 14498 19610
rect 14498 19558 14510 19610
rect 14510 19558 14524 19610
rect 14548 19558 14562 19610
rect 14562 19558 14574 19610
rect 14574 19558 14604 19610
rect 14628 19558 14638 19610
rect 14638 19558 14684 19610
rect 14388 19556 14444 19558
rect 14468 19556 14524 19558
rect 14548 19556 14604 19558
rect 14628 19556 14684 19558
rect 14370 19216 14426 19272
rect 14388 18522 14444 18524
rect 14468 18522 14524 18524
rect 14548 18522 14604 18524
rect 14628 18522 14684 18524
rect 14388 18470 14434 18522
rect 14434 18470 14444 18522
rect 14468 18470 14498 18522
rect 14498 18470 14510 18522
rect 14510 18470 14524 18522
rect 14548 18470 14562 18522
rect 14562 18470 14574 18522
rect 14574 18470 14604 18522
rect 14628 18470 14638 18522
rect 14638 18470 14684 18522
rect 14388 18468 14444 18470
rect 14468 18468 14524 18470
rect 14548 18468 14604 18470
rect 14628 18468 14684 18470
rect 14388 17434 14444 17436
rect 14468 17434 14524 17436
rect 14548 17434 14604 17436
rect 14628 17434 14684 17436
rect 14388 17382 14434 17434
rect 14434 17382 14444 17434
rect 14468 17382 14498 17434
rect 14498 17382 14510 17434
rect 14510 17382 14524 17434
rect 14548 17382 14562 17434
rect 14562 17382 14574 17434
rect 14574 17382 14604 17434
rect 14628 17382 14638 17434
rect 14638 17382 14684 17434
rect 14388 17380 14444 17382
rect 14468 17380 14524 17382
rect 14548 17380 14604 17382
rect 14628 17380 14684 17382
rect 14388 16346 14444 16348
rect 14468 16346 14524 16348
rect 14548 16346 14604 16348
rect 14628 16346 14684 16348
rect 14388 16294 14434 16346
rect 14434 16294 14444 16346
rect 14468 16294 14498 16346
rect 14498 16294 14510 16346
rect 14510 16294 14524 16346
rect 14548 16294 14562 16346
rect 14562 16294 14574 16346
rect 14574 16294 14604 16346
rect 14628 16294 14638 16346
rect 14638 16294 14684 16346
rect 14388 16292 14444 16294
rect 14468 16292 14524 16294
rect 14548 16292 14604 16294
rect 14628 16292 14684 16294
rect 14646 16088 14702 16144
rect 14388 15258 14444 15260
rect 14468 15258 14524 15260
rect 14548 15258 14604 15260
rect 14628 15258 14684 15260
rect 14388 15206 14434 15258
rect 14434 15206 14444 15258
rect 14468 15206 14498 15258
rect 14498 15206 14510 15258
rect 14510 15206 14524 15258
rect 14548 15206 14562 15258
rect 14562 15206 14574 15258
rect 14574 15206 14604 15258
rect 14628 15206 14638 15258
rect 14638 15206 14684 15258
rect 14388 15204 14444 15206
rect 14468 15204 14524 15206
rect 14548 15204 14604 15206
rect 14628 15204 14684 15206
rect 14370 14764 14372 14784
rect 14372 14764 14424 14784
rect 14424 14764 14426 14784
rect 14370 14728 14426 14764
rect 14388 14170 14444 14172
rect 14468 14170 14524 14172
rect 14548 14170 14604 14172
rect 14628 14170 14684 14172
rect 14388 14118 14434 14170
rect 14434 14118 14444 14170
rect 14468 14118 14498 14170
rect 14498 14118 14510 14170
rect 14510 14118 14524 14170
rect 14548 14118 14562 14170
rect 14562 14118 14574 14170
rect 14574 14118 14604 14170
rect 14628 14118 14638 14170
rect 14638 14118 14684 14170
rect 14388 14116 14444 14118
rect 14468 14116 14524 14118
rect 14548 14116 14604 14118
rect 14628 14116 14684 14118
rect 14370 13640 14426 13696
rect 14388 13082 14444 13084
rect 14468 13082 14524 13084
rect 14548 13082 14604 13084
rect 14628 13082 14684 13084
rect 14388 13030 14434 13082
rect 14434 13030 14444 13082
rect 14468 13030 14498 13082
rect 14498 13030 14510 13082
rect 14510 13030 14524 13082
rect 14548 13030 14562 13082
rect 14562 13030 14574 13082
rect 14574 13030 14604 13082
rect 14628 13030 14638 13082
rect 14638 13030 14684 13082
rect 14388 13028 14444 13030
rect 14468 13028 14524 13030
rect 14548 13028 14604 13030
rect 14628 13028 14684 13030
rect 14388 11994 14444 11996
rect 14468 11994 14524 11996
rect 14548 11994 14604 11996
rect 14628 11994 14684 11996
rect 14388 11942 14434 11994
rect 14434 11942 14444 11994
rect 14468 11942 14498 11994
rect 14498 11942 14510 11994
rect 14510 11942 14524 11994
rect 14548 11942 14562 11994
rect 14562 11942 14574 11994
rect 14574 11942 14604 11994
rect 14628 11942 14638 11994
rect 14638 11942 14684 11994
rect 14388 11940 14444 11942
rect 14468 11940 14524 11942
rect 14548 11940 14604 11942
rect 14628 11940 14684 11942
rect 14388 10906 14444 10908
rect 14468 10906 14524 10908
rect 14548 10906 14604 10908
rect 14628 10906 14684 10908
rect 14388 10854 14434 10906
rect 14434 10854 14444 10906
rect 14468 10854 14498 10906
rect 14498 10854 14510 10906
rect 14510 10854 14524 10906
rect 14548 10854 14562 10906
rect 14562 10854 14574 10906
rect 14574 10854 14604 10906
rect 14628 10854 14638 10906
rect 14638 10854 14684 10906
rect 14388 10852 14444 10854
rect 14468 10852 14524 10854
rect 14548 10852 14604 10854
rect 14628 10852 14684 10854
rect 14388 9818 14444 9820
rect 14468 9818 14524 9820
rect 14548 9818 14604 9820
rect 14628 9818 14684 9820
rect 14388 9766 14434 9818
rect 14434 9766 14444 9818
rect 14468 9766 14498 9818
rect 14498 9766 14510 9818
rect 14510 9766 14524 9818
rect 14548 9766 14562 9818
rect 14562 9766 14574 9818
rect 14574 9766 14604 9818
rect 14628 9766 14638 9818
rect 14638 9766 14684 9818
rect 14388 9764 14444 9766
rect 14468 9764 14524 9766
rect 14548 9764 14604 9766
rect 14628 9764 14684 9766
rect 14002 9324 14004 9344
rect 14004 9324 14056 9344
rect 14056 9324 14058 9344
rect 14002 9288 14058 9324
rect 14186 8472 14242 8528
rect 15014 35944 15070 36000
rect 14922 30232 14978 30288
rect 15014 29688 15070 29744
rect 15014 26152 15070 26208
rect 14922 23024 14978 23080
rect 14922 22888 14978 22944
rect 15014 20712 15070 20768
rect 15014 18536 15070 18592
rect 15014 17176 15070 17232
rect 15014 16768 15070 16824
rect 15014 16360 15070 16416
rect 15014 14184 15070 14240
rect 14388 8730 14444 8732
rect 14468 8730 14524 8732
rect 14548 8730 14604 8732
rect 14628 8730 14684 8732
rect 14388 8678 14434 8730
rect 14434 8678 14444 8730
rect 14468 8678 14498 8730
rect 14498 8678 14510 8730
rect 14510 8678 14524 8730
rect 14548 8678 14562 8730
rect 14562 8678 14574 8730
rect 14574 8678 14604 8730
rect 14628 8678 14638 8730
rect 14638 8678 14684 8730
rect 14388 8676 14444 8678
rect 14468 8676 14524 8678
rect 14548 8676 14604 8678
rect 14628 8676 14684 8678
rect 14388 7642 14444 7644
rect 14468 7642 14524 7644
rect 14548 7642 14604 7644
rect 14628 7642 14684 7644
rect 14388 7590 14434 7642
rect 14434 7590 14444 7642
rect 14468 7590 14498 7642
rect 14498 7590 14510 7642
rect 14510 7590 14524 7642
rect 14548 7590 14562 7642
rect 14562 7590 14574 7642
rect 14574 7590 14604 7642
rect 14628 7590 14638 7642
rect 14638 7590 14684 7642
rect 14388 7588 14444 7590
rect 14468 7588 14524 7590
rect 14548 7588 14604 7590
rect 14628 7588 14684 7590
rect 13450 6432 13506 6488
rect 13634 5616 13690 5672
rect 13726 5208 13782 5264
rect 14388 6554 14444 6556
rect 14468 6554 14524 6556
rect 14548 6554 14604 6556
rect 14628 6554 14684 6556
rect 14388 6502 14434 6554
rect 14434 6502 14444 6554
rect 14468 6502 14498 6554
rect 14498 6502 14510 6554
rect 14510 6502 14524 6554
rect 14548 6502 14562 6554
rect 14562 6502 14574 6554
rect 14574 6502 14604 6554
rect 14628 6502 14638 6554
rect 14638 6502 14684 6554
rect 14388 6500 14444 6502
rect 14468 6500 14524 6502
rect 14548 6500 14604 6502
rect 14628 6500 14684 6502
rect 14388 5466 14444 5468
rect 14468 5466 14524 5468
rect 14548 5466 14604 5468
rect 14628 5466 14684 5468
rect 14388 5414 14434 5466
rect 14434 5414 14444 5466
rect 14468 5414 14498 5466
rect 14498 5414 14510 5466
rect 14510 5414 14524 5466
rect 14548 5414 14562 5466
rect 14562 5414 14574 5466
rect 14574 5414 14604 5466
rect 14628 5414 14638 5466
rect 14638 5414 14684 5466
rect 14388 5412 14444 5414
rect 14468 5412 14524 5414
rect 14548 5412 14604 5414
rect 14628 5412 14684 5414
rect 13910 4936 13966 4992
rect 14388 4378 14444 4380
rect 14468 4378 14524 4380
rect 14548 4378 14604 4380
rect 14628 4378 14684 4380
rect 14388 4326 14434 4378
rect 14434 4326 14444 4378
rect 14468 4326 14498 4378
rect 14498 4326 14510 4378
rect 14510 4326 14524 4378
rect 14548 4326 14562 4378
rect 14562 4326 14574 4378
rect 14574 4326 14604 4378
rect 14628 4326 14638 4378
rect 14638 4326 14684 4378
rect 14388 4324 14444 4326
rect 14468 4324 14524 4326
rect 14548 4324 14604 4326
rect 14628 4324 14684 4326
rect 14388 3290 14444 3292
rect 14468 3290 14524 3292
rect 14548 3290 14604 3292
rect 14628 3290 14684 3292
rect 14388 3238 14434 3290
rect 14434 3238 14444 3290
rect 14468 3238 14498 3290
rect 14498 3238 14510 3290
rect 14510 3238 14524 3290
rect 14548 3238 14562 3290
rect 14562 3238 14574 3290
rect 14574 3238 14604 3290
rect 14628 3238 14638 3290
rect 14638 3238 14684 3290
rect 14388 3236 14444 3238
rect 14468 3236 14524 3238
rect 14548 3236 14604 3238
rect 14628 3236 14684 3238
rect 9351 2746 9407 2748
rect 9431 2746 9487 2748
rect 9511 2746 9567 2748
rect 9591 2746 9647 2748
rect 9351 2694 9397 2746
rect 9397 2694 9407 2746
rect 9431 2694 9461 2746
rect 9461 2694 9473 2746
rect 9473 2694 9487 2746
rect 9511 2694 9525 2746
rect 9525 2694 9537 2746
rect 9537 2694 9567 2746
rect 9591 2694 9601 2746
rect 9601 2694 9647 2746
rect 9351 2692 9407 2694
rect 9431 2692 9487 2694
rect 9511 2692 9567 2694
rect 9591 2692 9647 2694
rect 12709 2746 12765 2748
rect 12789 2746 12845 2748
rect 12869 2746 12925 2748
rect 12949 2746 13005 2748
rect 12709 2694 12755 2746
rect 12755 2694 12765 2746
rect 12789 2694 12819 2746
rect 12819 2694 12831 2746
rect 12831 2694 12845 2746
rect 12869 2694 12883 2746
rect 12883 2694 12895 2746
rect 12895 2694 12925 2746
rect 12949 2694 12959 2746
rect 12959 2694 13005 2746
rect 12709 2692 12765 2694
rect 12789 2692 12845 2694
rect 12869 2692 12925 2694
rect 12949 2692 13005 2694
rect 10874 2624 10930 2680
rect 9402 2488 9458 2544
rect 11030 2202 11086 2204
rect 11110 2202 11166 2204
rect 11190 2202 11246 2204
rect 11270 2202 11326 2204
rect 11030 2150 11076 2202
rect 11076 2150 11086 2202
rect 11110 2150 11140 2202
rect 11140 2150 11152 2202
rect 11152 2150 11166 2202
rect 11190 2150 11204 2202
rect 11204 2150 11216 2202
rect 11216 2150 11246 2202
rect 11270 2150 11280 2202
rect 11280 2150 11326 2202
rect 11030 2148 11086 2150
rect 11110 2148 11166 2150
rect 11190 2148 11246 2150
rect 11270 2148 11326 2150
rect 14388 2202 14444 2204
rect 14468 2202 14524 2204
rect 14548 2202 14604 2204
rect 14628 2202 14684 2204
rect 14388 2150 14434 2202
rect 14434 2150 14444 2202
rect 14468 2150 14498 2202
rect 14498 2150 14510 2202
rect 14510 2150 14524 2202
rect 14548 2150 14562 2202
rect 14562 2150 14574 2202
rect 14574 2150 14604 2202
rect 14628 2150 14638 2202
rect 14638 2150 14684 2202
rect 14388 2148 14444 2150
rect 14468 2148 14524 2150
rect 14548 2148 14604 2150
rect 14628 2148 14684 2150
rect 10138 1944 10194 2000
rect 9351 1658 9407 1660
rect 9431 1658 9487 1660
rect 9511 1658 9567 1660
rect 9591 1658 9647 1660
rect 9351 1606 9397 1658
rect 9397 1606 9407 1658
rect 9431 1606 9461 1658
rect 9461 1606 9473 1658
rect 9473 1606 9487 1658
rect 9511 1606 9525 1658
rect 9525 1606 9537 1658
rect 9537 1606 9567 1658
rect 9591 1606 9601 1658
rect 9601 1606 9647 1658
rect 9351 1604 9407 1606
rect 9431 1604 9487 1606
rect 9511 1604 9567 1606
rect 9591 1604 9647 1606
rect 12709 1658 12765 1660
rect 12789 1658 12845 1660
rect 12869 1658 12925 1660
rect 12949 1658 13005 1660
rect 12709 1606 12755 1658
rect 12755 1606 12765 1658
rect 12789 1606 12819 1658
rect 12819 1606 12831 1658
rect 12831 1606 12845 1658
rect 12869 1606 12883 1658
rect 12883 1606 12895 1658
rect 12895 1606 12925 1658
rect 12949 1606 12959 1658
rect 12959 1606 13005 1658
rect 12709 1604 12765 1606
rect 12789 1604 12845 1606
rect 12869 1604 12925 1606
rect 12949 1604 13005 1606
rect 4618 1300 4620 1320
rect 4620 1300 4672 1320
rect 4672 1300 4674 1320
rect 4618 1264 4674 1300
rect 5170 1300 5172 1320
rect 5172 1300 5224 1320
rect 5224 1300 5226 1320
rect 5170 1264 5226 1300
rect 6642 1300 6644 1320
rect 6644 1300 6696 1320
rect 6696 1300 6698 1320
rect 4314 1114 4370 1116
rect 4394 1114 4450 1116
rect 4474 1114 4530 1116
rect 4554 1114 4610 1116
rect 4314 1062 4360 1114
rect 4360 1062 4370 1114
rect 4394 1062 4424 1114
rect 4424 1062 4436 1114
rect 4436 1062 4450 1114
rect 4474 1062 4488 1114
rect 4488 1062 4500 1114
rect 4500 1062 4530 1114
rect 4554 1062 4564 1114
rect 4564 1062 4610 1114
rect 4314 1060 4370 1062
rect 4394 1060 4450 1062
rect 4474 1060 4530 1062
rect 4554 1060 4610 1062
rect 6642 1264 6698 1300
rect 7672 1114 7728 1116
rect 7752 1114 7808 1116
rect 7832 1114 7888 1116
rect 7912 1114 7968 1116
rect 7672 1062 7718 1114
rect 7718 1062 7728 1114
rect 7752 1062 7782 1114
rect 7782 1062 7794 1114
rect 7794 1062 7808 1114
rect 7832 1062 7846 1114
rect 7846 1062 7858 1114
rect 7858 1062 7888 1114
rect 7912 1062 7922 1114
rect 7922 1062 7968 1114
rect 7672 1060 7728 1062
rect 7752 1060 7808 1062
rect 7832 1060 7888 1062
rect 7912 1060 7968 1062
rect 11030 1114 11086 1116
rect 11110 1114 11166 1116
rect 11190 1114 11246 1116
rect 11270 1114 11326 1116
rect 11030 1062 11076 1114
rect 11076 1062 11086 1114
rect 11110 1062 11140 1114
rect 11140 1062 11152 1114
rect 11152 1062 11166 1114
rect 11190 1062 11204 1114
rect 11204 1062 11216 1114
rect 11216 1062 11246 1114
rect 11270 1062 11280 1114
rect 11280 1062 11326 1114
rect 11030 1060 11086 1062
rect 11110 1060 11166 1062
rect 11190 1060 11246 1062
rect 11270 1060 11326 1062
rect 13818 1264 13874 1320
rect 14830 8744 14886 8800
rect 14830 7656 14886 7712
rect 15198 27240 15254 27296
rect 15382 28600 15438 28656
rect 15382 27512 15438 27568
rect 15290 21800 15346 21856
rect 15198 21392 15254 21448
rect 15290 18264 15346 18320
rect 15382 16496 15438 16552
rect 15290 15952 15346 16008
rect 15382 14592 15438 14648
rect 15290 9560 15346 9616
rect 14830 5616 14886 5672
rect 14388 1114 14444 1116
rect 14468 1114 14524 1116
rect 14548 1114 14604 1116
rect 14628 1114 14684 1116
rect 14388 1062 14434 1114
rect 14434 1062 14444 1114
rect 14468 1062 14498 1114
rect 14498 1062 14510 1114
rect 14510 1062 14524 1114
rect 14548 1062 14562 1114
rect 14562 1062 14574 1114
rect 14574 1062 14604 1114
rect 14628 1062 14638 1114
rect 14638 1062 14684 1114
rect 14388 1060 14444 1062
rect 14468 1060 14524 1062
rect 14548 1060 14604 1062
rect 14628 1060 14684 1062
<< metal3 >>
rect 4304 43552 4620 43553
rect 4304 43488 4310 43552
rect 4374 43488 4390 43552
rect 4454 43488 4470 43552
rect 4534 43488 4550 43552
rect 4614 43488 4620 43552
rect 4304 43487 4620 43488
rect 7662 43552 7978 43553
rect 7662 43488 7668 43552
rect 7732 43488 7748 43552
rect 7812 43488 7828 43552
rect 7892 43488 7908 43552
rect 7972 43488 7978 43552
rect 7662 43487 7978 43488
rect 11020 43552 11336 43553
rect 11020 43488 11026 43552
rect 11090 43488 11106 43552
rect 11170 43488 11186 43552
rect 11250 43488 11266 43552
rect 11330 43488 11336 43552
rect 11020 43487 11336 43488
rect 14378 43552 14694 43553
rect 14378 43488 14384 43552
rect 14448 43488 14464 43552
rect 14528 43488 14544 43552
rect 14608 43488 14624 43552
rect 14688 43488 14694 43552
rect 14378 43487 14694 43488
rect 2625 43008 2941 43009
rect 2625 42944 2631 43008
rect 2695 42944 2711 43008
rect 2775 42944 2791 43008
rect 2855 42944 2871 43008
rect 2935 42944 2941 43008
rect 2625 42943 2941 42944
rect 5983 43008 6299 43009
rect 5983 42944 5989 43008
rect 6053 42944 6069 43008
rect 6133 42944 6149 43008
rect 6213 42944 6229 43008
rect 6293 42944 6299 43008
rect 5983 42943 6299 42944
rect 9341 43008 9657 43009
rect 9341 42944 9347 43008
rect 9411 42944 9427 43008
rect 9491 42944 9507 43008
rect 9571 42944 9587 43008
rect 9651 42944 9657 43008
rect 9341 42943 9657 42944
rect 12699 43008 13015 43009
rect 12699 42944 12705 43008
rect 12769 42944 12785 43008
rect 12849 42944 12865 43008
rect 12929 42944 12945 43008
rect 13009 42944 13015 43008
rect 12699 42943 13015 42944
rect 3918 42740 3924 42804
rect 3988 42802 3994 42804
rect 10041 42802 10107 42805
rect 3988 42800 10107 42802
rect 3988 42744 10046 42800
rect 10102 42744 10107 42800
rect 3988 42742 10107 42744
rect 3988 42740 3994 42742
rect 10041 42739 10107 42742
rect 3734 42604 3740 42668
rect 3804 42666 3810 42668
rect 7925 42666 7991 42669
rect 3804 42664 7991 42666
rect 3804 42608 7930 42664
rect 7986 42608 7991 42664
rect 3804 42606 7991 42608
rect 3804 42604 3810 42606
rect 7925 42603 7991 42606
rect 4304 42464 4620 42465
rect 4304 42400 4310 42464
rect 4374 42400 4390 42464
rect 4454 42400 4470 42464
rect 4534 42400 4550 42464
rect 4614 42400 4620 42464
rect 4304 42399 4620 42400
rect 7662 42464 7978 42465
rect 7662 42400 7668 42464
rect 7732 42400 7748 42464
rect 7812 42400 7828 42464
rect 7892 42400 7908 42464
rect 7972 42400 7978 42464
rect 7662 42399 7978 42400
rect 11020 42464 11336 42465
rect 11020 42400 11026 42464
rect 11090 42400 11106 42464
rect 11170 42400 11186 42464
rect 11250 42400 11266 42464
rect 11330 42400 11336 42464
rect 11020 42399 11336 42400
rect 14378 42464 14694 42465
rect 14378 42400 14384 42464
rect 14448 42400 14464 42464
rect 14528 42400 14544 42464
rect 14608 42400 14624 42464
rect 14688 42400 14694 42464
rect 14378 42399 14694 42400
rect 2262 42060 2268 42124
rect 2332 42122 2338 42124
rect 8661 42122 8727 42125
rect 2332 42120 8727 42122
rect 2332 42064 8666 42120
rect 8722 42064 8727 42120
rect 2332 42062 8727 42064
rect 2332 42060 2338 42062
rect 8661 42059 8727 42062
rect 2625 41920 2941 41921
rect 2625 41856 2631 41920
rect 2695 41856 2711 41920
rect 2775 41856 2791 41920
rect 2855 41856 2871 41920
rect 2935 41856 2941 41920
rect 2625 41855 2941 41856
rect 5983 41920 6299 41921
rect 5983 41856 5989 41920
rect 6053 41856 6069 41920
rect 6133 41856 6149 41920
rect 6213 41856 6229 41920
rect 6293 41856 6299 41920
rect 5983 41855 6299 41856
rect 9341 41920 9657 41921
rect 9341 41856 9347 41920
rect 9411 41856 9427 41920
rect 9491 41856 9507 41920
rect 9571 41856 9587 41920
rect 9651 41856 9657 41920
rect 9341 41855 9657 41856
rect 12699 41920 13015 41921
rect 12699 41856 12705 41920
rect 12769 41856 12785 41920
rect 12849 41856 12865 41920
rect 12929 41856 12945 41920
rect 13009 41856 13015 41920
rect 12699 41855 13015 41856
rect 2078 41652 2084 41716
rect 2148 41714 2154 41716
rect 7189 41714 7255 41717
rect 2148 41712 7255 41714
rect 2148 41656 7194 41712
rect 7250 41656 7255 41712
rect 2148 41654 7255 41656
rect 2148 41652 2154 41654
rect 7189 41651 7255 41654
rect 4245 41578 4311 41581
rect 4838 41578 4844 41580
rect 4245 41576 4844 41578
rect 4245 41520 4250 41576
rect 4306 41520 4844 41576
rect 4245 41518 4844 41520
rect 4245 41515 4311 41518
rect 4838 41516 4844 41518
rect 4908 41516 4914 41580
rect 13813 41578 13879 41581
rect 14958 41578 14964 41580
rect 13813 41576 14964 41578
rect 13813 41520 13818 41576
rect 13874 41520 14964 41576
rect 13813 41518 14964 41520
rect 13813 41515 13879 41518
rect 14958 41516 14964 41518
rect 15028 41516 15034 41580
rect 1393 41442 1459 41445
rect 1526 41442 1532 41444
rect 1393 41440 1532 41442
rect 1393 41384 1398 41440
rect 1454 41384 1532 41440
rect 1393 41382 1532 41384
rect 1393 41379 1459 41382
rect 1526 41380 1532 41382
rect 1596 41380 1602 41444
rect 4889 41442 4955 41445
rect 5206 41442 5212 41444
rect 4889 41440 5212 41442
rect 4889 41384 4894 41440
rect 4950 41384 5212 41440
rect 4889 41382 5212 41384
rect 4889 41379 4955 41382
rect 5206 41380 5212 41382
rect 5276 41380 5282 41444
rect 6453 41442 6519 41445
rect 6678 41442 6684 41444
rect 6453 41440 6684 41442
rect 6453 41384 6458 41440
rect 6514 41384 6684 41440
rect 6453 41382 6684 41384
rect 6453 41379 6519 41382
rect 6678 41380 6684 41382
rect 6748 41380 6754 41444
rect 4304 41376 4620 41377
rect 4304 41312 4310 41376
rect 4374 41312 4390 41376
rect 4454 41312 4470 41376
rect 4534 41312 4550 41376
rect 4614 41312 4620 41376
rect 4304 41311 4620 41312
rect 7662 41376 7978 41377
rect 7662 41312 7668 41376
rect 7732 41312 7748 41376
rect 7812 41312 7828 41376
rect 7892 41312 7908 41376
rect 7972 41312 7978 41376
rect 7662 41311 7978 41312
rect 11020 41376 11336 41377
rect 11020 41312 11026 41376
rect 11090 41312 11106 41376
rect 11170 41312 11186 41376
rect 11250 41312 11266 41376
rect 11330 41312 11336 41376
rect 11020 41311 11336 41312
rect 14378 41376 14694 41377
rect 14378 41312 14384 41376
rect 14448 41312 14464 41376
rect 14528 41312 14544 41376
rect 14608 41312 14624 41376
rect 14688 41312 14694 41376
rect 14378 41311 14694 41312
rect 2625 40832 2941 40833
rect 2625 40768 2631 40832
rect 2695 40768 2711 40832
rect 2775 40768 2791 40832
rect 2855 40768 2871 40832
rect 2935 40768 2941 40832
rect 2625 40767 2941 40768
rect 5983 40832 6299 40833
rect 5983 40768 5989 40832
rect 6053 40768 6069 40832
rect 6133 40768 6149 40832
rect 6213 40768 6229 40832
rect 6293 40768 6299 40832
rect 5983 40767 6299 40768
rect 9341 40832 9657 40833
rect 9341 40768 9347 40832
rect 9411 40768 9427 40832
rect 9491 40768 9507 40832
rect 9571 40768 9587 40832
rect 9651 40768 9657 40832
rect 9341 40767 9657 40768
rect 12699 40832 13015 40833
rect 12699 40768 12705 40832
rect 12769 40768 12785 40832
rect 12849 40768 12865 40832
rect 12929 40768 12945 40832
rect 13009 40768 13015 40832
rect 12699 40767 13015 40768
rect -300 40626 160 40656
rect 749 40626 815 40629
rect -300 40624 815 40626
rect -300 40568 754 40624
rect 810 40568 815 40624
rect -300 40566 815 40568
rect -300 40536 160 40566
rect 749 40563 815 40566
rect 4304 40288 4620 40289
rect 4304 40224 4310 40288
rect 4374 40224 4390 40288
rect 4454 40224 4470 40288
rect 4534 40224 4550 40288
rect 4614 40224 4620 40288
rect 4304 40223 4620 40224
rect 7662 40288 7978 40289
rect 7662 40224 7668 40288
rect 7732 40224 7748 40288
rect 7812 40224 7828 40288
rect 7892 40224 7908 40288
rect 7972 40224 7978 40288
rect 7662 40223 7978 40224
rect 11020 40288 11336 40289
rect 11020 40224 11026 40288
rect 11090 40224 11106 40288
rect 11170 40224 11186 40288
rect 11250 40224 11266 40288
rect 11330 40224 11336 40288
rect 11020 40223 11336 40224
rect 14378 40288 14694 40289
rect 14378 40224 14384 40288
rect 14448 40224 14464 40288
rect 14528 40224 14544 40288
rect 14608 40224 14624 40288
rect 14688 40224 14694 40288
rect 14378 40223 14694 40224
rect 1485 39944 1551 39949
rect 1485 39888 1490 39944
rect 1546 39888 1551 39944
rect 1485 39883 1551 39888
rect -300 39810 160 39840
rect 1488 39810 1548 39883
rect -300 39750 1548 39810
rect -300 39720 160 39750
rect 2625 39744 2941 39745
rect 2625 39680 2631 39744
rect 2695 39680 2711 39744
rect 2775 39680 2791 39744
rect 2855 39680 2871 39744
rect 2935 39680 2941 39744
rect 2625 39679 2941 39680
rect 5983 39744 6299 39745
rect 5983 39680 5989 39744
rect 6053 39680 6069 39744
rect 6133 39680 6149 39744
rect 6213 39680 6229 39744
rect 6293 39680 6299 39744
rect 5983 39679 6299 39680
rect 9341 39744 9657 39745
rect 9341 39680 9347 39744
rect 9411 39680 9427 39744
rect 9491 39680 9507 39744
rect 9571 39680 9587 39744
rect 9651 39680 9657 39744
rect 9341 39679 9657 39680
rect 12699 39744 13015 39745
rect 12699 39680 12705 39744
rect 12769 39680 12785 39744
rect 12849 39680 12865 39744
rect 12929 39680 12945 39744
rect 13009 39680 13015 39744
rect 12699 39679 13015 39680
rect 14089 39538 14155 39541
rect 15540 39538 16000 39568
rect 14089 39536 16000 39538
rect 14089 39480 14094 39536
rect 14150 39480 16000 39536
rect 14089 39478 16000 39480
rect 14089 39475 14155 39478
rect 15540 39448 16000 39478
rect 14825 39266 14891 39269
rect 15540 39266 16000 39296
rect 14825 39264 16000 39266
rect 14825 39208 14830 39264
rect 14886 39208 16000 39264
rect 14825 39206 16000 39208
rect 14825 39203 14891 39206
rect 4304 39200 4620 39201
rect 4304 39136 4310 39200
rect 4374 39136 4390 39200
rect 4454 39136 4470 39200
rect 4534 39136 4550 39200
rect 4614 39136 4620 39200
rect 4304 39135 4620 39136
rect 7662 39200 7978 39201
rect 7662 39136 7668 39200
rect 7732 39136 7748 39200
rect 7812 39136 7828 39200
rect 7892 39136 7908 39200
rect 7972 39136 7978 39200
rect 7662 39135 7978 39136
rect 11020 39200 11336 39201
rect 11020 39136 11026 39200
rect 11090 39136 11106 39200
rect 11170 39136 11186 39200
rect 11250 39136 11266 39200
rect 11330 39136 11336 39200
rect 11020 39135 11336 39136
rect 14378 39200 14694 39201
rect 14378 39136 14384 39200
rect 14448 39136 14464 39200
rect 14528 39136 14544 39200
rect 14608 39136 14624 39200
rect 14688 39136 14694 39200
rect 15540 39176 16000 39206
rect 14378 39135 14694 39136
rect -300 38994 160 39024
rect 749 38994 815 38997
rect -300 38992 815 38994
rect -300 38936 754 38992
rect 810 38936 815 38992
rect -300 38934 815 38936
rect -300 38904 160 38934
rect 749 38931 815 38934
rect 14273 38994 14339 38997
rect 15540 38994 16000 39024
rect 14273 38992 16000 38994
rect 14273 38936 14278 38992
rect 14334 38936 16000 38992
rect 14273 38934 16000 38936
rect 14273 38931 14339 38934
rect 15540 38904 16000 38934
rect 13905 38722 13971 38725
rect 15540 38722 16000 38752
rect 13905 38720 16000 38722
rect 13905 38664 13910 38720
rect 13966 38664 16000 38720
rect 13905 38662 16000 38664
rect 13905 38659 13971 38662
rect 2625 38656 2941 38657
rect 2625 38592 2631 38656
rect 2695 38592 2711 38656
rect 2775 38592 2791 38656
rect 2855 38592 2871 38656
rect 2935 38592 2941 38656
rect 2625 38591 2941 38592
rect 5983 38656 6299 38657
rect 5983 38592 5989 38656
rect 6053 38592 6069 38656
rect 6133 38592 6149 38656
rect 6213 38592 6229 38656
rect 6293 38592 6299 38656
rect 5983 38591 6299 38592
rect 9341 38656 9657 38657
rect 9341 38592 9347 38656
rect 9411 38592 9427 38656
rect 9491 38592 9507 38656
rect 9571 38592 9587 38656
rect 9651 38592 9657 38656
rect 9341 38591 9657 38592
rect 12699 38656 13015 38657
rect 12699 38592 12705 38656
rect 12769 38592 12785 38656
rect 12849 38592 12865 38656
rect 12929 38592 12945 38656
rect 13009 38592 13015 38656
rect 15540 38632 16000 38662
rect 12699 38591 13015 38592
rect 13353 38450 13419 38453
rect 15540 38450 16000 38480
rect 13353 38448 16000 38450
rect 13353 38392 13358 38448
rect 13414 38392 16000 38448
rect 13353 38390 16000 38392
rect 13353 38387 13419 38390
rect 15540 38360 16000 38390
rect -300 38178 160 38208
rect 749 38178 815 38181
rect -300 38176 815 38178
rect -300 38120 754 38176
rect 810 38120 815 38176
rect -300 38118 815 38120
rect -300 38088 160 38118
rect 749 38115 815 38118
rect 14825 38178 14891 38181
rect 15540 38178 16000 38208
rect 14825 38176 16000 38178
rect 14825 38120 14830 38176
rect 14886 38120 16000 38176
rect 14825 38118 16000 38120
rect 14825 38115 14891 38118
rect 4304 38112 4620 38113
rect 4304 38048 4310 38112
rect 4374 38048 4390 38112
rect 4454 38048 4470 38112
rect 4534 38048 4550 38112
rect 4614 38048 4620 38112
rect 4304 38047 4620 38048
rect 7662 38112 7978 38113
rect 7662 38048 7668 38112
rect 7732 38048 7748 38112
rect 7812 38048 7828 38112
rect 7892 38048 7908 38112
rect 7972 38048 7978 38112
rect 7662 38047 7978 38048
rect 11020 38112 11336 38113
rect 11020 38048 11026 38112
rect 11090 38048 11106 38112
rect 11170 38048 11186 38112
rect 11250 38048 11266 38112
rect 11330 38048 11336 38112
rect 11020 38047 11336 38048
rect 14378 38112 14694 38113
rect 14378 38048 14384 38112
rect 14448 38048 14464 38112
rect 14528 38048 14544 38112
rect 14608 38048 14624 38112
rect 14688 38048 14694 38112
rect 15540 38088 16000 38118
rect 14378 38047 14694 38048
rect 14273 37906 14339 37909
rect 15540 37906 16000 37936
rect 14273 37904 16000 37906
rect 14273 37848 14278 37904
rect 14334 37848 16000 37904
rect 14273 37846 16000 37848
rect 14273 37843 14339 37846
rect 15540 37816 16000 37846
rect 14365 37634 14431 37637
rect 15540 37634 16000 37664
rect 14365 37632 16000 37634
rect 14365 37576 14370 37632
rect 14426 37576 16000 37632
rect 14365 37574 16000 37576
rect 14365 37571 14431 37574
rect 2625 37568 2941 37569
rect 2625 37504 2631 37568
rect 2695 37504 2711 37568
rect 2775 37504 2791 37568
rect 2855 37504 2871 37568
rect 2935 37504 2941 37568
rect 2625 37503 2941 37504
rect 5983 37568 6299 37569
rect 5983 37504 5989 37568
rect 6053 37504 6069 37568
rect 6133 37504 6149 37568
rect 6213 37504 6229 37568
rect 6293 37504 6299 37568
rect 5983 37503 6299 37504
rect 9341 37568 9657 37569
rect 9341 37504 9347 37568
rect 9411 37504 9427 37568
rect 9491 37504 9507 37568
rect 9571 37504 9587 37568
rect 9651 37504 9657 37568
rect 9341 37503 9657 37504
rect 12699 37568 13015 37569
rect 12699 37504 12705 37568
rect 12769 37504 12785 37568
rect 12849 37504 12865 37568
rect 12929 37504 12945 37568
rect 13009 37504 13015 37568
rect 15540 37544 16000 37574
rect 12699 37503 13015 37504
rect -300 37362 160 37392
rect 749 37362 815 37365
rect 10409 37364 10475 37365
rect 10358 37362 10364 37364
rect -300 37360 815 37362
rect -300 37304 754 37360
rect 810 37304 815 37360
rect -300 37302 815 37304
rect 10318 37302 10364 37362
rect 10428 37360 10475 37364
rect 10470 37304 10475 37360
rect -300 37272 160 37302
rect 749 37299 815 37302
rect 10358 37300 10364 37302
rect 10428 37300 10475 37304
rect 10409 37299 10475 37300
rect 11789 37364 11855 37365
rect 11789 37360 11836 37364
rect 11900 37362 11906 37364
rect 14181 37362 14247 37365
rect 15540 37362 16000 37392
rect 11789 37304 11794 37360
rect 11789 37300 11836 37304
rect 11900 37302 11946 37362
rect 14181 37360 16000 37362
rect 14181 37304 14186 37360
rect 14242 37304 16000 37360
rect 14181 37302 16000 37304
rect 11900 37300 11906 37302
rect 11789 37299 11855 37300
rect 14181 37299 14247 37302
rect 15540 37272 16000 37302
rect 11697 37226 11763 37229
rect 12341 37226 12407 37229
rect 11697 37224 12407 37226
rect 11697 37168 11702 37224
rect 11758 37168 12346 37224
rect 12402 37168 12407 37224
rect 11697 37166 12407 37168
rect 11697 37163 11763 37166
rect 12341 37163 12407 37166
rect 14230 37166 14842 37226
rect 13353 37090 13419 37093
rect 14230 37090 14290 37166
rect 13353 37088 14290 37090
rect 13353 37032 13358 37088
rect 13414 37032 14290 37088
rect 13353 37030 14290 37032
rect 14782 37090 14842 37166
rect 15540 37090 16000 37120
rect 14782 37030 16000 37090
rect 13353 37027 13419 37030
rect 4304 37024 4620 37025
rect 4304 36960 4310 37024
rect 4374 36960 4390 37024
rect 4454 36960 4470 37024
rect 4534 36960 4550 37024
rect 4614 36960 4620 37024
rect 4304 36959 4620 36960
rect 7662 37024 7978 37025
rect 7662 36960 7668 37024
rect 7732 36960 7748 37024
rect 7812 36960 7828 37024
rect 7892 36960 7908 37024
rect 7972 36960 7978 37024
rect 7662 36959 7978 36960
rect 11020 37024 11336 37025
rect 11020 36960 11026 37024
rect 11090 36960 11106 37024
rect 11170 36960 11186 37024
rect 11250 36960 11266 37024
rect 11330 36960 11336 37024
rect 11020 36959 11336 36960
rect 14378 37024 14694 37025
rect 14378 36960 14384 37024
rect 14448 36960 14464 37024
rect 14528 36960 14544 37024
rect 14608 36960 14624 37024
rect 14688 36960 14694 37024
rect 15540 37000 16000 37030
rect 14378 36959 14694 36960
rect 11421 36954 11487 36957
rect 12709 36954 12775 36957
rect 11421 36952 12775 36954
rect 11421 36896 11426 36952
rect 11482 36896 12714 36952
rect 12770 36896 12775 36952
rect 11421 36894 12775 36896
rect 11421 36891 11487 36894
rect 12709 36891 12775 36894
rect 13721 36818 13787 36821
rect 15540 36818 16000 36848
rect 13721 36816 16000 36818
rect 13721 36760 13726 36816
rect 13782 36760 16000 36816
rect 13721 36758 16000 36760
rect 13721 36755 13787 36758
rect 15540 36728 16000 36758
rect -300 36546 160 36576
rect 749 36546 815 36549
rect -300 36544 815 36546
rect -300 36488 754 36544
rect 810 36488 815 36544
rect -300 36486 815 36488
rect -300 36456 160 36486
rect 749 36483 815 36486
rect 13629 36546 13695 36549
rect 15540 36546 16000 36576
rect 13629 36544 16000 36546
rect 13629 36488 13634 36544
rect 13690 36488 16000 36544
rect 13629 36486 16000 36488
rect 13629 36483 13695 36486
rect 2625 36480 2941 36481
rect 2625 36416 2631 36480
rect 2695 36416 2711 36480
rect 2775 36416 2791 36480
rect 2855 36416 2871 36480
rect 2935 36416 2941 36480
rect 2625 36415 2941 36416
rect 5983 36480 6299 36481
rect 5983 36416 5989 36480
rect 6053 36416 6069 36480
rect 6133 36416 6149 36480
rect 6213 36416 6229 36480
rect 6293 36416 6299 36480
rect 5983 36415 6299 36416
rect 9341 36480 9657 36481
rect 9341 36416 9347 36480
rect 9411 36416 9427 36480
rect 9491 36416 9507 36480
rect 9571 36416 9587 36480
rect 9651 36416 9657 36480
rect 9341 36415 9657 36416
rect 12699 36480 13015 36481
rect 12699 36416 12705 36480
rect 12769 36416 12785 36480
rect 12849 36416 12865 36480
rect 12929 36416 12945 36480
rect 13009 36416 13015 36480
rect 15540 36456 16000 36486
rect 12699 36415 13015 36416
rect 14181 36274 14247 36277
rect 15540 36274 16000 36304
rect 14181 36272 16000 36274
rect 14181 36216 14186 36272
rect 14242 36216 16000 36272
rect 14181 36214 16000 36216
rect 14181 36211 14247 36214
rect 15540 36184 16000 36214
rect 15009 36002 15075 36005
rect 15540 36002 16000 36032
rect 15009 36000 16000 36002
rect 15009 35944 15014 36000
rect 15070 35944 16000 36000
rect 15009 35942 16000 35944
rect 15009 35939 15075 35942
rect 4304 35936 4620 35937
rect 4304 35872 4310 35936
rect 4374 35872 4390 35936
rect 4454 35872 4470 35936
rect 4534 35872 4550 35936
rect 4614 35872 4620 35936
rect 4304 35871 4620 35872
rect 7662 35936 7978 35937
rect 7662 35872 7668 35936
rect 7732 35872 7748 35936
rect 7812 35872 7828 35936
rect 7892 35872 7908 35936
rect 7972 35872 7978 35936
rect 7662 35871 7978 35872
rect 11020 35936 11336 35937
rect 11020 35872 11026 35936
rect 11090 35872 11106 35936
rect 11170 35872 11186 35936
rect 11250 35872 11266 35936
rect 11330 35872 11336 35936
rect 11020 35871 11336 35872
rect 14378 35936 14694 35937
rect 14378 35872 14384 35936
rect 14448 35872 14464 35936
rect 14528 35872 14544 35936
rect 14608 35872 14624 35936
rect 14688 35872 14694 35936
rect 15540 35912 16000 35942
rect 14378 35871 14694 35872
rect 1485 35864 1551 35869
rect 1485 35808 1490 35864
rect 1546 35808 1551 35864
rect 1485 35803 1551 35808
rect -300 35730 160 35760
rect 1488 35730 1548 35803
rect -300 35670 1548 35730
rect 12617 35730 12683 35733
rect 15540 35730 16000 35760
rect 12617 35728 16000 35730
rect 12617 35672 12622 35728
rect 12678 35672 16000 35728
rect 12617 35670 16000 35672
rect -300 35640 160 35670
rect 12617 35667 12683 35670
rect 15540 35640 16000 35670
rect 6453 35594 6519 35597
rect 12709 35594 12775 35597
rect 6453 35592 12775 35594
rect 6453 35536 6458 35592
rect 6514 35536 12714 35592
rect 12770 35536 12775 35592
rect 6453 35534 12775 35536
rect 6453 35531 6519 35534
rect 12709 35531 12775 35534
rect 13169 35458 13235 35461
rect 15540 35458 16000 35488
rect 13169 35456 16000 35458
rect 13169 35400 13174 35456
rect 13230 35400 16000 35456
rect 13169 35398 16000 35400
rect 13169 35395 13235 35398
rect 2625 35392 2941 35393
rect 2625 35328 2631 35392
rect 2695 35328 2711 35392
rect 2775 35328 2791 35392
rect 2855 35328 2871 35392
rect 2935 35328 2941 35392
rect 2625 35327 2941 35328
rect 5983 35392 6299 35393
rect 5983 35328 5989 35392
rect 6053 35328 6069 35392
rect 6133 35328 6149 35392
rect 6213 35328 6229 35392
rect 6293 35328 6299 35392
rect 5983 35327 6299 35328
rect 9341 35392 9657 35393
rect 9341 35328 9347 35392
rect 9411 35328 9427 35392
rect 9491 35328 9507 35392
rect 9571 35328 9587 35392
rect 9651 35328 9657 35392
rect 9341 35327 9657 35328
rect 12699 35392 13015 35393
rect 12699 35328 12705 35392
rect 12769 35328 12785 35392
rect 12849 35328 12865 35392
rect 12929 35328 12945 35392
rect 13009 35328 13015 35392
rect 15540 35368 16000 35398
rect 12699 35327 13015 35328
rect 13997 35186 14063 35189
rect 15540 35186 16000 35216
rect 13997 35184 16000 35186
rect 13997 35128 14002 35184
rect 14058 35128 16000 35184
rect 13997 35126 16000 35128
rect 13997 35123 14063 35126
rect 15540 35096 16000 35126
rect 13721 35050 13787 35053
rect 13721 35048 14842 35050
rect 13721 34992 13726 35048
rect 13782 34992 14842 35048
rect 13721 34990 14842 34992
rect 13721 34987 13787 34990
rect -300 34914 160 34944
rect 749 34914 815 34917
rect -300 34912 815 34914
rect -300 34856 754 34912
rect 810 34856 815 34912
rect -300 34854 815 34856
rect 14782 34914 14842 34990
rect 15540 34914 16000 34944
rect 14782 34854 16000 34914
rect -300 34824 160 34854
rect 749 34851 815 34854
rect 4304 34848 4620 34849
rect 4304 34784 4310 34848
rect 4374 34784 4390 34848
rect 4454 34784 4470 34848
rect 4534 34784 4550 34848
rect 4614 34784 4620 34848
rect 4304 34783 4620 34784
rect 7662 34848 7978 34849
rect 7662 34784 7668 34848
rect 7732 34784 7748 34848
rect 7812 34784 7828 34848
rect 7892 34784 7908 34848
rect 7972 34784 7978 34848
rect 7662 34783 7978 34784
rect 11020 34848 11336 34849
rect 11020 34784 11026 34848
rect 11090 34784 11106 34848
rect 11170 34784 11186 34848
rect 11250 34784 11266 34848
rect 11330 34784 11336 34848
rect 11020 34783 11336 34784
rect 14378 34848 14694 34849
rect 14378 34784 14384 34848
rect 14448 34784 14464 34848
rect 14528 34784 14544 34848
rect 14608 34784 14624 34848
rect 14688 34784 14694 34848
rect 15540 34824 16000 34854
rect 14378 34783 14694 34784
rect 5717 34642 5783 34645
rect 6494 34642 6500 34644
rect 5717 34640 6500 34642
rect 5717 34584 5722 34640
rect 5778 34584 6500 34640
rect 5717 34582 6500 34584
rect 5717 34579 5783 34582
rect 6494 34580 6500 34582
rect 6564 34580 6570 34644
rect 12566 34580 12572 34644
rect 12636 34642 12642 34644
rect 13077 34642 13143 34645
rect 12636 34640 13143 34642
rect 12636 34584 13082 34640
rect 13138 34584 13143 34640
rect 12636 34582 13143 34584
rect 12636 34580 12642 34582
rect 13077 34579 13143 34582
rect 13537 34642 13603 34645
rect 15540 34642 16000 34672
rect 13537 34640 16000 34642
rect 13537 34584 13542 34640
rect 13598 34584 16000 34640
rect 13537 34582 16000 34584
rect 13537 34579 13603 34582
rect 15540 34552 16000 34582
rect 1393 34506 1459 34509
rect 798 34504 1459 34506
rect 798 34448 1398 34504
rect 1454 34448 1459 34504
rect 798 34446 1459 34448
rect -300 34098 160 34128
rect 798 34098 858 34446
rect 1393 34443 1459 34446
rect 13445 34370 13511 34373
rect 15540 34370 16000 34400
rect 13445 34368 16000 34370
rect 13445 34312 13450 34368
rect 13506 34312 16000 34368
rect 13445 34310 16000 34312
rect 13445 34307 13511 34310
rect 2625 34304 2941 34305
rect 2625 34240 2631 34304
rect 2695 34240 2711 34304
rect 2775 34240 2791 34304
rect 2855 34240 2871 34304
rect 2935 34240 2941 34304
rect 2625 34239 2941 34240
rect 5983 34304 6299 34305
rect 5983 34240 5989 34304
rect 6053 34240 6069 34304
rect 6133 34240 6149 34304
rect 6213 34240 6229 34304
rect 6293 34240 6299 34304
rect 5983 34239 6299 34240
rect 9341 34304 9657 34305
rect 9341 34240 9347 34304
rect 9411 34240 9427 34304
rect 9491 34240 9507 34304
rect 9571 34240 9587 34304
rect 9651 34240 9657 34304
rect 9341 34239 9657 34240
rect 12699 34304 13015 34305
rect 12699 34240 12705 34304
rect 12769 34240 12785 34304
rect 12849 34240 12865 34304
rect 12929 34240 12945 34304
rect 13009 34240 13015 34304
rect 15540 34280 16000 34310
rect 12699 34239 13015 34240
rect 13261 34234 13327 34237
rect 13721 34234 13787 34237
rect 13261 34232 13787 34234
rect 13261 34176 13266 34232
rect 13322 34176 13726 34232
rect 13782 34176 13787 34232
rect 13261 34174 13787 34176
rect 13261 34171 13327 34174
rect 13721 34171 13787 34174
rect -300 34038 858 34098
rect 11329 34098 11395 34101
rect 15540 34098 16000 34128
rect 11329 34096 16000 34098
rect 11329 34040 11334 34096
rect 11390 34040 16000 34096
rect 11329 34038 16000 34040
rect -300 34008 160 34038
rect 11329 34035 11395 34038
rect 15540 34008 16000 34038
rect 9857 33962 9923 33965
rect 10174 33962 10180 33964
rect 9857 33960 10180 33962
rect 9857 33904 9862 33960
rect 9918 33904 10180 33960
rect 9857 33902 10180 33904
rect 9857 33899 9923 33902
rect 10174 33900 10180 33902
rect 10244 33900 10250 33964
rect 10726 33900 10732 33964
rect 10796 33962 10802 33964
rect 12065 33962 12131 33965
rect 10796 33960 12131 33962
rect 10796 33904 12070 33960
rect 12126 33904 12131 33960
rect 10796 33902 12131 33904
rect 10796 33900 10802 33902
rect 12065 33899 12131 33902
rect 13721 33962 13787 33965
rect 13721 33960 14842 33962
rect 13721 33904 13726 33960
rect 13782 33904 14842 33960
rect 13721 33902 14842 33904
rect 13721 33899 13787 33902
rect 14782 33826 14842 33902
rect 15540 33826 16000 33856
rect 14782 33766 16000 33826
rect 4304 33760 4620 33761
rect 4304 33696 4310 33760
rect 4374 33696 4390 33760
rect 4454 33696 4470 33760
rect 4534 33696 4550 33760
rect 4614 33696 4620 33760
rect 4304 33695 4620 33696
rect 7662 33760 7978 33761
rect 7662 33696 7668 33760
rect 7732 33696 7748 33760
rect 7812 33696 7828 33760
rect 7892 33696 7908 33760
rect 7972 33696 7978 33760
rect 7662 33695 7978 33696
rect 11020 33760 11336 33761
rect 11020 33696 11026 33760
rect 11090 33696 11106 33760
rect 11170 33696 11186 33760
rect 11250 33696 11266 33760
rect 11330 33696 11336 33760
rect 11020 33695 11336 33696
rect 14378 33760 14694 33761
rect 14378 33696 14384 33760
rect 14448 33696 14464 33760
rect 14528 33696 14544 33760
rect 14608 33696 14624 33760
rect 14688 33696 14694 33760
rect 15540 33736 16000 33766
rect 14378 33695 14694 33696
rect 13629 33554 13695 33557
rect 15540 33554 16000 33584
rect 13629 33552 16000 33554
rect 13629 33496 13634 33552
rect 13690 33496 16000 33552
rect 13629 33494 16000 33496
rect 13629 33491 13695 33494
rect 15540 33464 16000 33494
rect -300 33282 160 33312
rect 749 33282 815 33285
rect -300 33280 815 33282
rect -300 33224 754 33280
rect 810 33224 815 33280
rect -300 33222 815 33224
rect -300 33192 160 33222
rect 749 33219 815 33222
rect 14089 33282 14155 33285
rect 15540 33282 16000 33312
rect 14089 33280 16000 33282
rect 14089 33224 14094 33280
rect 14150 33224 16000 33280
rect 14089 33222 16000 33224
rect 14089 33219 14155 33222
rect 2625 33216 2941 33217
rect 2625 33152 2631 33216
rect 2695 33152 2711 33216
rect 2775 33152 2791 33216
rect 2855 33152 2871 33216
rect 2935 33152 2941 33216
rect 2625 33151 2941 33152
rect 5983 33216 6299 33217
rect 5983 33152 5989 33216
rect 6053 33152 6069 33216
rect 6133 33152 6149 33216
rect 6213 33152 6229 33216
rect 6293 33152 6299 33216
rect 5983 33151 6299 33152
rect 9341 33216 9657 33217
rect 9341 33152 9347 33216
rect 9411 33152 9427 33216
rect 9491 33152 9507 33216
rect 9571 33152 9587 33216
rect 9651 33152 9657 33216
rect 9341 33151 9657 33152
rect 12699 33216 13015 33217
rect 12699 33152 12705 33216
rect 12769 33152 12785 33216
rect 12849 33152 12865 33216
rect 12929 33152 12945 33216
rect 13009 33152 13015 33216
rect 15540 33192 16000 33222
rect 12699 33151 13015 33152
rect 13353 33146 13419 33149
rect 13353 33144 14474 33146
rect 13353 33088 13358 33144
rect 13414 33088 14474 33144
rect 13353 33086 14474 33088
rect 13353 33083 13419 33086
rect 12341 33010 12407 33013
rect 12566 33010 12572 33012
rect 12341 33008 12572 33010
rect 12341 32952 12346 33008
rect 12402 32952 12572 33008
rect 12341 32950 12572 32952
rect 12341 32947 12407 32950
rect 12566 32948 12572 32950
rect 12636 32948 12642 33012
rect 13905 33010 13971 33013
rect 14414 33010 14474 33086
rect 15540 33010 16000 33040
rect 13905 33008 14290 33010
rect 13905 32952 13910 33008
rect 13966 32952 14290 33008
rect 13905 32950 14290 32952
rect 14414 32950 16000 33010
rect 13905 32947 13971 32950
rect 10174 32812 10180 32876
rect 10244 32874 10250 32876
rect 10961 32874 11027 32877
rect 10244 32872 11027 32874
rect 10244 32816 10966 32872
rect 11022 32816 11027 32872
rect 10244 32814 11027 32816
rect 10244 32812 10250 32814
rect 10961 32811 11027 32814
rect 11237 32874 11303 32877
rect 13445 32874 13511 32877
rect 11237 32872 13511 32874
rect 11237 32816 11242 32872
rect 11298 32816 13450 32872
rect 13506 32816 13511 32872
rect 11237 32814 13511 32816
rect 14230 32874 14290 32950
rect 15540 32920 16000 32950
rect 14230 32814 14842 32874
rect 11237 32811 11303 32814
rect 13445 32811 13511 32814
rect 14782 32738 14842 32814
rect 15540 32738 16000 32768
rect 14782 32678 16000 32738
rect 4304 32672 4620 32673
rect 4304 32608 4310 32672
rect 4374 32608 4390 32672
rect 4454 32608 4470 32672
rect 4534 32608 4550 32672
rect 4614 32608 4620 32672
rect 4304 32607 4620 32608
rect 7662 32672 7978 32673
rect 7662 32608 7668 32672
rect 7732 32608 7748 32672
rect 7812 32608 7828 32672
rect 7892 32608 7908 32672
rect 7972 32608 7978 32672
rect 7662 32607 7978 32608
rect 11020 32672 11336 32673
rect 11020 32608 11026 32672
rect 11090 32608 11106 32672
rect 11170 32608 11186 32672
rect 11250 32608 11266 32672
rect 11330 32608 11336 32672
rect 11020 32607 11336 32608
rect 14378 32672 14694 32673
rect 14378 32608 14384 32672
rect 14448 32608 14464 32672
rect 14528 32608 14544 32672
rect 14608 32608 14624 32672
rect 14688 32608 14694 32672
rect 15540 32648 16000 32678
rect 14378 32607 14694 32608
rect -300 32466 160 32496
rect 749 32466 815 32469
rect -300 32464 815 32466
rect -300 32408 754 32464
rect 810 32408 815 32464
rect -300 32406 815 32408
rect -300 32376 160 32406
rect 749 32403 815 32406
rect 12893 32466 12959 32469
rect 15540 32466 16000 32496
rect 12893 32464 16000 32466
rect 12893 32408 12898 32464
rect 12954 32408 16000 32464
rect 12893 32406 16000 32408
rect 12893 32403 12959 32406
rect 15540 32376 16000 32406
rect 12249 32330 12315 32333
rect 12249 32328 14106 32330
rect 12249 32272 12254 32328
rect 12310 32272 14106 32328
rect 12249 32270 14106 32272
rect 12249 32267 12315 32270
rect 14046 32194 14106 32270
rect 15540 32194 16000 32224
rect 14046 32134 16000 32194
rect 2625 32128 2941 32129
rect 2625 32064 2631 32128
rect 2695 32064 2711 32128
rect 2775 32064 2791 32128
rect 2855 32064 2871 32128
rect 2935 32064 2941 32128
rect 2625 32063 2941 32064
rect 5983 32128 6299 32129
rect 5983 32064 5989 32128
rect 6053 32064 6069 32128
rect 6133 32064 6149 32128
rect 6213 32064 6229 32128
rect 6293 32064 6299 32128
rect 5983 32063 6299 32064
rect 9341 32128 9657 32129
rect 9341 32064 9347 32128
rect 9411 32064 9427 32128
rect 9491 32064 9507 32128
rect 9571 32064 9587 32128
rect 9651 32064 9657 32128
rect 9341 32063 9657 32064
rect 12699 32128 13015 32129
rect 12699 32064 12705 32128
rect 12769 32064 12785 32128
rect 12849 32064 12865 32128
rect 12929 32064 12945 32128
rect 13009 32064 13015 32128
rect 15540 32104 16000 32134
rect 12699 32063 13015 32064
rect 14181 32060 14247 32061
rect 14181 32056 14228 32060
rect 14292 32058 14298 32060
rect 14181 32000 14186 32056
rect 14181 31996 14228 32000
rect 14292 31998 14338 32058
rect 14292 31996 14298 31998
rect 14181 31995 14247 31996
rect 13445 31920 13511 31925
rect 13445 31864 13450 31920
rect 13506 31864 13511 31920
rect 13445 31859 13511 31864
rect 13629 31922 13695 31925
rect 15540 31922 16000 31952
rect 13629 31920 16000 31922
rect 13629 31864 13634 31920
rect 13690 31864 16000 31920
rect 13629 31862 16000 31864
rect 13629 31859 13695 31862
rect 13448 31786 13508 31859
rect 15540 31832 16000 31862
rect 13448 31726 14842 31786
rect -300 31650 160 31680
rect 1393 31650 1459 31653
rect -300 31648 1459 31650
rect -300 31592 1398 31648
rect 1454 31592 1459 31648
rect -300 31590 1459 31592
rect 14782 31650 14842 31726
rect 15540 31650 16000 31680
rect 14782 31590 16000 31650
rect -300 31560 160 31590
rect 1393 31587 1459 31590
rect 4304 31584 4620 31585
rect 4304 31520 4310 31584
rect 4374 31520 4390 31584
rect 4454 31520 4470 31584
rect 4534 31520 4550 31584
rect 4614 31520 4620 31584
rect 4304 31519 4620 31520
rect 7662 31584 7978 31585
rect 7662 31520 7668 31584
rect 7732 31520 7748 31584
rect 7812 31520 7828 31584
rect 7892 31520 7908 31584
rect 7972 31520 7978 31584
rect 7662 31519 7978 31520
rect 11020 31584 11336 31585
rect 11020 31520 11026 31584
rect 11090 31520 11106 31584
rect 11170 31520 11186 31584
rect 11250 31520 11266 31584
rect 11330 31520 11336 31584
rect 11020 31519 11336 31520
rect 14378 31584 14694 31585
rect 14378 31520 14384 31584
rect 14448 31520 14464 31584
rect 14528 31520 14544 31584
rect 14608 31520 14624 31584
rect 14688 31520 14694 31584
rect 15540 31560 16000 31590
rect 14378 31519 14694 31520
rect 13261 31378 13327 31381
rect 13261 31376 13370 31378
rect 13261 31320 13266 31376
rect 13322 31320 13370 31376
rect 13261 31315 13370 31320
rect 14222 31316 14228 31380
rect 14292 31378 14298 31380
rect 15540 31378 16000 31408
rect 14292 31318 16000 31378
rect 14292 31316 14298 31318
rect 12985 31242 13051 31245
rect 12985 31240 13186 31242
rect 12985 31184 12990 31240
rect 13046 31184 13186 31240
rect 12985 31182 13186 31184
rect 12985 31179 13051 31182
rect 2625 31040 2941 31041
rect 2625 30976 2631 31040
rect 2695 30976 2711 31040
rect 2775 30976 2791 31040
rect 2855 30976 2871 31040
rect 2935 30976 2941 31040
rect 2625 30975 2941 30976
rect 5983 31040 6299 31041
rect 5983 30976 5989 31040
rect 6053 30976 6069 31040
rect 6133 30976 6149 31040
rect 6213 30976 6229 31040
rect 6293 30976 6299 31040
rect 5983 30975 6299 30976
rect 9341 31040 9657 31041
rect 9341 30976 9347 31040
rect 9411 30976 9427 31040
rect 9491 30976 9507 31040
rect 9571 30976 9587 31040
rect 9651 30976 9657 31040
rect 9341 30975 9657 30976
rect 12699 31040 13015 31041
rect 12699 30976 12705 31040
rect 12769 30976 12785 31040
rect 12849 30976 12865 31040
rect 12929 30976 12945 31040
rect 13009 30976 13015 31040
rect 12699 30975 13015 30976
rect 11789 30970 11855 30973
rect 12525 30970 12591 30973
rect 11789 30968 12591 30970
rect 11789 30912 11794 30968
rect 11850 30912 12530 30968
rect 12586 30912 12591 30968
rect 11789 30910 12591 30912
rect 13126 30970 13186 31182
rect 13310 31106 13370 31315
rect 15540 31288 16000 31318
rect 15540 31106 16000 31136
rect 13310 31046 16000 31106
rect 15540 31016 16000 31046
rect 13126 30910 15026 30970
rect 11789 30907 11855 30910
rect 12525 30907 12591 30910
rect -300 30834 160 30864
rect 749 30834 815 30837
rect -300 30832 815 30834
rect -300 30776 754 30832
rect 810 30776 815 30832
rect -300 30774 815 30776
rect -300 30744 160 30774
rect 749 30771 815 30774
rect 10174 30772 10180 30836
rect 10244 30834 10250 30836
rect 10317 30834 10383 30837
rect 10244 30832 10383 30834
rect 10244 30776 10322 30832
rect 10378 30776 10383 30832
rect 10244 30774 10383 30776
rect 10244 30772 10250 30774
rect 10317 30771 10383 30774
rect 12249 30834 12315 30837
rect 14966 30834 15026 30910
rect 15540 30834 16000 30864
rect 12249 30832 14842 30834
rect 12249 30776 12254 30832
rect 12310 30776 14842 30832
rect 12249 30774 14842 30776
rect 14966 30774 16000 30834
rect 12249 30771 12315 30774
rect 11789 30698 11855 30701
rect 13486 30698 13492 30700
rect 11789 30696 13492 30698
rect 11789 30640 11794 30696
rect 11850 30640 13492 30696
rect 11789 30638 13492 30640
rect 11789 30635 11855 30638
rect 13486 30636 13492 30638
rect 13556 30636 13562 30700
rect 14782 30562 14842 30774
rect 15540 30744 16000 30774
rect 15540 30562 16000 30592
rect 14782 30502 16000 30562
rect 4304 30496 4620 30497
rect 4304 30432 4310 30496
rect 4374 30432 4390 30496
rect 4454 30432 4470 30496
rect 4534 30432 4550 30496
rect 4614 30432 4620 30496
rect 4304 30431 4620 30432
rect 7662 30496 7978 30497
rect 7662 30432 7668 30496
rect 7732 30432 7748 30496
rect 7812 30432 7828 30496
rect 7892 30432 7908 30496
rect 7972 30432 7978 30496
rect 7662 30431 7978 30432
rect 11020 30496 11336 30497
rect 11020 30432 11026 30496
rect 11090 30432 11106 30496
rect 11170 30432 11186 30496
rect 11250 30432 11266 30496
rect 11330 30432 11336 30496
rect 11020 30431 11336 30432
rect 14378 30496 14694 30497
rect 14378 30432 14384 30496
rect 14448 30432 14464 30496
rect 14528 30432 14544 30496
rect 14608 30432 14624 30496
rect 14688 30432 14694 30496
rect 15540 30472 16000 30502
rect 14378 30431 14694 30432
rect 11881 30428 11947 30429
rect 11830 30364 11836 30428
rect 11900 30426 11947 30428
rect 11900 30424 11992 30426
rect 11942 30368 11992 30424
rect 11900 30366 11992 30368
rect 11900 30364 11947 30366
rect 11881 30363 11947 30364
rect 14089 30290 14155 30293
rect 14917 30290 14983 30293
rect 15540 30290 16000 30320
rect 14089 30288 14842 30290
rect 14089 30232 14094 30288
rect 14150 30232 14842 30288
rect 14089 30230 14842 30232
rect 14089 30227 14155 30230
rect -300 30018 160 30048
rect 749 30018 815 30021
rect -300 30016 815 30018
rect -300 29960 754 30016
rect 810 29960 815 30016
rect -300 29958 815 29960
rect 14782 30018 14842 30230
rect 14917 30288 16000 30290
rect 14917 30232 14922 30288
rect 14978 30232 16000 30288
rect 14917 30230 16000 30232
rect 14917 30227 14983 30230
rect 15540 30200 16000 30230
rect 15540 30018 16000 30048
rect 14782 29958 16000 30018
rect -300 29928 160 29958
rect 749 29955 815 29958
rect 2625 29952 2941 29953
rect 2625 29888 2631 29952
rect 2695 29888 2711 29952
rect 2775 29888 2791 29952
rect 2855 29888 2871 29952
rect 2935 29888 2941 29952
rect 2625 29887 2941 29888
rect 5983 29952 6299 29953
rect 5983 29888 5989 29952
rect 6053 29888 6069 29952
rect 6133 29888 6149 29952
rect 6213 29888 6229 29952
rect 6293 29888 6299 29952
rect 5983 29887 6299 29888
rect 9341 29952 9657 29953
rect 9341 29888 9347 29952
rect 9411 29888 9427 29952
rect 9491 29888 9507 29952
rect 9571 29888 9587 29952
rect 9651 29888 9657 29952
rect 9341 29887 9657 29888
rect 12699 29952 13015 29953
rect 12699 29888 12705 29952
rect 12769 29888 12785 29952
rect 12849 29888 12865 29952
rect 12929 29888 12945 29952
rect 13009 29888 13015 29952
rect 15540 29928 16000 29958
rect 12699 29887 13015 29888
rect 15009 29746 15075 29749
rect 15540 29746 16000 29776
rect 15009 29744 16000 29746
rect 15009 29688 15014 29744
rect 15070 29688 16000 29744
rect 15009 29686 16000 29688
rect 15009 29683 15075 29686
rect 15540 29656 16000 29686
rect 12525 29610 12591 29613
rect 12525 29608 14842 29610
rect 12525 29552 12530 29608
rect 12586 29552 14842 29608
rect 12525 29550 14842 29552
rect 12525 29547 12591 29550
rect 14782 29474 14842 29550
rect 15540 29474 16000 29504
rect 14782 29414 16000 29474
rect 4304 29408 4620 29409
rect 4304 29344 4310 29408
rect 4374 29344 4390 29408
rect 4454 29344 4470 29408
rect 4534 29344 4550 29408
rect 4614 29344 4620 29408
rect 4304 29343 4620 29344
rect 7662 29408 7978 29409
rect 7662 29344 7668 29408
rect 7732 29344 7748 29408
rect 7812 29344 7828 29408
rect 7892 29344 7908 29408
rect 7972 29344 7978 29408
rect 7662 29343 7978 29344
rect 11020 29408 11336 29409
rect 11020 29344 11026 29408
rect 11090 29344 11106 29408
rect 11170 29344 11186 29408
rect 11250 29344 11266 29408
rect 11330 29344 11336 29408
rect 11020 29343 11336 29344
rect 14378 29408 14694 29409
rect 14378 29344 14384 29408
rect 14448 29344 14464 29408
rect 14528 29344 14544 29408
rect 14608 29344 14624 29408
rect 14688 29344 14694 29408
rect 15540 29384 16000 29414
rect 14378 29343 14694 29344
rect -300 29202 160 29232
rect 749 29202 815 29205
rect -300 29200 815 29202
rect -300 29144 754 29200
rect 810 29144 815 29200
rect -300 29142 815 29144
rect -300 29112 160 29142
rect 749 29139 815 29142
rect 11053 29202 11119 29205
rect 11462 29202 11468 29204
rect 11053 29200 11468 29202
rect 11053 29144 11058 29200
rect 11114 29144 11468 29200
rect 11053 29142 11468 29144
rect 11053 29139 11119 29142
rect 11462 29140 11468 29142
rect 11532 29140 11538 29204
rect 11605 29202 11671 29205
rect 15540 29202 16000 29232
rect 11605 29200 16000 29202
rect 11605 29144 11610 29200
rect 11666 29144 16000 29200
rect 11605 29142 16000 29144
rect 11605 29139 11671 29142
rect 15540 29112 16000 29142
rect 1761 29066 1827 29069
rect 6913 29066 6979 29069
rect 9121 29068 9187 29069
rect 1761 29064 6979 29066
rect 1761 29008 1766 29064
rect 1822 29008 6918 29064
rect 6974 29008 6979 29064
rect 1761 29006 6979 29008
rect 1761 29003 1827 29006
rect 6913 29003 6979 29006
rect 9070 29004 9076 29068
rect 9140 29066 9187 29068
rect 9140 29064 9232 29066
rect 9182 29008 9232 29064
rect 9140 29006 9232 29008
rect 9140 29004 9187 29006
rect 9121 29003 9187 29004
rect 12249 28930 12315 28933
rect 12382 28930 12388 28932
rect 12249 28928 12388 28930
rect 12249 28872 12254 28928
rect 12310 28872 12388 28928
rect 12249 28870 12388 28872
rect 12249 28867 12315 28870
rect 12382 28868 12388 28870
rect 12452 28868 12458 28932
rect 15540 28930 16000 28960
rect 13908 28870 16000 28930
rect 2625 28864 2941 28865
rect 2625 28800 2631 28864
rect 2695 28800 2711 28864
rect 2775 28800 2791 28864
rect 2855 28800 2871 28864
rect 2935 28800 2941 28864
rect 2625 28799 2941 28800
rect 5983 28864 6299 28865
rect 5983 28800 5989 28864
rect 6053 28800 6069 28864
rect 6133 28800 6149 28864
rect 6213 28800 6229 28864
rect 6293 28800 6299 28864
rect 5983 28799 6299 28800
rect 9341 28864 9657 28865
rect 9341 28800 9347 28864
rect 9411 28800 9427 28864
rect 9491 28800 9507 28864
rect 9571 28800 9587 28864
rect 9651 28800 9657 28864
rect 9341 28799 9657 28800
rect 12699 28864 13015 28865
rect 12699 28800 12705 28864
rect 12769 28800 12785 28864
rect 12849 28800 12865 28864
rect 12929 28800 12945 28864
rect 13009 28800 13015 28864
rect 12699 28799 13015 28800
rect 11973 28796 12039 28797
rect 11973 28792 12020 28796
rect 12084 28794 12090 28796
rect 12249 28794 12315 28797
rect 12525 28794 12591 28797
rect 11973 28736 11978 28792
rect 11973 28732 12020 28736
rect 12084 28734 12130 28794
rect 12249 28792 12591 28794
rect 12249 28736 12254 28792
rect 12310 28736 12530 28792
rect 12586 28736 12591 28792
rect 12249 28734 12591 28736
rect 12084 28732 12090 28734
rect 11973 28731 12039 28732
rect 12249 28731 12315 28734
rect 12525 28731 12591 28734
rect 11421 28658 11487 28661
rect 13908 28658 13968 28870
rect 15540 28840 16000 28870
rect 11421 28656 13968 28658
rect 11421 28600 11426 28656
rect 11482 28600 13968 28656
rect 11421 28598 13968 28600
rect 15377 28658 15443 28661
rect 15540 28658 16000 28688
rect 15377 28656 16000 28658
rect 15377 28600 15382 28656
rect 15438 28600 16000 28656
rect 15377 28598 16000 28600
rect 11421 28595 11487 28598
rect 15377 28595 15443 28598
rect 15540 28568 16000 28598
rect 1577 28522 1643 28525
rect 6821 28522 6887 28525
rect 7189 28522 7255 28525
rect 1577 28520 7255 28522
rect 1577 28464 1582 28520
rect 1638 28464 6826 28520
rect 6882 28464 7194 28520
rect 7250 28464 7255 28520
rect 1577 28462 7255 28464
rect 1577 28459 1643 28462
rect 6821 28459 6887 28462
rect 7189 28459 7255 28462
rect 10685 28522 10751 28525
rect 12709 28522 12775 28525
rect 10685 28520 12775 28522
rect 10685 28464 10690 28520
rect 10746 28464 12714 28520
rect 12770 28464 12775 28520
rect 10685 28462 12775 28464
rect 10685 28459 10751 28462
rect 12709 28459 12775 28462
rect 13445 28522 13511 28525
rect 13445 28520 14842 28522
rect 13445 28464 13450 28520
rect 13506 28464 14842 28520
rect 13445 28462 14842 28464
rect 13445 28459 13511 28462
rect -300 28386 160 28416
rect 749 28386 815 28389
rect -300 28384 815 28386
rect -300 28328 754 28384
rect 810 28328 815 28384
rect -300 28326 815 28328
rect 14782 28386 14842 28462
rect 15540 28386 16000 28416
rect 14782 28326 16000 28386
rect -300 28296 160 28326
rect 749 28323 815 28326
rect 4304 28320 4620 28321
rect 4304 28256 4310 28320
rect 4374 28256 4390 28320
rect 4454 28256 4470 28320
rect 4534 28256 4550 28320
rect 4614 28256 4620 28320
rect 4304 28255 4620 28256
rect 7662 28320 7978 28321
rect 7662 28256 7668 28320
rect 7732 28256 7748 28320
rect 7812 28256 7828 28320
rect 7892 28256 7908 28320
rect 7972 28256 7978 28320
rect 7662 28255 7978 28256
rect 11020 28320 11336 28321
rect 11020 28256 11026 28320
rect 11090 28256 11106 28320
rect 11170 28256 11186 28320
rect 11250 28256 11266 28320
rect 11330 28256 11336 28320
rect 11020 28255 11336 28256
rect 14378 28320 14694 28321
rect 14378 28256 14384 28320
rect 14448 28256 14464 28320
rect 14528 28256 14544 28320
rect 14608 28256 14624 28320
rect 14688 28256 14694 28320
rect 15540 28296 16000 28326
rect 14378 28255 14694 28256
rect 14038 28250 14044 28252
rect 11470 28190 14044 28250
rect 8385 28114 8451 28117
rect 8518 28114 8524 28116
rect 8385 28112 8524 28114
rect 8385 28056 8390 28112
rect 8446 28056 8524 28112
rect 8385 28054 8524 28056
rect 8385 28051 8451 28054
rect 8518 28052 8524 28054
rect 8588 28052 8594 28116
rect 8937 28114 9003 28117
rect 10041 28114 10107 28117
rect 11470 28114 11530 28190
rect 14038 28188 14044 28190
rect 14108 28188 14114 28252
rect 8937 28112 11530 28114
rect 8937 28056 8942 28112
rect 8998 28056 10046 28112
rect 10102 28056 11530 28112
rect 8937 28054 11530 28056
rect 12341 28114 12407 28117
rect 14273 28114 14339 28117
rect 15540 28114 16000 28144
rect 12341 28112 12450 28114
rect 12341 28056 12346 28112
rect 12402 28056 12450 28112
rect 8937 28051 9003 28054
rect 10041 28051 10107 28054
rect 12341 28051 12450 28056
rect 14273 28112 16000 28114
rect 14273 28056 14278 28112
rect 14334 28056 16000 28112
rect 14273 28054 16000 28056
rect 14273 28051 14339 28054
rect 4061 27978 4127 27981
rect 9673 27978 9739 27981
rect 4061 27976 9739 27978
rect 4061 27920 4066 27976
rect 4122 27920 9678 27976
rect 9734 27920 9739 27976
rect 4061 27918 9739 27920
rect 12390 27978 12450 28051
rect 15540 28024 16000 28054
rect 12390 27918 14842 27978
rect 4061 27915 4127 27918
rect 9673 27915 9739 27918
rect 7925 27842 7991 27845
rect 8937 27842 9003 27845
rect 11973 27844 12039 27845
rect 11973 27842 12020 27844
rect 7925 27840 9003 27842
rect 7925 27784 7930 27840
rect 7986 27784 8942 27840
rect 8998 27784 9003 27840
rect 7925 27782 9003 27784
rect 11928 27840 12020 27842
rect 11928 27784 11978 27840
rect 11928 27782 12020 27784
rect 7925 27779 7991 27782
rect 8937 27779 9003 27782
rect 11973 27780 12020 27782
rect 12084 27780 12090 27844
rect 14782 27842 14842 27918
rect 15540 27842 16000 27872
rect 14782 27782 16000 27842
rect 11973 27779 12039 27780
rect 2625 27776 2941 27777
rect 2625 27712 2631 27776
rect 2695 27712 2711 27776
rect 2775 27712 2791 27776
rect 2855 27712 2871 27776
rect 2935 27712 2941 27776
rect 2625 27711 2941 27712
rect 5983 27776 6299 27777
rect 5983 27712 5989 27776
rect 6053 27712 6069 27776
rect 6133 27712 6149 27776
rect 6213 27712 6229 27776
rect 6293 27712 6299 27776
rect 5983 27711 6299 27712
rect 9341 27776 9657 27777
rect 9341 27712 9347 27776
rect 9411 27712 9427 27776
rect 9491 27712 9507 27776
rect 9571 27712 9587 27776
rect 9651 27712 9657 27776
rect 9341 27711 9657 27712
rect 12699 27776 13015 27777
rect 12699 27712 12705 27776
rect 12769 27712 12785 27776
rect 12849 27712 12865 27776
rect 12929 27712 12945 27776
rect 13009 27712 13015 27776
rect 15540 27752 16000 27782
rect 12699 27711 13015 27712
rect 8886 27644 8892 27708
rect 8956 27706 8962 27708
rect 9029 27706 9095 27709
rect 8956 27704 9095 27706
rect 8956 27648 9034 27704
rect 9090 27648 9095 27704
rect 8956 27646 9095 27648
rect 8956 27644 8962 27646
rect 9029 27643 9095 27646
rect 12014 27644 12020 27708
rect 12084 27706 12090 27708
rect 12341 27706 12407 27709
rect 12084 27704 12407 27706
rect 12084 27648 12346 27704
rect 12402 27648 12407 27704
rect 12084 27646 12407 27648
rect 12084 27644 12090 27646
rect 12341 27643 12407 27646
rect 13445 27706 13511 27709
rect 14222 27706 14228 27708
rect 13445 27704 14228 27706
rect 13445 27648 13450 27704
rect 13506 27648 14228 27704
rect 13445 27646 14228 27648
rect 13445 27643 13511 27646
rect 14222 27644 14228 27646
rect 14292 27644 14298 27708
rect -300 27570 160 27600
rect 1393 27570 1459 27573
rect -300 27568 1459 27570
rect -300 27512 1398 27568
rect 1454 27512 1459 27568
rect -300 27510 1459 27512
rect -300 27480 160 27510
rect 1393 27507 1459 27510
rect 10685 27570 10751 27573
rect 13905 27570 13971 27573
rect 10685 27568 13971 27570
rect 10685 27512 10690 27568
rect 10746 27512 13910 27568
rect 13966 27512 13971 27568
rect 10685 27510 13971 27512
rect 10685 27507 10751 27510
rect 13905 27507 13971 27510
rect 15377 27570 15443 27573
rect 15540 27570 16000 27600
rect 15377 27568 16000 27570
rect 15377 27512 15382 27568
rect 15438 27512 16000 27568
rect 15377 27510 16000 27512
rect 15377 27507 15443 27510
rect 15540 27480 16000 27510
rect 11881 27434 11947 27437
rect 12525 27434 12591 27437
rect 11881 27432 12591 27434
rect 11881 27376 11886 27432
rect 11942 27376 12530 27432
rect 12586 27376 12591 27432
rect 11881 27374 12591 27376
rect 11881 27371 11947 27374
rect 4304 27232 4620 27233
rect 4304 27168 4310 27232
rect 4374 27168 4390 27232
rect 4454 27168 4470 27232
rect 4534 27168 4550 27232
rect 4614 27168 4620 27232
rect 4304 27167 4620 27168
rect 7662 27232 7978 27233
rect 7662 27168 7668 27232
rect 7732 27168 7748 27232
rect 7812 27168 7828 27232
rect 7892 27168 7908 27232
rect 7972 27168 7978 27232
rect 7662 27167 7978 27168
rect 11020 27232 11336 27233
rect 11020 27168 11026 27232
rect 11090 27168 11106 27232
rect 11170 27168 11186 27232
rect 11250 27168 11266 27232
rect 11330 27168 11336 27232
rect 11020 27167 11336 27168
rect 12390 27162 12450 27374
rect 12525 27371 12591 27374
rect 15193 27298 15259 27301
rect 15540 27298 16000 27328
rect 15193 27296 16000 27298
rect 15193 27240 15198 27296
rect 15254 27240 16000 27296
rect 15193 27238 16000 27240
rect 15193 27235 15259 27238
rect 14378 27232 14694 27233
rect 14378 27168 14384 27232
rect 14448 27168 14464 27232
rect 14528 27168 14544 27232
rect 14608 27168 14624 27232
rect 14688 27168 14694 27232
rect 15540 27208 16000 27238
rect 14378 27167 14694 27168
rect 12566 27162 12572 27164
rect 12390 27102 12572 27162
rect 12566 27100 12572 27102
rect 12636 27100 12642 27164
rect 12065 27026 12131 27029
rect 15540 27026 16000 27056
rect 12065 27024 16000 27026
rect 12065 26968 12070 27024
rect 12126 26968 16000 27024
rect 12065 26966 16000 26968
rect 12065 26963 12131 26966
rect 15540 26936 16000 26966
rect 11605 26890 11671 26893
rect 11605 26888 13968 26890
rect 11605 26832 11610 26888
rect 11666 26832 13968 26888
rect 11605 26830 13968 26832
rect 11605 26827 11671 26830
rect -300 26754 160 26784
rect 749 26754 815 26757
rect -300 26752 815 26754
rect -300 26696 754 26752
rect 810 26696 815 26752
rect -300 26694 815 26696
rect -300 26664 160 26694
rect 749 26691 815 26694
rect 11605 26754 11671 26757
rect 11830 26754 11836 26756
rect 11605 26752 11836 26754
rect 11605 26696 11610 26752
rect 11666 26696 11836 26752
rect 11605 26694 11836 26696
rect 11605 26691 11671 26694
rect 11830 26692 11836 26694
rect 11900 26692 11906 26756
rect 13908 26754 13968 26830
rect 15540 26754 16000 26784
rect 13908 26694 16000 26754
rect 2625 26688 2941 26689
rect 2625 26624 2631 26688
rect 2695 26624 2711 26688
rect 2775 26624 2791 26688
rect 2855 26624 2871 26688
rect 2935 26624 2941 26688
rect 2625 26623 2941 26624
rect 5983 26688 6299 26689
rect 5983 26624 5989 26688
rect 6053 26624 6069 26688
rect 6133 26624 6149 26688
rect 6213 26624 6229 26688
rect 6293 26624 6299 26688
rect 5983 26623 6299 26624
rect 9341 26688 9657 26689
rect 9341 26624 9347 26688
rect 9411 26624 9427 26688
rect 9491 26624 9507 26688
rect 9571 26624 9587 26688
rect 9651 26624 9657 26688
rect 9341 26623 9657 26624
rect 12699 26688 13015 26689
rect 12699 26624 12705 26688
rect 12769 26624 12785 26688
rect 12849 26624 12865 26688
rect 12929 26624 12945 26688
rect 13009 26624 13015 26688
rect 15540 26664 16000 26694
rect 12699 26623 13015 26624
rect 9857 26482 9923 26485
rect 12893 26482 12959 26485
rect 9857 26480 12959 26482
rect 9857 26424 9862 26480
rect 9918 26424 12898 26480
rect 12954 26424 12959 26480
rect 9857 26422 12959 26424
rect 9857 26419 9923 26422
rect 12893 26419 12959 26422
rect 13997 26482 14063 26485
rect 15540 26482 16000 26512
rect 13997 26480 16000 26482
rect 13997 26424 14002 26480
rect 14058 26424 16000 26480
rect 13997 26422 16000 26424
rect 13997 26419 14063 26422
rect 15540 26392 16000 26422
rect 7281 26346 7347 26349
rect 7414 26346 7420 26348
rect 7281 26344 7420 26346
rect 7281 26288 7286 26344
rect 7342 26288 7420 26344
rect 7281 26286 7420 26288
rect 7281 26283 7347 26286
rect 7414 26284 7420 26286
rect 7484 26284 7490 26348
rect 1485 26210 1551 26213
rect 798 26208 1551 26210
rect 798 26152 1490 26208
rect 1546 26152 1551 26208
rect 798 26150 1551 26152
rect -300 25938 160 25968
rect 798 25938 858 26150
rect 1485 26147 1551 26150
rect 15009 26210 15075 26213
rect 15540 26210 16000 26240
rect 15009 26208 16000 26210
rect 15009 26152 15014 26208
rect 15070 26152 16000 26208
rect 15009 26150 16000 26152
rect 15009 26147 15075 26150
rect 4304 26144 4620 26145
rect 4304 26080 4310 26144
rect 4374 26080 4390 26144
rect 4454 26080 4470 26144
rect 4534 26080 4550 26144
rect 4614 26080 4620 26144
rect 4304 26079 4620 26080
rect 7662 26144 7978 26145
rect 7662 26080 7668 26144
rect 7732 26080 7748 26144
rect 7812 26080 7828 26144
rect 7892 26080 7908 26144
rect 7972 26080 7978 26144
rect 7662 26079 7978 26080
rect 11020 26144 11336 26145
rect 11020 26080 11026 26144
rect 11090 26080 11106 26144
rect 11170 26080 11186 26144
rect 11250 26080 11266 26144
rect 11330 26080 11336 26144
rect 11020 26079 11336 26080
rect 14378 26144 14694 26145
rect 14378 26080 14384 26144
rect 14448 26080 14464 26144
rect 14528 26080 14544 26144
rect 14608 26080 14624 26144
rect 14688 26080 14694 26144
rect 15540 26120 16000 26150
rect 14378 26079 14694 26080
rect -300 25878 858 25938
rect 10041 25938 10107 25941
rect 12433 25940 12499 25941
rect 10358 25938 10364 25940
rect 10041 25936 10364 25938
rect 10041 25880 10046 25936
rect 10102 25880 10364 25936
rect 10041 25878 10364 25880
rect -300 25848 160 25878
rect 10041 25875 10107 25878
rect 10358 25876 10364 25878
rect 10428 25876 10434 25940
rect 12382 25876 12388 25940
rect 12452 25938 12499 25940
rect 13721 25938 13787 25941
rect 15540 25938 16000 25968
rect 12452 25936 12544 25938
rect 12494 25880 12544 25936
rect 12452 25878 12544 25880
rect 13721 25936 16000 25938
rect 13721 25880 13726 25936
rect 13782 25880 16000 25936
rect 13721 25878 16000 25880
rect 12452 25876 12499 25878
rect 12433 25875 12499 25876
rect 13721 25875 13787 25878
rect 15540 25848 16000 25878
rect 13813 25666 13879 25669
rect 15540 25666 16000 25696
rect 13813 25664 16000 25666
rect 13813 25608 13818 25664
rect 13874 25608 16000 25664
rect 13813 25606 16000 25608
rect 13813 25603 13879 25606
rect 2625 25600 2941 25601
rect 2625 25536 2631 25600
rect 2695 25536 2711 25600
rect 2775 25536 2791 25600
rect 2855 25536 2871 25600
rect 2935 25536 2941 25600
rect 2625 25535 2941 25536
rect 5983 25600 6299 25601
rect 5983 25536 5989 25600
rect 6053 25536 6069 25600
rect 6133 25536 6149 25600
rect 6213 25536 6229 25600
rect 6293 25536 6299 25600
rect 5983 25535 6299 25536
rect 9341 25600 9657 25601
rect 9341 25536 9347 25600
rect 9411 25536 9427 25600
rect 9491 25536 9507 25600
rect 9571 25536 9587 25600
rect 9651 25536 9657 25600
rect 9341 25535 9657 25536
rect 12699 25600 13015 25601
rect 12699 25536 12705 25600
rect 12769 25536 12785 25600
rect 12849 25536 12865 25600
rect 12929 25536 12945 25600
rect 13009 25536 13015 25600
rect 15540 25576 16000 25606
rect 12699 25535 13015 25536
rect 10726 25332 10732 25396
rect 10796 25394 10802 25396
rect 11421 25394 11487 25397
rect 10796 25392 11487 25394
rect 10796 25336 11426 25392
rect 11482 25336 11487 25392
rect 10796 25334 11487 25336
rect 10796 25332 10802 25334
rect 11421 25331 11487 25334
rect 11881 25394 11947 25397
rect 15540 25394 16000 25424
rect 11881 25392 16000 25394
rect 11881 25336 11886 25392
rect 11942 25336 16000 25392
rect 11881 25334 16000 25336
rect 11881 25331 11947 25334
rect 15540 25304 16000 25334
rect 9673 25258 9739 25261
rect 10961 25258 11027 25261
rect 9673 25256 11027 25258
rect 9673 25200 9678 25256
rect 9734 25200 10966 25256
rect 11022 25200 11027 25256
rect 9673 25198 11027 25200
rect 9673 25195 9739 25198
rect 10961 25195 11027 25198
rect 14181 25258 14247 25261
rect 14181 25256 14842 25258
rect 14181 25200 14186 25256
rect 14242 25200 14842 25256
rect 14181 25198 14842 25200
rect 14181 25195 14247 25198
rect -300 25122 160 25152
rect 749 25122 815 25125
rect -300 25120 815 25122
rect -300 25064 754 25120
rect 810 25064 815 25120
rect -300 25062 815 25064
rect 14782 25122 14842 25198
rect 15540 25122 16000 25152
rect 14782 25062 16000 25122
rect -300 25032 160 25062
rect 749 25059 815 25062
rect 4304 25056 4620 25057
rect 4304 24992 4310 25056
rect 4374 24992 4390 25056
rect 4454 24992 4470 25056
rect 4534 24992 4550 25056
rect 4614 24992 4620 25056
rect 4304 24991 4620 24992
rect 7662 25056 7978 25057
rect 7662 24992 7668 25056
rect 7732 24992 7748 25056
rect 7812 24992 7828 25056
rect 7892 24992 7908 25056
rect 7972 24992 7978 25056
rect 7662 24991 7978 24992
rect 11020 25056 11336 25057
rect 11020 24992 11026 25056
rect 11090 24992 11106 25056
rect 11170 24992 11186 25056
rect 11250 24992 11266 25056
rect 11330 24992 11336 25056
rect 11020 24991 11336 24992
rect 14378 25056 14694 25057
rect 14378 24992 14384 25056
rect 14448 24992 14464 25056
rect 14528 24992 14544 25056
rect 14608 24992 14624 25056
rect 14688 24992 14694 25056
rect 15540 25032 16000 25062
rect 14378 24991 14694 24992
rect 12801 24986 12867 24989
rect 13670 24986 13676 24988
rect 12801 24984 13676 24986
rect 12801 24928 12806 24984
rect 12862 24928 13676 24984
rect 12801 24926 13676 24928
rect 12801 24923 12867 24926
rect 13670 24924 13676 24926
rect 13740 24924 13746 24988
rect 13997 24850 14063 24853
rect 15540 24850 16000 24880
rect 13997 24848 16000 24850
rect 13997 24792 14002 24848
rect 14058 24792 16000 24848
rect 13997 24790 16000 24792
rect 13997 24787 14063 24790
rect 15540 24760 16000 24790
rect 13445 24578 13511 24581
rect 15540 24578 16000 24608
rect 13445 24576 16000 24578
rect 13445 24520 13450 24576
rect 13506 24520 16000 24576
rect 13445 24518 16000 24520
rect 13445 24515 13511 24518
rect 2625 24512 2941 24513
rect 2625 24448 2631 24512
rect 2695 24448 2711 24512
rect 2775 24448 2791 24512
rect 2855 24448 2871 24512
rect 2935 24448 2941 24512
rect 2625 24447 2941 24448
rect 5983 24512 6299 24513
rect 5983 24448 5989 24512
rect 6053 24448 6069 24512
rect 6133 24448 6149 24512
rect 6213 24448 6229 24512
rect 6293 24448 6299 24512
rect 5983 24447 6299 24448
rect 9341 24512 9657 24513
rect 9341 24448 9347 24512
rect 9411 24448 9427 24512
rect 9491 24448 9507 24512
rect 9571 24448 9587 24512
rect 9651 24448 9657 24512
rect 9341 24447 9657 24448
rect 12699 24512 13015 24513
rect 12699 24448 12705 24512
rect 12769 24448 12785 24512
rect 12849 24448 12865 24512
rect 12929 24448 12945 24512
rect 13009 24448 13015 24512
rect 15540 24488 16000 24518
rect 12699 24447 13015 24448
rect -300 24306 160 24336
rect 749 24306 815 24309
rect -300 24304 815 24306
rect -300 24248 754 24304
rect 810 24248 815 24304
rect -300 24246 815 24248
rect -300 24216 160 24246
rect 749 24243 815 24246
rect 13997 24306 14063 24309
rect 15540 24306 16000 24336
rect 13997 24304 16000 24306
rect 13997 24248 14002 24304
rect 14058 24248 16000 24304
rect 13997 24246 16000 24248
rect 13997 24243 14063 24246
rect 15540 24216 16000 24246
rect 10041 24170 10107 24173
rect 10726 24170 10732 24172
rect 10041 24168 10732 24170
rect 10041 24112 10046 24168
rect 10102 24112 10732 24168
rect 10041 24110 10732 24112
rect 10041 24107 10107 24110
rect 10726 24108 10732 24110
rect 10796 24108 10802 24172
rect 11421 24170 11487 24173
rect 11421 24168 14842 24170
rect 11421 24112 11426 24168
rect 11482 24112 14842 24168
rect 11421 24110 14842 24112
rect 11421 24107 11487 24110
rect 14782 24034 14842 24110
rect 15540 24034 16000 24064
rect 14782 23974 16000 24034
rect 4304 23968 4620 23969
rect 4304 23904 4310 23968
rect 4374 23904 4390 23968
rect 4454 23904 4470 23968
rect 4534 23904 4550 23968
rect 4614 23904 4620 23968
rect 4304 23903 4620 23904
rect 7662 23968 7978 23969
rect 7662 23904 7668 23968
rect 7732 23904 7748 23968
rect 7812 23904 7828 23968
rect 7892 23904 7908 23968
rect 7972 23904 7978 23968
rect 7662 23903 7978 23904
rect 11020 23968 11336 23969
rect 11020 23904 11026 23968
rect 11090 23904 11106 23968
rect 11170 23904 11186 23968
rect 11250 23904 11266 23968
rect 11330 23904 11336 23968
rect 11020 23903 11336 23904
rect 14378 23968 14694 23969
rect 14378 23904 14384 23968
rect 14448 23904 14464 23968
rect 14528 23904 14544 23968
rect 14608 23904 14624 23968
rect 14688 23904 14694 23968
rect 15540 23944 16000 23974
rect 14378 23903 14694 23904
rect 14273 23762 14339 23765
rect 15540 23762 16000 23792
rect 14273 23760 16000 23762
rect 14273 23704 14278 23760
rect 14334 23704 16000 23760
rect 14273 23702 16000 23704
rect 14273 23699 14339 23702
rect 15540 23672 16000 23702
rect 7557 23626 7623 23629
rect 8150 23626 8156 23628
rect 7557 23624 8156 23626
rect 7557 23568 7562 23624
rect 7618 23568 8156 23624
rect 7557 23566 8156 23568
rect 7557 23563 7623 23566
rect 8150 23564 8156 23566
rect 8220 23564 8226 23628
rect 8518 23564 8524 23628
rect 8588 23626 8594 23628
rect 8661 23626 8727 23629
rect 8588 23624 8727 23626
rect 8588 23568 8666 23624
rect 8722 23568 8727 23624
rect 8588 23566 8727 23568
rect 8588 23564 8594 23566
rect 8661 23563 8727 23566
rect 9673 23626 9739 23629
rect 10225 23626 10291 23629
rect 12249 23626 12315 23629
rect 9673 23624 12315 23626
rect 9673 23568 9678 23624
rect 9734 23568 10230 23624
rect 10286 23568 12254 23624
rect 12310 23568 12315 23624
rect 9673 23566 12315 23568
rect 9673 23563 9739 23566
rect 10225 23563 10291 23566
rect 12249 23563 12315 23566
rect -300 23490 160 23520
rect 749 23490 815 23493
rect -300 23488 815 23490
rect -300 23432 754 23488
rect 810 23432 815 23488
rect -300 23430 815 23432
rect -300 23400 160 23430
rect 749 23427 815 23430
rect 13813 23490 13879 23493
rect 15540 23490 16000 23520
rect 13813 23488 16000 23490
rect 13813 23432 13818 23488
rect 13874 23432 16000 23488
rect 13813 23430 16000 23432
rect 13813 23427 13879 23430
rect 2625 23424 2941 23425
rect 2625 23360 2631 23424
rect 2695 23360 2711 23424
rect 2775 23360 2791 23424
rect 2855 23360 2871 23424
rect 2935 23360 2941 23424
rect 2625 23359 2941 23360
rect 5983 23424 6299 23425
rect 5983 23360 5989 23424
rect 6053 23360 6069 23424
rect 6133 23360 6149 23424
rect 6213 23360 6229 23424
rect 6293 23360 6299 23424
rect 5983 23359 6299 23360
rect 9341 23424 9657 23425
rect 9341 23360 9347 23424
rect 9411 23360 9427 23424
rect 9491 23360 9507 23424
rect 9571 23360 9587 23424
rect 9651 23360 9657 23424
rect 9341 23359 9657 23360
rect 12699 23424 13015 23425
rect 12699 23360 12705 23424
rect 12769 23360 12785 23424
rect 12849 23360 12865 23424
rect 12929 23360 12945 23424
rect 13009 23360 13015 23424
rect 15540 23400 16000 23430
rect 12699 23359 13015 23360
rect 11605 23218 11671 23221
rect 13169 23218 13235 23221
rect 11605 23216 13235 23218
rect 11605 23160 11610 23216
rect 11666 23160 13174 23216
rect 13230 23160 13235 23216
rect 11605 23158 13235 23160
rect 11605 23155 11671 23158
rect 13169 23155 13235 23158
rect 13721 23218 13787 23221
rect 15540 23218 16000 23248
rect 13721 23216 16000 23218
rect 13721 23160 13726 23216
rect 13782 23160 16000 23216
rect 13721 23158 16000 23160
rect 13721 23155 13787 23158
rect 15540 23128 16000 23158
rect 11605 23082 11671 23085
rect 14917 23082 14983 23085
rect 11605 23080 14983 23082
rect 11605 23024 11610 23080
rect 11666 23024 14922 23080
rect 14978 23024 14983 23080
rect 11605 23022 14983 23024
rect 11605 23019 11671 23022
rect 14917 23019 14983 23022
rect 14917 22946 14983 22949
rect 15540 22946 16000 22976
rect 14917 22944 16000 22946
rect 14917 22888 14922 22944
rect 14978 22888 16000 22944
rect 14917 22886 16000 22888
rect 14917 22883 14983 22886
rect 4304 22880 4620 22881
rect 4304 22816 4310 22880
rect 4374 22816 4390 22880
rect 4454 22816 4470 22880
rect 4534 22816 4550 22880
rect 4614 22816 4620 22880
rect 4304 22815 4620 22816
rect 7662 22880 7978 22881
rect 7662 22816 7668 22880
rect 7732 22816 7748 22880
rect 7812 22816 7828 22880
rect 7892 22816 7908 22880
rect 7972 22816 7978 22880
rect 7662 22815 7978 22816
rect 11020 22880 11336 22881
rect 11020 22816 11026 22880
rect 11090 22816 11106 22880
rect 11170 22816 11186 22880
rect 11250 22816 11266 22880
rect 11330 22816 11336 22880
rect 11020 22815 11336 22816
rect 14378 22880 14694 22881
rect 14378 22816 14384 22880
rect 14448 22816 14464 22880
rect 14528 22816 14544 22880
rect 14608 22816 14624 22880
rect 14688 22816 14694 22880
rect 15540 22856 16000 22886
rect 14378 22815 14694 22816
rect -300 22674 160 22704
rect 749 22674 815 22677
rect -300 22672 815 22674
rect -300 22616 754 22672
rect 810 22616 815 22672
rect -300 22614 815 22616
rect -300 22584 160 22614
rect 749 22611 815 22614
rect 14273 22674 14339 22677
rect 15540 22674 16000 22704
rect 14273 22672 16000 22674
rect 14273 22616 14278 22672
rect 14334 22616 16000 22672
rect 14273 22614 16000 22616
rect 14273 22611 14339 22614
rect 15540 22584 16000 22614
rect 8702 22476 8708 22540
rect 8772 22538 8778 22540
rect 9029 22538 9095 22541
rect 8772 22536 9095 22538
rect 8772 22480 9034 22536
rect 9090 22480 9095 22536
rect 8772 22478 9095 22480
rect 8772 22476 8778 22478
rect 9029 22475 9095 22478
rect 9765 22540 9831 22541
rect 9765 22536 9812 22540
rect 9876 22538 9882 22540
rect 10593 22538 10659 22541
rect 15326 22538 15332 22540
rect 9765 22480 9770 22536
rect 9765 22476 9812 22480
rect 9876 22478 9922 22538
rect 10593 22536 15332 22538
rect 10593 22480 10598 22536
rect 10654 22480 15332 22536
rect 10593 22478 15332 22480
rect 9876 22476 9882 22478
rect 9765 22475 9831 22476
rect 10593 22475 10659 22478
rect 15326 22476 15332 22478
rect 15396 22476 15402 22540
rect 15540 22402 16000 22432
rect 14598 22342 16000 22402
rect 2625 22336 2941 22337
rect 2625 22272 2631 22336
rect 2695 22272 2711 22336
rect 2775 22272 2791 22336
rect 2855 22272 2871 22336
rect 2935 22272 2941 22336
rect 2625 22271 2941 22272
rect 5983 22336 6299 22337
rect 5983 22272 5989 22336
rect 6053 22272 6069 22336
rect 6133 22272 6149 22336
rect 6213 22272 6229 22336
rect 6293 22272 6299 22336
rect 5983 22271 6299 22272
rect 9341 22336 9657 22337
rect 9341 22272 9347 22336
rect 9411 22272 9427 22336
rect 9491 22272 9507 22336
rect 9571 22272 9587 22336
rect 9651 22272 9657 22336
rect 9341 22271 9657 22272
rect 12699 22336 13015 22337
rect 12699 22272 12705 22336
rect 12769 22272 12785 22336
rect 12849 22272 12865 22336
rect 12929 22272 12945 22336
rect 13009 22272 13015 22336
rect 12699 22271 13015 22272
rect 13721 22266 13787 22269
rect 14598 22266 14658 22342
rect 15540 22312 16000 22342
rect 13721 22264 14658 22266
rect 13721 22208 13726 22264
rect 13782 22208 14658 22264
rect 13721 22206 14658 22208
rect 13721 22203 13787 22206
rect 13813 22130 13879 22133
rect 15540 22130 16000 22160
rect 13813 22128 16000 22130
rect 13813 22072 13818 22128
rect 13874 22072 16000 22128
rect 13813 22070 16000 22072
rect 13813 22067 13879 22070
rect 15540 22040 16000 22070
rect 9397 21994 9463 21997
rect 13905 21994 13971 21997
rect 9397 21992 13971 21994
rect 9397 21936 9402 21992
rect 9458 21936 13910 21992
rect 13966 21936 13971 21992
rect 9397 21934 13971 21936
rect 9397 21931 9463 21934
rect 13905 21931 13971 21934
rect -300 21858 160 21888
rect 749 21858 815 21861
rect -300 21856 815 21858
rect -300 21800 754 21856
rect 810 21800 815 21856
rect -300 21798 815 21800
rect -300 21768 160 21798
rect 749 21795 815 21798
rect 7373 21860 7439 21861
rect 7373 21856 7420 21860
rect 7484 21858 7490 21860
rect 15285 21858 15351 21861
rect 15540 21858 16000 21888
rect 7373 21800 7378 21856
rect 7373 21796 7420 21800
rect 7484 21798 7530 21858
rect 15285 21856 16000 21858
rect 15285 21800 15290 21856
rect 15346 21800 16000 21856
rect 15285 21798 16000 21800
rect 7484 21796 7490 21798
rect 7373 21795 7439 21796
rect 15285 21795 15351 21798
rect 4304 21792 4620 21793
rect 4304 21728 4310 21792
rect 4374 21728 4390 21792
rect 4454 21728 4470 21792
rect 4534 21728 4550 21792
rect 4614 21728 4620 21792
rect 4304 21727 4620 21728
rect 7662 21792 7978 21793
rect 7662 21728 7668 21792
rect 7732 21728 7748 21792
rect 7812 21728 7828 21792
rect 7892 21728 7908 21792
rect 7972 21728 7978 21792
rect 7662 21727 7978 21728
rect 11020 21792 11336 21793
rect 11020 21728 11026 21792
rect 11090 21728 11106 21792
rect 11170 21728 11186 21792
rect 11250 21728 11266 21792
rect 11330 21728 11336 21792
rect 11020 21727 11336 21728
rect 14378 21792 14694 21793
rect 14378 21728 14384 21792
rect 14448 21728 14464 21792
rect 14528 21728 14544 21792
rect 14608 21728 14624 21792
rect 14688 21728 14694 21792
rect 15540 21768 16000 21798
rect 14378 21727 14694 21728
rect 4521 21586 4587 21589
rect 8569 21586 8635 21589
rect 4521 21584 8635 21586
rect 4521 21528 4526 21584
rect 4582 21528 8574 21584
rect 8630 21528 8635 21584
rect 4521 21526 8635 21528
rect 4521 21523 4587 21526
rect 8569 21523 8635 21526
rect 13721 21586 13787 21589
rect 15540 21586 16000 21616
rect 13721 21584 16000 21586
rect 13721 21528 13726 21584
rect 13782 21528 16000 21584
rect 13721 21526 16000 21528
rect 13721 21523 13787 21526
rect 15540 21496 16000 21526
rect 13353 21450 13419 21453
rect 15193 21452 15259 21453
rect 15142 21450 15148 21452
rect 12390 21448 13419 21450
rect 12390 21392 13358 21448
rect 13414 21392 13419 21448
rect 12390 21390 13419 21392
rect 15102 21390 15148 21450
rect 15212 21448 15259 21452
rect 15254 21392 15259 21448
rect 10041 21312 10107 21317
rect 10041 21256 10046 21312
rect 10102 21256 10107 21312
rect 10041 21251 10107 21256
rect 12249 21314 12315 21317
rect 12390 21314 12450 21390
rect 13353 21387 13419 21390
rect 15142 21388 15148 21390
rect 15212 21388 15259 21392
rect 15193 21387 15259 21388
rect 12249 21312 12450 21314
rect 12249 21256 12254 21312
rect 12310 21256 12450 21312
rect 12249 21254 12450 21256
rect 13997 21314 14063 21317
rect 15540 21314 16000 21344
rect 13997 21312 16000 21314
rect 13997 21256 14002 21312
rect 14058 21256 16000 21312
rect 13997 21254 16000 21256
rect 12249 21251 12315 21254
rect 13997 21251 14063 21254
rect 2625 21248 2941 21249
rect 2625 21184 2631 21248
rect 2695 21184 2711 21248
rect 2775 21184 2791 21248
rect 2855 21184 2871 21248
rect 2935 21184 2941 21248
rect 2625 21183 2941 21184
rect 5983 21248 6299 21249
rect 5983 21184 5989 21248
rect 6053 21184 6069 21248
rect 6133 21184 6149 21248
rect 6213 21184 6229 21248
rect 6293 21184 6299 21248
rect 5983 21183 6299 21184
rect 9341 21248 9657 21249
rect 9341 21184 9347 21248
rect 9411 21184 9427 21248
rect 9491 21184 9507 21248
rect 9571 21184 9587 21248
rect 9651 21184 9657 21248
rect 9341 21183 9657 21184
rect -300 21042 160 21072
rect 749 21042 815 21045
rect -300 21040 815 21042
rect -300 20984 754 21040
rect 810 20984 815 21040
rect -300 20982 815 20984
rect 10044 21042 10104 21251
rect 12699 21248 13015 21249
rect 12699 21184 12705 21248
rect 12769 21184 12785 21248
rect 12849 21184 12865 21248
rect 12929 21184 12945 21248
rect 13009 21184 13015 21248
rect 15540 21224 16000 21254
rect 12699 21183 13015 21184
rect 13261 21042 13327 21045
rect 10044 21040 13327 21042
rect 10044 20984 13266 21040
rect 13322 20984 13327 21040
rect 10044 20982 13327 20984
rect -300 20952 160 20982
rect 749 20979 815 20982
rect 13261 20979 13327 20982
rect 14089 21042 14155 21045
rect 15540 21042 16000 21072
rect 14089 21040 16000 21042
rect 14089 20984 14094 21040
rect 14150 20984 16000 21040
rect 14089 20982 16000 20984
rect 14089 20979 14155 20982
rect 15540 20952 16000 20982
rect 9673 20906 9739 20909
rect 9806 20906 9812 20908
rect 9673 20904 9812 20906
rect 9673 20848 9678 20904
rect 9734 20848 9812 20904
rect 9673 20846 9812 20848
rect 9673 20843 9739 20846
rect 9806 20844 9812 20846
rect 9876 20844 9882 20908
rect 6913 20770 6979 20773
rect 13813 20772 13879 20773
rect 7046 20770 7052 20772
rect 6913 20768 7052 20770
rect 6913 20712 6918 20768
rect 6974 20712 7052 20768
rect 6913 20710 7052 20712
rect 6913 20707 6979 20710
rect 7046 20708 7052 20710
rect 7116 20708 7122 20772
rect 13813 20768 13860 20772
rect 13924 20770 13930 20772
rect 15009 20770 15075 20773
rect 15540 20770 16000 20800
rect 13813 20712 13818 20768
rect 13813 20708 13860 20712
rect 13924 20710 13970 20770
rect 15009 20768 16000 20770
rect 15009 20712 15014 20768
rect 15070 20712 16000 20768
rect 15009 20710 16000 20712
rect 13924 20708 13930 20710
rect 13813 20707 13879 20708
rect 15009 20707 15075 20710
rect 4304 20704 4620 20705
rect 4304 20640 4310 20704
rect 4374 20640 4390 20704
rect 4454 20640 4470 20704
rect 4534 20640 4550 20704
rect 4614 20640 4620 20704
rect 4304 20639 4620 20640
rect 7662 20704 7978 20705
rect 7662 20640 7668 20704
rect 7732 20640 7748 20704
rect 7812 20640 7828 20704
rect 7892 20640 7908 20704
rect 7972 20640 7978 20704
rect 7662 20639 7978 20640
rect 11020 20704 11336 20705
rect 11020 20640 11026 20704
rect 11090 20640 11106 20704
rect 11170 20640 11186 20704
rect 11250 20640 11266 20704
rect 11330 20640 11336 20704
rect 11020 20639 11336 20640
rect 14378 20704 14694 20705
rect 14378 20640 14384 20704
rect 14448 20640 14464 20704
rect 14528 20640 14544 20704
rect 14608 20640 14624 20704
rect 14688 20640 14694 20704
rect 15540 20680 16000 20710
rect 14378 20639 14694 20640
rect 12157 20636 12223 20637
rect 12157 20632 12204 20636
rect 12268 20634 12274 20636
rect 12709 20634 12775 20637
rect 12157 20576 12162 20632
rect 12157 20572 12204 20576
rect 12268 20574 12314 20634
rect 12709 20632 14106 20634
rect 12709 20576 12714 20632
rect 12770 20576 14106 20632
rect 12709 20574 14106 20576
rect 12268 20572 12274 20574
rect 12157 20571 12223 20572
rect 12709 20571 12775 20574
rect 1526 20436 1532 20500
rect 1596 20498 1602 20500
rect 4153 20498 4219 20501
rect 1596 20496 4219 20498
rect 1596 20440 4158 20496
rect 4214 20440 4219 20496
rect 1596 20438 4219 20440
rect 1596 20436 1602 20438
rect 4153 20435 4219 20438
rect 6913 20498 6979 20501
rect 7925 20498 7991 20501
rect 6913 20496 7991 20498
rect 6913 20440 6918 20496
rect 6974 20440 7930 20496
rect 7986 20440 7991 20496
rect 6913 20438 7991 20440
rect 14046 20498 14106 20574
rect 15540 20498 16000 20528
rect 14046 20438 16000 20498
rect 6913 20435 6979 20438
rect 7925 20435 7991 20438
rect 15540 20408 16000 20438
rect 5441 20362 5507 20365
rect 11605 20362 11671 20365
rect 5441 20360 11671 20362
rect 5441 20304 5446 20360
rect 5502 20304 11610 20360
rect 11666 20304 11671 20360
rect 5441 20302 11671 20304
rect 5441 20299 5507 20302
rect 11605 20299 11671 20302
rect -300 20226 160 20256
rect 749 20226 815 20229
rect -300 20224 815 20226
rect -300 20168 754 20224
rect 810 20168 815 20224
rect -300 20166 815 20168
rect -300 20136 160 20166
rect 749 20163 815 20166
rect 14089 20226 14155 20229
rect 15540 20226 16000 20256
rect 14089 20224 16000 20226
rect 14089 20168 14094 20224
rect 14150 20168 16000 20224
rect 14089 20166 16000 20168
rect 14089 20163 14155 20166
rect 2625 20160 2941 20161
rect 2625 20096 2631 20160
rect 2695 20096 2711 20160
rect 2775 20096 2791 20160
rect 2855 20096 2871 20160
rect 2935 20096 2941 20160
rect 2625 20095 2941 20096
rect 5983 20160 6299 20161
rect 5983 20096 5989 20160
rect 6053 20096 6069 20160
rect 6133 20096 6149 20160
rect 6213 20096 6229 20160
rect 6293 20096 6299 20160
rect 5983 20095 6299 20096
rect 9341 20160 9657 20161
rect 9341 20096 9347 20160
rect 9411 20096 9427 20160
rect 9491 20096 9507 20160
rect 9571 20096 9587 20160
rect 9651 20096 9657 20160
rect 9341 20095 9657 20096
rect 12699 20160 13015 20161
rect 12699 20096 12705 20160
rect 12769 20096 12785 20160
rect 12849 20096 12865 20160
rect 12929 20096 12945 20160
rect 13009 20096 13015 20160
rect 15540 20136 16000 20166
rect 12699 20095 13015 20096
rect 7005 19954 7071 19957
rect 8937 19954 9003 19957
rect 7005 19952 9003 19954
rect 7005 19896 7010 19952
rect 7066 19896 8942 19952
rect 8998 19896 9003 19952
rect 7005 19894 9003 19896
rect 7005 19891 7071 19894
rect 8937 19891 9003 19894
rect 12617 19954 12683 19957
rect 15540 19954 16000 19984
rect 12617 19952 16000 19954
rect 12617 19896 12622 19952
rect 12678 19896 16000 19952
rect 12617 19894 16000 19896
rect 12617 19891 12683 19894
rect 15540 19864 16000 19894
rect 12157 19818 12223 19821
rect 12157 19816 14842 19818
rect 12157 19760 12162 19816
rect 12218 19760 14842 19816
rect 12157 19758 14842 19760
rect 12157 19755 12223 19758
rect 14782 19682 14842 19758
rect 15540 19682 16000 19712
rect 14782 19622 16000 19682
rect 4304 19616 4620 19617
rect 4304 19552 4310 19616
rect 4374 19552 4390 19616
rect 4454 19552 4470 19616
rect 4534 19552 4550 19616
rect 4614 19552 4620 19616
rect 4304 19551 4620 19552
rect 7662 19616 7978 19617
rect 7662 19552 7668 19616
rect 7732 19552 7748 19616
rect 7812 19552 7828 19616
rect 7892 19552 7908 19616
rect 7972 19552 7978 19616
rect 7662 19551 7978 19552
rect 11020 19616 11336 19617
rect 11020 19552 11026 19616
rect 11090 19552 11106 19616
rect 11170 19552 11186 19616
rect 11250 19552 11266 19616
rect 11330 19552 11336 19616
rect 11020 19551 11336 19552
rect 14378 19616 14694 19617
rect 14378 19552 14384 19616
rect 14448 19552 14464 19616
rect 14528 19552 14544 19616
rect 14608 19552 14624 19616
rect 14688 19552 14694 19616
rect 15540 19592 16000 19622
rect 14378 19551 14694 19552
rect -300 19410 160 19440
rect 749 19410 815 19413
rect -300 19408 815 19410
rect -300 19352 754 19408
rect 810 19352 815 19408
rect -300 19350 815 19352
rect -300 19320 160 19350
rect 749 19347 815 19350
rect 8293 19410 8359 19413
rect 9070 19410 9076 19412
rect 8293 19408 9076 19410
rect 8293 19352 8298 19408
rect 8354 19352 9076 19408
rect 8293 19350 9076 19352
rect 8293 19347 8359 19350
rect 9070 19348 9076 19350
rect 9140 19348 9146 19412
rect 9765 19410 9831 19413
rect 9990 19410 9996 19412
rect 9765 19408 9996 19410
rect 9765 19352 9770 19408
rect 9826 19352 9996 19408
rect 9765 19350 9996 19352
rect 9765 19347 9831 19350
rect 9990 19348 9996 19350
rect 10060 19348 10066 19412
rect 11237 19410 11303 19413
rect 15540 19410 16000 19440
rect 11237 19408 16000 19410
rect 11237 19352 11242 19408
rect 11298 19352 16000 19408
rect 11237 19350 16000 19352
rect 11237 19347 11303 19350
rect 15540 19320 16000 19350
rect 7005 19274 7071 19277
rect 7465 19274 7531 19277
rect 7005 19272 7531 19274
rect 7005 19216 7010 19272
rect 7066 19216 7470 19272
rect 7526 19216 7531 19272
rect 7005 19214 7531 19216
rect 7005 19211 7071 19214
rect 7465 19211 7531 19214
rect 8886 19212 8892 19276
rect 8956 19274 8962 19276
rect 9397 19274 9463 19277
rect 8956 19272 9463 19274
rect 8956 19216 9402 19272
rect 9458 19216 9463 19272
rect 8956 19214 9463 19216
rect 8956 19212 8962 19214
rect 9397 19211 9463 19214
rect 13670 19212 13676 19276
rect 13740 19274 13746 19276
rect 14365 19274 14431 19277
rect 13740 19272 14431 19274
rect 13740 19216 14370 19272
rect 14426 19216 14431 19272
rect 13740 19214 14431 19216
rect 13740 19212 13746 19214
rect 14365 19211 14431 19214
rect 6821 19138 6887 19141
rect 8845 19138 8911 19141
rect 6821 19136 8911 19138
rect 6821 19080 6826 19136
rect 6882 19080 8850 19136
rect 8906 19080 8911 19136
rect 6821 19078 8911 19080
rect 6821 19075 6887 19078
rect 8845 19075 8911 19078
rect 13997 19138 14063 19141
rect 15540 19138 16000 19168
rect 13997 19136 16000 19138
rect 13997 19080 14002 19136
rect 14058 19080 16000 19136
rect 13997 19078 16000 19080
rect 13997 19075 14063 19078
rect 2625 19072 2941 19073
rect 2625 19008 2631 19072
rect 2695 19008 2711 19072
rect 2775 19008 2791 19072
rect 2855 19008 2871 19072
rect 2935 19008 2941 19072
rect 2625 19007 2941 19008
rect 5983 19072 6299 19073
rect 5983 19008 5989 19072
rect 6053 19008 6069 19072
rect 6133 19008 6149 19072
rect 6213 19008 6229 19072
rect 6293 19008 6299 19072
rect 5983 19007 6299 19008
rect 9341 19072 9657 19073
rect 9341 19008 9347 19072
rect 9411 19008 9427 19072
rect 9491 19008 9507 19072
rect 9571 19008 9587 19072
rect 9651 19008 9657 19072
rect 9341 19007 9657 19008
rect 12699 19072 13015 19073
rect 12699 19008 12705 19072
rect 12769 19008 12785 19072
rect 12849 19008 12865 19072
rect 12929 19008 12945 19072
rect 13009 19008 13015 19072
rect 15540 19048 16000 19078
rect 12699 19007 13015 19008
rect 4981 18866 5047 18869
rect 7414 18866 7420 18868
rect 4981 18864 7420 18866
rect 4981 18808 4986 18864
rect 5042 18808 7420 18864
rect 4981 18806 7420 18808
rect 4981 18803 5047 18806
rect 7414 18804 7420 18806
rect 7484 18866 7490 18868
rect 10685 18866 10751 18869
rect 7484 18864 10751 18866
rect 7484 18808 10690 18864
rect 10746 18808 10751 18864
rect 7484 18806 10751 18808
rect 7484 18804 7490 18806
rect 10685 18803 10751 18806
rect 12065 18866 12131 18869
rect 15540 18866 16000 18896
rect 12065 18864 16000 18866
rect 12065 18808 12070 18864
rect 12126 18808 16000 18864
rect 12065 18806 16000 18808
rect 12065 18803 12131 18806
rect 15540 18776 16000 18806
rect 3693 18730 3759 18733
rect 7230 18730 7236 18732
rect 3693 18728 7236 18730
rect 3693 18672 3698 18728
rect 3754 18672 7236 18728
rect 3693 18670 7236 18672
rect 3693 18667 3759 18670
rect 7230 18668 7236 18670
rect 7300 18730 7306 18732
rect 7557 18730 7623 18733
rect 8201 18732 8267 18733
rect 8150 18730 8156 18732
rect 7300 18728 7623 18730
rect 7300 18672 7562 18728
rect 7618 18672 7623 18728
rect 7300 18670 7623 18672
rect 8110 18670 8156 18730
rect 8220 18728 8267 18732
rect 8262 18672 8267 18728
rect 7300 18668 7306 18670
rect 7557 18667 7623 18670
rect 8150 18668 8156 18670
rect 8220 18668 8267 18672
rect 8201 18667 8267 18668
rect -300 18594 160 18624
rect 749 18594 815 18597
rect -300 18592 815 18594
rect -300 18536 754 18592
rect 810 18536 815 18592
rect -300 18534 815 18536
rect -300 18504 160 18534
rect 749 18531 815 18534
rect 15009 18594 15075 18597
rect 15540 18594 16000 18624
rect 15009 18592 16000 18594
rect 15009 18536 15014 18592
rect 15070 18536 16000 18592
rect 15009 18534 16000 18536
rect 15009 18531 15075 18534
rect 4304 18528 4620 18529
rect 4304 18464 4310 18528
rect 4374 18464 4390 18528
rect 4454 18464 4470 18528
rect 4534 18464 4550 18528
rect 4614 18464 4620 18528
rect 4304 18463 4620 18464
rect 7662 18528 7978 18529
rect 7662 18464 7668 18528
rect 7732 18464 7748 18528
rect 7812 18464 7828 18528
rect 7892 18464 7908 18528
rect 7972 18464 7978 18528
rect 7662 18463 7978 18464
rect 11020 18528 11336 18529
rect 11020 18464 11026 18528
rect 11090 18464 11106 18528
rect 11170 18464 11186 18528
rect 11250 18464 11266 18528
rect 11330 18464 11336 18528
rect 11020 18463 11336 18464
rect 14378 18528 14694 18529
rect 14378 18464 14384 18528
rect 14448 18464 14464 18528
rect 14528 18464 14544 18528
rect 14608 18464 14624 18528
rect 14688 18464 14694 18528
rect 15540 18504 16000 18534
rect 14378 18463 14694 18464
rect 13302 18396 13308 18460
rect 13372 18458 13378 18460
rect 13445 18458 13511 18461
rect 13372 18456 13511 18458
rect 13372 18400 13450 18456
rect 13506 18400 13511 18456
rect 13372 18398 13511 18400
rect 13372 18396 13378 18398
rect 13445 18395 13511 18398
rect 3601 18322 3667 18325
rect 9070 18322 9076 18324
rect 3601 18320 9076 18322
rect 3601 18264 3606 18320
rect 3662 18264 9076 18320
rect 3601 18262 9076 18264
rect 3601 18259 3667 18262
rect 9070 18260 9076 18262
rect 9140 18260 9146 18324
rect 9857 18322 9923 18325
rect 12341 18324 12407 18325
rect 13445 18324 13511 18325
rect 11462 18322 11468 18324
rect 9857 18320 11468 18322
rect 9857 18264 9862 18320
rect 9918 18264 11468 18320
rect 9857 18262 11468 18264
rect 9857 18259 9923 18262
rect 11462 18260 11468 18262
rect 11532 18260 11538 18324
rect 12341 18322 12388 18324
rect 12296 18320 12388 18322
rect 12296 18264 12346 18320
rect 12296 18262 12388 18264
rect 12341 18260 12388 18262
rect 12452 18260 12458 18324
rect 13445 18322 13492 18324
rect 13400 18320 13492 18322
rect 13400 18264 13450 18320
rect 13400 18262 13492 18264
rect 13445 18260 13492 18262
rect 13556 18260 13562 18324
rect 15285 18322 15351 18325
rect 15540 18322 16000 18352
rect 15285 18320 16000 18322
rect 15285 18264 15290 18320
rect 15346 18264 16000 18320
rect 15285 18262 16000 18264
rect 12341 18259 12407 18260
rect 13445 18259 13511 18260
rect 15285 18259 15351 18262
rect 15540 18232 16000 18262
rect 8753 18186 8819 18189
rect 9857 18186 9923 18189
rect 8753 18184 9923 18186
rect 8753 18128 8758 18184
rect 8814 18128 9862 18184
rect 9918 18128 9923 18184
rect 8753 18126 9923 18128
rect 8753 18123 8819 18126
rect 9857 18123 9923 18126
rect 12341 18186 12407 18189
rect 12341 18184 14106 18186
rect 12341 18128 12346 18184
rect 12402 18128 14106 18184
rect 12341 18126 14106 18128
rect 12341 18123 12407 18126
rect 8017 18050 8083 18053
rect 8477 18050 8543 18053
rect 8017 18048 8543 18050
rect 8017 17992 8022 18048
rect 8078 17992 8482 18048
rect 8538 17992 8543 18048
rect 8017 17990 8543 17992
rect 14046 18050 14106 18126
rect 15540 18050 16000 18080
rect 14046 17990 16000 18050
rect 8017 17987 8083 17990
rect 8477 17987 8543 17990
rect 2625 17984 2941 17985
rect 2625 17920 2631 17984
rect 2695 17920 2711 17984
rect 2775 17920 2791 17984
rect 2855 17920 2871 17984
rect 2935 17920 2941 17984
rect 2625 17919 2941 17920
rect 5983 17984 6299 17985
rect 5983 17920 5989 17984
rect 6053 17920 6069 17984
rect 6133 17920 6149 17984
rect 6213 17920 6229 17984
rect 6293 17920 6299 17984
rect 5983 17919 6299 17920
rect 9341 17984 9657 17985
rect 9341 17920 9347 17984
rect 9411 17920 9427 17984
rect 9491 17920 9507 17984
rect 9571 17920 9587 17984
rect 9651 17920 9657 17984
rect 9341 17919 9657 17920
rect 12699 17984 13015 17985
rect 12699 17920 12705 17984
rect 12769 17920 12785 17984
rect 12849 17920 12865 17984
rect 12929 17920 12945 17984
rect 13009 17920 13015 17984
rect 15540 17960 16000 17990
rect 12699 17919 13015 17920
rect 1485 17914 1551 17917
rect 798 17912 1551 17914
rect 798 17856 1490 17912
rect 1546 17856 1551 17912
rect 798 17854 1551 17856
rect -300 17778 160 17808
rect 798 17778 858 17854
rect 1485 17851 1551 17854
rect 9765 17916 9831 17917
rect 9765 17912 9812 17916
rect 9876 17914 9882 17916
rect 9765 17856 9770 17912
rect 9765 17852 9812 17856
rect 9876 17854 9922 17914
rect 9876 17852 9882 17854
rect 9765 17851 9831 17852
rect -300 17718 858 17778
rect 10501 17778 10567 17781
rect 15540 17778 16000 17808
rect 10501 17776 16000 17778
rect 10501 17720 10506 17776
rect 10562 17720 16000 17776
rect 10501 17718 16000 17720
rect -300 17688 160 17718
rect 10501 17715 10567 17718
rect 15540 17688 16000 17718
rect 6913 17642 6979 17645
rect 7046 17642 7052 17644
rect 6913 17640 7052 17642
rect 6913 17584 6918 17640
rect 6974 17584 7052 17640
rect 6913 17582 7052 17584
rect 6913 17579 6979 17582
rect 7046 17580 7052 17582
rect 7116 17580 7122 17644
rect 10869 17642 10935 17645
rect 10734 17640 10935 17642
rect 10734 17584 10874 17640
rect 10930 17584 10935 17640
rect 10734 17582 10935 17584
rect 4304 17440 4620 17441
rect 4304 17376 4310 17440
rect 4374 17376 4390 17440
rect 4454 17376 4470 17440
rect 4534 17376 4550 17440
rect 4614 17376 4620 17440
rect 4304 17375 4620 17376
rect 7662 17440 7978 17441
rect 7662 17376 7668 17440
rect 7732 17376 7748 17440
rect 7812 17376 7828 17440
rect 7892 17376 7908 17440
rect 7972 17376 7978 17440
rect 7662 17375 7978 17376
rect 10734 17373 10794 17582
rect 10869 17579 10935 17582
rect 11697 17642 11763 17645
rect 12065 17642 12131 17645
rect 11697 17640 12131 17642
rect 11697 17584 11702 17640
rect 11758 17584 12070 17640
rect 12126 17584 12131 17640
rect 11697 17582 12131 17584
rect 11697 17579 11763 17582
rect 12065 17579 12131 17582
rect 14038 17580 14044 17644
rect 14108 17580 14114 17644
rect 12985 17506 13051 17509
rect 14046 17506 14106 17580
rect 15540 17506 16000 17536
rect 12985 17504 14106 17506
rect 12985 17448 12990 17504
rect 13046 17448 14106 17504
rect 12985 17446 14106 17448
rect 14782 17446 16000 17506
rect 12985 17443 13051 17446
rect 11020 17440 11336 17441
rect 11020 17376 11026 17440
rect 11090 17376 11106 17440
rect 11170 17376 11186 17440
rect 11250 17376 11266 17440
rect 11330 17376 11336 17440
rect 11020 17375 11336 17376
rect 14378 17440 14694 17441
rect 14378 17376 14384 17440
rect 14448 17376 14464 17440
rect 14528 17376 14544 17440
rect 14608 17376 14624 17440
rect 14688 17376 14694 17440
rect 14378 17375 14694 17376
rect 10734 17368 10843 17373
rect 10734 17312 10782 17368
rect 10838 17312 10843 17368
rect 10734 17310 10843 17312
rect 10777 17307 10843 17310
rect 13537 17370 13603 17373
rect 14222 17370 14228 17372
rect 13537 17368 14228 17370
rect 13537 17312 13542 17368
rect 13598 17312 14228 17368
rect 13537 17310 14228 17312
rect 13537 17307 13603 17310
rect 14222 17308 14228 17310
rect 14292 17308 14298 17372
rect 11697 17234 11763 17237
rect 2730 17232 11763 17234
rect 2730 17176 11702 17232
rect 11758 17176 11763 17232
rect 2730 17174 11763 17176
rect 2405 17098 2471 17101
rect 2730 17098 2790 17174
rect 11697 17171 11763 17174
rect 11881 17234 11947 17237
rect 14782 17234 14842 17446
rect 15540 17416 16000 17446
rect 11881 17232 14842 17234
rect 11881 17176 11886 17232
rect 11942 17176 14842 17232
rect 11881 17174 14842 17176
rect 15009 17234 15075 17237
rect 15540 17234 16000 17264
rect 15009 17232 16000 17234
rect 15009 17176 15014 17232
rect 15070 17176 16000 17232
rect 15009 17174 16000 17176
rect 11881 17171 11947 17174
rect 15009 17171 15075 17174
rect 15540 17144 16000 17174
rect 2405 17096 2790 17098
rect 2405 17040 2410 17096
rect 2466 17040 2790 17096
rect 2405 17038 2790 17040
rect 3969 17098 4035 17101
rect 10358 17098 10364 17100
rect 3969 17096 10364 17098
rect 3969 17040 3974 17096
rect 4030 17040 10364 17096
rect 3969 17038 10364 17040
rect 2405 17035 2471 17038
rect 3969 17035 4035 17038
rect 10358 17036 10364 17038
rect 10428 17036 10434 17100
rect 11145 17098 11211 17101
rect 11145 17096 14106 17098
rect 11145 17040 11150 17096
rect 11206 17040 14106 17096
rect 11145 17038 14106 17040
rect 11145 17035 11211 17038
rect -300 16962 160 16992
rect 749 16962 815 16965
rect -300 16960 815 16962
rect -300 16904 754 16960
rect 810 16904 815 16960
rect -300 16902 815 16904
rect 14046 16962 14106 17038
rect 15540 16962 16000 16992
rect 14046 16902 16000 16962
rect -300 16872 160 16902
rect 749 16899 815 16902
rect 2625 16896 2941 16897
rect 2625 16832 2631 16896
rect 2695 16832 2711 16896
rect 2775 16832 2791 16896
rect 2855 16832 2871 16896
rect 2935 16832 2941 16896
rect 2625 16831 2941 16832
rect 5983 16896 6299 16897
rect 5983 16832 5989 16896
rect 6053 16832 6069 16896
rect 6133 16832 6149 16896
rect 6213 16832 6229 16896
rect 6293 16832 6299 16896
rect 5983 16831 6299 16832
rect 9341 16896 9657 16897
rect 9341 16832 9347 16896
rect 9411 16832 9427 16896
rect 9491 16832 9507 16896
rect 9571 16832 9587 16896
rect 9651 16832 9657 16896
rect 9341 16831 9657 16832
rect 12699 16896 13015 16897
rect 12699 16832 12705 16896
rect 12769 16832 12785 16896
rect 12849 16832 12865 16896
rect 12929 16832 12945 16896
rect 13009 16832 13015 16896
rect 15540 16872 16000 16902
rect 12699 16831 13015 16832
rect 15009 16826 15075 16829
rect 13862 16824 15075 16826
rect 13862 16768 15014 16824
rect 15070 16768 15075 16824
rect 13862 16766 15075 16768
rect 11145 16690 11211 16693
rect 13862 16690 13922 16766
rect 15009 16763 15075 16766
rect 11145 16688 13922 16690
rect 11145 16632 11150 16688
rect 11206 16632 13922 16688
rect 11145 16630 13922 16632
rect 13997 16690 14063 16693
rect 15540 16690 16000 16720
rect 13997 16688 16000 16690
rect 13997 16632 14002 16688
rect 14058 16632 16000 16688
rect 13997 16630 16000 16632
rect 11145 16627 11211 16630
rect 13997 16627 14063 16630
rect 15540 16600 16000 16630
rect 9673 16554 9739 16557
rect 10726 16554 10732 16556
rect 9673 16552 10732 16554
rect 9673 16496 9678 16552
rect 9734 16496 10732 16552
rect 9673 16494 10732 16496
rect 9673 16491 9739 16494
rect 10726 16492 10732 16494
rect 10796 16492 10802 16556
rect 13486 16492 13492 16556
rect 13556 16554 13562 16556
rect 13629 16554 13695 16557
rect 15377 16554 15443 16557
rect 13556 16552 13695 16554
rect 13556 16496 13634 16552
rect 13690 16496 13695 16552
rect 13556 16494 13695 16496
rect 13556 16492 13562 16494
rect 13629 16491 13695 16494
rect 13816 16552 15443 16554
rect 13816 16496 15382 16552
rect 15438 16496 15443 16552
rect 13816 16494 15443 16496
rect 11605 16418 11671 16421
rect 13816 16418 13876 16494
rect 15377 16491 15443 16494
rect 11605 16416 13876 16418
rect 11605 16360 11610 16416
rect 11666 16360 13876 16416
rect 11605 16358 13876 16360
rect 15009 16418 15075 16421
rect 15540 16418 16000 16448
rect 15009 16416 16000 16418
rect 15009 16360 15014 16416
rect 15070 16360 16000 16416
rect 15009 16358 16000 16360
rect 11605 16355 11671 16358
rect 15009 16355 15075 16358
rect 4304 16352 4620 16353
rect 4304 16288 4310 16352
rect 4374 16288 4390 16352
rect 4454 16288 4470 16352
rect 4534 16288 4550 16352
rect 4614 16288 4620 16352
rect 4304 16287 4620 16288
rect 7662 16352 7978 16353
rect 7662 16288 7668 16352
rect 7732 16288 7748 16352
rect 7812 16288 7828 16352
rect 7892 16288 7908 16352
rect 7972 16288 7978 16352
rect 7662 16287 7978 16288
rect 11020 16352 11336 16353
rect 11020 16288 11026 16352
rect 11090 16288 11106 16352
rect 11170 16288 11186 16352
rect 11250 16288 11266 16352
rect 11330 16288 11336 16352
rect 11020 16287 11336 16288
rect 14378 16352 14694 16353
rect 14378 16288 14384 16352
rect 14448 16288 14464 16352
rect 14528 16288 14544 16352
rect 14608 16288 14624 16352
rect 14688 16288 14694 16352
rect 15540 16328 16000 16358
rect 14378 16287 14694 16288
rect -300 16146 160 16176
rect 749 16146 815 16149
rect -300 16144 815 16146
rect -300 16088 754 16144
rect 810 16088 815 16144
rect -300 16086 815 16088
rect -300 16056 160 16086
rect 749 16083 815 16086
rect 14641 16146 14707 16149
rect 15540 16146 16000 16176
rect 14641 16144 16000 16146
rect 14641 16088 14646 16144
rect 14702 16088 16000 16144
rect 14641 16086 16000 16088
rect 14641 16083 14707 16086
rect 15540 16056 16000 16086
rect 15285 16012 15351 16013
rect 15285 16010 15332 16012
rect 15240 16008 15332 16010
rect 15240 15952 15290 16008
rect 15240 15950 15332 15952
rect 15285 15948 15332 15950
rect 15396 15948 15402 16012
rect 15285 15947 15351 15948
rect 7230 15812 7236 15876
rect 7300 15874 7306 15876
rect 7557 15874 7623 15877
rect 7300 15872 7623 15874
rect 7300 15816 7562 15872
rect 7618 15816 7623 15872
rect 7300 15814 7623 15816
rect 7300 15812 7306 15814
rect 7557 15811 7623 15814
rect 13077 15874 13143 15877
rect 15540 15874 16000 15904
rect 13077 15872 16000 15874
rect 13077 15816 13082 15872
rect 13138 15816 16000 15872
rect 13077 15814 16000 15816
rect 13077 15811 13143 15814
rect 2625 15808 2941 15809
rect 2625 15744 2631 15808
rect 2695 15744 2711 15808
rect 2775 15744 2791 15808
rect 2855 15744 2871 15808
rect 2935 15744 2941 15808
rect 2625 15743 2941 15744
rect 5983 15808 6299 15809
rect 5983 15744 5989 15808
rect 6053 15744 6069 15808
rect 6133 15744 6149 15808
rect 6213 15744 6229 15808
rect 6293 15744 6299 15808
rect 5983 15743 6299 15744
rect 9341 15808 9657 15809
rect 9341 15744 9347 15808
rect 9411 15744 9427 15808
rect 9491 15744 9507 15808
rect 9571 15744 9587 15808
rect 9651 15744 9657 15808
rect 9341 15743 9657 15744
rect 12699 15808 13015 15809
rect 12699 15744 12705 15808
rect 12769 15744 12785 15808
rect 12849 15744 12865 15808
rect 12929 15744 12945 15808
rect 13009 15744 13015 15808
rect 15540 15784 16000 15814
rect 12699 15743 13015 15744
rect 9673 15602 9739 15605
rect 10726 15602 10732 15604
rect 9673 15600 10732 15602
rect 9673 15544 9678 15600
rect 9734 15544 10732 15600
rect 9673 15542 10732 15544
rect 9673 15539 9739 15542
rect 10726 15540 10732 15542
rect 10796 15602 10802 15604
rect 11053 15602 11119 15605
rect 10796 15600 11119 15602
rect 10796 15544 11058 15600
rect 11114 15544 11119 15600
rect 10796 15542 11119 15544
rect 10796 15540 10802 15542
rect 11053 15539 11119 15542
rect 11462 15540 11468 15604
rect 11532 15602 11538 15604
rect 12065 15602 12131 15605
rect 11532 15600 12131 15602
rect 11532 15544 12070 15600
rect 12126 15544 12131 15600
rect 11532 15542 12131 15544
rect 11532 15540 11538 15542
rect 12065 15539 12131 15542
rect 13813 15602 13879 15605
rect 15540 15602 16000 15632
rect 13813 15600 16000 15602
rect 13813 15544 13818 15600
rect 13874 15544 16000 15600
rect 13813 15542 16000 15544
rect 13813 15539 13879 15542
rect 15540 15512 16000 15542
rect 9990 15404 9996 15468
rect 10060 15466 10066 15468
rect 11697 15466 11763 15469
rect 10060 15464 11763 15466
rect 10060 15408 11702 15464
rect 11758 15408 11763 15464
rect 10060 15406 11763 15408
rect 10060 15404 10066 15406
rect 11697 15403 11763 15406
rect 13724 15406 14842 15466
rect -300 15330 160 15360
rect 13724 15333 13784 15406
rect 749 15330 815 15333
rect -300 15328 815 15330
rect -300 15272 754 15328
rect 810 15272 815 15328
rect -300 15270 815 15272
rect -300 15240 160 15270
rect 749 15267 815 15270
rect 13721 15328 13787 15333
rect 13721 15272 13726 15328
rect 13782 15272 13787 15328
rect 13721 15267 13787 15272
rect 14782 15330 14842 15406
rect 15540 15330 16000 15360
rect 14782 15270 16000 15330
rect 4304 15264 4620 15265
rect 4304 15200 4310 15264
rect 4374 15200 4390 15264
rect 4454 15200 4470 15264
rect 4534 15200 4550 15264
rect 4614 15200 4620 15264
rect 4304 15199 4620 15200
rect 7662 15264 7978 15265
rect 7662 15200 7668 15264
rect 7732 15200 7748 15264
rect 7812 15200 7828 15264
rect 7892 15200 7908 15264
rect 7972 15200 7978 15264
rect 7662 15199 7978 15200
rect 11020 15264 11336 15265
rect 11020 15200 11026 15264
rect 11090 15200 11106 15264
rect 11170 15200 11186 15264
rect 11250 15200 11266 15264
rect 11330 15200 11336 15264
rect 11020 15199 11336 15200
rect 14378 15264 14694 15265
rect 14378 15200 14384 15264
rect 14448 15200 14464 15264
rect 14528 15200 14544 15264
rect 14608 15200 14624 15264
rect 14688 15200 14694 15264
rect 15540 15240 16000 15270
rect 14378 15199 14694 15200
rect 12157 15194 12223 15197
rect 14089 15194 14155 15197
rect 12157 15192 14155 15194
rect 12157 15136 12162 15192
rect 12218 15136 14094 15192
rect 14150 15136 14155 15192
rect 12157 15134 14155 15136
rect 12157 15131 12223 15134
rect 14089 15131 14155 15134
rect 9857 15058 9923 15061
rect 12525 15058 12591 15061
rect 13118 15058 13124 15060
rect 9857 15056 13124 15058
rect 9857 15000 9862 15056
rect 9918 15000 12530 15056
rect 12586 15000 13124 15056
rect 9857 14998 13124 15000
rect 9857 14995 9923 14998
rect 12525 14995 12591 14998
rect 13118 14996 13124 14998
rect 13188 14996 13194 15060
rect 13905 15058 13971 15061
rect 15540 15058 16000 15088
rect 13905 15056 16000 15058
rect 13905 15000 13910 15056
rect 13966 15000 16000 15056
rect 13905 14998 16000 15000
rect 13905 14995 13971 14998
rect 15540 14968 16000 14998
rect 10777 14922 10843 14925
rect 15142 14922 15148 14924
rect 10777 14920 15148 14922
rect 10777 14864 10782 14920
rect 10838 14864 15148 14920
rect 10777 14862 15148 14864
rect 10777 14859 10843 14862
rect 15142 14860 15148 14862
rect 15212 14860 15218 14924
rect 9765 14786 9831 14789
rect 10317 14786 10383 14789
rect 9765 14784 10383 14786
rect 9765 14728 9770 14784
rect 9826 14728 10322 14784
rect 10378 14728 10383 14784
rect 9765 14726 10383 14728
rect 9765 14723 9831 14726
rect 10317 14723 10383 14726
rect 14365 14786 14431 14789
rect 15540 14786 16000 14816
rect 14365 14784 16000 14786
rect 14365 14728 14370 14784
rect 14426 14728 16000 14784
rect 14365 14726 16000 14728
rect 14365 14723 14431 14726
rect 2625 14720 2941 14721
rect 2625 14656 2631 14720
rect 2695 14656 2711 14720
rect 2775 14656 2791 14720
rect 2855 14656 2871 14720
rect 2935 14656 2941 14720
rect 2625 14655 2941 14656
rect 5983 14720 6299 14721
rect 5983 14656 5989 14720
rect 6053 14656 6069 14720
rect 6133 14656 6149 14720
rect 6213 14656 6229 14720
rect 6293 14656 6299 14720
rect 5983 14655 6299 14656
rect 9341 14720 9657 14721
rect 9341 14656 9347 14720
rect 9411 14656 9427 14720
rect 9491 14656 9507 14720
rect 9571 14656 9587 14720
rect 9651 14656 9657 14720
rect 9341 14655 9657 14656
rect 12699 14720 13015 14721
rect 12699 14656 12705 14720
rect 12769 14656 12785 14720
rect 12849 14656 12865 14720
rect 12929 14656 12945 14720
rect 13009 14656 13015 14720
rect 15540 14696 16000 14726
rect 12699 14655 13015 14656
rect 10174 14588 10180 14652
rect 10244 14650 10250 14652
rect 10317 14650 10383 14653
rect 11053 14650 11119 14653
rect 10244 14648 11119 14650
rect 10244 14592 10322 14648
rect 10378 14592 11058 14648
rect 11114 14592 11119 14648
rect 10244 14590 11119 14592
rect 10244 14588 10250 14590
rect 10317 14587 10383 14590
rect 11053 14587 11119 14590
rect 11881 14650 11947 14653
rect 12433 14650 12499 14653
rect 11881 14648 12499 14650
rect 11881 14592 11886 14648
rect 11942 14592 12438 14648
rect 12494 14592 12499 14648
rect 11881 14590 12499 14592
rect 11881 14587 11947 14590
rect 12433 14587 12499 14590
rect 14222 14588 14228 14652
rect 14292 14650 14298 14652
rect 15377 14650 15443 14653
rect 14292 14648 15443 14650
rect 14292 14592 15382 14648
rect 15438 14592 15443 14648
rect 14292 14590 15443 14592
rect 14292 14588 14298 14590
rect 15377 14587 15443 14590
rect -300 14514 160 14544
rect 841 14514 907 14517
rect -300 14512 907 14514
rect -300 14456 846 14512
rect 902 14456 907 14512
rect -300 14454 907 14456
rect -300 14424 160 14454
rect 841 14451 907 14454
rect 10593 14514 10659 14517
rect 11145 14514 11211 14517
rect 11973 14514 12039 14517
rect 10593 14512 12039 14514
rect 10593 14456 10598 14512
rect 10654 14456 11150 14512
rect 11206 14456 11978 14512
rect 12034 14456 12039 14512
rect 10593 14454 12039 14456
rect 10593 14451 10659 14454
rect 11145 14451 11211 14454
rect 11973 14451 12039 14454
rect 12985 14514 13051 14517
rect 13302 14514 13308 14516
rect 12985 14512 13308 14514
rect 12985 14456 12990 14512
rect 13046 14456 13308 14512
rect 12985 14454 13308 14456
rect 12985 14451 13051 14454
rect 13302 14452 13308 14454
rect 13372 14452 13378 14516
rect 15540 14514 16000 14544
rect 14000 14454 16000 14514
rect 13854 14378 13860 14380
rect 9676 14318 13860 14378
rect 9676 14245 9736 14318
rect 13854 14316 13860 14318
rect 13924 14316 13930 14380
rect 9673 14240 9739 14245
rect 9673 14184 9678 14240
rect 9734 14184 9739 14240
rect 9673 14179 9739 14184
rect 11697 14242 11763 14245
rect 14000 14242 14060 14454
rect 15540 14424 16000 14454
rect 11697 14240 14060 14242
rect 11697 14184 11702 14240
rect 11758 14184 14060 14240
rect 11697 14182 14060 14184
rect 15009 14242 15075 14245
rect 15540 14242 16000 14272
rect 15009 14240 16000 14242
rect 15009 14184 15014 14240
rect 15070 14184 16000 14240
rect 15009 14182 16000 14184
rect 11697 14179 11763 14182
rect 15009 14179 15075 14182
rect 4304 14176 4620 14177
rect 4304 14112 4310 14176
rect 4374 14112 4390 14176
rect 4454 14112 4470 14176
rect 4534 14112 4550 14176
rect 4614 14112 4620 14176
rect 4304 14111 4620 14112
rect 7662 14176 7978 14177
rect 7662 14112 7668 14176
rect 7732 14112 7748 14176
rect 7812 14112 7828 14176
rect 7892 14112 7908 14176
rect 7972 14112 7978 14176
rect 7662 14111 7978 14112
rect 11020 14176 11336 14177
rect 11020 14112 11026 14176
rect 11090 14112 11106 14176
rect 11170 14112 11186 14176
rect 11250 14112 11266 14176
rect 11330 14112 11336 14176
rect 11020 14111 11336 14112
rect 14378 14176 14694 14177
rect 14378 14112 14384 14176
rect 14448 14112 14464 14176
rect 14528 14112 14544 14176
rect 14608 14112 14624 14176
rect 14688 14112 14694 14176
rect 15540 14152 16000 14182
rect 14378 14111 14694 14112
rect 7649 13970 7715 13973
rect 11329 13970 11395 13973
rect 7649 13968 11395 13970
rect 7649 13912 7654 13968
rect 7710 13912 11334 13968
rect 11390 13912 11395 13968
rect 7649 13910 11395 13912
rect 7649 13907 7715 13910
rect 11329 13907 11395 13910
rect 12198 13908 12204 13972
rect 12268 13970 12274 13972
rect 12433 13970 12499 13973
rect 12268 13968 12499 13970
rect 12268 13912 12438 13968
rect 12494 13912 12499 13968
rect 12268 13910 12499 13912
rect 12268 13908 12274 13910
rect 12433 13907 12499 13910
rect 14089 13970 14155 13973
rect 15540 13970 16000 14000
rect 14089 13968 16000 13970
rect 14089 13912 14094 13968
rect 14150 13912 16000 13968
rect 14089 13910 16000 13912
rect 14089 13907 14155 13910
rect 15540 13880 16000 13910
rect -300 13698 160 13728
rect 1577 13698 1643 13701
rect -300 13696 1643 13698
rect -300 13640 1582 13696
rect 1638 13640 1643 13696
rect -300 13638 1643 13640
rect -300 13608 160 13638
rect 1577 13635 1643 13638
rect 7414 13636 7420 13700
rect 7484 13698 7490 13700
rect 7557 13698 7623 13701
rect 7484 13696 7623 13698
rect 7484 13640 7562 13696
rect 7618 13640 7623 13696
rect 7484 13638 7623 13640
rect 7484 13636 7490 13638
rect 7557 13635 7623 13638
rect 14365 13698 14431 13701
rect 15540 13698 16000 13728
rect 14365 13696 16000 13698
rect 14365 13640 14370 13696
rect 14426 13640 16000 13696
rect 14365 13638 16000 13640
rect 14365 13635 14431 13638
rect 2625 13632 2941 13633
rect 2625 13568 2631 13632
rect 2695 13568 2711 13632
rect 2775 13568 2791 13632
rect 2855 13568 2871 13632
rect 2935 13568 2941 13632
rect 2625 13567 2941 13568
rect 5983 13632 6299 13633
rect 5983 13568 5989 13632
rect 6053 13568 6069 13632
rect 6133 13568 6149 13632
rect 6213 13568 6229 13632
rect 6293 13568 6299 13632
rect 5983 13567 6299 13568
rect 9341 13632 9657 13633
rect 9341 13568 9347 13632
rect 9411 13568 9427 13632
rect 9491 13568 9507 13632
rect 9571 13568 9587 13632
rect 9651 13568 9657 13632
rect 9341 13567 9657 13568
rect 12699 13632 13015 13633
rect 12699 13568 12705 13632
rect 12769 13568 12785 13632
rect 12849 13568 12865 13632
rect 12929 13568 12945 13632
rect 13009 13568 13015 13632
rect 15540 13608 16000 13638
rect 12699 13567 13015 13568
rect 8886 13364 8892 13428
rect 8956 13426 8962 13428
rect 9397 13426 9463 13429
rect 8956 13424 9463 13426
rect 8956 13368 9402 13424
rect 9458 13368 9463 13424
rect 8956 13366 9463 13368
rect 8956 13364 8962 13366
rect 9397 13363 9463 13366
rect 13997 13426 14063 13429
rect 15540 13426 16000 13456
rect 13997 13424 16000 13426
rect 13997 13368 14002 13424
rect 14058 13368 16000 13424
rect 13997 13366 16000 13368
rect 13997 13363 14063 13366
rect 15540 13336 16000 13366
rect 8569 13290 8635 13293
rect 9029 13290 9095 13293
rect 8569 13288 9095 13290
rect 8569 13232 8574 13288
rect 8630 13232 9034 13288
rect 9090 13232 9095 13288
rect 8569 13230 9095 13232
rect 8569 13227 8635 13230
rect 9029 13227 9095 13230
rect 11237 13290 11303 13293
rect 11462 13290 11468 13292
rect 11237 13288 11468 13290
rect 11237 13232 11242 13288
rect 11298 13232 11468 13288
rect 11237 13230 11468 13232
rect 11237 13227 11303 13230
rect 11462 13228 11468 13230
rect 11532 13228 11538 13292
rect 13077 13290 13143 13293
rect 13077 13288 14842 13290
rect 13077 13232 13082 13288
rect 13138 13232 14842 13288
rect 13077 13230 14842 13232
rect 13077 13227 13143 13230
rect 14782 13154 14842 13230
rect 15540 13154 16000 13184
rect 14782 13094 16000 13154
rect 4304 13088 4620 13089
rect 4304 13024 4310 13088
rect 4374 13024 4390 13088
rect 4454 13024 4470 13088
rect 4534 13024 4550 13088
rect 4614 13024 4620 13088
rect 4304 13023 4620 13024
rect 7662 13088 7978 13089
rect 7662 13024 7668 13088
rect 7732 13024 7748 13088
rect 7812 13024 7828 13088
rect 7892 13024 7908 13088
rect 7972 13024 7978 13088
rect 7662 13023 7978 13024
rect 11020 13088 11336 13089
rect 11020 13024 11026 13088
rect 11090 13024 11106 13088
rect 11170 13024 11186 13088
rect 11250 13024 11266 13088
rect 11330 13024 11336 13088
rect 11020 13023 11336 13024
rect 14378 13088 14694 13089
rect 14378 13024 14384 13088
rect 14448 13024 14464 13088
rect 14528 13024 14544 13088
rect 14608 13024 14624 13088
rect 14688 13024 14694 13088
rect 15540 13064 16000 13094
rect 14378 13023 14694 13024
rect -300 12882 160 12912
rect 841 12882 907 12885
rect -300 12880 907 12882
rect -300 12824 846 12880
rect 902 12824 907 12880
rect -300 12822 907 12824
rect -300 12792 160 12822
rect 841 12819 907 12822
rect 12341 12882 12407 12885
rect 15540 12882 16000 12912
rect 12341 12880 16000 12882
rect 12341 12824 12346 12880
rect 12402 12824 16000 12880
rect 12341 12822 16000 12824
rect 12341 12819 12407 12822
rect 15540 12792 16000 12822
rect 12709 12746 12775 12749
rect 12436 12744 12775 12746
rect 12436 12688 12714 12744
rect 12770 12688 12775 12744
rect 12436 12686 12775 12688
rect 11329 12610 11395 12613
rect 12436 12610 12496 12686
rect 12709 12683 12775 12686
rect 15540 12610 16000 12640
rect 11329 12608 12496 12610
rect 11329 12552 11334 12608
rect 11390 12552 12496 12608
rect 11329 12550 12496 12552
rect 11329 12547 11395 12550
rect 2625 12544 2941 12545
rect 2625 12480 2631 12544
rect 2695 12480 2711 12544
rect 2775 12480 2791 12544
rect 2855 12480 2871 12544
rect 2935 12480 2941 12544
rect 2625 12479 2941 12480
rect 5983 12544 6299 12545
rect 5983 12480 5989 12544
rect 6053 12480 6069 12544
rect 6133 12480 6149 12544
rect 6213 12480 6229 12544
rect 6293 12480 6299 12544
rect 5983 12479 6299 12480
rect 9341 12544 9657 12545
rect 9341 12480 9347 12544
rect 9411 12480 9427 12544
rect 9491 12480 9507 12544
rect 9571 12480 9587 12544
rect 9651 12480 9657 12544
rect 9341 12479 9657 12480
rect 12436 12477 12496 12550
rect 13724 12550 16000 12610
rect 12699 12544 13015 12545
rect 12699 12480 12705 12544
rect 12769 12480 12785 12544
rect 12849 12480 12865 12544
rect 12929 12480 12945 12544
rect 13009 12480 13015 12544
rect 12699 12479 13015 12480
rect 13724 12477 13784 12550
rect 15540 12520 16000 12550
rect 12433 12472 12499 12477
rect 12433 12416 12438 12472
rect 12494 12416 12499 12472
rect 12433 12411 12499 12416
rect 13721 12472 13787 12477
rect 13721 12416 13726 12472
rect 13782 12416 13787 12472
rect 13721 12411 13787 12416
rect 9397 12338 9463 12341
rect 10225 12338 10291 12341
rect 9397 12336 10291 12338
rect 9397 12280 9402 12336
rect 9458 12280 10230 12336
rect 10286 12280 10291 12336
rect 9397 12278 10291 12280
rect 9397 12275 9463 12278
rect 10225 12275 10291 12278
rect 12157 12338 12223 12341
rect 15540 12338 16000 12368
rect 12157 12336 16000 12338
rect 12157 12280 12162 12336
rect 12218 12280 16000 12336
rect 12157 12278 16000 12280
rect 12157 12275 12223 12278
rect 15540 12248 16000 12278
rect 13445 12202 13511 12205
rect 13445 12200 13554 12202
rect 13445 12144 13450 12200
rect 13506 12144 13554 12200
rect 13445 12139 13554 12144
rect -300 12066 160 12096
rect 841 12066 907 12069
rect -300 12064 907 12066
rect -300 12008 846 12064
rect 902 12008 907 12064
rect -300 12006 907 12008
rect -300 11976 160 12006
rect 841 12003 907 12006
rect 11605 12066 11671 12069
rect 13494 12066 13554 12139
rect 14230 12142 14842 12202
rect 13721 12066 13787 12069
rect 11605 12064 13370 12066
rect 11605 12008 11610 12064
rect 11666 12008 13370 12064
rect 11605 12006 13370 12008
rect 13494 12064 13787 12066
rect 13494 12008 13726 12064
rect 13782 12008 13787 12064
rect 13494 12006 13787 12008
rect 11605 12003 11671 12006
rect 4304 12000 4620 12001
rect 4304 11936 4310 12000
rect 4374 11936 4390 12000
rect 4454 11936 4470 12000
rect 4534 11936 4550 12000
rect 4614 11936 4620 12000
rect 4304 11935 4620 11936
rect 7662 12000 7978 12001
rect 7662 11936 7668 12000
rect 7732 11936 7748 12000
rect 7812 11936 7828 12000
rect 7892 11936 7908 12000
rect 7972 11936 7978 12000
rect 7662 11935 7978 11936
rect 11020 12000 11336 12001
rect 11020 11936 11026 12000
rect 11090 11936 11106 12000
rect 11170 11936 11186 12000
rect 11250 11936 11266 12000
rect 11330 11936 11336 12000
rect 11020 11935 11336 11936
rect 13310 11930 13370 12006
rect 13721 12003 13787 12006
rect 14230 11930 14290 12142
rect 14782 12066 14842 12142
rect 15540 12066 16000 12096
rect 14782 12006 16000 12066
rect 14378 12000 14694 12001
rect 14378 11936 14384 12000
rect 14448 11936 14464 12000
rect 14528 11936 14544 12000
rect 14608 11936 14624 12000
rect 14688 11936 14694 12000
rect 15540 11976 16000 12006
rect 14378 11935 14694 11936
rect 13310 11870 14290 11930
rect 12065 11794 12131 11797
rect 15540 11794 16000 11824
rect 12065 11792 16000 11794
rect 12065 11736 12070 11792
rect 12126 11736 16000 11792
rect 12065 11734 16000 11736
rect 12065 11731 12131 11734
rect 15540 11704 16000 11734
rect 12065 11658 12131 11661
rect 12065 11656 14106 11658
rect 12065 11600 12070 11656
rect 12126 11600 14106 11656
rect 12065 11598 14106 11600
rect 12065 11595 12131 11598
rect 11881 11522 11947 11525
rect 12525 11522 12591 11525
rect 11881 11520 12591 11522
rect 11881 11464 11886 11520
rect 11942 11464 12530 11520
rect 12586 11464 12591 11520
rect 11881 11462 12591 11464
rect 14046 11522 14106 11598
rect 15540 11522 16000 11552
rect 14046 11462 16000 11522
rect 11881 11459 11947 11462
rect 12525 11459 12591 11462
rect 2625 11456 2941 11457
rect 2625 11392 2631 11456
rect 2695 11392 2711 11456
rect 2775 11392 2791 11456
rect 2855 11392 2871 11456
rect 2935 11392 2941 11456
rect 2625 11391 2941 11392
rect 5983 11456 6299 11457
rect 5983 11392 5989 11456
rect 6053 11392 6069 11456
rect 6133 11392 6149 11456
rect 6213 11392 6229 11456
rect 6293 11392 6299 11456
rect 5983 11391 6299 11392
rect 9341 11456 9657 11457
rect 9341 11392 9347 11456
rect 9411 11392 9427 11456
rect 9491 11392 9507 11456
rect 9571 11392 9587 11456
rect 9651 11392 9657 11456
rect 9341 11391 9657 11392
rect 12699 11456 13015 11457
rect 12699 11392 12705 11456
rect 12769 11392 12785 11456
rect 12849 11392 12865 11456
rect 12929 11392 12945 11456
rect 13009 11392 13015 11456
rect 15540 11432 16000 11462
rect 12699 11391 13015 11392
rect -300 11250 160 11280
rect 841 11250 907 11253
rect -300 11248 907 11250
rect -300 11192 846 11248
rect 902 11192 907 11248
rect -300 11190 907 11192
rect -300 11160 160 11190
rect 841 11187 907 11190
rect 8845 11250 8911 11253
rect 11789 11250 11855 11253
rect 15540 11250 16000 11280
rect 8845 11248 8954 11250
rect 8845 11192 8850 11248
rect 8906 11192 8954 11248
rect 8845 11187 8954 11192
rect 11789 11248 16000 11250
rect 11789 11192 11794 11248
rect 11850 11192 16000 11248
rect 11789 11190 16000 11192
rect 11789 11187 11855 11190
rect 3734 11052 3740 11116
rect 3804 11114 3810 11116
rect 7465 11114 7531 11117
rect 3804 11112 7531 11114
rect 3804 11056 7470 11112
rect 7526 11056 7531 11112
rect 3804 11054 7531 11056
rect 3804 11052 3810 11054
rect 7465 11051 7531 11054
rect 8894 10978 8954 11187
rect 15540 11160 16000 11190
rect 10317 11114 10383 11117
rect 12709 11114 12775 11117
rect 10317 11112 12775 11114
rect 10317 11056 10322 11112
rect 10378 11056 12714 11112
rect 12770 11056 12775 11112
rect 10317 11054 12775 11056
rect 10317 11051 10383 11054
rect 12709 11051 12775 11054
rect 14230 11054 14842 11114
rect 9029 10978 9095 10981
rect 8894 10976 9095 10978
rect 8894 10920 9034 10976
rect 9090 10920 9095 10976
rect 8894 10918 9095 10920
rect 9029 10915 9095 10918
rect 11973 10978 12039 10981
rect 14230 10978 14290 11054
rect 11973 10976 14290 10978
rect 11973 10920 11978 10976
rect 12034 10920 14290 10976
rect 11973 10918 14290 10920
rect 14782 10978 14842 11054
rect 15540 10978 16000 11008
rect 14782 10918 16000 10978
rect 11973 10915 12039 10918
rect 4304 10912 4620 10913
rect 4304 10848 4310 10912
rect 4374 10848 4390 10912
rect 4454 10848 4470 10912
rect 4534 10848 4550 10912
rect 4614 10848 4620 10912
rect 4304 10847 4620 10848
rect 7662 10912 7978 10913
rect 7662 10848 7668 10912
rect 7732 10848 7748 10912
rect 7812 10848 7828 10912
rect 7892 10848 7908 10912
rect 7972 10848 7978 10912
rect 7662 10847 7978 10848
rect 11020 10912 11336 10913
rect 11020 10848 11026 10912
rect 11090 10848 11106 10912
rect 11170 10848 11186 10912
rect 11250 10848 11266 10912
rect 11330 10848 11336 10912
rect 11020 10847 11336 10848
rect 14378 10912 14694 10913
rect 14378 10848 14384 10912
rect 14448 10848 14464 10912
rect 14528 10848 14544 10912
rect 14608 10848 14624 10912
rect 14688 10848 14694 10912
rect 15540 10888 16000 10918
rect 14378 10847 14694 10848
rect 1853 10706 1919 10709
rect 8201 10706 8267 10709
rect 1853 10704 8267 10706
rect 1853 10648 1858 10704
rect 1914 10648 8206 10704
rect 8262 10648 8267 10704
rect 1853 10646 8267 10648
rect 1853 10643 1919 10646
rect 8201 10643 8267 10646
rect 11462 10644 11468 10708
rect 11532 10706 11538 10708
rect 11881 10706 11947 10709
rect 11532 10704 11947 10706
rect 11532 10648 11886 10704
rect 11942 10648 11947 10704
rect 11532 10646 11947 10648
rect 11532 10644 11538 10646
rect 11881 10643 11947 10646
rect 12341 10706 12407 10709
rect 15540 10706 16000 10736
rect 12341 10704 16000 10706
rect 12341 10648 12346 10704
rect 12402 10648 16000 10704
rect 12341 10646 16000 10648
rect 12341 10643 12407 10646
rect 15540 10616 16000 10646
rect 3877 10570 3943 10573
rect 9397 10570 9463 10573
rect 3877 10568 9463 10570
rect 3877 10512 3882 10568
rect 3938 10512 9402 10568
rect 9458 10512 9463 10568
rect 3877 10510 9463 10512
rect 3877 10507 3943 10510
rect 9397 10507 9463 10510
rect 12341 10570 12407 10573
rect 12566 10570 12572 10572
rect 12341 10568 12572 10570
rect 12341 10512 12346 10568
rect 12402 10512 12572 10568
rect 12341 10510 12572 10512
rect 12341 10507 12407 10510
rect 12566 10508 12572 10510
rect 12636 10508 12642 10572
rect -300 10434 160 10464
rect 841 10434 907 10437
rect -300 10432 907 10434
rect -300 10376 846 10432
rect 902 10376 907 10432
rect -300 10374 907 10376
rect -300 10344 160 10374
rect 841 10371 907 10374
rect 14089 10434 14155 10437
rect 15540 10434 16000 10464
rect 14089 10432 16000 10434
rect 14089 10376 14094 10432
rect 14150 10376 16000 10432
rect 14089 10374 16000 10376
rect 14089 10371 14155 10374
rect 2625 10368 2941 10369
rect 2625 10304 2631 10368
rect 2695 10304 2711 10368
rect 2775 10304 2791 10368
rect 2855 10304 2871 10368
rect 2935 10304 2941 10368
rect 2625 10303 2941 10304
rect 5983 10368 6299 10369
rect 5983 10304 5989 10368
rect 6053 10304 6069 10368
rect 6133 10304 6149 10368
rect 6213 10304 6229 10368
rect 6293 10304 6299 10368
rect 5983 10303 6299 10304
rect 9341 10368 9657 10369
rect 9341 10304 9347 10368
rect 9411 10304 9427 10368
rect 9491 10304 9507 10368
rect 9571 10304 9587 10368
rect 9651 10304 9657 10368
rect 9341 10303 9657 10304
rect 12699 10368 13015 10369
rect 12699 10304 12705 10368
rect 12769 10304 12785 10368
rect 12849 10304 12865 10368
rect 12929 10304 12945 10368
rect 13009 10304 13015 10368
rect 15540 10344 16000 10374
rect 12699 10303 13015 10304
rect 11605 10162 11671 10165
rect 12433 10162 12499 10165
rect 11605 10160 12499 10162
rect 11605 10104 11610 10160
rect 11666 10104 12438 10160
rect 12494 10104 12499 10160
rect 11605 10102 12499 10104
rect 11605 10099 11671 10102
rect 12433 10099 12499 10102
rect 13997 10162 14063 10165
rect 15540 10162 16000 10192
rect 13997 10160 16000 10162
rect 13997 10104 14002 10160
rect 14058 10104 16000 10160
rect 13997 10102 16000 10104
rect 13997 10099 14063 10102
rect 15540 10072 16000 10102
rect 10133 10026 10199 10029
rect 10409 10026 10475 10029
rect 10133 10024 10475 10026
rect 10133 9968 10138 10024
rect 10194 9968 10414 10024
rect 10470 9968 10475 10024
rect 10133 9966 10475 9968
rect 10133 9963 10199 9966
rect 10409 9963 10475 9966
rect 14230 9966 14842 10026
rect 13629 9890 13695 9893
rect 14230 9890 14290 9966
rect 13629 9888 14290 9890
rect 13629 9832 13634 9888
rect 13690 9832 14290 9888
rect 13629 9830 14290 9832
rect 14782 9890 14842 9966
rect 15540 9890 16000 9920
rect 14782 9830 16000 9890
rect 13629 9827 13695 9830
rect 4304 9824 4620 9825
rect 4304 9760 4310 9824
rect 4374 9760 4390 9824
rect 4454 9760 4470 9824
rect 4534 9760 4550 9824
rect 4614 9760 4620 9824
rect 4304 9759 4620 9760
rect 7662 9824 7978 9825
rect 7662 9760 7668 9824
rect 7732 9760 7748 9824
rect 7812 9760 7828 9824
rect 7892 9760 7908 9824
rect 7972 9760 7978 9824
rect 7662 9759 7978 9760
rect 11020 9824 11336 9825
rect 11020 9760 11026 9824
rect 11090 9760 11106 9824
rect 11170 9760 11186 9824
rect 11250 9760 11266 9824
rect 11330 9760 11336 9824
rect 11020 9759 11336 9760
rect 14378 9824 14694 9825
rect 14378 9760 14384 9824
rect 14448 9760 14464 9824
rect 14528 9760 14544 9824
rect 14608 9760 14624 9824
rect 14688 9760 14694 9824
rect 15540 9800 16000 9830
rect 14378 9759 14694 9760
rect 13118 9692 13124 9756
rect 13188 9754 13194 9756
rect 13261 9754 13327 9757
rect 13188 9752 13327 9754
rect 13188 9696 13266 9752
rect 13322 9696 13327 9752
rect 13188 9694 13327 9696
rect 13188 9692 13194 9694
rect 13261 9691 13327 9694
rect -300 9618 160 9648
rect 2773 9618 2839 9621
rect -300 9616 2839 9618
rect -300 9560 2778 9616
rect 2834 9560 2839 9616
rect -300 9558 2839 9560
rect -300 9528 160 9558
rect 2773 9555 2839 9558
rect 12433 9618 12499 9621
rect 13077 9618 13143 9621
rect 12433 9616 13143 9618
rect 12433 9560 12438 9616
rect 12494 9560 13082 9616
rect 13138 9560 13143 9616
rect 12433 9558 13143 9560
rect 12433 9555 12499 9558
rect 13077 9555 13143 9558
rect 13261 9618 13327 9621
rect 13721 9618 13787 9621
rect 13261 9616 13787 9618
rect 13261 9560 13266 9616
rect 13322 9560 13726 9616
rect 13782 9560 13787 9616
rect 13261 9558 13787 9560
rect 13261 9555 13327 9558
rect 13721 9555 13787 9558
rect 15285 9618 15351 9621
rect 15540 9618 16000 9648
rect 15285 9616 16000 9618
rect 15285 9560 15290 9616
rect 15346 9560 16000 9616
rect 15285 9558 16000 9560
rect 15285 9555 15351 9558
rect 15540 9528 16000 9558
rect 9581 9482 9647 9485
rect 10726 9482 10732 9484
rect 9581 9480 10732 9482
rect 9581 9424 9586 9480
rect 9642 9424 10732 9480
rect 9581 9422 10732 9424
rect 9581 9419 9647 9422
rect 10726 9420 10732 9422
rect 10796 9482 10802 9484
rect 11605 9482 11671 9485
rect 10796 9480 11671 9482
rect 10796 9424 11610 9480
rect 11666 9424 11671 9480
rect 10796 9422 11671 9424
rect 10796 9420 10802 9422
rect 11605 9419 11671 9422
rect 10133 9348 10199 9349
rect 10133 9346 10180 9348
rect 10088 9344 10180 9346
rect 10088 9288 10138 9344
rect 10088 9286 10180 9288
rect 10133 9284 10180 9286
rect 10244 9284 10250 9348
rect 10501 9346 10567 9349
rect 11421 9346 11487 9349
rect 10501 9344 11487 9346
rect 10501 9288 10506 9344
rect 10562 9288 11426 9344
rect 11482 9288 11487 9344
rect 10501 9286 11487 9288
rect 10133 9283 10199 9284
rect 10501 9283 10567 9286
rect 11421 9283 11487 9286
rect 13997 9346 14063 9349
rect 15540 9346 16000 9376
rect 13997 9344 16000 9346
rect 13997 9288 14002 9344
rect 14058 9288 16000 9344
rect 13997 9286 16000 9288
rect 13997 9283 14063 9286
rect 2625 9280 2941 9281
rect 2625 9216 2631 9280
rect 2695 9216 2711 9280
rect 2775 9216 2791 9280
rect 2855 9216 2871 9280
rect 2935 9216 2941 9280
rect 2625 9215 2941 9216
rect 5983 9280 6299 9281
rect 5983 9216 5989 9280
rect 6053 9216 6069 9280
rect 6133 9216 6149 9280
rect 6213 9216 6229 9280
rect 6293 9216 6299 9280
rect 5983 9215 6299 9216
rect 9341 9280 9657 9281
rect 9341 9216 9347 9280
rect 9411 9216 9427 9280
rect 9491 9216 9507 9280
rect 9571 9216 9587 9280
rect 9651 9216 9657 9280
rect 9341 9215 9657 9216
rect 12699 9280 13015 9281
rect 12699 9216 12705 9280
rect 12769 9216 12785 9280
rect 12849 9216 12865 9280
rect 12929 9216 12945 9280
rect 13009 9216 13015 9280
rect 15540 9256 16000 9286
rect 12699 9215 13015 9216
rect 11237 9074 11303 9077
rect 15540 9074 16000 9104
rect 11237 9072 16000 9074
rect 11237 9016 11242 9072
rect 11298 9016 16000 9072
rect 11237 9014 16000 9016
rect 11237 9011 11303 9014
rect 15540 8984 16000 9014
rect -300 8802 160 8832
rect 841 8802 907 8805
rect -300 8800 907 8802
rect -300 8744 846 8800
rect 902 8744 907 8800
rect -300 8742 907 8744
rect -300 8712 160 8742
rect 841 8739 907 8742
rect 8477 8802 8543 8805
rect 8886 8802 8892 8804
rect 8477 8800 8892 8802
rect 8477 8744 8482 8800
rect 8538 8744 8892 8800
rect 8477 8742 8892 8744
rect 8477 8739 8543 8742
rect 8886 8740 8892 8742
rect 8956 8740 8962 8804
rect 14825 8802 14891 8805
rect 15540 8802 16000 8832
rect 14825 8800 16000 8802
rect 14825 8744 14830 8800
rect 14886 8744 16000 8800
rect 14825 8742 16000 8744
rect 14825 8739 14891 8742
rect 4304 8736 4620 8737
rect 4304 8672 4310 8736
rect 4374 8672 4390 8736
rect 4454 8672 4470 8736
rect 4534 8672 4550 8736
rect 4614 8672 4620 8736
rect 4304 8671 4620 8672
rect 7662 8736 7978 8737
rect 7662 8672 7668 8736
rect 7732 8672 7748 8736
rect 7812 8672 7828 8736
rect 7892 8672 7908 8736
rect 7972 8672 7978 8736
rect 7662 8671 7978 8672
rect 11020 8736 11336 8737
rect 11020 8672 11026 8736
rect 11090 8672 11106 8736
rect 11170 8672 11186 8736
rect 11250 8672 11266 8736
rect 11330 8672 11336 8736
rect 11020 8671 11336 8672
rect 14378 8736 14694 8737
rect 14378 8672 14384 8736
rect 14448 8672 14464 8736
rect 14528 8672 14544 8736
rect 14608 8672 14624 8736
rect 14688 8672 14694 8736
rect 15540 8712 16000 8742
rect 14378 8671 14694 8672
rect 9857 8668 9923 8669
rect 9806 8604 9812 8668
rect 9876 8666 9923 8668
rect 9876 8664 9968 8666
rect 9918 8608 9968 8664
rect 9876 8606 9968 8608
rect 9876 8604 9923 8606
rect 9857 8603 9923 8604
rect 5901 8530 5967 8533
rect 11329 8530 11395 8533
rect 5901 8528 11395 8530
rect 5901 8472 5906 8528
rect 5962 8472 11334 8528
rect 11390 8472 11395 8528
rect 5901 8470 11395 8472
rect 5901 8467 5967 8470
rect 11329 8467 11395 8470
rect 14181 8530 14247 8533
rect 15540 8530 16000 8560
rect 14181 8528 16000 8530
rect 14181 8472 14186 8528
rect 14242 8472 16000 8528
rect 14181 8470 16000 8472
rect 14181 8467 14247 8470
rect 15540 8440 16000 8470
rect 1669 8258 1735 8261
rect 15540 8258 16000 8288
rect 798 8256 1735 8258
rect 798 8200 1674 8256
rect 1730 8200 1735 8256
rect 798 8198 1735 8200
rect -300 7986 160 8016
rect 798 7986 858 8198
rect 1669 8195 1735 8198
rect 14046 8198 16000 8258
rect 2625 8192 2941 8193
rect 2625 8128 2631 8192
rect 2695 8128 2711 8192
rect 2775 8128 2791 8192
rect 2855 8128 2871 8192
rect 2935 8128 2941 8192
rect 2625 8127 2941 8128
rect 5983 8192 6299 8193
rect 5983 8128 5989 8192
rect 6053 8128 6069 8192
rect 6133 8128 6149 8192
rect 6213 8128 6229 8192
rect 6293 8128 6299 8192
rect 5983 8127 6299 8128
rect 9341 8192 9657 8193
rect 9341 8128 9347 8192
rect 9411 8128 9427 8192
rect 9491 8128 9507 8192
rect 9571 8128 9587 8192
rect 9651 8128 9657 8192
rect 9341 8127 9657 8128
rect 12699 8192 13015 8193
rect 12699 8128 12705 8192
rect 12769 8128 12785 8192
rect 12849 8128 12865 8192
rect 12929 8128 12945 8192
rect 13009 8128 13015 8192
rect 12699 8127 13015 8128
rect 8017 8122 8083 8125
rect 8150 8122 8156 8124
rect 8017 8120 8156 8122
rect 8017 8064 8022 8120
rect 8078 8064 8156 8120
rect 8017 8062 8156 8064
rect 8017 8059 8083 8062
rect 8150 8060 8156 8062
rect 8220 8060 8226 8124
rect -300 7926 858 7986
rect 7097 7986 7163 7989
rect 9857 7986 9923 7989
rect 7097 7984 9923 7986
rect 7097 7928 7102 7984
rect 7158 7928 9862 7984
rect 9918 7928 9923 7984
rect 7097 7926 9923 7928
rect -300 7896 160 7926
rect 7097 7923 7163 7926
rect 9857 7923 9923 7926
rect 11237 7986 11303 7989
rect 14046 7986 14106 8198
rect 15540 8168 16000 8198
rect 15540 7986 16000 8016
rect 11237 7984 14106 7986
rect 11237 7928 11242 7984
rect 11298 7928 14106 7984
rect 11237 7926 14106 7928
rect 14230 7926 16000 7986
rect 11237 7923 11303 7926
rect 7189 7850 7255 7853
rect 7649 7850 7715 7853
rect 9673 7850 9739 7853
rect 7189 7848 9739 7850
rect 7189 7792 7194 7848
rect 7250 7792 7654 7848
rect 7710 7792 9678 7848
rect 9734 7792 9739 7848
rect 7189 7790 9739 7792
rect 7189 7787 7255 7790
rect 7649 7787 7715 7790
rect 9673 7787 9739 7790
rect 11145 7850 11211 7853
rect 14230 7850 14290 7926
rect 15540 7896 16000 7926
rect 11145 7848 14290 7850
rect 11145 7792 11150 7848
rect 11206 7792 14290 7848
rect 11145 7790 14290 7792
rect 11145 7787 11211 7790
rect 8886 7652 8892 7716
rect 8956 7714 8962 7716
rect 9489 7714 9555 7717
rect 10777 7714 10843 7717
rect 8956 7712 10843 7714
rect 8956 7656 9494 7712
rect 9550 7656 10782 7712
rect 10838 7656 10843 7712
rect 8956 7654 10843 7656
rect 8956 7652 8962 7654
rect 9489 7651 9555 7654
rect 10777 7651 10843 7654
rect 14825 7714 14891 7717
rect 15540 7714 16000 7744
rect 14825 7712 16000 7714
rect 14825 7656 14830 7712
rect 14886 7656 16000 7712
rect 14825 7654 16000 7656
rect 14825 7651 14891 7654
rect 4304 7648 4620 7649
rect 4304 7584 4310 7648
rect 4374 7584 4390 7648
rect 4454 7584 4470 7648
rect 4534 7584 4550 7648
rect 4614 7584 4620 7648
rect 4304 7583 4620 7584
rect 7662 7648 7978 7649
rect 7662 7584 7668 7648
rect 7732 7584 7748 7648
rect 7812 7584 7828 7648
rect 7892 7584 7908 7648
rect 7972 7584 7978 7648
rect 7662 7583 7978 7584
rect 11020 7648 11336 7649
rect 11020 7584 11026 7648
rect 11090 7584 11106 7648
rect 11170 7584 11186 7648
rect 11250 7584 11266 7648
rect 11330 7584 11336 7648
rect 11020 7583 11336 7584
rect 14378 7648 14694 7649
rect 14378 7584 14384 7648
rect 14448 7584 14464 7648
rect 14528 7584 14544 7648
rect 14608 7584 14624 7648
rect 14688 7584 14694 7648
rect 15540 7624 16000 7654
rect 14378 7583 14694 7584
rect 8109 7578 8175 7581
rect 9305 7578 9371 7581
rect 8109 7576 9371 7578
rect 8109 7520 8114 7576
rect 8170 7520 9310 7576
rect 9366 7520 9371 7576
rect 8109 7518 9371 7520
rect 8109 7515 8175 7518
rect 9305 7515 9371 7518
rect 9627 7474 9693 7479
rect 7281 7442 7347 7445
rect 9489 7442 9555 7445
rect 7281 7440 9555 7442
rect 7281 7384 7286 7440
rect 7342 7384 9494 7440
rect 9550 7384 9555 7440
rect 9627 7418 9632 7474
rect 9688 7418 9693 7474
rect 9627 7413 9693 7418
rect 9765 7442 9831 7445
rect 10777 7442 10843 7445
rect 9765 7440 10843 7442
rect 7281 7382 9555 7384
rect 7281 7379 7347 7382
rect 9489 7379 9555 7382
rect 9630 7309 9690 7413
rect 9765 7384 9770 7440
rect 9826 7384 10782 7440
rect 10838 7384 10843 7440
rect 9765 7382 10843 7384
rect 9765 7379 9831 7382
rect 10777 7379 10843 7382
rect 11697 7442 11763 7445
rect 15540 7442 16000 7472
rect 11697 7440 16000 7442
rect 11697 7384 11702 7440
rect 11758 7384 16000 7440
rect 11697 7382 16000 7384
rect 11697 7379 11763 7382
rect 15540 7352 16000 7382
rect 5165 7306 5231 7309
rect 5165 7304 9138 7306
rect 5165 7248 5170 7304
rect 5226 7248 9138 7304
rect 5165 7246 9138 7248
rect 9630 7304 9739 7309
rect 9630 7248 9678 7304
rect 9734 7248 9739 7304
rect 9630 7246 9739 7248
rect 5165 7243 5231 7246
rect -300 7170 160 7200
rect 841 7170 907 7173
rect -300 7168 907 7170
rect -300 7112 846 7168
rect 902 7112 907 7168
rect -300 7110 907 7112
rect -300 7080 160 7110
rect 841 7107 907 7110
rect 2625 7104 2941 7105
rect 2625 7040 2631 7104
rect 2695 7040 2711 7104
rect 2775 7040 2791 7104
rect 2855 7040 2871 7104
rect 2935 7040 2941 7104
rect 2625 7039 2941 7040
rect 5983 7104 6299 7105
rect 5983 7040 5989 7104
rect 6053 7040 6069 7104
rect 6133 7040 6149 7104
rect 6213 7040 6229 7104
rect 6293 7040 6299 7104
rect 5983 7039 6299 7040
rect 9078 6898 9138 7246
rect 9673 7243 9739 7246
rect 12065 7306 12131 7309
rect 12065 7304 14106 7306
rect 12065 7248 12070 7304
rect 12126 7248 14106 7304
rect 12065 7246 14106 7248
rect 12065 7243 12131 7246
rect 14046 7170 14106 7246
rect 15540 7170 16000 7200
rect 14046 7110 16000 7170
rect 9341 7104 9657 7105
rect 9341 7040 9347 7104
rect 9411 7040 9427 7104
rect 9491 7040 9507 7104
rect 9571 7040 9587 7104
rect 9651 7040 9657 7104
rect 9341 7039 9657 7040
rect 12699 7104 13015 7105
rect 12699 7040 12705 7104
rect 12769 7040 12785 7104
rect 12849 7040 12865 7104
rect 12929 7040 12945 7104
rect 13009 7040 13015 7104
rect 15540 7080 16000 7110
rect 12699 7039 13015 7040
rect 9765 7034 9831 7037
rect 9765 7032 12634 7034
rect 9765 6976 9770 7032
rect 9826 6976 12634 7032
rect 9765 6974 12634 6976
rect 9765 6971 9831 6974
rect 9305 6898 9371 6901
rect 9078 6896 9371 6898
rect 9078 6840 9310 6896
rect 9366 6840 9371 6896
rect 9078 6838 9371 6840
rect 12574 6898 12634 6974
rect 15540 6898 16000 6928
rect 12574 6838 16000 6898
rect 9305 6835 9371 6838
rect 15540 6808 16000 6838
rect 9765 6764 9831 6765
rect 9765 6760 9812 6764
rect 9876 6762 9882 6764
rect 11697 6762 11763 6765
rect 9765 6704 9770 6760
rect 9765 6700 9812 6704
rect 9876 6702 9922 6762
rect 11697 6760 14842 6762
rect 11697 6704 11702 6760
rect 11758 6704 14842 6760
rect 11697 6702 14842 6704
rect 9876 6700 9882 6702
rect 9765 6699 9831 6700
rect 11697 6699 11763 6702
rect 14782 6626 14842 6702
rect 15540 6626 16000 6656
rect 14782 6566 16000 6626
rect 4304 6560 4620 6561
rect 4304 6496 4310 6560
rect 4374 6496 4390 6560
rect 4454 6496 4470 6560
rect 4534 6496 4550 6560
rect 4614 6496 4620 6560
rect 4304 6495 4620 6496
rect 7662 6560 7978 6561
rect 7662 6496 7668 6560
rect 7732 6496 7748 6560
rect 7812 6496 7828 6560
rect 7892 6496 7908 6560
rect 7972 6496 7978 6560
rect 7662 6495 7978 6496
rect 11020 6560 11336 6561
rect 11020 6496 11026 6560
rect 11090 6496 11106 6560
rect 11170 6496 11186 6560
rect 11250 6496 11266 6560
rect 11330 6496 11336 6560
rect 11020 6495 11336 6496
rect 14378 6560 14694 6561
rect 14378 6496 14384 6560
rect 14448 6496 14464 6560
rect 14528 6496 14544 6560
rect 14608 6496 14624 6560
rect 14688 6496 14694 6560
rect 15540 6536 16000 6566
rect 14378 6495 14694 6496
rect 13445 6490 13511 6493
rect 12068 6488 13511 6490
rect 12068 6432 13450 6488
rect 13506 6432 13511 6488
rect 12068 6430 13511 6432
rect -300 6354 160 6384
rect 841 6354 907 6357
rect -300 6352 907 6354
rect -300 6296 846 6352
rect 902 6296 907 6352
rect -300 6294 907 6296
rect -300 6264 160 6294
rect 841 6291 907 6294
rect 10317 6354 10383 6357
rect 12068 6354 12128 6430
rect 13445 6427 13511 6430
rect 10317 6352 12128 6354
rect 10317 6296 10322 6352
rect 10378 6296 12128 6352
rect 10317 6294 12128 6296
rect 12249 6354 12315 6357
rect 15540 6354 16000 6384
rect 12249 6352 16000 6354
rect 12249 6296 12254 6352
rect 12310 6296 16000 6352
rect 12249 6294 16000 6296
rect 10317 6291 10383 6294
rect 12249 6291 12315 6294
rect 15540 6264 16000 6294
rect 8201 6220 8267 6221
rect 8150 6218 8156 6220
rect 8074 6158 8156 6218
rect 8220 6218 8267 6220
rect 12525 6218 12591 6221
rect 8220 6216 12591 6218
rect 8262 6160 12530 6216
rect 12586 6160 12591 6216
rect 8150 6156 8156 6158
rect 8220 6158 12591 6160
rect 8220 6156 8267 6158
rect 8201 6155 8267 6156
rect 12525 6155 12591 6158
rect 15540 6082 16000 6112
rect 14046 6022 16000 6082
rect 2625 6016 2941 6017
rect 2625 5952 2631 6016
rect 2695 5952 2711 6016
rect 2775 5952 2791 6016
rect 2855 5952 2871 6016
rect 2935 5952 2941 6016
rect 2625 5951 2941 5952
rect 5983 6016 6299 6017
rect 5983 5952 5989 6016
rect 6053 5952 6069 6016
rect 6133 5952 6149 6016
rect 6213 5952 6229 6016
rect 6293 5952 6299 6016
rect 5983 5951 6299 5952
rect 9341 6016 9657 6017
rect 9341 5952 9347 6016
rect 9411 5952 9427 6016
rect 9491 5952 9507 6016
rect 9571 5952 9587 6016
rect 9651 5952 9657 6016
rect 9341 5951 9657 5952
rect 12699 6016 13015 6017
rect 12699 5952 12705 6016
rect 12769 5952 12785 6016
rect 12849 5952 12865 6016
rect 12929 5952 12945 6016
rect 13009 5952 13015 6016
rect 12699 5951 13015 5952
rect 12341 5810 12407 5813
rect 14046 5810 14106 6022
rect 15540 5992 16000 6022
rect 15540 5810 16000 5840
rect 12341 5808 14106 5810
rect 12341 5752 12346 5808
rect 12402 5752 14106 5808
rect 12341 5750 14106 5752
rect 14598 5750 16000 5810
rect 12341 5747 12407 5750
rect 8293 5674 8359 5677
rect 12433 5674 12499 5677
rect 8293 5672 12499 5674
rect 8293 5616 8298 5672
rect 8354 5616 12438 5672
rect 12494 5616 12499 5672
rect 8293 5614 12499 5616
rect 8293 5611 8359 5614
rect 12433 5611 12499 5614
rect 13629 5674 13695 5677
rect 14598 5674 14658 5750
rect 15540 5720 16000 5750
rect 13629 5672 14658 5674
rect 13629 5616 13634 5672
rect 13690 5616 14658 5672
rect 13629 5614 14658 5616
rect 14825 5674 14891 5677
rect 14958 5674 14964 5676
rect 14825 5672 14964 5674
rect 14825 5616 14830 5672
rect 14886 5616 14964 5672
rect 14825 5614 14964 5616
rect 13629 5611 13695 5614
rect 14825 5611 14891 5614
rect 14958 5612 14964 5614
rect 15028 5612 15034 5676
rect -300 5538 160 5568
rect 1577 5538 1643 5541
rect 15540 5538 16000 5568
rect -300 5536 1643 5538
rect -300 5480 1582 5536
rect 1638 5480 1643 5536
rect -300 5478 1643 5480
rect -300 5448 160 5478
rect 1577 5475 1643 5478
rect 14782 5478 16000 5538
rect 4304 5472 4620 5473
rect 4304 5408 4310 5472
rect 4374 5408 4390 5472
rect 4454 5408 4470 5472
rect 4534 5408 4550 5472
rect 4614 5408 4620 5472
rect 4304 5407 4620 5408
rect 7662 5472 7978 5473
rect 7662 5408 7668 5472
rect 7732 5408 7748 5472
rect 7812 5408 7828 5472
rect 7892 5408 7908 5472
rect 7972 5408 7978 5472
rect 7662 5407 7978 5408
rect 11020 5472 11336 5473
rect 11020 5408 11026 5472
rect 11090 5408 11106 5472
rect 11170 5408 11186 5472
rect 11250 5408 11266 5472
rect 11330 5408 11336 5472
rect 11020 5407 11336 5408
rect 14378 5472 14694 5473
rect 14378 5408 14384 5472
rect 14448 5408 14464 5472
rect 14528 5408 14544 5472
rect 14608 5408 14624 5472
rect 14688 5408 14694 5472
rect 14378 5407 14694 5408
rect 13721 5266 13787 5269
rect 14782 5266 14842 5478
rect 15540 5448 16000 5478
rect 15540 5266 16000 5296
rect 13721 5264 14842 5266
rect 13721 5208 13726 5264
rect 13782 5208 14842 5264
rect 13721 5206 14842 5208
rect 14920 5206 16000 5266
rect 13721 5203 13787 5206
rect 11973 5130 12039 5133
rect 14920 5130 14980 5206
rect 15540 5176 16000 5206
rect 11973 5128 14980 5130
rect 11973 5072 11978 5128
rect 12034 5072 14980 5128
rect 11973 5070 14980 5072
rect 11973 5067 12039 5070
rect 13905 4994 13971 4997
rect 15540 4994 16000 5024
rect 13905 4992 16000 4994
rect 13905 4936 13910 4992
rect 13966 4936 16000 4992
rect 13905 4934 16000 4936
rect 13905 4931 13971 4934
rect 2625 4928 2941 4929
rect 2625 4864 2631 4928
rect 2695 4864 2711 4928
rect 2775 4864 2791 4928
rect 2855 4864 2871 4928
rect 2935 4864 2941 4928
rect 2625 4863 2941 4864
rect 5983 4928 6299 4929
rect 5983 4864 5989 4928
rect 6053 4864 6069 4928
rect 6133 4864 6149 4928
rect 6213 4864 6229 4928
rect 6293 4864 6299 4928
rect 5983 4863 6299 4864
rect 9341 4928 9657 4929
rect 9341 4864 9347 4928
rect 9411 4864 9427 4928
rect 9491 4864 9507 4928
rect 9571 4864 9587 4928
rect 9651 4864 9657 4928
rect 9341 4863 9657 4864
rect 12699 4928 13015 4929
rect 12699 4864 12705 4928
rect 12769 4864 12785 4928
rect 12849 4864 12865 4928
rect 12929 4864 12945 4928
rect 13009 4864 13015 4928
rect 15540 4904 16000 4934
rect 12699 4863 13015 4864
rect -300 4722 160 4752
rect 841 4722 907 4725
rect -300 4720 907 4722
rect -300 4664 846 4720
rect 902 4664 907 4720
rect -300 4662 907 4664
rect -300 4632 160 4662
rect 841 4659 907 4662
rect 4304 4384 4620 4385
rect 4304 4320 4310 4384
rect 4374 4320 4390 4384
rect 4454 4320 4470 4384
rect 4534 4320 4550 4384
rect 4614 4320 4620 4384
rect 4304 4319 4620 4320
rect 7662 4384 7978 4385
rect 7662 4320 7668 4384
rect 7732 4320 7748 4384
rect 7812 4320 7828 4384
rect 7892 4320 7908 4384
rect 7972 4320 7978 4384
rect 7662 4319 7978 4320
rect 11020 4384 11336 4385
rect 11020 4320 11026 4384
rect 11090 4320 11106 4384
rect 11170 4320 11186 4384
rect 11250 4320 11266 4384
rect 11330 4320 11336 4384
rect 11020 4319 11336 4320
rect 14378 4384 14694 4385
rect 14378 4320 14384 4384
rect 14448 4320 14464 4384
rect 14528 4320 14544 4384
rect 14608 4320 14624 4384
rect 14688 4320 14694 4384
rect 14378 4319 14694 4320
rect -300 3906 160 3936
rect 749 3906 815 3909
rect -300 3904 815 3906
rect -300 3848 754 3904
rect 810 3848 815 3904
rect -300 3846 815 3848
rect -300 3816 160 3846
rect 749 3843 815 3846
rect 2625 3840 2941 3841
rect 2625 3776 2631 3840
rect 2695 3776 2711 3840
rect 2775 3776 2791 3840
rect 2855 3776 2871 3840
rect 2935 3776 2941 3840
rect 2625 3775 2941 3776
rect 5983 3840 6299 3841
rect 5983 3776 5989 3840
rect 6053 3776 6069 3840
rect 6133 3776 6149 3840
rect 6213 3776 6229 3840
rect 6293 3776 6299 3840
rect 5983 3775 6299 3776
rect 9341 3840 9657 3841
rect 9341 3776 9347 3840
rect 9411 3776 9427 3840
rect 9491 3776 9507 3840
rect 9571 3776 9587 3840
rect 9651 3776 9657 3840
rect 9341 3775 9657 3776
rect 12699 3840 13015 3841
rect 12699 3776 12705 3840
rect 12769 3776 12785 3840
rect 12849 3776 12865 3840
rect 12929 3776 12945 3840
rect 13009 3776 13015 3840
rect 12699 3775 13015 3776
rect 4304 3296 4620 3297
rect 4304 3232 4310 3296
rect 4374 3232 4390 3296
rect 4454 3232 4470 3296
rect 4534 3232 4550 3296
rect 4614 3232 4620 3296
rect 4304 3231 4620 3232
rect 7662 3296 7978 3297
rect 7662 3232 7668 3296
rect 7732 3232 7748 3296
rect 7812 3232 7828 3296
rect 7892 3232 7908 3296
rect 7972 3232 7978 3296
rect 7662 3231 7978 3232
rect 11020 3296 11336 3297
rect 11020 3232 11026 3296
rect 11090 3232 11106 3296
rect 11170 3232 11186 3296
rect 11250 3232 11266 3296
rect 11330 3232 11336 3296
rect 11020 3231 11336 3232
rect 14378 3296 14694 3297
rect 14378 3232 14384 3296
rect 14448 3232 14464 3296
rect 14528 3232 14544 3296
rect 14608 3232 14624 3296
rect 14688 3232 14694 3296
rect 14378 3231 14694 3232
rect 2625 2752 2941 2753
rect 2625 2688 2631 2752
rect 2695 2688 2711 2752
rect 2775 2688 2791 2752
rect 2855 2688 2871 2752
rect 2935 2688 2941 2752
rect 2625 2687 2941 2688
rect 5983 2752 6299 2753
rect 5983 2688 5989 2752
rect 6053 2688 6069 2752
rect 6133 2688 6149 2752
rect 6213 2688 6229 2752
rect 6293 2688 6299 2752
rect 5983 2687 6299 2688
rect 9341 2752 9657 2753
rect 9341 2688 9347 2752
rect 9411 2688 9427 2752
rect 9491 2688 9507 2752
rect 9571 2688 9587 2752
rect 9651 2688 9657 2752
rect 9341 2687 9657 2688
rect 12699 2752 13015 2753
rect 12699 2688 12705 2752
rect 12769 2688 12785 2752
rect 12849 2688 12865 2752
rect 12929 2688 12945 2752
rect 13009 2688 13015 2752
rect 12699 2687 13015 2688
rect 6637 2684 6703 2685
rect 6637 2682 6684 2684
rect 6592 2680 6684 2682
rect 6592 2624 6642 2680
rect 6592 2622 6684 2624
rect 6637 2620 6684 2622
rect 6748 2620 6754 2684
rect 10358 2620 10364 2684
rect 10428 2682 10434 2684
rect 10869 2682 10935 2685
rect 10428 2680 10935 2682
rect 10428 2624 10874 2680
rect 10930 2624 10935 2680
rect 10428 2622 10935 2624
rect 10428 2620 10434 2622
rect 6637 2619 6703 2620
rect 10869 2619 10935 2622
rect 2078 2484 2084 2548
rect 2148 2546 2154 2548
rect 7189 2546 7255 2549
rect 2148 2544 7255 2546
rect 2148 2488 7194 2544
rect 7250 2488 7255 2544
rect 2148 2486 7255 2488
rect 2148 2484 2154 2486
rect 7189 2483 7255 2486
rect 9070 2484 9076 2548
rect 9140 2546 9146 2548
rect 9397 2546 9463 2549
rect 9140 2544 9463 2546
rect 9140 2488 9402 2544
rect 9458 2488 9463 2544
rect 9140 2486 9463 2488
rect 9140 2484 9146 2486
rect 9397 2483 9463 2486
rect 2262 2348 2268 2412
rect 2332 2410 2338 2412
rect 8661 2410 8727 2413
rect 2332 2408 8727 2410
rect 2332 2352 8666 2408
rect 8722 2352 8727 2408
rect 2332 2350 8727 2352
rect 2332 2348 2338 2350
rect 8661 2347 8727 2350
rect 4304 2208 4620 2209
rect 4304 2144 4310 2208
rect 4374 2144 4390 2208
rect 4454 2144 4470 2208
rect 4534 2144 4550 2208
rect 4614 2144 4620 2208
rect 4304 2143 4620 2144
rect 7662 2208 7978 2209
rect 7662 2144 7668 2208
rect 7732 2144 7748 2208
rect 7812 2144 7828 2208
rect 7892 2144 7908 2208
rect 7972 2144 7978 2208
rect 7662 2143 7978 2144
rect 11020 2208 11336 2209
rect 11020 2144 11026 2208
rect 11090 2144 11106 2208
rect 11170 2144 11186 2208
rect 11250 2144 11266 2208
rect 11330 2144 11336 2208
rect 11020 2143 11336 2144
rect 14378 2208 14694 2209
rect 14378 2144 14384 2208
rect 14448 2144 14464 2208
rect 14528 2144 14544 2208
rect 14608 2144 14624 2208
rect 14688 2144 14694 2208
rect 14378 2143 14694 2144
rect 3918 1940 3924 2004
rect 3988 2002 3994 2004
rect 10133 2002 10199 2005
rect 3988 2000 10199 2002
rect 3988 1944 10138 2000
rect 10194 1944 10199 2000
rect 3988 1942 10199 1944
rect 3988 1940 3994 1942
rect 10133 1939 10199 1942
rect 2625 1664 2941 1665
rect 2625 1600 2631 1664
rect 2695 1600 2711 1664
rect 2775 1600 2791 1664
rect 2855 1600 2871 1664
rect 2935 1600 2941 1664
rect 2625 1599 2941 1600
rect 5983 1664 6299 1665
rect 5983 1600 5989 1664
rect 6053 1600 6069 1664
rect 6133 1600 6149 1664
rect 6213 1600 6229 1664
rect 6293 1600 6299 1664
rect 5983 1599 6299 1600
rect 9341 1664 9657 1665
rect 9341 1600 9347 1664
rect 9411 1600 9427 1664
rect 9491 1600 9507 1664
rect 9571 1600 9587 1664
rect 9651 1600 9657 1664
rect 9341 1599 9657 1600
rect 12699 1664 13015 1665
rect 12699 1600 12705 1664
rect 12769 1600 12785 1664
rect 12849 1600 12865 1664
rect 12929 1600 12945 1664
rect 13009 1600 13015 1664
rect 12699 1599 13015 1600
rect 4613 1322 4679 1325
rect 5165 1324 5231 1325
rect 4838 1322 4844 1324
rect 4613 1320 4844 1322
rect 4613 1264 4618 1320
rect 4674 1264 4844 1320
rect 4613 1262 4844 1264
rect 4613 1259 4679 1262
rect 4838 1260 4844 1262
rect 4908 1260 4914 1324
rect 5165 1322 5212 1324
rect 5120 1320 5212 1322
rect 5120 1264 5170 1320
rect 5120 1262 5212 1264
rect 5165 1260 5212 1262
rect 5276 1260 5282 1324
rect 6494 1260 6500 1324
rect 6564 1322 6570 1324
rect 6637 1322 6703 1325
rect 6564 1320 6703 1322
rect 6564 1264 6642 1320
rect 6698 1264 6703 1320
rect 6564 1262 6703 1264
rect 6564 1260 6570 1262
rect 5165 1259 5231 1260
rect 6637 1259 6703 1262
rect 8702 1260 8708 1324
rect 8772 1322 8778 1324
rect 13813 1322 13879 1325
rect 8772 1320 13879 1322
rect 8772 1264 13818 1320
rect 13874 1264 13879 1320
rect 8772 1262 13879 1264
rect 8772 1260 8778 1262
rect 13813 1259 13879 1262
rect 4304 1120 4620 1121
rect 4304 1056 4310 1120
rect 4374 1056 4390 1120
rect 4454 1056 4470 1120
rect 4534 1056 4550 1120
rect 4614 1056 4620 1120
rect 4304 1055 4620 1056
rect 7662 1120 7978 1121
rect 7662 1056 7668 1120
rect 7732 1056 7748 1120
rect 7812 1056 7828 1120
rect 7892 1056 7908 1120
rect 7972 1056 7978 1120
rect 7662 1055 7978 1056
rect 11020 1120 11336 1121
rect 11020 1056 11026 1120
rect 11090 1056 11106 1120
rect 11170 1056 11186 1120
rect 11250 1056 11266 1120
rect 11330 1056 11336 1120
rect 11020 1055 11336 1056
rect 14378 1120 14694 1121
rect 14378 1056 14384 1120
rect 14448 1056 14464 1120
rect 14528 1056 14544 1120
rect 14608 1056 14624 1120
rect 14688 1056 14694 1120
rect 14378 1055 14694 1056
<< via3 >>
rect 4310 43548 4374 43552
rect 4310 43492 4314 43548
rect 4314 43492 4370 43548
rect 4370 43492 4374 43548
rect 4310 43488 4374 43492
rect 4390 43548 4454 43552
rect 4390 43492 4394 43548
rect 4394 43492 4450 43548
rect 4450 43492 4454 43548
rect 4390 43488 4454 43492
rect 4470 43548 4534 43552
rect 4470 43492 4474 43548
rect 4474 43492 4530 43548
rect 4530 43492 4534 43548
rect 4470 43488 4534 43492
rect 4550 43548 4614 43552
rect 4550 43492 4554 43548
rect 4554 43492 4610 43548
rect 4610 43492 4614 43548
rect 4550 43488 4614 43492
rect 7668 43548 7732 43552
rect 7668 43492 7672 43548
rect 7672 43492 7728 43548
rect 7728 43492 7732 43548
rect 7668 43488 7732 43492
rect 7748 43548 7812 43552
rect 7748 43492 7752 43548
rect 7752 43492 7808 43548
rect 7808 43492 7812 43548
rect 7748 43488 7812 43492
rect 7828 43548 7892 43552
rect 7828 43492 7832 43548
rect 7832 43492 7888 43548
rect 7888 43492 7892 43548
rect 7828 43488 7892 43492
rect 7908 43548 7972 43552
rect 7908 43492 7912 43548
rect 7912 43492 7968 43548
rect 7968 43492 7972 43548
rect 7908 43488 7972 43492
rect 11026 43548 11090 43552
rect 11026 43492 11030 43548
rect 11030 43492 11086 43548
rect 11086 43492 11090 43548
rect 11026 43488 11090 43492
rect 11106 43548 11170 43552
rect 11106 43492 11110 43548
rect 11110 43492 11166 43548
rect 11166 43492 11170 43548
rect 11106 43488 11170 43492
rect 11186 43548 11250 43552
rect 11186 43492 11190 43548
rect 11190 43492 11246 43548
rect 11246 43492 11250 43548
rect 11186 43488 11250 43492
rect 11266 43548 11330 43552
rect 11266 43492 11270 43548
rect 11270 43492 11326 43548
rect 11326 43492 11330 43548
rect 11266 43488 11330 43492
rect 14384 43548 14448 43552
rect 14384 43492 14388 43548
rect 14388 43492 14444 43548
rect 14444 43492 14448 43548
rect 14384 43488 14448 43492
rect 14464 43548 14528 43552
rect 14464 43492 14468 43548
rect 14468 43492 14524 43548
rect 14524 43492 14528 43548
rect 14464 43488 14528 43492
rect 14544 43548 14608 43552
rect 14544 43492 14548 43548
rect 14548 43492 14604 43548
rect 14604 43492 14608 43548
rect 14544 43488 14608 43492
rect 14624 43548 14688 43552
rect 14624 43492 14628 43548
rect 14628 43492 14684 43548
rect 14684 43492 14688 43548
rect 14624 43488 14688 43492
rect 2631 43004 2695 43008
rect 2631 42948 2635 43004
rect 2635 42948 2691 43004
rect 2691 42948 2695 43004
rect 2631 42944 2695 42948
rect 2711 43004 2775 43008
rect 2711 42948 2715 43004
rect 2715 42948 2771 43004
rect 2771 42948 2775 43004
rect 2711 42944 2775 42948
rect 2791 43004 2855 43008
rect 2791 42948 2795 43004
rect 2795 42948 2851 43004
rect 2851 42948 2855 43004
rect 2791 42944 2855 42948
rect 2871 43004 2935 43008
rect 2871 42948 2875 43004
rect 2875 42948 2931 43004
rect 2931 42948 2935 43004
rect 2871 42944 2935 42948
rect 5989 43004 6053 43008
rect 5989 42948 5993 43004
rect 5993 42948 6049 43004
rect 6049 42948 6053 43004
rect 5989 42944 6053 42948
rect 6069 43004 6133 43008
rect 6069 42948 6073 43004
rect 6073 42948 6129 43004
rect 6129 42948 6133 43004
rect 6069 42944 6133 42948
rect 6149 43004 6213 43008
rect 6149 42948 6153 43004
rect 6153 42948 6209 43004
rect 6209 42948 6213 43004
rect 6149 42944 6213 42948
rect 6229 43004 6293 43008
rect 6229 42948 6233 43004
rect 6233 42948 6289 43004
rect 6289 42948 6293 43004
rect 6229 42944 6293 42948
rect 9347 43004 9411 43008
rect 9347 42948 9351 43004
rect 9351 42948 9407 43004
rect 9407 42948 9411 43004
rect 9347 42944 9411 42948
rect 9427 43004 9491 43008
rect 9427 42948 9431 43004
rect 9431 42948 9487 43004
rect 9487 42948 9491 43004
rect 9427 42944 9491 42948
rect 9507 43004 9571 43008
rect 9507 42948 9511 43004
rect 9511 42948 9567 43004
rect 9567 42948 9571 43004
rect 9507 42944 9571 42948
rect 9587 43004 9651 43008
rect 9587 42948 9591 43004
rect 9591 42948 9647 43004
rect 9647 42948 9651 43004
rect 9587 42944 9651 42948
rect 12705 43004 12769 43008
rect 12705 42948 12709 43004
rect 12709 42948 12765 43004
rect 12765 42948 12769 43004
rect 12705 42944 12769 42948
rect 12785 43004 12849 43008
rect 12785 42948 12789 43004
rect 12789 42948 12845 43004
rect 12845 42948 12849 43004
rect 12785 42944 12849 42948
rect 12865 43004 12929 43008
rect 12865 42948 12869 43004
rect 12869 42948 12925 43004
rect 12925 42948 12929 43004
rect 12865 42944 12929 42948
rect 12945 43004 13009 43008
rect 12945 42948 12949 43004
rect 12949 42948 13005 43004
rect 13005 42948 13009 43004
rect 12945 42944 13009 42948
rect 3924 42740 3988 42804
rect 3740 42604 3804 42668
rect 4310 42460 4374 42464
rect 4310 42404 4314 42460
rect 4314 42404 4370 42460
rect 4370 42404 4374 42460
rect 4310 42400 4374 42404
rect 4390 42460 4454 42464
rect 4390 42404 4394 42460
rect 4394 42404 4450 42460
rect 4450 42404 4454 42460
rect 4390 42400 4454 42404
rect 4470 42460 4534 42464
rect 4470 42404 4474 42460
rect 4474 42404 4530 42460
rect 4530 42404 4534 42460
rect 4470 42400 4534 42404
rect 4550 42460 4614 42464
rect 4550 42404 4554 42460
rect 4554 42404 4610 42460
rect 4610 42404 4614 42460
rect 4550 42400 4614 42404
rect 7668 42460 7732 42464
rect 7668 42404 7672 42460
rect 7672 42404 7728 42460
rect 7728 42404 7732 42460
rect 7668 42400 7732 42404
rect 7748 42460 7812 42464
rect 7748 42404 7752 42460
rect 7752 42404 7808 42460
rect 7808 42404 7812 42460
rect 7748 42400 7812 42404
rect 7828 42460 7892 42464
rect 7828 42404 7832 42460
rect 7832 42404 7888 42460
rect 7888 42404 7892 42460
rect 7828 42400 7892 42404
rect 7908 42460 7972 42464
rect 7908 42404 7912 42460
rect 7912 42404 7968 42460
rect 7968 42404 7972 42460
rect 7908 42400 7972 42404
rect 11026 42460 11090 42464
rect 11026 42404 11030 42460
rect 11030 42404 11086 42460
rect 11086 42404 11090 42460
rect 11026 42400 11090 42404
rect 11106 42460 11170 42464
rect 11106 42404 11110 42460
rect 11110 42404 11166 42460
rect 11166 42404 11170 42460
rect 11106 42400 11170 42404
rect 11186 42460 11250 42464
rect 11186 42404 11190 42460
rect 11190 42404 11246 42460
rect 11246 42404 11250 42460
rect 11186 42400 11250 42404
rect 11266 42460 11330 42464
rect 11266 42404 11270 42460
rect 11270 42404 11326 42460
rect 11326 42404 11330 42460
rect 11266 42400 11330 42404
rect 14384 42460 14448 42464
rect 14384 42404 14388 42460
rect 14388 42404 14444 42460
rect 14444 42404 14448 42460
rect 14384 42400 14448 42404
rect 14464 42460 14528 42464
rect 14464 42404 14468 42460
rect 14468 42404 14524 42460
rect 14524 42404 14528 42460
rect 14464 42400 14528 42404
rect 14544 42460 14608 42464
rect 14544 42404 14548 42460
rect 14548 42404 14604 42460
rect 14604 42404 14608 42460
rect 14544 42400 14608 42404
rect 14624 42460 14688 42464
rect 14624 42404 14628 42460
rect 14628 42404 14684 42460
rect 14684 42404 14688 42460
rect 14624 42400 14688 42404
rect 2268 42060 2332 42124
rect 2631 41916 2695 41920
rect 2631 41860 2635 41916
rect 2635 41860 2691 41916
rect 2691 41860 2695 41916
rect 2631 41856 2695 41860
rect 2711 41916 2775 41920
rect 2711 41860 2715 41916
rect 2715 41860 2771 41916
rect 2771 41860 2775 41916
rect 2711 41856 2775 41860
rect 2791 41916 2855 41920
rect 2791 41860 2795 41916
rect 2795 41860 2851 41916
rect 2851 41860 2855 41916
rect 2791 41856 2855 41860
rect 2871 41916 2935 41920
rect 2871 41860 2875 41916
rect 2875 41860 2931 41916
rect 2931 41860 2935 41916
rect 2871 41856 2935 41860
rect 5989 41916 6053 41920
rect 5989 41860 5993 41916
rect 5993 41860 6049 41916
rect 6049 41860 6053 41916
rect 5989 41856 6053 41860
rect 6069 41916 6133 41920
rect 6069 41860 6073 41916
rect 6073 41860 6129 41916
rect 6129 41860 6133 41916
rect 6069 41856 6133 41860
rect 6149 41916 6213 41920
rect 6149 41860 6153 41916
rect 6153 41860 6209 41916
rect 6209 41860 6213 41916
rect 6149 41856 6213 41860
rect 6229 41916 6293 41920
rect 6229 41860 6233 41916
rect 6233 41860 6289 41916
rect 6289 41860 6293 41916
rect 6229 41856 6293 41860
rect 9347 41916 9411 41920
rect 9347 41860 9351 41916
rect 9351 41860 9407 41916
rect 9407 41860 9411 41916
rect 9347 41856 9411 41860
rect 9427 41916 9491 41920
rect 9427 41860 9431 41916
rect 9431 41860 9487 41916
rect 9487 41860 9491 41916
rect 9427 41856 9491 41860
rect 9507 41916 9571 41920
rect 9507 41860 9511 41916
rect 9511 41860 9567 41916
rect 9567 41860 9571 41916
rect 9507 41856 9571 41860
rect 9587 41916 9651 41920
rect 9587 41860 9591 41916
rect 9591 41860 9647 41916
rect 9647 41860 9651 41916
rect 9587 41856 9651 41860
rect 12705 41916 12769 41920
rect 12705 41860 12709 41916
rect 12709 41860 12765 41916
rect 12765 41860 12769 41916
rect 12705 41856 12769 41860
rect 12785 41916 12849 41920
rect 12785 41860 12789 41916
rect 12789 41860 12845 41916
rect 12845 41860 12849 41916
rect 12785 41856 12849 41860
rect 12865 41916 12929 41920
rect 12865 41860 12869 41916
rect 12869 41860 12925 41916
rect 12925 41860 12929 41916
rect 12865 41856 12929 41860
rect 12945 41916 13009 41920
rect 12945 41860 12949 41916
rect 12949 41860 13005 41916
rect 13005 41860 13009 41916
rect 12945 41856 13009 41860
rect 2084 41652 2148 41716
rect 4844 41516 4908 41580
rect 14964 41516 15028 41580
rect 1532 41380 1596 41444
rect 5212 41380 5276 41444
rect 6684 41380 6748 41444
rect 4310 41372 4374 41376
rect 4310 41316 4314 41372
rect 4314 41316 4370 41372
rect 4370 41316 4374 41372
rect 4310 41312 4374 41316
rect 4390 41372 4454 41376
rect 4390 41316 4394 41372
rect 4394 41316 4450 41372
rect 4450 41316 4454 41372
rect 4390 41312 4454 41316
rect 4470 41372 4534 41376
rect 4470 41316 4474 41372
rect 4474 41316 4530 41372
rect 4530 41316 4534 41372
rect 4470 41312 4534 41316
rect 4550 41372 4614 41376
rect 4550 41316 4554 41372
rect 4554 41316 4610 41372
rect 4610 41316 4614 41372
rect 4550 41312 4614 41316
rect 7668 41372 7732 41376
rect 7668 41316 7672 41372
rect 7672 41316 7728 41372
rect 7728 41316 7732 41372
rect 7668 41312 7732 41316
rect 7748 41372 7812 41376
rect 7748 41316 7752 41372
rect 7752 41316 7808 41372
rect 7808 41316 7812 41372
rect 7748 41312 7812 41316
rect 7828 41372 7892 41376
rect 7828 41316 7832 41372
rect 7832 41316 7888 41372
rect 7888 41316 7892 41372
rect 7828 41312 7892 41316
rect 7908 41372 7972 41376
rect 7908 41316 7912 41372
rect 7912 41316 7968 41372
rect 7968 41316 7972 41372
rect 7908 41312 7972 41316
rect 11026 41372 11090 41376
rect 11026 41316 11030 41372
rect 11030 41316 11086 41372
rect 11086 41316 11090 41372
rect 11026 41312 11090 41316
rect 11106 41372 11170 41376
rect 11106 41316 11110 41372
rect 11110 41316 11166 41372
rect 11166 41316 11170 41372
rect 11106 41312 11170 41316
rect 11186 41372 11250 41376
rect 11186 41316 11190 41372
rect 11190 41316 11246 41372
rect 11246 41316 11250 41372
rect 11186 41312 11250 41316
rect 11266 41372 11330 41376
rect 11266 41316 11270 41372
rect 11270 41316 11326 41372
rect 11326 41316 11330 41372
rect 11266 41312 11330 41316
rect 14384 41372 14448 41376
rect 14384 41316 14388 41372
rect 14388 41316 14444 41372
rect 14444 41316 14448 41372
rect 14384 41312 14448 41316
rect 14464 41372 14528 41376
rect 14464 41316 14468 41372
rect 14468 41316 14524 41372
rect 14524 41316 14528 41372
rect 14464 41312 14528 41316
rect 14544 41372 14608 41376
rect 14544 41316 14548 41372
rect 14548 41316 14604 41372
rect 14604 41316 14608 41372
rect 14544 41312 14608 41316
rect 14624 41372 14688 41376
rect 14624 41316 14628 41372
rect 14628 41316 14684 41372
rect 14684 41316 14688 41372
rect 14624 41312 14688 41316
rect 2631 40828 2695 40832
rect 2631 40772 2635 40828
rect 2635 40772 2691 40828
rect 2691 40772 2695 40828
rect 2631 40768 2695 40772
rect 2711 40828 2775 40832
rect 2711 40772 2715 40828
rect 2715 40772 2771 40828
rect 2771 40772 2775 40828
rect 2711 40768 2775 40772
rect 2791 40828 2855 40832
rect 2791 40772 2795 40828
rect 2795 40772 2851 40828
rect 2851 40772 2855 40828
rect 2791 40768 2855 40772
rect 2871 40828 2935 40832
rect 2871 40772 2875 40828
rect 2875 40772 2931 40828
rect 2931 40772 2935 40828
rect 2871 40768 2935 40772
rect 5989 40828 6053 40832
rect 5989 40772 5993 40828
rect 5993 40772 6049 40828
rect 6049 40772 6053 40828
rect 5989 40768 6053 40772
rect 6069 40828 6133 40832
rect 6069 40772 6073 40828
rect 6073 40772 6129 40828
rect 6129 40772 6133 40828
rect 6069 40768 6133 40772
rect 6149 40828 6213 40832
rect 6149 40772 6153 40828
rect 6153 40772 6209 40828
rect 6209 40772 6213 40828
rect 6149 40768 6213 40772
rect 6229 40828 6293 40832
rect 6229 40772 6233 40828
rect 6233 40772 6289 40828
rect 6289 40772 6293 40828
rect 6229 40768 6293 40772
rect 9347 40828 9411 40832
rect 9347 40772 9351 40828
rect 9351 40772 9407 40828
rect 9407 40772 9411 40828
rect 9347 40768 9411 40772
rect 9427 40828 9491 40832
rect 9427 40772 9431 40828
rect 9431 40772 9487 40828
rect 9487 40772 9491 40828
rect 9427 40768 9491 40772
rect 9507 40828 9571 40832
rect 9507 40772 9511 40828
rect 9511 40772 9567 40828
rect 9567 40772 9571 40828
rect 9507 40768 9571 40772
rect 9587 40828 9651 40832
rect 9587 40772 9591 40828
rect 9591 40772 9647 40828
rect 9647 40772 9651 40828
rect 9587 40768 9651 40772
rect 12705 40828 12769 40832
rect 12705 40772 12709 40828
rect 12709 40772 12765 40828
rect 12765 40772 12769 40828
rect 12705 40768 12769 40772
rect 12785 40828 12849 40832
rect 12785 40772 12789 40828
rect 12789 40772 12845 40828
rect 12845 40772 12849 40828
rect 12785 40768 12849 40772
rect 12865 40828 12929 40832
rect 12865 40772 12869 40828
rect 12869 40772 12925 40828
rect 12925 40772 12929 40828
rect 12865 40768 12929 40772
rect 12945 40828 13009 40832
rect 12945 40772 12949 40828
rect 12949 40772 13005 40828
rect 13005 40772 13009 40828
rect 12945 40768 13009 40772
rect 4310 40284 4374 40288
rect 4310 40228 4314 40284
rect 4314 40228 4370 40284
rect 4370 40228 4374 40284
rect 4310 40224 4374 40228
rect 4390 40284 4454 40288
rect 4390 40228 4394 40284
rect 4394 40228 4450 40284
rect 4450 40228 4454 40284
rect 4390 40224 4454 40228
rect 4470 40284 4534 40288
rect 4470 40228 4474 40284
rect 4474 40228 4530 40284
rect 4530 40228 4534 40284
rect 4470 40224 4534 40228
rect 4550 40284 4614 40288
rect 4550 40228 4554 40284
rect 4554 40228 4610 40284
rect 4610 40228 4614 40284
rect 4550 40224 4614 40228
rect 7668 40284 7732 40288
rect 7668 40228 7672 40284
rect 7672 40228 7728 40284
rect 7728 40228 7732 40284
rect 7668 40224 7732 40228
rect 7748 40284 7812 40288
rect 7748 40228 7752 40284
rect 7752 40228 7808 40284
rect 7808 40228 7812 40284
rect 7748 40224 7812 40228
rect 7828 40284 7892 40288
rect 7828 40228 7832 40284
rect 7832 40228 7888 40284
rect 7888 40228 7892 40284
rect 7828 40224 7892 40228
rect 7908 40284 7972 40288
rect 7908 40228 7912 40284
rect 7912 40228 7968 40284
rect 7968 40228 7972 40284
rect 7908 40224 7972 40228
rect 11026 40284 11090 40288
rect 11026 40228 11030 40284
rect 11030 40228 11086 40284
rect 11086 40228 11090 40284
rect 11026 40224 11090 40228
rect 11106 40284 11170 40288
rect 11106 40228 11110 40284
rect 11110 40228 11166 40284
rect 11166 40228 11170 40284
rect 11106 40224 11170 40228
rect 11186 40284 11250 40288
rect 11186 40228 11190 40284
rect 11190 40228 11246 40284
rect 11246 40228 11250 40284
rect 11186 40224 11250 40228
rect 11266 40284 11330 40288
rect 11266 40228 11270 40284
rect 11270 40228 11326 40284
rect 11326 40228 11330 40284
rect 11266 40224 11330 40228
rect 14384 40284 14448 40288
rect 14384 40228 14388 40284
rect 14388 40228 14444 40284
rect 14444 40228 14448 40284
rect 14384 40224 14448 40228
rect 14464 40284 14528 40288
rect 14464 40228 14468 40284
rect 14468 40228 14524 40284
rect 14524 40228 14528 40284
rect 14464 40224 14528 40228
rect 14544 40284 14608 40288
rect 14544 40228 14548 40284
rect 14548 40228 14604 40284
rect 14604 40228 14608 40284
rect 14544 40224 14608 40228
rect 14624 40284 14688 40288
rect 14624 40228 14628 40284
rect 14628 40228 14684 40284
rect 14684 40228 14688 40284
rect 14624 40224 14688 40228
rect 2631 39740 2695 39744
rect 2631 39684 2635 39740
rect 2635 39684 2691 39740
rect 2691 39684 2695 39740
rect 2631 39680 2695 39684
rect 2711 39740 2775 39744
rect 2711 39684 2715 39740
rect 2715 39684 2771 39740
rect 2771 39684 2775 39740
rect 2711 39680 2775 39684
rect 2791 39740 2855 39744
rect 2791 39684 2795 39740
rect 2795 39684 2851 39740
rect 2851 39684 2855 39740
rect 2791 39680 2855 39684
rect 2871 39740 2935 39744
rect 2871 39684 2875 39740
rect 2875 39684 2931 39740
rect 2931 39684 2935 39740
rect 2871 39680 2935 39684
rect 5989 39740 6053 39744
rect 5989 39684 5993 39740
rect 5993 39684 6049 39740
rect 6049 39684 6053 39740
rect 5989 39680 6053 39684
rect 6069 39740 6133 39744
rect 6069 39684 6073 39740
rect 6073 39684 6129 39740
rect 6129 39684 6133 39740
rect 6069 39680 6133 39684
rect 6149 39740 6213 39744
rect 6149 39684 6153 39740
rect 6153 39684 6209 39740
rect 6209 39684 6213 39740
rect 6149 39680 6213 39684
rect 6229 39740 6293 39744
rect 6229 39684 6233 39740
rect 6233 39684 6289 39740
rect 6289 39684 6293 39740
rect 6229 39680 6293 39684
rect 9347 39740 9411 39744
rect 9347 39684 9351 39740
rect 9351 39684 9407 39740
rect 9407 39684 9411 39740
rect 9347 39680 9411 39684
rect 9427 39740 9491 39744
rect 9427 39684 9431 39740
rect 9431 39684 9487 39740
rect 9487 39684 9491 39740
rect 9427 39680 9491 39684
rect 9507 39740 9571 39744
rect 9507 39684 9511 39740
rect 9511 39684 9567 39740
rect 9567 39684 9571 39740
rect 9507 39680 9571 39684
rect 9587 39740 9651 39744
rect 9587 39684 9591 39740
rect 9591 39684 9647 39740
rect 9647 39684 9651 39740
rect 9587 39680 9651 39684
rect 12705 39740 12769 39744
rect 12705 39684 12709 39740
rect 12709 39684 12765 39740
rect 12765 39684 12769 39740
rect 12705 39680 12769 39684
rect 12785 39740 12849 39744
rect 12785 39684 12789 39740
rect 12789 39684 12845 39740
rect 12845 39684 12849 39740
rect 12785 39680 12849 39684
rect 12865 39740 12929 39744
rect 12865 39684 12869 39740
rect 12869 39684 12925 39740
rect 12925 39684 12929 39740
rect 12865 39680 12929 39684
rect 12945 39740 13009 39744
rect 12945 39684 12949 39740
rect 12949 39684 13005 39740
rect 13005 39684 13009 39740
rect 12945 39680 13009 39684
rect 4310 39196 4374 39200
rect 4310 39140 4314 39196
rect 4314 39140 4370 39196
rect 4370 39140 4374 39196
rect 4310 39136 4374 39140
rect 4390 39196 4454 39200
rect 4390 39140 4394 39196
rect 4394 39140 4450 39196
rect 4450 39140 4454 39196
rect 4390 39136 4454 39140
rect 4470 39196 4534 39200
rect 4470 39140 4474 39196
rect 4474 39140 4530 39196
rect 4530 39140 4534 39196
rect 4470 39136 4534 39140
rect 4550 39196 4614 39200
rect 4550 39140 4554 39196
rect 4554 39140 4610 39196
rect 4610 39140 4614 39196
rect 4550 39136 4614 39140
rect 7668 39196 7732 39200
rect 7668 39140 7672 39196
rect 7672 39140 7728 39196
rect 7728 39140 7732 39196
rect 7668 39136 7732 39140
rect 7748 39196 7812 39200
rect 7748 39140 7752 39196
rect 7752 39140 7808 39196
rect 7808 39140 7812 39196
rect 7748 39136 7812 39140
rect 7828 39196 7892 39200
rect 7828 39140 7832 39196
rect 7832 39140 7888 39196
rect 7888 39140 7892 39196
rect 7828 39136 7892 39140
rect 7908 39196 7972 39200
rect 7908 39140 7912 39196
rect 7912 39140 7968 39196
rect 7968 39140 7972 39196
rect 7908 39136 7972 39140
rect 11026 39196 11090 39200
rect 11026 39140 11030 39196
rect 11030 39140 11086 39196
rect 11086 39140 11090 39196
rect 11026 39136 11090 39140
rect 11106 39196 11170 39200
rect 11106 39140 11110 39196
rect 11110 39140 11166 39196
rect 11166 39140 11170 39196
rect 11106 39136 11170 39140
rect 11186 39196 11250 39200
rect 11186 39140 11190 39196
rect 11190 39140 11246 39196
rect 11246 39140 11250 39196
rect 11186 39136 11250 39140
rect 11266 39196 11330 39200
rect 11266 39140 11270 39196
rect 11270 39140 11326 39196
rect 11326 39140 11330 39196
rect 11266 39136 11330 39140
rect 14384 39196 14448 39200
rect 14384 39140 14388 39196
rect 14388 39140 14444 39196
rect 14444 39140 14448 39196
rect 14384 39136 14448 39140
rect 14464 39196 14528 39200
rect 14464 39140 14468 39196
rect 14468 39140 14524 39196
rect 14524 39140 14528 39196
rect 14464 39136 14528 39140
rect 14544 39196 14608 39200
rect 14544 39140 14548 39196
rect 14548 39140 14604 39196
rect 14604 39140 14608 39196
rect 14544 39136 14608 39140
rect 14624 39196 14688 39200
rect 14624 39140 14628 39196
rect 14628 39140 14684 39196
rect 14684 39140 14688 39196
rect 14624 39136 14688 39140
rect 2631 38652 2695 38656
rect 2631 38596 2635 38652
rect 2635 38596 2691 38652
rect 2691 38596 2695 38652
rect 2631 38592 2695 38596
rect 2711 38652 2775 38656
rect 2711 38596 2715 38652
rect 2715 38596 2771 38652
rect 2771 38596 2775 38652
rect 2711 38592 2775 38596
rect 2791 38652 2855 38656
rect 2791 38596 2795 38652
rect 2795 38596 2851 38652
rect 2851 38596 2855 38652
rect 2791 38592 2855 38596
rect 2871 38652 2935 38656
rect 2871 38596 2875 38652
rect 2875 38596 2931 38652
rect 2931 38596 2935 38652
rect 2871 38592 2935 38596
rect 5989 38652 6053 38656
rect 5989 38596 5993 38652
rect 5993 38596 6049 38652
rect 6049 38596 6053 38652
rect 5989 38592 6053 38596
rect 6069 38652 6133 38656
rect 6069 38596 6073 38652
rect 6073 38596 6129 38652
rect 6129 38596 6133 38652
rect 6069 38592 6133 38596
rect 6149 38652 6213 38656
rect 6149 38596 6153 38652
rect 6153 38596 6209 38652
rect 6209 38596 6213 38652
rect 6149 38592 6213 38596
rect 6229 38652 6293 38656
rect 6229 38596 6233 38652
rect 6233 38596 6289 38652
rect 6289 38596 6293 38652
rect 6229 38592 6293 38596
rect 9347 38652 9411 38656
rect 9347 38596 9351 38652
rect 9351 38596 9407 38652
rect 9407 38596 9411 38652
rect 9347 38592 9411 38596
rect 9427 38652 9491 38656
rect 9427 38596 9431 38652
rect 9431 38596 9487 38652
rect 9487 38596 9491 38652
rect 9427 38592 9491 38596
rect 9507 38652 9571 38656
rect 9507 38596 9511 38652
rect 9511 38596 9567 38652
rect 9567 38596 9571 38652
rect 9507 38592 9571 38596
rect 9587 38652 9651 38656
rect 9587 38596 9591 38652
rect 9591 38596 9647 38652
rect 9647 38596 9651 38652
rect 9587 38592 9651 38596
rect 12705 38652 12769 38656
rect 12705 38596 12709 38652
rect 12709 38596 12765 38652
rect 12765 38596 12769 38652
rect 12705 38592 12769 38596
rect 12785 38652 12849 38656
rect 12785 38596 12789 38652
rect 12789 38596 12845 38652
rect 12845 38596 12849 38652
rect 12785 38592 12849 38596
rect 12865 38652 12929 38656
rect 12865 38596 12869 38652
rect 12869 38596 12925 38652
rect 12925 38596 12929 38652
rect 12865 38592 12929 38596
rect 12945 38652 13009 38656
rect 12945 38596 12949 38652
rect 12949 38596 13005 38652
rect 13005 38596 13009 38652
rect 12945 38592 13009 38596
rect 4310 38108 4374 38112
rect 4310 38052 4314 38108
rect 4314 38052 4370 38108
rect 4370 38052 4374 38108
rect 4310 38048 4374 38052
rect 4390 38108 4454 38112
rect 4390 38052 4394 38108
rect 4394 38052 4450 38108
rect 4450 38052 4454 38108
rect 4390 38048 4454 38052
rect 4470 38108 4534 38112
rect 4470 38052 4474 38108
rect 4474 38052 4530 38108
rect 4530 38052 4534 38108
rect 4470 38048 4534 38052
rect 4550 38108 4614 38112
rect 4550 38052 4554 38108
rect 4554 38052 4610 38108
rect 4610 38052 4614 38108
rect 4550 38048 4614 38052
rect 7668 38108 7732 38112
rect 7668 38052 7672 38108
rect 7672 38052 7728 38108
rect 7728 38052 7732 38108
rect 7668 38048 7732 38052
rect 7748 38108 7812 38112
rect 7748 38052 7752 38108
rect 7752 38052 7808 38108
rect 7808 38052 7812 38108
rect 7748 38048 7812 38052
rect 7828 38108 7892 38112
rect 7828 38052 7832 38108
rect 7832 38052 7888 38108
rect 7888 38052 7892 38108
rect 7828 38048 7892 38052
rect 7908 38108 7972 38112
rect 7908 38052 7912 38108
rect 7912 38052 7968 38108
rect 7968 38052 7972 38108
rect 7908 38048 7972 38052
rect 11026 38108 11090 38112
rect 11026 38052 11030 38108
rect 11030 38052 11086 38108
rect 11086 38052 11090 38108
rect 11026 38048 11090 38052
rect 11106 38108 11170 38112
rect 11106 38052 11110 38108
rect 11110 38052 11166 38108
rect 11166 38052 11170 38108
rect 11106 38048 11170 38052
rect 11186 38108 11250 38112
rect 11186 38052 11190 38108
rect 11190 38052 11246 38108
rect 11246 38052 11250 38108
rect 11186 38048 11250 38052
rect 11266 38108 11330 38112
rect 11266 38052 11270 38108
rect 11270 38052 11326 38108
rect 11326 38052 11330 38108
rect 11266 38048 11330 38052
rect 14384 38108 14448 38112
rect 14384 38052 14388 38108
rect 14388 38052 14444 38108
rect 14444 38052 14448 38108
rect 14384 38048 14448 38052
rect 14464 38108 14528 38112
rect 14464 38052 14468 38108
rect 14468 38052 14524 38108
rect 14524 38052 14528 38108
rect 14464 38048 14528 38052
rect 14544 38108 14608 38112
rect 14544 38052 14548 38108
rect 14548 38052 14604 38108
rect 14604 38052 14608 38108
rect 14544 38048 14608 38052
rect 14624 38108 14688 38112
rect 14624 38052 14628 38108
rect 14628 38052 14684 38108
rect 14684 38052 14688 38108
rect 14624 38048 14688 38052
rect 2631 37564 2695 37568
rect 2631 37508 2635 37564
rect 2635 37508 2691 37564
rect 2691 37508 2695 37564
rect 2631 37504 2695 37508
rect 2711 37564 2775 37568
rect 2711 37508 2715 37564
rect 2715 37508 2771 37564
rect 2771 37508 2775 37564
rect 2711 37504 2775 37508
rect 2791 37564 2855 37568
rect 2791 37508 2795 37564
rect 2795 37508 2851 37564
rect 2851 37508 2855 37564
rect 2791 37504 2855 37508
rect 2871 37564 2935 37568
rect 2871 37508 2875 37564
rect 2875 37508 2931 37564
rect 2931 37508 2935 37564
rect 2871 37504 2935 37508
rect 5989 37564 6053 37568
rect 5989 37508 5993 37564
rect 5993 37508 6049 37564
rect 6049 37508 6053 37564
rect 5989 37504 6053 37508
rect 6069 37564 6133 37568
rect 6069 37508 6073 37564
rect 6073 37508 6129 37564
rect 6129 37508 6133 37564
rect 6069 37504 6133 37508
rect 6149 37564 6213 37568
rect 6149 37508 6153 37564
rect 6153 37508 6209 37564
rect 6209 37508 6213 37564
rect 6149 37504 6213 37508
rect 6229 37564 6293 37568
rect 6229 37508 6233 37564
rect 6233 37508 6289 37564
rect 6289 37508 6293 37564
rect 6229 37504 6293 37508
rect 9347 37564 9411 37568
rect 9347 37508 9351 37564
rect 9351 37508 9407 37564
rect 9407 37508 9411 37564
rect 9347 37504 9411 37508
rect 9427 37564 9491 37568
rect 9427 37508 9431 37564
rect 9431 37508 9487 37564
rect 9487 37508 9491 37564
rect 9427 37504 9491 37508
rect 9507 37564 9571 37568
rect 9507 37508 9511 37564
rect 9511 37508 9567 37564
rect 9567 37508 9571 37564
rect 9507 37504 9571 37508
rect 9587 37564 9651 37568
rect 9587 37508 9591 37564
rect 9591 37508 9647 37564
rect 9647 37508 9651 37564
rect 9587 37504 9651 37508
rect 12705 37564 12769 37568
rect 12705 37508 12709 37564
rect 12709 37508 12765 37564
rect 12765 37508 12769 37564
rect 12705 37504 12769 37508
rect 12785 37564 12849 37568
rect 12785 37508 12789 37564
rect 12789 37508 12845 37564
rect 12845 37508 12849 37564
rect 12785 37504 12849 37508
rect 12865 37564 12929 37568
rect 12865 37508 12869 37564
rect 12869 37508 12925 37564
rect 12925 37508 12929 37564
rect 12865 37504 12929 37508
rect 12945 37564 13009 37568
rect 12945 37508 12949 37564
rect 12949 37508 13005 37564
rect 13005 37508 13009 37564
rect 12945 37504 13009 37508
rect 10364 37360 10428 37364
rect 10364 37304 10414 37360
rect 10414 37304 10428 37360
rect 10364 37300 10428 37304
rect 11836 37360 11900 37364
rect 11836 37304 11850 37360
rect 11850 37304 11900 37360
rect 11836 37300 11900 37304
rect 4310 37020 4374 37024
rect 4310 36964 4314 37020
rect 4314 36964 4370 37020
rect 4370 36964 4374 37020
rect 4310 36960 4374 36964
rect 4390 37020 4454 37024
rect 4390 36964 4394 37020
rect 4394 36964 4450 37020
rect 4450 36964 4454 37020
rect 4390 36960 4454 36964
rect 4470 37020 4534 37024
rect 4470 36964 4474 37020
rect 4474 36964 4530 37020
rect 4530 36964 4534 37020
rect 4470 36960 4534 36964
rect 4550 37020 4614 37024
rect 4550 36964 4554 37020
rect 4554 36964 4610 37020
rect 4610 36964 4614 37020
rect 4550 36960 4614 36964
rect 7668 37020 7732 37024
rect 7668 36964 7672 37020
rect 7672 36964 7728 37020
rect 7728 36964 7732 37020
rect 7668 36960 7732 36964
rect 7748 37020 7812 37024
rect 7748 36964 7752 37020
rect 7752 36964 7808 37020
rect 7808 36964 7812 37020
rect 7748 36960 7812 36964
rect 7828 37020 7892 37024
rect 7828 36964 7832 37020
rect 7832 36964 7888 37020
rect 7888 36964 7892 37020
rect 7828 36960 7892 36964
rect 7908 37020 7972 37024
rect 7908 36964 7912 37020
rect 7912 36964 7968 37020
rect 7968 36964 7972 37020
rect 7908 36960 7972 36964
rect 11026 37020 11090 37024
rect 11026 36964 11030 37020
rect 11030 36964 11086 37020
rect 11086 36964 11090 37020
rect 11026 36960 11090 36964
rect 11106 37020 11170 37024
rect 11106 36964 11110 37020
rect 11110 36964 11166 37020
rect 11166 36964 11170 37020
rect 11106 36960 11170 36964
rect 11186 37020 11250 37024
rect 11186 36964 11190 37020
rect 11190 36964 11246 37020
rect 11246 36964 11250 37020
rect 11186 36960 11250 36964
rect 11266 37020 11330 37024
rect 11266 36964 11270 37020
rect 11270 36964 11326 37020
rect 11326 36964 11330 37020
rect 11266 36960 11330 36964
rect 14384 37020 14448 37024
rect 14384 36964 14388 37020
rect 14388 36964 14444 37020
rect 14444 36964 14448 37020
rect 14384 36960 14448 36964
rect 14464 37020 14528 37024
rect 14464 36964 14468 37020
rect 14468 36964 14524 37020
rect 14524 36964 14528 37020
rect 14464 36960 14528 36964
rect 14544 37020 14608 37024
rect 14544 36964 14548 37020
rect 14548 36964 14604 37020
rect 14604 36964 14608 37020
rect 14544 36960 14608 36964
rect 14624 37020 14688 37024
rect 14624 36964 14628 37020
rect 14628 36964 14684 37020
rect 14684 36964 14688 37020
rect 14624 36960 14688 36964
rect 2631 36476 2695 36480
rect 2631 36420 2635 36476
rect 2635 36420 2691 36476
rect 2691 36420 2695 36476
rect 2631 36416 2695 36420
rect 2711 36476 2775 36480
rect 2711 36420 2715 36476
rect 2715 36420 2771 36476
rect 2771 36420 2775 36476
rect 2711 36416 2775 36420
rect 2791 36476 2855 36480
rect 2791 36420 2795 36476
rect 2795 36420 2851 36476
rect 2851 36420 2855 36476
rect 2791 36416 2855 36420
rect 2871 36476 2935 36480
rect 2871 36420 2875 36476
rect 2875 36420 2931 36476
rect 2931 36420 2935 36476
rect 2871 36416 2935 36420
rect 5989 36476 6053 36480
rect 5989 36420 5993 36476
rect 5993 36420 6049 36476
rect 6049 36420 6053 36476
rect 5989 36416 6053 36420
rect 6069 36476 6133 36480
rect 6069 36420 6073 36476
rect 6073 36420 6129 36476
rect 6129 36420 6133 36476
rect 6069 36416 6133 36420
rect 6149 36476 6213 36480
rect 6149 36420 6153 36476
rect 6153 36420 6209 36476
rect 6209 36420 6213 36476
rect 6149 36416 6213 36420
rect 6229 36476 6293 36480
rect 6229 36420 6233 36476
rect 6233 36420 6289 36476
rect 6289 36420 6293 36476
rect 6229 36416 6293 36420
rect 9347 36476 9411 36480
rect 9347 36420 9351 36476
rect 9351 36420 9407 36476
rect 9407 36420 9411 36476
rect 9347 36416 9411 36420
rect 9427 36476 9491 36480
rect 9427 36420 9431 36476
rect 9431 36420 9487 36476
rect 9487 36420 9491 36476
rect 9427 36416 9491 36420
rect 9507 36476 9571 36480
rect 9507 36420 9511 36476
rect 9511 36420 9567 36476
rect 9567 36420 9571 36476
rect 9507 36416 9571 36420
rect 9587 36476 9651 36480
rect 9587 36420 9591 36476
rect 9591 36420 9647 36476
rect 9647 36420 9651 36476
rect 9587 36416 9651 36420
rect 12705 36476 12769 36480
rect 12705 36420 12709 36476
rect 12709 36420 12765 36476
rect 12765 36420 12769 36476
rect 12705 36416 12769 36420
rect 12785 36476 12849 36480
rect 12785 36420 12789 36476
rect 12789 36420 12845 36476
rect 12845 36420 12849 36476
rect 12785 36416 12849 36420
rect 12865 36476 12929 36480
rect 12865 36420 12869 36476
rect 12869 36420 12925 36476
rect 12925 36420 12929 36476
rect 12865 36416 12929 36420
rect 12945 36476 13009 36480
rect 12945 36420 12949 36476
rect 12949 36420 13005 36476
rect 13005 36420 13009 36476
rect 12945 36416 13009 36420
rect 4310 35932 4374 35936
rect 4310 35876 4314 35932
rect 4314 35876 4370 35932
rect 4370 35876 4374 35932
rect 4310 35872 4374 35876
rect 4390 35932 4454 35936
rect 4390 35876 4394 35932
rect 4394 35876 4450 35932
rect 4450 35876 4454 35932
rect 4390 35872 4454 35876
rect 4470 35932 4534 35936
rect 4470 35876 4474 35932
rect 4474 35876 4530 35932
rect 4530 35876 4534 35932
rect 4470 35872 4534 35876
rect 4550 35932 4614 35936
rect 4550 35876 4554 35932
rect 4554 35876 4610 35932
rect 4610 35876 4614 35932
rect 4550 35872 4614 35876
rect 7668 35932 7732 35936
rect 7668 35876 7672 35932
rect 7672 35876 7728 35932
rect 7728 35876 7732 35932
rect 7668 35872 7732 35876
rect 7748 35932 7812 35936
rect 7748 35876 7752 35932
rect 7752 35876 7808 35932
rect 7808 35876 7812 35932
rect 7748 35872 7812 35876
rect 7828 35932 7892 35936
rect 7828 35876 7832 35932
rect 7832 35876 7888 35932
rect 7888 35876 7892 35932
rect 7828 35872 7892 35876
rect 7908 35932 7972 35936
rect 7908 35876 7912 35932
rect 7912 35876 7968 35932
rect 7968 35876 7972 35932
rect 7908 35872 7972 35876
rect 11026 35932 11090 35936
rect 11026 35876 11030 35932
rect 11030 35876 11086 35932
rect 11086 35876 11090 35932
rect 11026 35872 11090 35876
rect 11106 35932 11170 35936
rect 11106 35876 11110 35932
rect 11110 35876 11166 35932
rect 11166 35876 11170 35932
rect 11106 35872 11170 35876
rect 11186 35932 11250 35936
rect 11186 35876 11190 35932
rect 11190 35876 11246 35932
rect 11246 35876 11250 35932
rect 11186 35872 11250 35876
rect 11266 35932 11330 35936
rect 11266 35876 11270 35932
rect 11270 35876 11326 35932
rect 11326 35876 11330 35932
rect 11266 35872 11330 35876
rect 14384 35932 14448 35936
rect 14384 35876 14388 35932
rect 14388 35876 14444 35932
rect 14444 35876 14448 35932
rect 14384 35872 14448 35876
rect 14464 35932 14528 35936
rect 14464 35876 14468 35932
rect 14468 35876 14524 35932
rect 14524 35876 14528 35932
rect 14464 35872 14528 35876
rect 14544 35932 14608 35936
rect 14544 35876 14548 35932
rect 14548 35876 14604 35932
rect 14604 35876 14608 35932
rect 14544 35872 14608 35876
rect 14624 35932 14688 35936
rect 14624 35876 14628 35932
rect 14628 35876 14684 35932
rect 14684 35876 14688 35932
rect 14624 35872 14688 35876
rect 2631 35388 2695 35392
rect 2631 35332 2635 35388
rect 2635 35332 2691 35388
rect 2691 35332 2695 35388
rect 2631 35328 2695 35332
rect 2711 35388 2775 35392
rect 2711 35332 2715 35388
rect 2715 35332 2771 35388
rect 2771 35332 2775 35388
rect 2711 35328 2775 35332
rect 2791 35388 2855 35392
rect 2791 35332 2795 35388
rect 2795 35332 2851 35388
rect 2851 35332 2855 35388
rect 2791 35328 2855 35332
rect 2871 35388 2935 35392
rect 2871 35332 2875 35388
rect 2875 35332 2931 35388
rect 2931 35332 2935 35388
rect 2871 35328 2935 35332
rect 5989 35388 6053 35392
rect 5989 35332 5993 35388
rect 5993 35332 6049 35388
rect 6049 35332 6053 35388
rect 5989 35328 6053 35332
rect 6069 35388 6133 35392
rect 6069 35332 6073 35388
rect 6073 35332 6129 35388
rect 6129 35332 6133 35388
rect 6069 35328 6133 35332
rect 6149 35388 6213 35392
rect 6149 35332 6153 35388
rect 6153 35332 6209 35388
rect 6209 35332 6213 35388
rect 6149 35328 6213 35332
rect 6229 35388 6293 35392
rect 6229 35332 6233 35388
rect 6233 35332 6289 35388
rect 6289 35332 6293 35388
rect 6229 35328 6293 35332
rect 9347 35388 9411 35392
rect 9347 35332 9351 35388
rect 9351 35332 9407 35388
rect 9407 35332 9411 35388
rect 9347 35328 9411 35332
rect 9427 35388 9491 35392
rect 9427 35332 9431 35388
rect 9431 35332 9487 35388
rect 9487 35332 9491 35388
rect 9427 35328 9491 35332
rect 9507 35388 9571 35392
rect 9507 35332 9511 35388
rect 9511 35332 9567 35388
rect 9567 35332 9571 35388
rect 9507 35328 9571 35332
rect 9587 35388 9651 35392
rect 9587 35332 9591 35388
rect 9591 35332 9647 35388
rect 9647 35332 9651 35388
rect 9587 35328 9651 35332
rect 12705 35388 12769 35392
rect 12705 35332 12709 35388
rect 12709 35332 12765 35388
rect 12765 35332 12769 35388
rect 12705 35328 12769 35332
rect 12785 35388 12849 35392
rect 12785 35332 12789 35388
rect 12789 35332 12845 35388
rect 12845 35332 12849 35388
rect 12785 35328 12849 35332
rect 12865 35388 12929 35392
rect 12865 35332 12869 35388
rect 12869 35332 12925 35388
rect 12925 35332 12929 35388
rect 12865 35328 12929 35332
rect 12945 35388 13009 35392
rect 12945 35332 12949 35388
rect 12949 35332 13005 35388
rect 13005 35332 13009 35388
rect 12945 35328 13009 35332
rect 4310 34844 4374 34848
rect 4310 34788 4314 34844
rect 4314 34788 4370 34844
rect 4370 34788 4374 34844
rect 4310 34784 4374 34788
rect 4390 34844 4454 34848
rect 4390 34788 4394 34844
rect 4394 34788 4450 34844
rect 4450 34788 4454 34844
rect 4390 34784 4454 34788
rect 4470 34844 4534 34848
rect 4470 34788 4474 34844
rect 4474 34788 4530 34844
rect 4530 34788 4534 34844
rect 4470 34784 4534 34788
rect 4550 34844 4614 34848
rect 4550 34788 4554 34844
rect 4554 34788 4610 34844
rect 4610 34788 4614 34844
rect 4550 34784 4614 34788
rect 7668 34844 7732 34848
rect 7668 34788 7672 34844
rect 7672 34788 7728 34844
rect 7728 34788 7732 34844
rect 7668 34784 7732 34788
rect 7748 34844 7812 34848
rect 7748 34788 7752 34844
rect 7752 34788 7808 34844
rect 7808 34788 7812 34844
rect 7748 34784 7812 34788
rect 7828 34844 7892 34848
rect 7828 34788 7832 34844
rect 7832 34788 7888 34844
rect 7888 34788 7892 34844
rect 7828 34784 7892 34788
rect 7908 34844 7972 34848
rect 7908 34788 7912 34844
rect 7912 34788 7968 34844
rect 7968 34788 7972 34844
rect 7908 34784 7972 34788
rect 11026 34844 11090 34848
rect 11026 34788 11030 34844
rect 11030 34788 11086 34844
rect 11086 34788 11090 34844
rect 11026 34784 11090 34788
rect 11106 34844 11170 34848
rect 11106 34788 11110 34844
rect 11110 34788 11166 34844
rect 11166 34788 11170 34844
rect 11106 34784 11170 34788
rect 11186 34844 11250 34848
rect 11186 34788 11190 34844
rect 11190 34788 11246 34844
rect 11246 34788 11250 34844
rect 11186 34784 11250 34788
rect 11266 34844 11330 34848
rect 11266 34788 11270 34844
rect 11270 34788 11326 34844
rect 11326 34788 11330 34844
rect 11266 34784 11330 34788
rect 14384 34844 14448 34848
rect 14384 34788 14388 34844
rect 14388 34788 14444 34844
rect 14444 34788 14448 34844
rect 14384 34784 14448 34788
rect 14464 34844 14528 34848
rect 14464 34788 14468 34844
rect 14468 34788 14524 34844
rect 14524 34788 14528 34844
rect 14464 34784 14528 34788
rect 14544 34844 14608 34848
rect 14544 34788 14548 34844
rect 14548 34788 14604 34844
rect 14604 34788 14608 34844
rect 14544 34784 14608 34788
rect 14624 34844 14688 34848
rect 14624 34788 14628 34844
rect 14628 34788 14684 34844
rect 14684 34788 14688 34844
rect 14624 34784 14688 34788
rect 6500 34580 6564 34644
rect 12572 34580 12636 34644
rect 2631 34300 2695 34304
rect 2631 34244 2635 34300
rect 2635 34244 2691 34300
rect 2691 34244 2695 34300
rect 2631 34240 2695 34244
rect 2711 34300 2775 34304
rect 2711 34244 2715 34300
rect 2715 34244 2771 34300
rect 2771 34244 2775 34300
rect 2711 34240 2775 34244
rect 2791 34300 2855 34304
rect 2791 34244 2795 34300
rect 2795 34244 2851 34300
rect 2851 34244 2855 34300
rect 2791 34240 2855 34244
rect 2871 34300 2935 34304
rect 2871 34244 2875 34300
rect 2875 34244 2931 34300
rect 2931 34244 2935 34300
rect 2871 34240 2935 34244
rect 5989 34300 6053 34304
rect 5989 34244 5993 34300
rect 5993 34244 6049 34300
rect 6049 34244 6053 34300
rect 5989 34240 6053 34244
rect 6069 34300 6133 34304
rect 6069 34244 6073 34300
rect 6073 34244 6129 34300
rect 6129 34244 6133 34300
rect 6069 34240 6133 34244
rect 6149 34300 6213 34304
rect 6149 34244 6153 34300
rect 6153 34244 6209 34300
rect 6209 34244 6213 34300
rect 6149 34240 6213 34244
rect 6229 34300 6293 34304
rect 6229 34244 6233 34300
rect 6233 34244 6289 34300
rect 6289 34244 6293 34300
rect 6229 34240 6293 34244
rect 9347 34300 9411 34304
rect 9347 34244 9351 34300
rect 9351 34244 9407 34300
rect 9407 34244 9411 34300
rect 9347 34240 9411 34244
rect 9427 34300 9491 34304
rect 9427 34244 9431 34300
rect 9431 34244 9487 34300
rect 9487 34244 9491 34300
rect 9427 34240 9491 34244
rect 9507 34300 9571 34304
rect 9507 34244 9511 34300
rect 9511 34244 9567 34300
rect 9567 34244 9571 34300
rect 9507 34240 9571 34244
rect 9587 34300 9651 34304
rect 9587 34244 9591 34300
rect 9591 34244 9647 34300
rect 9647 34244 9651 34300
rect 9587 34240 9651 34244
rect 12705 34300 12769 34304
rect 12705 34244 12709 34300
rect 12709 34244 12765 34300
rect 12765 34244 12769 34300
rect 12705 34240 12769 34244
rect 12785 34300 12849 34304
rect 12785 34244 12789 34300
rect 12789 34244 12845 34300
rect 12845 34244 12849 34300
rect 12785 34240 12849 34244
rect 12865 34300 12929 34304
rect 12865 34244 12869 34300
rect 12869 34244 12925 34300
rect 12925 34244 12929 34300
rect 12865 34240 12929 34244
rect 12945 34300 13009 34304
rect 12945 34244 12949 34300
rect 12949 34244 13005 34300
rect 13005 34244 13009 34300
rect 12945 34240 13009 34244
rect 10180 33900 10244 33964
rect 10732 33900 10796 33964
rect 4310 33756 4374 33760
rect 4310 33700 4314 33756
rect 4314 33700 4370 33756
rect 4370 33700 4374 33756
rect 4310 33696 4374 33700
rect 4390 33756 4454 33760
rect 4390 33700 4394 33756
rect 4394 33700 4450 33756
rect 4450 33700 4454 33756
rect 4390 33696 4454 33700
rect 4470 33756 4534 33760
rect 4470 33700 4474 33756
rect 4474 33700 4530 33756
rect 4530 33700 4534 33756
rect 4470 33696 4534 33700
rect 4550 33756 4614 33760
rect 4550 33700 4554 33756
rect 4554 33700 4610 33756
rect 4610 33700 4614 33756
rect 4550 33696 4614 33700
rect 7668 33756 7732 33760
rect 7668 33700 7672 33756
rect 7672 33700 7728 33756
rect 7728 33700 7732 33756
rect 7668 33696 7732 33700
rect 7748 33756 7812 33760
rect 7748 33700 7752 33756
rect 7752 33700 7808 33756
rect 7808 33700 7812 33756
rect 7748 33696 7812 33700
rect 7828 33756 7892 33760
rect 7828 33700 7832 33756
rect 7832 33700 7888 33756
rect 7888 33700 7892 33756
rect 7828 33696 7892 33700
rect 7908 33756 7972 33760
rect 7908 33700 7912 33756
rect 7912 33700 7968 33756
rect 7968 33700 7972 33756
rect 7908 33696 7972 33700
rect 11026 33756 11090 33760
rect 11026 33700 11030 33756
rect 11030 33700 11086 33756
rect 11086 33700 11090 33756
rect 11026 33696 11090 33700
rect 11106 33756 11170 33760
rect 11106 33700 11110 33756
rect 11110 33700 11166 33756
rect 11166 33700 11170 33756
rect 11106 33696 11170 33700
rect 11186 33756 11250 33760
rect 11186 33700 11190 33756
rect 11190 33700 11246 33756
rect 11246 33700 11250 33756
rect 11186 33696 11250 33700
rect 11266 33756 11330 33760
rect 11266 33700 11270 33756
rect 11270 33700 11326 33756
rect 11326 33700 11330 33756
rect 11266 33696 11330 33700
rect 14384 33756 14448 33760
rect 14384 33700 14388 33756
rect 14388 33700 14444 33756
rect 14444 33700 14448 33756
rect 14384 33696 14448 33700
rect 14464 33756 14528 33760
rect 14464 33700 14468 33756
rect 14468 33700 14524 33756
rect 14524 33700 14528 33756
rect 14464 33696 14528 33700
rect 14544 33756 14608 33760
rect 14544 33700 14548 33756
rect 14548 33700 14604 33756
rect 14604 33700 14608 33756
rect 14544 33696 14608 33700
rect 14624 33756 14688 33760
rect 14624 33700 14628 33756
rect 14628 33700 14684 33756
rect 14684 33700 14688 33756
rect 14624 33696 14688 33700
rect 2631 33212 2695 33216
rect 2631 33156 2635 33212
rect 2635 33156 2691 33212
rect 2691 33156 2695 33212
rect 2631 33152 2695 33156
rect 2711 33212 2775 33216
rect 2711 33156 2715 33212
rect 2715 33156 2771 33212
rect 2771 33156 2775 33212
rect 2711 33152 2775 33156
rect 2791 33212 2855 33216
rect 2791 33156 2795 33212
rect 2795 33156 2851 33212
rect 2851 33156 2855 33212
rect 2791 33152 2855 33156
rect 2871 33212 2935 33216
rect 2871 33156 2875 33212
rect 2875 33156 2931 33212
rect 2931 33156 2935 33212
rect 2871 33152 2935 33156
rect 5989 33212 6053 33216
rect 5989 33156 5993 33212
rect 5993 33156 6049 33212
rect 6049 33156 6053 33212
rect 5989 33152 6053 33156
rect 6069 33212 6133 33216
rect 6069 33156 6073 33212
rect 6073 33156 6129 33212
rect 6129 33156 6133 33212
rect 6069 33152 6133 33156
rect 6149 33212 6213 33216
rect 6149 33156 6153 33212
rect 6153 33156 6209 33212
rect 6209 33156 6213 33212
rect 6149 33152 6213 33156
rect 6229 33212 6293 33216
rect 6229 33156 6233 33212
rect 6233 33156 6289 33212
rect 6289 33156 6293 33212
rect 6229 33152 6293 33156
rect 9347 33212 9411 33216
rect 9347 33156 9351 33212
rect 9351 33156 9407 33212
rect 9407 33156 9411 33212
rect 9347 33152 9411 33156
rect 9427 33212 9491 33216
rect 9427 33156 9431 33212
rect 9431 33156 9487 33212
rect 9487 33156 9491 33212
rect 9427 33152 9491 33156
rect 9507 33212 9571 33216
rect 9507 33156 9511 33212
rect 9511 33156 9567 33212
rect 9567 33156 9571 33212
rect 9507 33152 9571 33156
rect 9587 33212 9651 33216
rect 9587 33156 9591 33212
rect 9591 33156 9647 33212
rect 9647 33156 9651 33212
rect 9587 33152 9651 33156
rect 12705 33212 12769 33216
rect 12705 33156 12709 33212
rect 12709 33156 12765 33212
rect 12765 33156 12769 33212
rect 12705 33152 12769 33156
rect 12785 33212 12849 33216
rect 12785 33156 12789 33212
rect 12789 33156 12845 33212
rect 12845 33156 12849 33212
rect 12785 33152 12849 33156
rect 12865 33212 12929 33216
rect 12865 33156 12869 33212
rect 12869 33156 12925 33212
rect 12925 33156 12929 33212
rect 12865 33152 12929 33156
rect 12945 33212 13009 33216
rect 12945 33156 12949 33212
rect 12949 33156 13005 33212
rect 13005 33156 13009 33212
rect 12945 33152 13009 33156
rect 12572 32948 12636 33012
rect 10180 32812 10244 32876
rect 4310 32668 4374 32672
rect 4310 32612 4314 32668
rect 4314 32612 4370 32668
rect 4370 32612 4374 32668
rect 4310 32608 4374 32612
rect 4390 32668 4454 32672
rect 4390 32612 4394 32668
rect 4394 32612 4450 32668
rect 4450 32612 4454 32668
rect 4390 32608 4454 32612
rect 4470 32668 4534 32672
rect 4470 32612 4474 32668
rect 4474 32612 4530 32668
rect 4530 32612 4534 32668
rect 4470 32608 4534 32612
rect 4550 32668 4614 32672
rect 4550 32612 4554 32668
rect 4554 32612 4610 32668
rect 4610 32612 4614 32668
rect 4550 32608 4614 32612
rect 7668 32668 7732 32672
rect 7668 32612 7672 32668
rect 7672 32612 7728 32668
rect 7728 32612 7732 32668
rect 7668 32608 7732 32612
rect 7748 32668 7812 32672
rect 7748 32612 7752 32668
rect 7752 32612 7808 32668
rect 7808 32612 7812 32668
rect 7748 32608 7812 32612
rect 7828 32668 7892 32672
rect 7828 32612 7832 32668
rect 7832 32612 7888 32668
rect 7888 32612 7892 32668
rect 7828 32608 7892 32612
rect 7908 32668 7972 32672
rect 7908 32612 7912 32668
rect 7912 32612 7968 32668
rect 7968 32612 7972 32668
rect 7908 32608 7972 32612
rect 11026 32668 11090 32672
rect 11026 32612 11030 32668
rect 11030 32612 11086 32668
rect 11086 32612 11090 32668
rect 11026 32608 11090 32612
rect 11106 32668 11170 32672
rect 11106 32612 11110 32668
rect 11110 32612 11166 32668
rect 11166 32612 11170 32668
rect 11106 32608 11170 32612
rect 11186 32668 11250 32672
rect 11186 32612 11190 32668
rect 11190 32612 11246 32668
rect 11246 32612 11250 32668
rect 11186 32608 11250 32612
rect 11266 32668 11330 32672
rect 11266 32612 11270 32668
rect 11270 32612 11326 32668
rect 11326 32612 11330 32668
rect 11266 32608 11330 32612
rect 14384 32668 14448 32672
rect 14384 32612 14388 32668
rect 14388 32612 14444 32668
rect 14444 32612 14448 32668
rect 14384 32608 14448 32612
rect 14464 32668 14528 32672
rect 14464 32612 14468 32668
rect 14468 32612 14524 32668
rect 14524 32612 14528 32668
rect 14464 32608 14528 32612
rect 14544 32668 14608 32672
rect 14544 32612 14548 32668
rect 14548 32612 14604 32668
rect 14604 32612 14608 32668
rect 14544 32608 14608 32612
rect 14624 32668 14688 32672
rect 14624 32612 14628 32668
rect 14628 32612 14684 32668
rect 14684 32612 14688 32668
rect 14624 32608 14688 32612
rect 2631 32124 2695 32128
rect 2631 32068 2635 32124
rect 2635 32068 2691 32124
rect 2691 32068 2695 32124
rect 2631 32064 2695 32068
rect 2711 32124 2775 32128
rect 2711 32068 2715 32124
rect 2715 32068 2771 32124
rect 2771 32068 2775 32124
rect 2711 32064 2775 32068
rect 2791 32124 2855 32128
rect 2791 32068 2795 32124
rect 2795 32068 2851 32124
rect 2851 32068 2855 32124
rect 2791 32064 2855 32068
rect 2871 32124 2935 32128
rect 2871 32068 2875 32124
rect 2875 32068 2931 32124
rect 2931 32068 2935 32124
rect 2871 32064 2935 32068
rect 5989 32124 6053 32128
rect 5989 32068 5993 32124
rect 5993 32068 6049 32124
rect 6049 32068 6053 32124
rect 5989 32064 6053 32068
rect 6069 32124 6133 32128
rect 6069 32068 6073 32124
rect 6073 32068 6129 32124
rect 6129 32068 6133 32124
rect 6069 32064 6133 32068
rect 6149 32124 6213 32128
rect 6149 32068 6153 32124
rect 6153 32068 6209 32124
rect 6209 32068 6213 32124
rect 6149 32064 6213 32068
rect 6229 32124 6293 32128
rect 6229 32068 6233 32124
rect 6233 32068 6289 32124
rect 6289 32068 6293 32124
rect 6229 32064 6293 32068
rect 9347 32124 9411 32128
rect 9347 32068 9351 32124
rect 9351 32068 9407 32124
rect 9407 32068 9411 32124
rect 9347 32064 9411 32068
rect 9427 32124 9491 32128
rect 9427 32068 9431 32124
rect 9431 32068 9487 32124
rect 9487 32068 9491 32124
rect 9427 32064 9491 32068
rect 9507 32124 9571 32128
rect 9507 32068 9511 32124
rect 9511 32068 9567 32124
rect 9567 32068 9571 32124
rect 9507 32064 9571 32068
rect 9587 32124 9651 32128
rect 9587 32068 9591 32124
rect 9591 32068 9647 32124
rect 9647 32068 9651 32124
rect 9587 32064 9651 32068
rect 12705 32124 12769 32128
rect 12705 32068 12709 32124
rect 12709 32068 12765 32124
rect 12765 32068 12769 32124
rect 12705 32064 12769 32068
rect 12785 32124 12849 32128
rect 12785 32068 12789 32124
rect 12789 32068 12845 32124
rect 12845 32068 12849 32124
rect 12785 32064 12849 32068
rect 12865 32124 12929 32128
rect 12865 32068 12869 32124
rect 12869 32068 12925 32124
rect 12925 32068 12929 32124
rect 12865 32064 12929 32068
rect 12945 32124 13009 32128
rect 12945 32068 12949 32124
rect 12949 32068 13005 32124
rect 13005 32068 13009 32124
rect 12945 32064 13009 32068
rect 14228 32056 14292 32060
rect 14228 32000 14242 32056
rect 14242 32000 14292 32056
rect 14228 31996 14292 32000
rect 4310 31580 4374 31584
rect 4310 31524 4314 31580
rect 4314 31524 4370 31580
rect 4370 31524 4374 31580
rect 4310 31520 4374 31524
rect 4390 31580 4454 31584
rect 4390 31524 4394 31580
rect 4394 31524 4450 31580
rect 4450 31524 4454 31580
rect 4390 31520 4454 31524
rect 4470 31580 4534 31584
rect 4470 31524 4474 31580
rect 4474 31524 4530 31580
rect 4530 31524 4534 31580
rect 4470 31520 4534 31524
rect 4550 31580 4614 31584
rect 4550 31524 4554 31580
rect 4554 31524 4610 31580
rect 4610 31524 4614 31580
rect 4550 31520 4614 31524
rect 7668 31580 7732 31584
rect 7668 31524 7672 31580
rect 7672 31524 7728 31580
rect 7728 31524 7732 31580
rect 7668 31520 7732 31524
rect 7748 31580 7812 31584
rect 7748 31524 7752 31580
rect 7752 31524 7808 31580
rect 7808 31524 7812 31580
rect 7748 31520 7812 31524
rect 7828 31580 7892 31584
rect 7828 31524 7832 31580
rect 7832 31524 7888 31580
rect 7888 31524 7892 31580
rect 7828 31520 7892 31524
rect 7908 31580 7972 31584
rect 7908 31524 7912 31580
rect 7912 31524 7968 31580
rect 7968 31524 7972 31580
rect 7908 31520 7972 31524
rect 11026 31580 11090 31584
rect 11026 31524 11030 31580
rect 11030 31524 11086 31580
rect 11086 31524 11090 31580
rect 11026 31520 11090 31524
rect 11106 31580 11170 31584
rect 11106 31524 11110 31580
rect 11110 31524 11166 31580
rect 11166 31524 11170 31580
rect 11106 31520 11170 31524
rect 11186 31580 11250 31584
rect 11186 31524 11190 31580
rect 11190 31524 11246 31580
rect 11246 31524 11250 31580
rect 11186 31520 11250 31524
rect 11266 31580 11330 31584
rect 11266 31524 11270 31580
rect 11270 31524 11326 31580
rect 11326 31524 11330 31580
rect 11266 31520 11330 31524
rect 14384 31580 14448 31584
rect 14384 31524 14388 31580
rect 14388 31524 14444 31580
rect 14444 31524 14448 31580
rect 14384 31520 14448 31524
rect 14464 31580 14528 31584
rect 14464 31524 14468 31580
rect 14468 31524 14524 31580
rect 14524 31524 14528 31580
rect 14464 31520 14528 31524
rect 14544 31580 14608 31584
rect 14544 31524 14548 31580
rect 14548 31524 14604 31580
rect 14604 31524 14608 31580
rect 14544 31520 14608 31524
rect 14624 31580 14688 31584
rect 14624 31524 14628 31580
rect 14628 31524 14684 31580
rect 14684 31524 14688 31580
rect 14624 31520 14688 31524
rect 14228 31316 14292 31380
rect 2631 31036 2695 31040
rect 2631 30980 2635 31036
rect 2635 30980 2691 31036
rect 2691 30980 2695 31036
rect 2631 30976 2695 30980
rect 2711 31036 2775 31040
rect 2711 30980 2715 31036
rect 2715 30980 2771 31036
rect 2771 30980 2775 31036
rect 2711 30976 2775 30980
rect 2791 31036 2855 31040
rect 2791 30980 2795 31036
rect 2795 30980 2851 31036
rect 2851 30980 2855 31036
rect 2791 30976 2855 30980
rect 2871 31036 2935 31040
rect 2871 30980 2875 31036
rect 2875 30980 2931 31036
rect 2931 30980 2935 31036
rect 2871 30976 2935 30980
rect 5989 31036 6053 31040
rect 5989 30980 5993 31036
rect 5993 30980 6049 31036
rect 6049 30980 6053 31036
rect 5989 30976 6053 30980
rect 6069 31036 6133 31040
rect 6069 30980 6073 31036
rect 6073 30980 6129 31036
rect 6129 30980 6133 31036
rect 6069 30976 6133 30980
rect 6149 31036 6213 31040
rect 6149 30980 6153 31036
rect 6153 30980 6209 31036
rect 6209 30980 6213 31036
rect 6149 30976 6213 30980
rect 6229 31036 6293 31040
rect 6229 30980 6233 31036
rect 6233 30980 6289 31036
rect 6289 30980 6293 31036
rect 6229 30976 6293 30980
rect 9347 31036 9411 31040
rect 9347 30980 9351 31036
rect 9351 30980 9407 31036
rect 9407 30980 9411 31036
rect 9347 30976 9411 30980
rect 9427 31036 9491 31040
rect 9427 30980 9431 31036
rect 9431 30980 9487 31036
rect 9487 30980 9491 31036
rect 9427 30976 9491 30980
rect 9507 31036 9571 31040
rect 9507 30980 9511 31036
rect 9511 30980 9567 31036
rect 9567 30980 9571 31036
rect 9507 30976 9571 30980
rect 9587 31036 9651 31040
rect 9587 30980 9591 31036
rect 9591 30980 9647 31036
rect 9647 30980 9651 31036
rect 9587 30976 9651 30980
rect 12705 31036 12769 31040
rect 12705 30980 12709 31036
rect 12709 30980 12765 31036
rect 12765 30980 12769 31036
rect 12705 30976 12769 30980
rect 12785 31036 12849 31040
rect 12785 30980 12789 31036
rect 12789 30980 12845 31036
rect 12845 30980 12849 31036
rect 12785 30976 12849 30980
rect 12865 31036 12929 31040
rect 12865 30980 12869 31036
rect 12869 30980 12925 31036
rect 12925 30980 12929 31036
rect 12865 30976 12929 30980
rect 12945 31036 13009 31040
rect 12945 30980 12949 31036
rect 12949 30980 13005 31036
rect 13005 30980 13009 31036
rect 12945 30976 13009 30980
rect 10180 30772 10244 30836
rect 13492 30636 13556 30700
rect 4310 30492 4374 30496
rect 4310 30436 4314 30492
rect 4314 30436 4370 30492
rect 4370 30436 4374 30492
rect 4310 30432 4374 30436
rect 4390 30492 4454 30496
rect 4390 30436 4394 30492
rect 4394 30436 4450 30492
rect 4450 30436 4454 30492
rect 4390 30432 4454 30436
rect 4470 30492 4534 30496
rect 4470 30436 4474 30492
rect 4474 30436 4530 30492
rect 4530 30436 4534 30492
rect 4470 30432 4534 30436
rect 4550 30492 4614 30496
rect 4550 30436 4554 30492
rect 4554 30436 4610 30492
rect 4610 30436 4614 30492
rect 4550 30432 4614 30436
rect 7668 30492 7732 30496
rect 7668 30436 7672 30492
rect 7672 30436 7728 30492
rect 7728 30436 7732 30492
rect 7668 30432 7732 30436
rect 7748 30492 7812 30496
rect 7748 30436 7752 30492
rect 7752 30436 7808 30492
rect 7808 30436 7812 30492
rect 7748 30432 7812 30436
rect 7828 30492 7892 30496
rect 7828 30436 7832 30492
rect 7832 30436 7888 30492
rect 7888 30436 7892 30492
rect 7828 30432 7892 30436
rect 7908 30492 7972 30496
rect 7908 30436 7912 30492
rect 7912 30436 7968 30492
rect 7968 30436 7972 30492
rect 7908 30432 7972 30436
rect 11026 30492 11090 30496
rect 11026 30436 11030 30492
rect 11030 30436 11086 30492
rect 11086 30436 11090 30492
rect 11026 30432 11090 30436
rect 11106 30492 11170 30496
rect 11106 30436 11110 30492
rect 11110 30436 11166 30492
rect 11166 30436 11170 30492
rect 11106 30432 11170 30436
rect 11186 30492 11250 30496
rect 11186 30436 11190 30492
rect 11190 30436 11246 30492
rect 11246 30436 11250 30492
rect 11186 30432 11250 30436
rect 11266 30492 11330 30496
rect 11266 30436 11270 30492
rect 11270 30436 11326 30492
rect 11326 30436 11330 30492
rect 11266 30432 11330 30436
rect 14384 30492 14448 30496
rect 14384 30436 14388 30492
rect 14388 30436 14444 30492
rect 14444 30436 14448 30492
rect 14384 30432 14448 30436
rect 14464 30492 14528 30496
rect 14464 30436 14468 30492
rect 14468 30436 14524 30492
rect 14524 30436 14528 30492
rect 14464 30432 14528 30436
rect 14544 30492 14608 30496
rect 14544 30436 14548 30492
rect 14548 30436 14604 30492
rect 14604 30436 14608 30492
rect 14544 30432 14608 30436
rect 14624 30492 14688 30496
rect 14624 30436 14628 30492
rect 14628 30436 14684 30492
rect 14684 30436 14688 30492
rect 14624 30432 14688 30436
rect 11836 30424 11900 30428
rect 11836 30368 11886 30424
rect 11886 30368 11900 30424
rect 11836 30364 11900 30368
rect 2631 29948 2695 29952
rect 2631 29892 2635 29948
rect 2635 29892 2691 29948
rect 2691 29892 2695 29948
rect 2631 29888 2695 29892
rect 2711 29948 2775 29952
rect 2711 29892 2715 29948
rect 2715 29892 2771 29948
rect 2771 29892 2775 29948
rect 2711 29888 2775 29892
rect 2791 29948 2855 29952
rect 2791 29892 2795 29948
rect 2795 29892 2851 29948
rect 2851 29892 2855 29948
rect 2791 29888 2855 29892
rect 2871 29948 2935 29952
rect 2871 29892 2875 29948
rect 2875 29892 2931 29948
rect 2931 29892 2935 29948
rect 2871 29888 2935 29892
rect 5989 29948 6053 29952
rect 5989 29892 5993 29948
rect 5993 29892 6049 29948
rect 6049 29892 6053 29948
rect 5989 29888 6053 29892
rect 6069 29948 6133 29952
rect 6069 29892 6073 29948
rect 6073 29892 6129 29948
rect 6129 29892 6133 29948
rect 6069 29888 6133 29892
rect 6149 29948 6213 29952
rect 6149 29892 6153 29948
rect 6153 29892 6209 29948
rect 6209 29892 6213 29948
rect 6149 29888 6213 29892
rect 6229 29948 6293 29952
rect 6229 29892 6233 29948
rect 6233 29892 6289 29948
rect 6289 29892 6293 29948
rect 6229 29888 6293 29892
rect 9347 29948 9411 29952
rect 9347 29892 9351 29948
rect 9351 29892 9407 29948
rect 9407 29892 9411 29948
rect 9347 29888 9411 29892
rect 9427 29948 9491 29952
rect 9427 29892 9431 29948
rect 9431 29892 9487 29948
rect 9487 29892 9491 29948
rect 9427 29888 9491 29892
rect 9507 29948 9571 29952
rect 9507 29892 9511 29948
rect 9511 29892 9567 29948
rect 9567 29892 9571 29948
rect 9507 29888 9571 29892
rect 9587 29948 9651 29952
rect 9587 29892 9591 29948
rect 9591 29892 9647 29948
rect 9647 29892 9651 29948
rect 9587 29888 9651 29892
rect 12705 29948 12769 29952
rect 12705 29892 12709 29948
rect 12709 29892 12765 29948
rect 12765 29892 12769 29948
rect 12705 29888 12769 29892
rect 12785 29948 12849 29952
rect 12785 29892 12789 29948
rect 12789 29892 12845 29948
rect 12845 29892 12849 29948
rect 12785 29888 12849 29892
rect 12865 29948 12929 29952
rect 12865 29892 12869 29948
rect 12869 29892 12925 29948
rect 12925 29892 12929 29948
rect 12865 29888 12929 29892
rect 12945 29948 13009 29952
rect 12945 29892 12949 29948
rect 12949 29892 13005 29948
rect 13005 29892 13009 29948
rect 12945 29888 13009 29892
rect 4310 29404 4374 29408
rect 4310 29348 4314 29404
rect 4314 29348 4370 29404
rect 4370 29348 4374 29404
rect 4310 29344 4374 29348
rect 4390 29404 4454 29408
rect 4390 29348 4394 29404
rect 4394 29348 4450 29404
rect 4450 29348 4454 29404
rect 4390 29344 4454 29348
rect 4470 29404 4534 29408
rect 4470 29348 4474 29404
rect 4474 29348 4530 29404
rect 4530 29348 4534 29404
rect 4470 29344 4534 29348
rect 4550 29404 4614 29408
rect 4550 29348 4554 29404
rect 4554 29348 4610 29404
rect 4610 29348 4614 29404
rect 4550 29344 4614 29348
rect 7668 29404 7732 29408
rect 7668 29348 7672 29404
rect 7672 29348 7728 29404
rect 7728 29348 7732 29404
rect 7668 29344 7732 29348
rect 7748 29404 7812 29408
rect 7748 29348 7752 29404
rect 7752 29348 7808 29404
rect 7808 29348 7812 29404
rect 7748 29344 7812 29348
rect 7828 29404 7892 29408
rect 7828 29348 7832 29404
rect 7832 29348 7888 29404
rect 7888 29348 7892 29404
rect 7828 29344 7892 29348
rect 7908 29404 7972 29408
rect 7908 29348 7912 29404
rect 7912 29348 7968 29404
rect 7968 29348 7972 29404
rect 7908 29344 7972 29348
rect 11026 29404 11090 29408
rect 11026 29348 11030 29404
rect 11030 29348 11086 29404
rect 11086 29348 11090 29404
rect 11026 29344 11090 29348
rect 11106 29404 11170 29408
rect 11106 29348 11110 29404
rect 11110 29348 11166 29404
rect 11166 29348 11170 29404
rect 11106 29344 11170 29348
rect 11186 29404 11250 29408
rect 11186 29348 11190 29404
rect 11190 29348 11246 29404
rect 11246 29348 11250 29404
rect 11186 29344 11250 29348
rect 11266 29404 11330 29408
rect 11266 29348 11270 29404
rect 11270 29348 11326 29404
rect 11326 29348 11330 29404
rect 11266 29344 11330 29348
rect 14384 29404 14448 29408
rect 14384 29348 14388 29404
rect 14388 29348 14444 29404
rect 14444 29348 14448 29404
rect 14384 29344 14448 29348
rect 14464 29404 14528 29408
rect 14464 29348 14468 29404
rect 14468 29348 14524 29404
rect 14524 29348 14528 29404
rect 14464 29344 14528 29348
rect 14544 29404 14608 29408
rect 14544 29348 14548 29404
rect 14548 29348 14604 29404
rect 14604 29348 14608 29404
rect 14544 29344 14608 29348
rect 14624 29404 14688 29408
rect 14624 29348 14628 29404
rect 14628 29348 14684 29404
rect 14684 29348 14688 29404
rect 14624 29344 14688 29348
rect 11468 29140 11532 29204
rect 9076 29064 9140 29068
rect 9076 29008 9126 29064
rect 9126 29008 9140 29064
rect 9076 29004 9140 29008
rect 12388 28868 12452 28932
rect 2631 28860 2695 28864
rect 2631 28804 2635 28860
rect 2635 28804 2691 28860
rect 2691 28804 2695 28860
rect 2631 28800 2695 28804
rect 2711 28860 2775 28864
rect 2711 28804 2715 28860
rect 2715 28804 2771 28860
rect 2771 28804 2775 28860
rect 2711 28800 2775 28804
rect 2791 28860 2855 28864
rect 2791 28804 2795 28860
rect 2795 28804 2851 28860
rect 2851 28804 2855 28860
rect 2791 28800 2855 28804
rect 2871 28860 2935 28864
rect 2871 28804 2875 28860
rect 2875 28804 2931 28860
rect 2931 28804 2935 28860
rect 2871 28800 2935 28804
rect 5989 28860 6053 28864
rect 5989 28804 5993 28860
rect 5993 28804 6049 28860
rect 6049 28804 6053 28860
rect 5989 28800 6053 28804
rect 6069 28860 6133 28864
rect 6069 28804 6073 28860
rect 6073 28804 6129 28860
rect 6129 28804 6133 28860
rect 6069 28800 6133 28804
rect 6149 28860 6213 28864
rect 6149 28804 6153 28860
rect 6153 28804 6209 28860
rect 6209 28804 6213 28860
rect 6149 28800 6213 28804
rect 6229 28860 6293 28864
rect 6229 28804 6233 28860
rect 6233 28804 6289 28860
rect 6289 28804 6293 28860
rect 6229 28800 6293 28804
rect 9347 28860 9411 28864
rect 9347 28804 9351 28860
rect 9351 28804 9407 28860
rect 9407 28804 9411 28860
rect 9347 28800 9411 28804
rect 9427 28860 9491 28864
rect 9427 28804 9431 28860
rect 9431 28804 9487 28860
rect 9487 28804 9491 28860
rect 9427 28800 9491 28804
rect 9507 28860 9571 28864
rect 9507 28804 9511 28860
rect 9511 28804 9567 28860
rect 9567 28804 9571 28860
rect 9507 28800 9571 28804
rect 9587 28860 9651 28864
rect 9587 28804 9591 28860
rect 9591 28804 9647 28860
rect 9647 28804 9651 28860
rect 9587 28800 9651 28804
rect 12705 28860 12769 28864
rect 12705 28804 12709 28860
rect 12709 28804 12765 28860
rect 12765 28804 12769 28860
rect 12705 28800 12769 28804
rect 12785 28860 12849 28864
rect 12785 28804 12789 28860
rect 12789 28804 12845 28860
rect 12845 28804 12849 28860
rect 12785 28800 12849 28804
rect 12865 28860 12929 28864
rect 12865 28804 12869 28860
rect 12869 28804 12925 28860
rect 12925 28804 12929 28860
rect 12865 28800 12929 28804
rect 12945 28860 13009 28864
rect 12945 28804 12949 28860
rect 12949 28804 13005 28860
rect 13005 28804 13009 28860
rect 12945 28800 13009 28804
rect 12020 28792 12084 28796
rect 12020 28736 12034 28792
rect 12034 28736 12084 28792
rect 12020 28732 12084 28736
rect 4310 28316 4374 28320
rect 4310 28260 4314 28316
rect 4314 28260 4370 28316
rect 4370 28260 4374 28316
rect 4310 28256 4374 28260
rect 4390 28316 4454 28320
rect 4390 28260 4394 28316
rect 4394 28260 4450 28316
rect 4450 28260 4454 28316
rect 4390 28256 4454 28260
rect 4470 28316 4534 28320
rect 4470 28260 4474 28316
rect 4474 28260 4530 28316
rect 4530 28260 4534 28316
rect 4470 28256 4534 28260
rect 4550 28316 4614 28320
rect 4550 28260 4554 28316
rect 4554 28260 4610 28316
rect 4610 28260 4614 28316
rect 4550 28256 4614 28260
rect 7668 28316 7732 28320
rect 7668 28260 7672 28316
rect 7672 28260 7728 28316
rect 7728 28260 7732 28316
rect 7668 28256 7732 28260
rect 7748 28316 7812 28320
rect 7748 28260 7752 28316
rect 7752 28260 7808 28316
rect 7808 28260 7812 28316
rect 7748 28256 7812 28260
rect 7828 28316 7892 28320
rect 7828 28260 7832 28316
rect 7832 28260 7888 28316
rect 7888 28260 7892 28316
rect 7828 28256 7892 28260
rect 7908 28316 7972 28320
rect 7908 28260 7912 28316
rect 7912 28260 7968 28316
rect 7968 28260 7972 28316
rect 7908 28256 7972 28260
rect 11026 28316 11090 28320
rect 11026 28260 11030 28316
rect 11030 28260 11086 28316
rect 11086 28260 11090 28316
rect 11026 28256 11090 28260
rect 11106 28316 11170 28320
rect 11106 28260 11110 28316
rect 11110 28260 11166 28316
rect 11166 28260 11170 28316
rect 11106 28256 11170 28260
rect 11186 28316 11250 28320
rect 11186 28260 11190 28316
rect 11190 28260 11246 28316
rect 11246 28260 11250 28316
rect 11186 28256 11250 28260
rect 11266 28316 11330 28320
rect 11266 28260 11270 28316
rect 11270 28260 11326 28316
rect 11326 28260 11330 28316
rect 11266 28256 11330 28260
rect 14384 28316 14448 28320
rect 14384 28260 14388 28316
rect 14388 28260 14444 28316
rect 14444 28260 14448 28316
rect 14384 28256 14448 28260
rect 14464 28316 14528 28320
rect 14464 28260 14468 28316
rect 14468 28260 14524 28316
rect 14524 28260 14528 28316
rect 14464 28256 14528 28260
rect 14544 28316 14608 28320
rect 14544 28260 14548 28316
rect 14548 28260 14604 28316
rect 14604 28260 14608 28316
rect 14544 28256 14608 28260
rect 14624 28316 14688 28320
rect 14624 28260 14628 28316
rect 14628 28260 14684 28316
rect 14684 28260 14688 28316
rect 14624 28256 14688 28260
rect 8524 28052 8588 28116
rect 14044 28188 14108 28252
rect 12020 27840 12084 27844
rect 12020 27784 12034 27840
rect 12034 27784 12084 27840
rect 12020 27780 12084 27784
rect 2631 27772 2695 27776
rect 2631 27716 2635 27772
rect 2635 27716 2691 27772
rect 2691 27716 2695 27772
rect 2631 27712 2695 27716
rect 2711 27772 2775 27776
rect 2711 27716 2715 27772
rect 2715 27716 2771 27772
rect 2771 27716 2775 27772
rect 2711 27712 2775 27716
rect 2791 27772 2855 27776
rect 2791 27716 2795 27772
rect 2795 27716 2851 27772
rect 2851 27716 2855 27772
rect 2791 27712 2855 27716
rect 2871 27772 2935 27776
rect 2871 27716 2875 27772
rect 2875 27716 2931 27772
rect 2931 27716 2935 27772
rect 2871 27712 2935 27716
rect 5989 27772 6053 27776
rect 5989 27716 5993 27772
rect 5993 27716 6049 27772
rect 6049 27716 6053 27772
rect 5989 27712 6053 27716
rect 6069 27772 6133 27776
rect 6069 27716 6073 27772
rect 6073 27716 6129 27772
rect 6129 27716 6133 27772
rect 6069 27712 6133 27716
rect 6149 27772 6213 27776
rect 6149 27716 6153 27772
rect 6153 27716 6209 27772
rect 6209 27716 6213 27772
rect 6149 27712 6213 27716
rect 6229 27772 6293 27776
rect 6229 27716 6233 27772
rect 6233 27716 6289 27772
rect 6289 27716 6293 27772
rect 6229 27712 6293 27716
rect 9347 27772 9411 27776
rect 9347 27716 9351 27772
rect 9351 27716 9407 27772
rect 9407 27716 9411 27772
rect 9347 27712 9411 27716
rect 9427 27772 9491 27776
rect 9427 27716 9431 27772
rect 9431 27716 9487 27772
rect 9487 27716 9491 27772
rect 9427 27712 9491 27716
rect 9507 27772 9571 27776
rect 9507 27716 9511 27772
rect 9511 27716 9567 27772
rect 9567 27716 9571 27772
rect 9507 27712 9571 27716
rect 9587 27772 9651 27776
rect 9587 27716 9591 27772
rect 9591 27716 9647 27772
rect 9647 27716 9651 27772
rect 9587 27712 9651 27716
rect 12705 27772 12769 27776
rect 12705 27716 12709 27772
rect 12709 27716 12765 27772
rect 12765 27716 12769 27772
rect 12705 27712 12769 27716
rect 12785 27772 12849 27776
rect 12785 27716 12789 27772
rect 12789 27716 12845 27772
rect 12845 27716 12849 27772
rect 12785 27712 12849 27716
rect 12865 27772 12929 27776
rect 12865 27716 12869 27772
rect 12869 27716 12925 27772
rect 12925 27716 12929 27772
rect 12865 27712 12929 27716
rect 12945 27772 13009 27776
rect 12945 27716 12949 27772
rect 12949 27716 13005 27772
rect 13005 27716 13009 27772
rect 12945 27712 13009 27716
rect 8892 27644 8956 27708
rect 12020 27644 12084 27708
rect 14228 27644 14292 27708
rect 4310 27228 4374 27232
rect 4310 27172 4314 27228
rect 4314 27172 4370 27228
rect 4370 27172 4374 27228
rect 4310 27168 4374 27172
rect 4390 27228 4454 27232
rect 4390 27172 4394 27228
rect 4394 27172 4450 27228
rect 4450 27172 4454 27228
rect 4390 27168 4454 27172
rect 4470 27228 4534 27232
rect 4470 27172 4474 27228
rect 4474 27172 4530 27228
rect 4530 27172 4534 27228
rect 4470 27168 4534 27172
rect 4550 27228 4614 27232
rect 4550 27172 4554 27228
rect 4554 27172 4610 27228
rect 4610 27172 4614 27228
rect 4550 27168 4614 27172
rect 7668 27228 7732 27232
rect 7668 27172 7672 27228
rect 7672 27172 7728 27228
rect 7728 27172 7732 27228
rect 7668 27168 7732 27172
rect 7748 27228 7812 27232
rect 7748 27172 7752 27228
rect 7752 27172 7808 27228
rect 7808 27172 7812 27228
rect 7748 27168 7812 27172
rect 7828 27228 7892 27232
rect 7828 27172 7832 27228
rect 7832 27172 7888 27228
rect 7888 27172 7892 27228
rect 7828 27168 7892 27172
rect 7908 27228 7972 27232
rect 7908 27172 7912 27228
rect 7912 27172 7968 27228
rect 7968 27172 7972 27228
rect 7908 27168 7972 27172
rect 11026 27228 11090 27232
rect 11026 27172 11030 27228
rect 11030 27172 11086 27228
rect 11086 27172 11090 27228
rect 11026 27168 11090 27172
rect 11106 27228 11170 27232
rect 11106 27172 11110 27228
rect 11110 27172 11166 27228
rect 11166 27172 11170 27228
rect 11106 27168 11170 27172
rect 11186 27228 11250 27232
rect 11186 27172 11190 27228
rect 11190 27172 11246 27228
rect 11246 27172 11250 27228
rect 11186 27168 11250 27172
rect 11266 27228 11330 27232
rect 11266 27172 11270 27228
rect 11270 27172 11326 27228
rect 11326 27172 11330 27228
rect 11266 27168 11330 27172
rect 14384 27228 14448 27232
rect 14384 27172 14388 27228
rect 14388 27172 14444 27228
rect 14444 27172 14448 27228
rect 14384 27168 14448 27172
rect 14464 27228 14528 27232
rect 14464 27172 14468 27228
rect 14468 27172 14524 27228
rect 14524 27172 14528 27228
rect 14464 27168 14528 27172
rect 14544 27228 14608 27232
rect 14544 27172 14548 27228
rect 14548 27172 14604 27228
rect 14604 27172 14608 27228
rect 14544 27168 14608 27172
rect 14624 27228 14688 27232
rect 14624 27172 14628 27228
rect 14628 27172 14684 27228
rect 14684 27172 14688 27228
rect 14624 27168 14688 27172
rect 12572 27100 12636 27164
rect 11836 26692 11900 26756
rect 2631 26684 2695 26688
rect 2631 26628 2635 26684
rect 2635 26628 2691 26684
rect 2691 26628 2695 26684
rect 2631 26624 2695 26628
rect 2711 26684 2775 26688
rect 2711 26628 2715 26684
rect 2715 26628 2771 26684
rect 2771 26628 2775 26684
rect 2711 26624 2775 26628
rect 2791 26684 2855 26688
rect 2791 26628 2795 26684
rect 2795 26628 2851 26684
rect 2851 26628 2855 26684
rect 2791 26624 2855 26628
rect 2871 26684 2935 26688
rect 2871 26628 2875 26684
rect 2875 26628 2931 26684
rect 2931 26628 2935 26684
rect 2871 26624 2935 26628
rect 5989 26684 6053 26688
rect 5989 26628 5993 26684
rect 5993 26628 6049 26684
rect 6049 26628 6053 26684
rect 5989 26624 6053 26628
rect 6069 26684 6133 26688
rect 6069 26628 6073 26684
rect 6073 26628 6129 26684
rect 6129 26628 6133 26684
rect 6069 26624 6133 26628
rect 6149 26684 6213 26688
rect 6149 26628 6153 26684
rect 6153 26628 6209 26684
rect 6209 26628 6213 26684
rect 6149 26624 6213 26628
rect 6229 26684 6293 26688
rect 6229 26628 6233 26684
rect 6233 26628 6289 26684
rect 6289 26628 6293 26684
rect 6229 26624 6293 26628
rect 9347 26684 9411 26688
rect 9347 26628 9351 26684
rect 9351 26628 9407 26684
rect 9407 26628 9411 26684
rect 9347 26624 9411 26628
rect 9427 26684 9491 26688
rect 9427 26628 9431 26684
rect 9431 26628 9487 26684
rect 9487 26628 9491 26684
rect 9427 26624 9491 26628
rect 9507 26684 9571 26688
rect 9507 26628 9511 26684
rect 9511 26628 9567 26684
rect 9567 26628 9571 26684
rect 9507 26624 9571 26628
rect 9587 26684 9651 26688
rect 9587 26628 9591 26684
rect 9591 26628 9647 26684
rect 9647 26628 9651 26684
rect 9587 26624 9651 26628
rect 12705 26684 12769 26688
rect 12705 26628 12709 26684
rect 12709 26628 12765 26684
rect 12765 26628 12769 26684
rect 12705 26624 12769 26628
rect 12785 26684 12849 26688
rect 12785 26628 12789 26684
rect 12789 26628 12845 26684
rect 12845 26628 12849 26684
rect 12785 26624 12849 26628
rect 12865 26684 12929 26688
rect 12865 26628 12869 26684
rect 12869 26628 12925 26684
rect 12925 26628 12929 26684
rect 12865 26624 12929 26628
rect 12945 26684 13009 26688
rect 12945 26628 12949 26684
rect 12949 26628 13005 26684
rect 13005 26628 13009 26684
rect 12945 26624 13009 26628
rect 7420 26284 7484 26348
rect 4310 26140 4374 26144
rect 4310 26084 4314 26140
rect 4314 26084 4370 26140
rect 4370 26084 4374 26140
rect 4310 26080 4374 26084
rect 4390 26140 4454 26144
rect 4390 26084 4394 26140
rect 4394 26084 4450 26140
rect 4450 26084 4454 26140
rect 4390 26080 4454 26084
rect 4470 26140 4534 26144
rect 4470 26084 4474 26140
rect 4474 26084 4530 26140
rect 4530 26084 4534 26140
rect 4470 26080 4534 26084
rect 4550 26140 4614 26144
rect 4550 26084 4554 26140
rect 4554 26084 4610 26140
rect 4610 26084 4614 26140
rect 4550 26080 4614 26084
rect 7668 26140 7732 26144
rect 7668 26084 7672 26140
rect 7672 26084 7728 26140
rect 7728 26084 7732 26140
rect 7668 26080 7732 26084
rect 7748 26140 7812 26144
rect 7748 26084 7752 26140
rect 7752 26084 7808 26140
rect 7808 26084 7812 26140
rect 7748 26080 7812 26084
rect 7828 26140 7892 26144
rect 7828 26084 7832 26140
rect 7832 26084 7888 26140
rect 7888 26084 7892 26140
rect 7828 26080 7892 26084
rect 7908 26140 7972 26144
rect 7908 26084 7912 26140
rect 7912 26084 7968 26140
rect 7968 26084 7972 26140
rect 7908 26080 7972 26084
rect 11026 26140 11090 26144
rect 11026 26084 11030 26140
rect 11030 26084 11086 26140
rect 11086 26084 11090 26140
rect 11026 26080 11090 26084
rect 11106 26140 11170 26144
rect 11106 26084 11110 26140
rect 11110 26084 11166 26140
rect 11166 26084 11170 26140
rect 11106 26080 11170 26084
rect 11186 26140 11250 26144
rect 11186 26084 11190 26140
rect 11190 26084 11246 26140
rect 11246 26084 11250 26140
rect 11186 26080 11250 26084
rect 11266 26140 11330 26144
rect 11266 26084 11270 26140
rect 11270 26084 11326 26140
rect 11326 26084 11330 26140
rect 11266 26080 11330 26084
rect 14384 26140 14448 26144
rect 14384 26084 14388 26140
rect 14388 26084 14444 26140
rect 14444 26084 14448 26140
rect 14384 26080 14448 26084
rect 14464 26140 14528 26144
rect 14464 26084 14468 26140
rect 14468 26084 14524 26140
rect 14524 26084 14528 26140
rect 14464 26080 14528 26084
rect 14544 26140 14608 26144
rect 14544 26084 14548 26140
rect 14548 26084 14604 26140
rect 14604 26084 14608 26140
rect 14544 26080 14608 26084
rect 14624 26140 14688 26144
rect 14624 26084 14628 26140
rect 14628 26084 14684 26140
rect 14684 26084 14688 26140
rect 14624 26080 14688 26084
rect 10364 25876 10428 25940
rect 12388 25936 12452 25940
rect 12388 25880 12438 25936
rect 12438 25880 12452 25936
rect 12388 25876 12452 25880
rect 2631 25596 2695 25600
rect 2631 25540 2635 25596
rect 2635 25540 2691 25596
rect 2691 25540 2695 25596
rect 2631 25536 2695 25540
rect 2711 25596 2775 25600
rect 2711 25540 2715 25596
rect 2715 25540 2771 25596
rect 2771 25540 2775 25596
rect 2711 25536 2775 25540
rect 2791 25596 2855 25600
rect 2791 25540 2795 25596
rect 2795 25540 2851 25596
rect 2851 25540 2855 25596
rect 2791 25536 2855 25540
rect 2871 25596 2935 25600
rect 2871 25540 2875 25596
rect 2875 25540 2931 25596
rect 2931 25540 2935 25596
rect 2871 25536 2935 25540
rect 5989 25596 6053 25600
rect 5989 25540 5993 25596
rect 5993 25540 6049 25596
rect 6049 25540 6053 25596
rect 5989 25536 6053 25540
rect 6069 25596 6133 25600
rect 6069 25540 6073 25596
rect 6073 25540 6129 25596
rect 6129 25540 6133 25596
rect 6069 25536 6133 25540
rect 6149 25596 6213 25600
rect 6149 25540 6153 25596
rect 6153 25540 6209 25596
rect 6209 25540 6213 25596
rect 6149 25536 6213 25540
rect 6229 25596 6293 25600
rect 6229 25540 6233 25596
rect 6233 25540 6289 25596
rect 6289 25540 6293 25596
rect 6229 25536 6293 25540
rect 9347 25596 9411 25600
rect 9347 25540 9351 25596
rect 9351 25540 9407 25596
rect 9407 25540 9411 25596
rect 9347 25536 9411 25540
rect 9427 25596 9491 25600
rect 9427 25540 9431 25596
rect 9431 25540 9487 25596
rect 9487 25540 9491 25596
rect 9427 25536 9491 25540
rect 9507 25596 9571 25600
rect 9507 25540 9511 25596
rect 9511 25540 9567 25596
rect 9567 25540 9571 25596
rect 9507 25536 9571 25540
rect 9587 25596 9651 25600
rect 9587 25540 9591 25596
rect 9591 25540 9647 25596
rect 9647 25540 9651 25596
rect 9587 25536 9651 25540
rect 12705 25596 12769 25600
rect 12705 25540 12709 25596
rect 12709 25540 12765 25596
rect 12765 25540 12769 25596
rect 12705 25536 12769 25540
rect 12785 25596 12849 25600
rect 12785 25540 12789 25596
rect 12789 25540 12845 25596
rect 12845 25540 12849 25596
rect 12785 25536 12849 25540
rect 12865 25596 12929 25600
rect 12865 25540 12869 25596
rect 12869 25540 12925 25596
rect 12925 25540 12929 25596
rect 12865 25536 12929 25540
rect 12945 25596 13009 25600
rect 12945 25540 12949 25596
rect 12949 25540 13005 25596
rect 13005 25540 13009 25596
rect 12945 25536 13009 25540
rect 10732 25332 10796 25396
rect 4310 25052 4374 25056
rect 4310 24996 4314 25052
rect 4314 24996 4370 25052
rect 4370 24996 4374 25052
rect 4310 24992 4374 24996
rect 4390 25052 4454 25056
rect 4390 24996 4394 25052
rect 4394 24996 4450 25052
rect 4450 24996 4454 25052
rect 4390 24992 4454 24996
rect 4470 25052 4534 25056
rect 4470 24996 4474 25052
rect 4474 24996 4530 25052
rect 4530 24996 4534 25052
rect 4470 24992 4534 24996
rect 4550 25052 4614 25056
rect 4550 24996 4554 25052
rect 4554 24996 4610 25052
rect 4610 24996 4614 25052
rect 4550 24992 4614 24996
rect 7668 25052 7732 25056
rect 7668 24996 7672 25052
rect 7672 24996 7728 25052
rect 7728 24996 7732 25052
rect 7668 24992 7732 24996
rect 7748 25052 7812 25056
rect 7748 24996 7752 25052
rect 7752 24996 7808 25052
rect 7808 24996 7812 25052
rect 7748 24992 7812 24996
rect 7828 25052 7892 25056
rect 7828 24996 7832 25052
rect 7832 24996 7888 25052
rect 7888 24996 7892 25052
rect 7828 24992 7892 24996
rect 7908 25052 7972 25056
rect 7908 24996 7912 25052
rect 7912 24996 7968 25052
rect 7968 24996 7972 25052
rect 7908 24992 7972 24996
rect 11026 25052 11090 25056
rect 11026 24996 11030 25052
rect 11030 24996 11086 25052
rect 11086 24996 11090 25052
rect 11026 24992 11090 24996
rect 11106 25052 11170 25056
rect 11106 24996 11110 25052
rect 11110 24996 11166 25052
rect 11166 24996 11170 25052
rect 11106 24992 11170 24996
rect 11186 25052 11250 25056
rect 11186 24996 11190 25052
rect 11190 24996 11246 25052
rect 11246 24996 11250 25052
rect 11186 24992 11250 24996
rect 11266 25052 11330 25056
rect 11266 24996 11270 25052
rect 11270 24996 11326 25052
rect 11326 24996 11330 25052
rect 11266 24992 11330 24996
rect 14384 25052 14448 25056
rect 14384 24996 14388 25052
rect 14388 24996 14444 25052
rect 14444 24996 14448 25052
rect 14384 24992 14448 24996
rect 14464 25052 14528 25056
rect 14464 24996 14468 25052
rect 14468 24996 14524 25052
rect 14524 24996 14528 25052
rect 14464 24992 14528 24996
rect 14544 25052 14608 25056
rect 14544 24996 14548 25052
rect 14548 24996 14604 25052
rect 14604 24996 14608 25052
rect 14544 24992 14608 24996
rect 14624 25052 14688 25056
rect 14624 24996 14628 25052
rect 14628 24996 14684 25052
rect 14684 24996 14688 25052
rect 14624 24992 14688 24996
rect 13676 24924 13740 24988
rect 2631 24508 2695 24512
rect 2631 24452 2635 24508
rect 2635 24452 2691 24508
rect 2691 24452 2695 24508
rect 2631 24448 2695 24452
rect 2711 24508 2775 24512
rect 2711 24452 2715 24508
rect 2715 24452 2771 24508
rect 2771 24452 2775 24508
rect 2711 24448 2775 24452
rect 2791 24508 2855 24512
rect 2791 24452 2795 24508
rect 2795 24452 2851 24508
rect 2851 24452 2855 24508
rect 2791 24448 2855 24452
rect 2871 24508 2935 24512
rect 2871 24452 2875 24508
rect 2875 24452 2931 24508
rect 2931 24452 2935 24508
rect 2871 24448 2935 24452
rect 5989 24508 6053 24512
rect 5989 24452 5993 24508
rect 5993 24452 6049 24508
rect 6049 24452 6053 24508
rect 5989 24448 6053 24452
rect 6069 24508 6133 24512
rect 6069 24452 6073 24508
rect 6073 24452 6129 24508
rect 6129 24452 6133 24508
rect 6069 24448 6133 24452
rect 6149 24508 6213 24512
rect 6149 24452 6153 24508
rect 6153 24452 6209 24508
rect 6209 24452 6213 24508
rect 6149 24448 6213 24452
rect 6229 24508 6293 24512
rect 6229 24452 6233 24508
rect 6233 24452 6289 24508
rect 6289 24452 6293 24508
rect 6229 24448 6293 24452
rect 9347 24508 9411 24512
rect 9347 24452 9351 24508
rect 9351 24452 9407 24508
rect 9407 24452 9411 24508
rect 9347 24448 9411 24452
rect 9427 24508 9491 24512
rect 9427 24452 9431 24508
rect 9431 24452 9487 24508
rect 9487 24452 9491 24508
rect 9427 24448 9491 24452
rect 9507 24508 9571 24512
rect 9507 24452 9511 24508
rect 9511 24452 9567 24508
rect 9567 24452 9571 24508
rect 9507 24448 9571 24452
rect 9587 24508 9651 24512
rect 9587 24452 9591 24508
rect 9591 24452 9647 24508
rect 9647 24452 9651 24508
rect 9587 24448 9651 24452
rect 12705 24508 12769 24512
rect 12705 24452 12709 24508
rect 12709 24452 12765 24508
rect 12765 24452 12769 24508
rect 12705 24448 12769 24452
rect 12785 24508 12849 24512
rect 12785 24452 12789 24508
rect 12789 24452 12845 24508
rect 12845 24452 12849 24508
rect 12785 24448 12849 24452
rect 12865 24508 12929 24512
rect 12865 24452 12869 24508
rect 12869 24452 12925 24508
rect 12925 24452 12929 24508
rect 12865 24448 12929 24452
rect 12945 24508 13009 24512
rect 12945 24452 12949 24508
rect 12949 24452 13005 24508
rect 13005 24452 13009 24508
rect 12945 24448 13009 24452
rect 10732 24108 10796 24172
rect 4310 23964 4374 23968
rect 4310 23908 4314 23964
rect 4314 23908 4370 23964
rect 4370 23908 4374 23964
rect 4310 23904 4374 23908
rect 4390 23964 4454 23968
rect 4390 23908 4394 23964
rect 4394 23908 4450 23964
rect 4450 23908 4454 23964
rect 4390 23904 4454 23908
rect 4470 23964 4534 23968
rect 4470 23908 4474 23964
rect 4474 23908 4530 23964
rect 4530 23908 4534 23964
rect 4470 23904 4534 23908
rect 4550 23964 4614 23968
rect 4550 23908 4554 23964
rect 4554 23908 4610 23964
rect 4610 23908 4614 23964
rect 4550 23904 4614 23908
rect 7668 23964 7732 23968
rect 7668 23908 7672 23964
rect 7672 23908 7728 23964
rect 7728 23908 7732 23964
rect 7668 23904 7732 23908
rect 7748 23964 7812 23968
rect 7748 23908 7752 23964
rect 7752 23908 7808 23964
rect 7808 23908 7812 23964
rect 7748 23904 7812 23908
rect 7828 23964 7892 23968
rect 7828 23908 7832 23964
rect 7832 23908 7888 23964
rect 7888 23908 7892 23964
rect 7828 23904 7892 23908
rect 7908 23964 7972 23968
rect 7908 23908 7912 23964
rect 7912 23908 7968 23964
rect 7968 23908 7972 23964
rect 7908 23904 7972 23908
rect 11026 23964 11090 23968
rect 11026 23908 11030 23964
rect 11030 23908 11086 23964
rect 11086 23908 11090 23964
rect 11026 23904 11090 23908
rect 11106 23964 11170 23968
rect 11106 23908 11110 23964
rect 11110 23908 11166 23964
rect 11166 23908 11170 23964
rect 11106 23904 11170 23908
rect 11186 23964 11250 23968
rect 11186 23908 11190 23964
rect 11190 23908 11246 23964
rect 11246 23908 11250 23964
rect 11186 23904 11250 23908
rect 11266 23964 11330 23968
rect 11266 23908 11270 23964
rect 11270 23908 11326 23964
rect 11326 23908 11330 23964
rect 11266 23904 11330 23908
rect 14384 23964 14448 23968
rect 14384 23908 14388 23964
rect 14388 23908 14444 23964
rect 14444 23908 14448 23964
rect 14384 23904 14448 23908
rect 14464 23964 14528 23968
rect 14464 23908 14468 23964
rect 14468 23908 14524 23964
rect 14524 23908 14528 23964
rect 14464 23904 14528 23908
rect 14544 23964 14608 23968
rect 14544 23908 14548 23964
rect 14548 23908 14604 23964
rect 14604 23908 14608 23964
rect 14544 23904 14608 23908
rect 14624 23964 14688 23968
rect 14624 23908 14628 23964
rect 14628 23908 14684 23964
rect 14684 23908 14688 23964
rect 14624 23904 14688 23908
rect 8156 23564 8220 23628
rect 8524 23564 8588 23628
rect 2631 23420 2695 23424
rect 2631 23364 2635 23420
rect 2635 23364 2691 23420
rect 2691 23364 2695 23420
rect 2631 23360 2695 23364
rect 2711 23420 2775 23424
rect 2711 23364 2715 23420
rect 2715 23364 2771 23420
rect 2771 23364 2775 23420
rect 2711 23360 2775 23364
rect 2791 23420 2855 23424
rect 2791 23364 2795 23420
rect 2795 23364 2851 23420
rect 2851 23364 2855 23420
rect 2791 23360 2855 23364
rect 2871 23420 2935 23424
rect 2871 23364 2875 23420
rect 2875 23364 2931 23420
rect 2931 23364 2935 23420
rect 2871 23360 2935 23364
rect 5989 23420 6053 23424
rect 5989 23364 5993 23420
rect 5993 23364 6049 23420
rect 6049 23364 6053 23420
rect 5989 23360 6053 23364
rect 6069 23420 6133 23424
rect 6069 23364 6073 23420
rect 6073 23364 6129 23420
rect 6129 23364 6133 23420
rect 6069 23360 6133 23364
rect 6149 23420 6213 23424
rect 6149 23364 6153 23420
rect 6153 23364 6209 23420
rect 6209 23364 6213 23420
rect 6149 23360 6213 23364
rect 6229 23420 6293 23424
rect 6229 23364 6233 23420
rect 6233 23364 6289 23420
rect 6289 23364 6293 23420
rect 6229 23360 6293 23364
rect 9347 23420 9411 23424
rect 9347 23364 9351 23420
rect 9351 23364 9407 23420
rect 9407 23364 9411 23420
rect 9347 23360 9411 23364
rect 9427 23420 9491 23424
rect 9427 23364 9431 23420
rect 9431 23364 9487 23420
rect 9487 23364 9491 23420
rect 9427 23360 9491 23364
rect 9507 23420 9571 23424
rect 9507 23364 9511 23420
rect 9511 23364 9567 23420
rect 9567 23364 9571 23420
rect 9507 23360 9571 23364
rect 9587 23420 9651 23424
rect 9587 23364 9591 23420
rect 9591 23364 9647 23420
rect 9647 23364 9651 23420
rect 9587 23360 9651 23364
rect 12705 23420 12769 23424
rect 12705 23364 12709 23420
rect 12709 23364 12765 23420
rect 12765 23364 12769 23420
rect 12705 23360 12769 23364
rect 12785 23420 12849 23424
rect 12785 23364 12789 23420
rect 12789 23364 12845 23420
rect 12845 23364 12849 23420
rect 12785 23360 12849 23364
rect 12865 23420 12929 23424
rect 12865 23364 12869 23420
rect 12869 23364 12925 23420
rect 12925 23364 12929 23420
rect 12865 23360 12929 23364
rect 12945 23420 13009 23424
rect 12945 23364 12949 23420
rect 12949 23364 13005 23420
rect 13005 23364 13009 23420
rect 12945 23360 13009 23364
rect 4310 22876 4374 22880
rect 4310 22820 4314 22876
rect 4314 22820 4370 22876
rect 4370 22820 4374 22876
rect 4310 22816 4374 22820
rect 4390 22876 4454 22880
rect 4390 22820 4394 22876
rect 4394 22820 4450 22876
rect 4450 22820 4454 22876
rect 4390 22816 4454 22820
rect 4470 22876 4534 22880
rect 4470 22820 4474 22876
rect 4474 22820 4530 22876
rect 4530 22820 4534 22876
rect 4470 22816 4534 22820
rect 4550 22876 4614 22880
rect 4550 22820 4554 22876
rect 4554 22820 4610 22876
rect 4610 22820 4614 22876
rect 4550 22816 4614 22820
rect 7668 22876 7732 22880
rect 7668 22820 7672 22876
rect 7672 22820 7728 22876
rect 7728 22820 7732 22876
rect 7668 22816 7732 22820
rect 7748 22876 7812 22880
rect 7748 22820 7752 22876
rect 7752 22820 7808 22876
rect 7808 22820 7812 22876
rect 7748 22816 7812 22820
rect 7828 22876 7892 22880
rect 7828 22820 7832 22876
rect 7832 22820 7888 22876
rect 7888 22820 7892 22876
rect 7828 22816 7892 22820
rect 7908 22876 7972 22880
rect 7908 22820 7912 22876
rect 7912 22820 7968 22876
rect 7968 22820 7972 22876
rect 7908 22816 7972 22820
rect 11026 22876 11090 22880
rect 11026 22820 11030 22876
rect 11030 22820 11086 22876
rect 11086 22820 11090 22876
rect 11026 22816 11090 22820
rect 11106 22876 11170 22880
rect 11106 22820 11110 22876
rect 11110 22820 11166 22876
rect 11166 22820 11170 22876
rect 11106 22816 11170 22820
rect 11186 22876 11250 22880
rect 11186 22820 11190 22876
rect 11190 22820 11246 22876
rect 11246 22820 11250 22876
rect 11186 22816 11250 22820
rect 11266 22876 11330 22880
rect 11266 22820 11270 22876
rect 11270 22820 11326 22876
rect 11326 22820 11330 22876
rect 11266 22816 11330 22820
rect 14384 22876 14448 22880
rect 14384 22820 14388 22876
rect 14388 22820 14444 22876
rect 14444 22820 14448 22876
rect 14384 22816 14448 22820
rect 14464 22876 14528 22880
rect 14464 22820 14468 22876
rect 14468 22820 14524 22876
rect 14524 22820 14528 22876
rect 14464 22816 14528 22820
rect 14544 22876 14608 22880
rect 14544 22820 14548 22876
rect 14548 22820 14604 22876
rect 14604 22820 14608 22876
rect 14544 22816 14608 22820
rect 14624 22876 14688 22880
rect 14624 22820 14628 22876
rect 14628 22820 14684 22876
rect 14684 22820 14688 22876
rect 14624 22816 14688 22820
rect 8708 22476 8772 22540
rect 9812 22536 9876 22540
rect 9812 22480 9826 22536
rect 9826 22480 9876 22536
rect 9812 22476 9876 22480
rect 15332 22476 15396 22540
rect 2631 22332 2695 22336
rect 2631 22276 2635 22332
rect 2635 22276 2691 22332
rect 2691 22276 2695 22332
rect 2631 22272 2695 22276
rect 2711 22332 2775 22336
rect 2711 22276 2715 22332
rect 2715 22276 2771 22332
rect 2771 22276 2775 22332
rect 2711 22272 2775 22276
rect 2791 22332 2855 22336
rect 2791 22276 2795 22332
rect 2795 22276 2851 22332
rect 2851 22276 2855 22332
rect 2791 22272 2855 22276
rect 2871 22332 2935 22336
rect 2871 22276 2875 22332
rect 2875 22276 2931 22332
rect 2931 22276 2935 22332
rect 2871 22272 2935 22276
rect 5989 22332 6053 22336
rect 5989 22276 5993 22332
rect 5993 22276 6049 22332
rect 6049 22276 6053 22332
rect 5989 22272 6053 22276
rect 6069 22332 6133 22336
rect 6069 22276 6073 22332
rect 6073 22276 6129 22332
rect 6129 22276 6133 22332
rect 6069 22272 6133 22276
rect 6149 22332 6213 22336
rect 6149 22276 6153 22332
rect 6153 22276 6209 22332
rect 6209 22276 6213 22332
rect 6149 22272 6213 22276
rect 6229 22332 6293 22336
rect 6229 22276 6233 22332
rect 6233 22276 6289 22332
rect 6289 22276 6293 22332
rect 6229 22272 6293 22276
rect 9347 22332 9411 22336
rect 9347 22276 9351 22332
rect 9351 22276 9407 22332
rect 9407 22276 9411 22332
rect 9347 22272 9411 22276
rect 9427 22332 9491 22336
rect 9427 22276 9431 22332
rect 9431 22276 9487 22332
rect 9487 22276 9491 22332
rect 9427 22272 9491 22276
rect 9507 22332 9571 22336
rect 9507 22276 9511 22332
rect 9511 22276 9567 22332
rect 9567 22276 9571 22332
rect 9507 22272 9571 22276
rect 9587 22332 9651 22336
rect 9587 22276 9591 22332
rect 9591 22276 9647 22332
rect 9647 22276 9651 22332
rect 9587 22272 9651 22276
rect 12705 22332 12769 22336
rect 12705 22276 12709 22332
rect 12709 22276 12765 22332
rect 12765 22276 12769 22332
rect 12705 22272 12769 22276
rect 12785 22332 12849 22336
rect 12785 22276 12789 22332
rect 12789 22276 12845 22332
rect 12845 22276 12849 22332
rect 12785 22272 12849 22276
rect 12865 22332 12929 22336
rect 12865 22276 12869 22332
rect 12869 22276 12925 22332
rect 12925 22276 12929 22332
rect 12865 22272 12929 22276
rect 12945 22332 13009 22336
rect 12945 22276 12949 22332
rect 12949 22276 13005 22332
rect 13005 22276 13009 22332
rect 12945 22272 13009 22276
rect 7420 21856 7484 21860
rect 7420 21800 7434 21856
rect 7434 21800 7484 21856
rect 7420 21796 7484 21800
rect 4310 21788 4374 21792
rect 4310 21732 4314 21788
rect 4314 21732 4370 21788
rect 4370 21732 4374 21788
rect 4310 21728 4374 21732
rect 4390 21788 4454 21792
rect 4390 21732 4394 21788
rect 4394 21732 4450 21788
rect 4450 21732 4454 21788
rect 4390 21728 4454 21732
rect 4470 21788 4534 21792
rect 4470 21732 4474 21788
rect 4474 21732 4530 21788
rect 4530 21732 4534 21788
rect 4470 21728 4534 21732
rect 4550 21788 4614 21792
rect 4550 21732 4554 21788
rect 4554 21732 4610 21788
rect 4610 21732 4614 21788
rect 4550 21728 4614 21732
rect 7668 21788 7732 21792
rect 7668 21732 7672 21788
rect 7672 21732 7728 21788
rect 7728 21732 7732 21788
rect 7668 21728 7732 21732
rect 7748 21788 7812 21792
rect 7748 21732 7752 21788
rect 7752 21732 7808 21788
rect 7808 21732 7812 21788
rect 7748 21728 7812 21732
rect 7828 21788 7892 21792
rect 7828 21732 7832 21788
rect 7832 21732 7888 21788
rect 7888 21732 7892 21788
rect 7828 21728 7892 21732
rect 7908 21788 7972 21792
rect 7908 21732 7912 21788
rect 7912 21732 7968 21788
rect 7968 21732 7972 21788
rect 7908 21728 7972 21732
rect 11026 21788 11090 21792
rect 11026 21732 11030 21788
rect 11030 21732 11086 21788
rect 11086 21732 11090 21788
rect 11026 21728 11090 21732
rect 11106 21788 11170 21792
rect 11106 21732 11110 21788
rect 11110 21732 11166 21788
rect 11166 21732 11170 21788
rect 11106 21728 11170 21732
rect 11186 21788 11250 21792
rect 11186 21732 11190 21788
rect 11190 21732 11246 21788
rect 11246 21732 11250 21788
rect 11186 21728 11250 21732
rect 11266 21788 11330 21792
rect 11266 21732 11270 21788
rect 11270 21732 11326 21788
rect 11326 21732 11330 21788
rect 11266 21728 11330 21732
rect 14384 21788 14448 21792
rect 14384 21732 14388 21788
rect 14388 21732 14444 21788
rect 14444 21732 14448 21788
rect 14384 21728 14448 21732
rect 14464 21788 14528 21792
rect 14464 21732 14468 21788
rect 14468 21732 14524 21788
rect 14524 21732 14528 21788
rect 14464 21728 14528 21732
rect 14544 21788 14608 21792
rect 14544 21732 14548 21788
rect 14548 21732 14604 21788
rect 14604 21732 14608 21788
rect 14544 21728 14608 21732
rect 14624 21788 14688 21792
rect 14624 21732 14628 21788
rect 14628 21732 14684 21788
rect 14684 21732 14688 21788
rect 14624 21728 14688 21732
rect 15148 21448 15212 21452
rect 15148 21392 15198 21448
rect 15198 21392 15212 21448
rect 15148 21388 15212 21392
rect 2631 21244 2695 21248
rect 2631 21188 2635 21244
rect 2635 21188 2691 21244
rect 2691 21188 2695 21244
rect 2631 21184 2695 21188
rect 2711 21244 2775 21248
rect 2711 21188 2715 21244
rect 2715 21188 2771 21244
rect 2771 21188 2775 21244
rect 2711 21184 2775 21188
rect 2791 21244 2855 21248
rect 2791 21188 2795 21244
rect 2795 21188 2851 21244
rect 2851 21188 2855 21244
rect 2791 21184 2855 21188
rect 2871 21244 2935 21248
rect 2871 21188 2875 21244
rect 2875 21188 2931 21244
rect 2931 21188 2935 21244
rect 2871 21184 2935 21188
rect 5989 21244 6053 21248
rect 5989 21188 5993 21244
rect 5993 21188 6049 21244
rect 6049 21188 6053 21244
rect 5989 21184 6053 21188
rect 6069 21244 6133 21248
rect 6069 21188 6073 21244
rect 6073 21188 6129 21244
rect 6129 21188 6133 21244
rect 6069 21184 6133 21188
rect 6149 21244 6213 21248
rect 6149 21188 6153 21244
rect 6153 21188 6209 21244
rect 6209 21188 6213 21244
rect 6149 21184 6213 21188
rect 6229 21244 6293 21248
rect 6229 21188 6233 21244
rect 6233 21188 6289 21244
rect 6289 21188 6293 21244
rect 6229 21184 6293 21188
rect 9347 21244 9411 21248
rect 9347 21188 9351 21244
rect 9351 21188 9407 21244
rect 9407 21188 9411 21244
rect 9347 21184 9411 21188
rect 9427 21244 9491 21248
rect 9427 21188 9431 21244
rect 9431 21188 9487 21244
rect 9487 21188 9491 21244
rect 9427 21184 9491 21188
rect 9507 21244 9571 21248
rect 9507 21188 9511 21244
rect 9511 21188 9567 21244
rect 9567 21188 9571 21244
rect 9507 21184 9571 21188
rect 9587 21244 9651 21248
rect 9587 21188 9591 21244
rect 9591 21188 9647 21244
rect 9647 21188 9651 21244
rect 9587 21184 9651 21188
rect 12705 21244 12769 21248
rect 12705 21188 12709 21244
rect 12709 21188 12765 21244
rect 12765 21188 12769 21244
rect 12705 21184 12769 21188
rect 12785 21244 12849 21248
rect 12785 21188 12789 21244
rect 12789 21188 12845 21244
rect 12845 21188 12849 21244
rect 12785 21184 12849 21188
rect 12865 21244 12929 21248
rect 12865 21188 12869 21244
rect 12869 21188 12925 21244
rect 12925 21188 12929 21244
rect 12865 21184 12929 21188
rect 12945 21244 13009 21248
rect 12945 21188 12949 21244
rect 12949 21188 13005 21244
rect 13005 21188 13009 21244
rect 12945 21184 13009 21188
rect 9812 20844 9876 20908
rect 7052 20708 7116 20772
rect 13860 20768 13924 20772
rect 13860 20712 13874 20768
rect 13874 20712 13924 20768
rect 13860 20708 13924 20712
rect 4310 20700 4374 20704
rect 4310 20644 4314 20700
rect 4314 20644 4370 20700
rect 4370 20644 4374 20700
rect 4310 20640 4374 20644
rect 4390 20700 4454 20704
rect 4390 20644 4394 20700
rect 4394 20644 4450 20700
rect 4450 20644 4454 20700
rect 4390 20640 4454 20644
rect 4470 20700 4534 20704
rect 4470 20644 4474 20700
rect 4474 20644 4530 20700
rect 4530 20644 4534 20700
rect 4470 20640 4534 20644
rect 4550 20700 4614 20704
rect 4550 20644 4554 20700
rect 4554 20644 4610 20700
rect 4610 20644 4614 20700
rect 4550 20640 4614 20644
rect 7668 20700 7732 20704
rect 7668 20644 7672 20700
rect 7672 20644 7728 20700
rect 7728 20644 7732 20700
rect 7668 20640 7732 20644
rect 7748 20700 7812 20704
rect 7748 20644 7752 20700
rect 7752 20644 7808 20700
rect 7808 20644 7812 20700
rect 7748 20640 7812 20644
rect 7828 20700 7892 20704
rect 7828 20644 7832 20700
rect 7832 20644 7888 20700
rect 7888 20644 7892 20700
rect 7828 20640 7892 20644
rect 7908 20700 7972 20704
rect 7908 20644 7912 20700
rect 7912 20644 7968 20700
rect 7968 20644 7972 20700
rect 7908 20640 7972 20644
rect 11026 20700 11090 20704
rect 11026 20644 11030 20700
rect 11030 20644 11086 20700
rect 11086 20644 11090 20700
rect 11026 20640 11090 20644
rect 11106 20700 11170 20704
rect 11106 20644 11110 20700
rect 11110 20644 11166 20700
rect 11166 20644 11170 20700
rect 11106 20640 11170 20644
rect 11186 20700 11250 20704
rect 11186 20644 11190 20700
rect 11190 20644 11246 20700
rect 11246 20644 11250 20700
rect 11186 20640 11250 20644
rect 11266 20700 11330 20704
rect 11266 20644 11270 20700
rect 11270 20644 11326 20700
rect 11326 20644 11330 20700
rect 11266 20640 11330 20644
rect 14384 20700 14448 20704
rect 14384 20644 14388 20700
rect 14388 20644 14444 20700
rect 14444 20644 14448 20700
rect 14384 20640 14448 20644
rect 14464 20700 14528 20704
rect 14464 20644 14468 20700
rect 14468 20644 14524 20700
rect 14524 20644 14528 20700
rect 14464 20640 14528 20644
rect 14544 20700 14608 20704
rect 14544 20644 14548 20700
rect 14548 20644 14604 20700
rect 14604 20644 14608 20700
rect 14544 20640 14608 20644
rect 14624 20700 14688 20704
rect 14624 20644 14628 20700
rect 14628 20644 14684 20700
rect 14684 20644 14688 20700
rect 14624 20640 14688 20644
rect 12204 20632 12268 20636
rect 12204 20576 12218 20632
rect 12218 20576 12268 20632
rect 12204 20572 12268 20576
rect 1532 20436 1596 20500
rect 2631 20156 2695 20160
rect 2631 20100 2635 20156
rect 2635 20100 2691 20156
rect 2691 20100 2695 20156
rect 2631 20096 2695 20100
rect 2711 20156 2775 20160
rect 2711 20100 2715 20156
rect 2715 20100 2771 20156
rect 2771 20100 2775 20156
rect 2711 20096 2775 20100
rect 2791 20156 2855 20160
rect 2791 20100 2795 20156
rect 2795 20100 2851 20156
rect 2851 20100 2855 20156
rect 2791 20096 2855 20100
rect 2871 20156 2935 20160
rect 2871 20100 2875 20156
rect 2875 20100 2931 20156
rect 2931 20100 2935 20156
rect 2871 20096 2935 20100
rect 5989 20156 6053 20160
rect 5989 20100 5993 20156
rect 5993 20100 6049 20156
rect 6049 20100 6053 20156
rect 5989 20096 6053 20100
rect 6069 20156 6133 20160
rect 6069 20100 6073 20156
rect 6073 20100 6129 20156
rect 6129 20100 6133 20156
rect 6069 20096 6133 20100
rect 6149 20156 6213 20160
rect 6149 20100 6153 20156
rect 6153 20100 6209 20156
rect 6209 20100 6213 20156
rect 6149 20096 6213 20100
rect 6229 20156 6293 20160
rect 6229 20100 6233 20156
rect 6233 20100 6289 20156
rect 6289 20100 6293 20156
rect 6229 20096 6293 20100
rect 9347 20156 9411 20160
rect 9347 20100 9351 20156
rect 9351 20100 9407 20156
rect 9407 20100 9411 20156
rect 9347 20096 9411 20100
rect 9427 20156 9491 20160
rect 9427 20100 9431 20156
rect 9431 20100 9487 20156
rect 9487 20100 9491 20156
rect 9427 20096 9491 20100
rect 9507 20156 9571 20160
rect 9507 20100 9511 20156
rect 9511 20100 9567 20156
rect 9567 20100 9571 20156
rect 9507 20096 9571 20100
rect 9587 20156 9651 20160
rect 9587 20100 9591 20156
rect 9591 20100 9647 20156
rect 9647 20100 9651 20156
rect 9587 20096 9651 20100
rect 12705 20156 12769 20160
rect 12705 20100 12709 20156
rect 12709 20100 12765 20156
rect 12765 20100 12769 20156
rect 12705 20096 12769 20100
rect 12785 20156 12849 20160
rect 12785 20100 12789 20156
rect 12789 20100 12845 20156
rect 12845 20100 12849 20156
rect 12785 20096 12849 20100
rect 12865 20156 12929 20160
rect 12865 20100 12869 20156
rect 12869 20100 12925 20156
rect 12925 20100 12929 20156
rect 12865 20096 12929 20100
rect 12945 20156 13009 20160
rect 12945 20100 12949 20156
rect 12949 20100 13005 20156
rect 13005 20100 13009 20156
rect 12945 20096 13009 20100
rect 4310 19612 4374 19616
rect 4310 19556 4314 19612
rect 4314 19556 4370 19612
rect 4370 19556 4374 19612
rect 4310 19552 4374 19556
rect 4390 19612 4454 19616
rect 4390 19556 4394 19612
rect 4394 19556 4450 19612
rect 4450 19556 4454 19612
rect 4390 19552 4454 19556
rect 4470 19612 4534 19616
rect 4470 19556 4474 19612
rect 4474 19556 4530 19612
rect 4530 19556 4534 19612
rect 4470 19552 4534 19556
rect 4550 19612 4614 19616
rect 4550 19556 4554 19612
rect 4554 19556 4610 19612
rect 4610 19556 4614 19612
rect 4550 19552 4614 19556
rect 7668 19612 7732 19616
rect 7668 19556 7672 19612
rect 7672 19556 7728 19612
rect 7728 19556 7732 19612
rect 7668 19552 7732 19556
rect 7748 19612 7812 19616
rect 7748 19556 7752 19612
rect 7752 19556 7808 19612
rect 7808 19556 7812 19612
rect 7748 19552 7812 19556
rect 7828 19612 7892 19616
rect 7828 19556 7832 19612
rect 7832 19556 7888 19612
rect 7888 19556 7892 19612
rect 7828 19552 7892 19556
rect 7908 19612 7972 19616
rect 7908 19556 7912 19612
rect 7912 19556 7968 19612
rect 7968 19556 7972 19612
rect 7908 19552 7972 19556
rect 11026 19612 11090 19616
rect 11026 19556 11030 19612
rect 11030 19556 11086 19612
rect 11086 19556 11090 19612
rect 11026 19552 11090 19556
rect 11106 19612 11170 19616
rect 11106 19556 11110 19612
rect 11110 19556 11166 19612
rect 11166 19556 11170 19612
rect 11106 19552 11170 19556
rect 11186 19612 11250 19616
rect 11186 19556 11190 19612
rect 11190 19556 11246 19612
rect 11246 19556 11250 19612
rect 11186 19552 11250 19556
rect 11266 19612 11330 19616
rect 11266 19556 11270 19612
rect 11270 19556 11326 19612
rect 11326 19556 11330 19612
rect 11266 19552 11330 19556
rect 14384 19612 14448 19616
rect 14384 19556 14388 19612
rect 14388 19556 14444 19612
rect 14444 19556 14448 19612
rect 14384 19552 14448 19556
rect 14464 19612 14528 19616
rect 14464 19556 14468 19612
rect 14468 19556 14524 19612
rect 14524 19556 14528 19612
rect 14464 19552 14528 19556
rect 14544 19612 14608 19616
rect 14544 19556 14548 19612
rect 14548 19556 14604 19612
rect 14604 19556 14608 19612
rect 14544 19552 14608 19556
rect 14624 19612 14688 19616
rect 14624 19556 14628 19612
rect 14628 19556 14684 19612
rect 14684 19556 14688 19612
rect 14624 19552 14688 19556
rect 9076 19348 9140 19412
rect 9996 19348 10060 19412
rect 8892 19212 8956 19276
rect 13676 19212 13740 19276
rect 2631 19068 2695 19072
rect 2631 19012 2635 19068
rect 2635 19012 2691 19068
rect 2691 19012 2695 19068
rect 2631 19008 2695 19012
rect 2711 19068 2775 19072
rect 2711 19012 2715 19068
rect 2715 19012 2771 19068
rect 2771 19012 2775 19068
rect 2711 19008 2775 19012
rect 2791 19068 2855 19072
rect 2791 19012 2795 19068
rect 2795 19012 2851 19068
rect 2851 19012 2855 19068
rect 2791 19008 2855 19012
rect 2871 19068 2935 19072
rect 2871 19012 2875 19068
rect 2875 19012 2931 19068
rect 2931 19012 2935 19068
rect 2871 19008 2935 19012
rect 5989 19068 6053 19072
rect 5989 19012 5993 19068
rect 5993 19012 6049 19068
rect 6049 19012 6053 19068
rect 5989 19008 6053 19012
rect 6069 19068 6133 19072
rect 6069 19012 6073 19068
rect 6073 19012 6129 19068
rect 6129 19012 6133 19068
rect 6069 19008 6133 19012
rect 6149 19068 6213 19072
rect 6149 19012 6153 19068
rect 6153 19012 6209 19068
rect 6209 19012 6213 19068
rect 6149 19008 6213 19012
rect 6229 19068 6293 19072
rect 6229 19012 6233 19068
rect 6233 19012 6289 19068
rect 6289 19012 6293 19068
rect 6229 19008 6293 19012
rect 9347 19068 9411 19072
rect 9347 19012 9351 19068
rect 9351 19012 9407 19068
rect 9407 19012 9411 19068
rect 9347 19008 9411 19012
rect 9427 19068 9491 19072
rect 9427 19012 9431 19068
rect 9431 19012 9487 19068
rect 9487 19012 9491 19068
rect 9427 19008 9491 19012
rect 9507 19068 9571 19072
rect 9507 19012 9511 19068
rect 9511 19012 9567 19068
rect 9567 19012 9571 19068
rect 9507 19008 9571 19012
rect 9587 19068 9651 19072
rect 9587 19012 9591 19068
rect 9591 19012 9647 19068
rect 9647 19012 9651 19068
rect 9587 19008 9651 19012
rect 12705 19068 12769 19072
rect 12705 19012 12709 19068
rect 12709 19012 12765 19068
rect 12765 19012 12769 19068
rect 12705 19008 12769 19012
rect 12785 19068 12849 19072
rect 12785 19012 12789 19068
rect 12789 19012 12845 19068
rect 12845 19012 12849 19068
rect 12785 19008 12849 19012
rect 12865 19068 12929 19072
rect 12865 19012 12869 19068
rect 12869 19012 12925 19068
rect 12925 19012 12929 19068
rect 12865 19008 12929 19012
rect 12945 19068 13009 19072
rect 12945 19012 12949 19068
rect 12949 19012 13005 19068
rect 13005 19012 13009 19068
rect 12945 19008 13009 19012
rect 7420 18804 7484 18868
rect 7236 18668 7300 18732
rect 8156 18728 8220 18732
rect 8156 18672 8206 18728
rect 8206 18672 8220 18728
rect 8156 18668 8220 18672
rect 4310 18524 4374 18528
rect 4310 18468 4314 18524
rect 4314 18468 4370 18524
rect 4370 18468 4374 18524
rect 4310 18464 4374 18468
rect 4390 18524 4454 18528
rect 4390 18468 4394 18524
rect 4394 18468 4450 18524
rect 4450 18468 4454 18524
rect 4390 18464 4454 18468
rect 4470 18524 4534 18528
rect 4470 18468 4474 18524
rect 4474 18468 4530 18524
rect 4530 18468 4534 18524
rect 4470 18464 4534 18468
rect 4550 18524 4614 18528
rect 4550 18468 4554 18524
rect 4554 18468 4610 18524
rect 4610 18468 4614 18524
rect 4550 18464 4614 18468
rect 7668 18524 7732 18528
rect 7668 18468 7672 18524
rect 7672 18468 7728 18524
rect 7728 18468 7732 18524
rect 7668 18464 7732 18468
rect 7748 18524 7812 18528
rect 7748 18468 7752 18524
rect 7752 18468 7808 18524
rect 7808 18468 7812 18524
rect 7748 18464 7812 18468
rect 7828 18524 7892 18528
rect 7828 18468 7832 18524
rect 7832 18468 7888 18524
rect 7888 18468 7892 18524
rect 7828 18464 7892 18468
rect 7908 18524 7972 18528
rect 7908 18468 7912 18524
rect 7912 18468 7968 18524
rect 7968 18468 7972 18524
rect 7908 18464 7972 18468
rect 11026 18524 11090 18528
rect 11026 18468 11030 18524
rect 11030 18468 11086 18524
rect 11086 18468 11090 18524
rect 11026 18464 11090 18468
rect 11106 18524 11170 18528
rect 11106 18468 11110 18524
rect 11110 18468 11166 18524
rect 11166 18468 11170 18524
rect 11106 18464 11170 18468
rect 11186 18524 11250 18528
rect 11186 18468 11190 18524
rect 11190 18468 11246 18524
rect 11246 18468 11250 18524
rect 11186 18464 11250 18468
rect 11266 18524 11330 18528
rect 11266 18468 11270 18524
rect 11270 18468 11326 18524
rect 11326 18468 11330 18524
rect 11266 18464 11330 18468
rect 14384 18524 14448 18528
rect 14384 18468 14388 18524
rect 14388 18468 14444 18524
rect 14444 18468 14448 18524
rect 14384 18464 14448 18468
rect 14464 18524 14528 18528
rect 14464 18468 14468 18524
rect 14468 18468 14524 18524
rect 14524 18468 14528 18524
rect 14464 18464 14528 18468
rect 14544 18524 14608 18528
rect 14544 18468 14548 18524
rect 14548 18468 14604 18524
rect 14604 18468 14608 18524
rect 14544 18464 14608 18468
rect 14624 18524 14688 18528
rect 14624 18468 14628 18524
rect 14628 18468 14684 18524
rect 14684 18468 14688 18524
rect 14624 18464 14688 18468
rect 13308 18396 13372 18460
rect 9076 18260 9140 18324
rect 11468 18260 11532 18324
rect 12388 18320 12452 18324
rect 12388 18264 12402 18320
rect 12402 18264 12452 18320
rect 12388 18260 12452 18264
rect 13492 18320 13556 18324
rect 13492 18264 13506 18320
rect 13506 18264 13556 18320
rect 13492 18260 13556 18264
rect 2631 17980 2695 17984
rect 2631 17924 2635 17980
rect 2635 17924 2691 17980
rect 2691 17924 2695 17980
rect 2631 17920 2695 17924
rect 2711 17980 2775 17984
rect 2711 17924 2715 17980
rect 2715 17924 2771 17980
rect 2771 17924 2775 17980
rect 2711 17920 2775 17924
rect 2791 17980 2855 17984
rect 2791 17924 2795 17980
rect 2795 17924 2851 17980
rect 2851 17924 2855 17980
rect 2791 17920 2855 17924
rect 2871 17980 2935 17984
rect 2871 17924 2875 17980
rect 2875 17924 2931 17980
rect 2931 17924 2935 17980
rect 2871 17920 2935 17924
rect 5989 17980 6053 17984
rect 5989 17924 5993 17980
rect 5993 17924 6049 17980
rect 6049 17924 6053 17980
rect 5989 17920 6053 17924
rect 6069 17980 6133 17984
rect 6069 17924 6073 17980
rect 6073 17924 6129 17980
rect 6129 17924 6133 17980
rect 6069 17920 6133 17924
rect 6149 17980 6213 17984
rect 6149 17924 6153 17980
rect 6153 17924 6209 17980
rect 6209 17924 6213 17980
rect 6149 17920 6213 17924
rect 6229 17980 6293 17984
rect 6229 17924 6233 17980
rect 6233 17924 6289 17980
rect 6289 17924 6293 17980
rect 6229 17920 6293 17924
rect 9347 17980 9411 17984
rect 9347 17924 9351 17980
rect 9351 17924 9407 17980
rect 9407 17924 9411 17980
rect 9347 17920 9411 17924
rect 9427 17980 9491 17984
rect 9427 17924 9431 17980
rect 9431 17924 9487 17980
rect 9487 17924 9491 17980
rect 9427 17920 9491 17924
rect 9507 17980 9571 17984
rect 9507 17924 9511 17980
rect 9511 17924 9567 17980
rect 9567 17924 9571 17980
rect 9507 17920 9571 17924
rect 9587 17980 9651 17984
rect 9587 17924 9591 17980
rect 9591 17924 9647 17980
rect 9647 17924 9651 17980
rect 9587 17920 9651 17924
rect 12705 17980 12769 17984
rect 12705 17924 12709 17980
rect 12709 17924 12765 17980
rect 12765 17924 12769 17980
rect 12705 17920 12769 17924
rect 12785 17980 12849 17984
rect 12785 17924 12789 17980
rect 12789 17924 12845 17980
rect 12845 17924 12849 17980
rect 12785 17920 12849 17924
rect 12865 17980 12929 17984
rect 12865 17924 12869 17980
rect 12869 17924 12925 17980
rect 12925 17924 12929 17980
rect 12865 17920 12929 17924
rect 12945 17980 13009 17984
rect 12945 17924 12949 17980
rect 12949 17924 13005 17980
rect 13005 17924 13009 17980
rect 12945 17920 13009 17924
rect 9812 17912 9876 17916
rect 9812 17856 9826 17912
rect 9826 17856 9876 17912
rect 9812 17852 9876 17856
rect 7052 17580 7116 17644
rect 4310 17436 4374 17440
rect 4310 17380 4314 17436
rect 4314 17380 4370 17436
rect 4370 17380 4374 17436
rect 4310 17376 4374 17380
rect 4390 17436 4454 17440
rect 4390 17380 4394 17436
rect 4394 17380 4450 17436
rect 4450 17380 4454 17436
rect 4390 17376 4454 17380
rect 4470 17436 4534 17440
rect 4470 17380 4474 17436
rect 4474 17380 4530 17436
rect 4530 17380 4534 17436
rect 4470 17376 4534 17380
rect 4550 17436 4614 17440
rect 4550 17380 4554 17436
rect 4554 17380 4610 17436
rect 4610 17380 4614 17436
rect 4550 17376 4614 17380
rect 7668 17436 7732 17440
rect 7668 17380 7672 17436
rect 7672 17380 7728 17436
rect 7728 17380 7732 17436
rect 7668 17376 7732 17380
rect 7748 17436 7812 17440
rect 7748 17380 7752 17436
rect 7752 17380 7808 17436
rect 7808 17380 7812 17436
rect 7748 17376 7812 17380
rect 7828 17436 7892 17440
rect 7828 17380 7832 17436
rect 7832 17380 7888 17436
rect 7888 17380 7892 17436
rect 7828 17376 7892 17380
rect 7908 17436 7972 17440
rect 7908 17380 7912 17436
rect 7912 17380 7968 17436
rect 7968 17380 7972 17436
rect 7908 17376 7972 17380
rect 14044 17580 14108 17644
rect 11026 17436 11090 17440
rect 11026 17380 11030 17436
rect 11030 17380 11086 17436
rect 11086 17380 11090 17436
rect 11026 17376 11090 17380
rect 11106 17436 11170 17440
rect 11106 17380 11110 17436
rect 11110 17380 11166 17436
rect 11166 17380 11170 17436
rect 11106 17376 11170 17380
rect 11186 17436 11250 17440
rect 11186 17380 11190 17436
rect 11190 17380 11246 17436
rect 11246 17380 11250 17436
rect 11186 17376 11250 17380
rect 11266 17436 11330 17440
rect 11266 17380 11270 17436
rect 11270 17380 11326 17436
rect 11326 17380 11330 17436
rect 11266 17376 11330 17380
rect 14384 17436 14448 17440
rect 14384 17380 14388 17436
rect 14388 17380 14444 17436
rect 14444 17380 14448 17436
rect 14384 17376 14448 17380
rect 14464 17436 14528 17440
rect 14464 17380 14468 17436
rect 14468 17380 14524 17436
rect 14524 17380 14528 17436
rect 14464 17376 14528 17380
rect 14544 17436 14608 17440
rect 14544 17380 14548 17436
rect 14548 17380 14604 17436
rect 14604 17380 14608 17436
rect 14544 17376 14608 17380
rect 14624 17436 14688 17440
rect 14624 17380 14628 17436
rect 14628 17380 14684 17436
rect 14684 17380 14688 17436
rect 14624 17376 14688 17380
rect 14228 17308 14292 17372
rect 10364 17036 10428 17100
rect 2631 16892 2695 16896
rect 2631 16836 2635 16892
rect 2635 16836 2691 16892
rect 2691 16836 2695 16892
rect 2631 16832 2695 16836
rect 2711 16892 2775 16896
rect 2711 16836 2715 16892
rect 2715 16836 2771 16892
rect 2771 16836 2775 16892
rect 2711 16832 2775 16836
rect 2791 16892 2855 16896
rect 2791 16836 2795 16892
rect 2795 16836 2851 16892
rect 2851 16836 2855 16892
rect 2791 16832 2855 16836
rect 2871 16892 2935 16896
rect 2871 16836 2875 16892
rect 2875 16836 2931 16892
rect 2931 16836 2935 16892
rect 2871 16832 2935 16836
rect 5989 16892 6053 16896
rect 5989 16836 5993 16892
rect 5993 16836 6049 16892
rect 6049 16836 6053 16892
rect 5989 16832 6053 16836
rect 6069 16892 6133 16896
rect 6069 16836 6073 16892
rect 6073 16836 6129 16892
rect 6129 16836 6133 16892
rect 6069 16832 6133 16836
rect 6149 16892 6213 16896
rect 6149 16836 6153 16892
rect 6153 16836 6209 16892
rect 6209 16836 6213 16892
rect 6149 16832 6213 16836
rect 6229 16892 6293 16896
rect 6229 16836 6233 16892
rect 6233 16836 6289 16892
rect 6289 16836 6293 16892
rect 6229 16832 6293 16836
rect 9347 16892 9411 16896
rect 9347 16836 9351 16892
rect 9351 16836 9407 16892
rect 9407 16836 9411 16892
rect 9347 16832 9411 16836
rect 9427 16892 9491 16896
rect 9427 16836 9431 16892
rect 9431 16836 9487 16892
rect 9487 16836 9491 16892
rect 9427 16832 9491 16836
rect 9507 16892 9571 16896
rect 9507 16836 9511 16892
rect 9511 16836 9567 16892
rect 9567 16836 9571 16892
rect 9507 16832 9571 16836
rect 9587 16892 9651 16896
rect 9587 16836 9591 16892
rect 9591 16836 9647 16892
rect 9647 16836 9651 16892
rect 9587 16832 9651 16836
rect 12705 16892 12769 16896
rect 12705 16836 12709 16892
rect 12709 16836 12765 16892
rect 12765 16836 12769 16892
rect 12705 16832 12769 16836
rect 12785 16892 12849 16896
rect 12785 16836 12789 16892
rect 12789 16836 12845 16892
rect 12845 16836 12849 16892
rect 12785 16832 12849 16836
rect 12865 16892 12929 16896
rect 12865 16836 12869 16892
rect 12869 16836 12925 16892
rect 12925 16836 12929 16892
rect 12865 16832 12929 16836
rect 12945 16892 13009 16896
rect 12945 16836 12949 16892
rect 12949 16836 13005 16892
rect 13005 16836 13009 16892
rect 12945 16832 13009 16836
rect 10732 16492 10796 16556
rect 13492 16492 13556 16556
rect 4310 16348 4374 16352
rect 4310 16292 4314 16348
rect 4314 16292 4370 16348
rect 4370 16292 4374 16348
rect 4310 16288 4374 16292
rect 4390 16348 4454 16352
rect 4390 16292 4394 16348
rect 4394 16292 4450 16348
rect 4450 16292 4454 16348
rect 4390 16288 4454 16292
rect 4470 16348 4534 16352
rect 4470 16292 4474 16348
rect 4474 16292 4530 16348
rect 4530 16292 4534 16348
rect 4470 16288 4534 16292
rect 4550 16348 4614 16352
rect 4550 16292 4554 16348
rect 4554 16292 4610 16348
rect 4610 16292 4614 16348
rect 4550 16288 4614 16292
rect 7668 16348 7732 16352
rect 7668 16292 7672 16348
rect 7672 16292 7728 16348
rect 7728 16292 7732 16348
rect 7668 16288 7732 16292
rect 7748 16348 7812 16352
rect 7748 16292 7752 16348
rect 7752 16292 7808 16348
rect 7808 16292 7812 16348
rect 7748 16288 7812 16292
rect 7828 16348 7892 16352
rect 7828 16292 7832 16348
rect 7832 16292 7888 16348
rect 7888 16292 7892 16348
rect 7828 16288 7892 16292
rect 7908 16348 7972 16352
rect 7908 16292 7912 16348
rect 7912 16292 7968 16348
rect 7968 16292 7972 16348
rect 7908 16288 7972 16292
rect 11026 16348 11090 16352
rect 11026 16292 11030 16348
rect 11030 16292 11086 16348
rect 11086 16292 11090 16348
rect 11026 16288 11090 16292
rect 11106 16348 11170 16352
rect 11106 16292 11110 16348
rect 11110 16292 11166 16348
rect 11166 16292 11170 16348
rect 11106 16288 11170 16292
rect 11186 16348 11250 16352
rect 11186 16292 11190 16348
rect 11190 16292 11246 16348
rect 11246 16292 11250 16348
rect 11186 16288 11250 16292
rect 11266 16348 11330 16352
rect 11266 16292 11270 16348
rect 11270 16292 11326 16348
rect 11326 16292 11330 16348
rect 11266 16288 11330 16292
rect 14384 16348 14448 16352
rect 14384 16292 14388 16348
rect 14388 16292 14444 16348
rect 14444 16292 14448 16348
rect 14384 16288 14448 16292
rect 14464 16348 14528 16352
rect 14464 16292 14468 16348
rect 14468 16292 14524 16348
rect 14524 16292 14528 16348
rect 14464 16288 14528 16292
rect 14544 16348 14608 16352
rect 14544 16292 14548 16348
rect 14548 16292 14604 16348
rect 14604 16292 14608 16348
rect 14544 16288 14608 16292
rect 14624 16348 14688 16352
rect 14624 16292 14628 16348
rect 14628 16292 14684 16348
rect 14684 16292 14688 16348
rect 14624 16288 14688 16292
rect 15332 16008 15396 16012
rect 15332 15952 15346 16008
rect 15346 15952 15396 16008
rect 15332 15948 15396 15952
rect 7236 15812 7300 15876
rect 2631 15804 2695 15808
rect 2631 15748 2635 15804
rect 2635 15748 2691 15804
rect 2691 15748 2695 15804
rect 2631 15744 2695 15748
rect 2711 15804 2775 15808
rect 2711 15748 2715 15804
rect 2715 15748 2771 15804
rect 2771 15748 2775 15804
rect 2711 15744 2775 15748
rect 2791 15804 2855 15808
rect 2791 15748 2795 15804
rect 2795 15748 2851 15804
rect 2851 15748 2855 15804
rect 2791 15744 2855 15748
rect 2871 15804 2935 15808
rect 2871 15748 2875 15804
rect 2875 15748 2931 15804
rect 2931 15748 2935 15804
rect 2871 15744 2935 15748
rect 5989 15804 6053 15808
rect 5989 15748 5993 15804
rect 5993 15748 6049 15804
rect 6049 15748 6053 15804
rect 5989 15744 6053 15748
rect 6069 15804 6133 15808
rect 6069 15748 6073 15804
rect 6073 15748 6129 15804
rect 6129 15748 6133 15804
rect 6069 15744 6133 15748
rect 6149 15804 6213 15808
rect 6149 15748 6153 15804
rect 6153 15748 6209 15804
rect 6209 15748 6213 15804
rect 6149 15744 6213 15748
rect 6229 15804 6293 15808
rect 6229 15748 6233 15804
rect 6233 15748 6289 15804
rect 6289 15748 6293 15804
rect 6229 15744 6293 15748
rect 9347 15804 9411 15808
rect 9347 15748 9351 15804
rect 9351 15748 9407 15804
rect 9407 15748 9411 15804
rect 9347 15744 9411 15748
rect 9427 15804 9491 15808
rect 9427 15748 9431 15804
rect 9431 15748 9487 15804
rect 9487 15748 9491 15804
rect 9427 15744 9491 15748
rect 9507 15804 9571 15808
rect 9507 15748 9511 15804
rect 9511 15748 9567 15804
rect 9567 15748 9571 15804
rect 9507 15744 9571 15748
rect 9587 15804 9651 15808
rect 9587 15748 9591 15804
rect 9591 15748 9647 15804
rect 9647 15748 9651 15804
rect 9587 15744 9651 15748
rect 12705 15804 12769 15808
rect 12705 15748 12709 15804
rect 12709 15748 12765 15804
rect 12765 15748 12769 15804
rect 12705 15744 12769 15748
rect 12785 15804 12849 15808
rect 12785 15748 12789 15804
rect 12789 15748 12845 15804
rect 12845 15748 12849 15804
rect 12785 15744 12849 15748
rect 12865 15804 12929 15808
rect 12865 15748 12869 15804
rect 12869 15748 12925 15804
rect 12925 15748 12929 15804
rect 12865 15744 12929 15748
rect 12945 15804 13009 15808
rect 12945 15748 12949 15804
rect 12949 15748 13005 15804
rect 13005 15748 13009 15804
rect 12945 15744 13009 15748
rect 10732 15540 10796 15604
rect 11468 15540 11532 15604
rect 9996 15404 10060 15468
rect 4310 15260 4374 15264
rect 4310 15204 4314 15260
rect 4314 15204 4370 15260
rect 4370 15204 4374 15260
rect 4310 15200 4374 15204
rect 4390 15260 4454 15264
rect 4390 15204 4394 15260
rect 4394 15204 4450 15260
rect 4450 15204 4454 15260
rect 4390 15200 4454 15204
rect 4470 15260 4534 15264
rect 4470 15204 4474 15260
rect 4474 15204 4530 15260
rect 4530 15204 4534 15260
rect 4470 15200 4534 15204
rect 4550 15260 4614 15264
rect 4550 15204 4554 15260
rect 4554 15204 4610 15260
rect 4610 15204 4614 15260
rect 4550 15200 4614 15204
rect 7668 15260 7732 15264
rect 7668 15204 7672 15260
rect 7672 15204 7728 15260
rect 7728 15204 7732 15260
rect 7668 15200 7732 15204
rect 7748 15260 7812 15264
rect 7748 15204 7752 15260
rect 7752 15204 7808 15260
rect 7808 15204 7812 15260
rect 7748 15200 7812 15204
rect 7828 15260 7892 15264
rect 7828 15204 7832 15260
rect 7832 15204 7888 15260
rect 7888 15204 7892 15260
rect 7828 15200 7892 15204
rect 7908 15260 7972 15264
rect 7908 15204 7912 15260
rect 7912 15204 7968 15260
rect 7968 15204 7972 15260
rect 7908 15200 7972 15204
rect 11026 15260 11090 15264
rect 11026 15204 11030 15260
rect 11030 15204 11086 15260
rect 11086 15204 11090 15260
rect 11026 15200 11090 15204
rect 11106 15260 11170 15264
rect 11106 15204 11110 15260
rect 11110 15204 11166 15260
rect 11166 15204 11170 15260
rect 11106 15200 11170 15204
rect 11186 15260 11250 15264
rect 11186 15204 11190 15260
rect 11190 15204 11246 15260
rect 11246 15204 11250 15260
rect 11186 15200 11250 15204
rect 11266 15260 11330 15264
rect 11266 15204 11270 15260
rect 11270 15204 11326 15260
rect 11326 15204 11330 15260
rect 11266 15200 11330 15204
rect 14384 15260 14448 15264
rect 14384 15204 14388 15260
rect 14388 15204 14444 15260
rect 14444 15204 14448 15260
rect 14384 15200 14448 15204
rect 14464 15260 14528 15264
rect 14464 15204 14468 15260
rect 14468 15204 14524 15260
rect 14524 15204 14528 15260
rect 14464 15200 14528 15204
rect 14544 15260 14608 15264
rect 14544 15204 14548 15260
rect 14548 15204 14604 15260
rect 14604 15204 14608 15260
rect 14544 15200 14608 15204
rect 14624 15260 14688 15264
rect 14624 15204 14628 15260
rect 14628 15204 14684 15260
rect 14684 15204 14688 15260
rect 14624 15200 14688 15204
rect 13124 14996 13188 15060
rect 15148 14860 15212 14924
rect 2631 14716 2695 14720
rect 2631 14660 2635 14716
rect 2635 14660 2691 14716
rect 2691 14660 2695 14716
rect 2631 14656 2695 14660
rect 2711 14716 2775 14720
rect 2711 14660 2715 14716
rect 2715 14660 2771 14716
rect 2771 14660 2775 14716
rect 2711 14656 2775 14660
rect 2791 14716 2855 14720
rect 2791 14660 2795 14716
rect 2795 14660 2851 14716
rect 2851 14660 2855 14716
rect 2791 14656 2855 14660
rect 2871 14716 2935 14720
rect 2871 14660 2875 14716
rect 2875 14660 2931 14716
rect 2931 14660 2935 14716
rect 2871 14656 2935 14660
rect 5989 14716 6053 14720
rect 5989 14660 5993 14716
rect 5993 14660 6049 14716
rect 6049 14660 6053 14716
rect 5989 14656 6053 14660
rect 6069 14716 6133 14720
rect 6069 14660 6073 14716
rect 6073 14660 6129 14716
rect 6129 14660 6133 14716
rect 6069 14656 6133 14660
rect 6149 14716 6213 14720
rect 6149 14660 6153 14716
rect 6153 14660 6209 14716
rect 6209 14660 6213 14716
rect 6149 14656 6213 14660
rect 6229 14716 6293 14720
rect 6229 14660 6233 14716
rect 6233 14660 6289 14716
rect 6289 14660 6293 14716
rect 6229 14656 6293 14660
rect 9347 14716 9411 14720
rect 9347 14660 9351 14716
rect 9351 14660 9407 14716
rect 9407 14660 9411 14716
rect 9347 14656 9411 14660
rect 9427 14716 9491 14720
rect 9427 14660 9431 14716
rect 9431 14660 9487 14716
rect 9487 14660 9491 14716
rect 9427 14656 9491 14660
rect 9507 14716 9571 14720
rect 9507 14660 9511 14716
rect 9511 14660 9567 14716
rect 9567 14660 9571 14716
rect 9507 14656 9571 14660
rect 9587 14716 9651 14720
rect 9587 14660 9591 14716
rect 9591 14660 9647 14716
rect 9647 14660 9651 14716
rect 9587 14656 9651 14660
rect 12705 14716 12769 14720
rect 12705 14660 12709 14716
rect 12709 14660 12765 14716
rect 12765 14660 12769 14716
rect 12705 14656 12769 14660
rect 12785 14716 12849 14720
rect 12785 14660 12789 14716
rect 12789 14660 12845 14716
rect 12845 14660 12849 14716
rect 12785 14656 12849 14660
rect 12865 14716 12929 14720
rect 12865 14660 12869 14716
rect 12869 14660 12925 14716
rect 12925 14660 12929 14716
rect 12865 14656 12929 14660
rect 12945 14716 13009 14720
rect 12945 14660 12949 14716
rect 12949 14660 13005 14716
rect 13005 14660 13009 14716
rect 12945 14656 13009 14660
rect 10180 14588 10244 14652
rect 14228 14588 14292 14652
rect 13308 14452 13372 14516
rect 13860 14316 13924 14380
rect 4310 14172 4374 14176
rect 4310 14116 4314 14172
rect 4314 14116 4370 14172
rect 4370 14116 4374 14172
rect 4310 14112 4374 14116
rect 4390 14172 4454 14176
rect 4390 14116 4394 14172
rect 4394 14116 4450 14172
rect 4450 14116 4454 14172
rect 4390 14112 4454 14116
rect 4470 14172 4534 14176
rect 4470 14116 4474 14172
rect 4474 14116 4530 14172
rect 4530 14116 4534 14172
rect 4470 14112 4534 14116
rect 4550 14172 4614 14176
rect 4550 14116 4554 14172
rect 4554 14116 4610 14172
rect 4610 14116 4614 14172
rect 4550 14112 4614 14116
rect 7668 14172 7732 14176
rect 7668 14116 7672 14172
rect 7672 14116 7728 14172
rect 7728 14116 7732 14172
rect 7668 14112 7732 14116
rect 7748 14172 7812 14176
rect 7748 14116 7752 14172
rect 7752 14116 7808 14172
rect 7808 14116 7812 14172
rect 7748 14112 7812 14116
rect 7828 14172 7892 14176
rect 7828 14116 7832 14172
rect 7832 14116 7888 14172
rect 7888 14116 7892 14172
rect 7828 14112 7892 14116
rect 7908 14172 7972 14176
rect 7908 14116 7912 14172
rect 7912 14116 7968 14172
rect 7968 14116 7972 14172
rect 7908 14112 7972 14116
rect 11026 14172 11090 14176
rect 11026 14116 11030 14172
rect 11030 14116 11086 14172
rect 11086 14116 11090 14172
rect 11026 14112 11090 14116
rect 11106 14172 11170 14176
rect 11106 14116 11110 14172
rect 11110 14116 11166 14172
rect 11166 14116 11170 14172
rect 11106 14112 11170 14116
rect 11186 14172 11250 14176
rect 11186 14116 11190 14172
rect 11190 14116 11246 14172
rect 11246 14116 11250 14172
rect 11186 14112 11250 14116
rect 11266 14172 11330 14176
rect 11266 14116 11270 14172
rect 11270 14116 11326 14172
rect 11326 14116 11330 14172
rect 11266 14112 11330 14116
rect 14384 14172 14448 14176
rect 14384 14116 14388 14172
rect 14388 14116 14444 14172
rect 14444 14116 14448 14172
rect 14384 14112 14448 14116
rect 14464 14172 14528 14176
rect 14464 14116 14468 14172
rect 14468 14116 14524 14172
rect 14524 14116 14528 14172
rect 14464 14112 14528 14116
rect 14544 14172 14608 14176
rect 14544 14116 14548 14172
rect 14548 14116 14604 14172
rect 14604 14116 14608 14172
rect 14544 14112 14608 14116
rect 14624 14172 14688 14176
rect 14624 14116 14628 14172
rect 14628 14116 14684 14172
rect 14684 14116 14688 14172
rect 14624 14112 14688 14116
rect 12204 13908 12268 13972
rect 7420 13636 7484 13700
rect 2631 13628 2695 13632
rect 2631 13572 2635 13628
rect 2635 13572 2691 13628
rect 2691 13572 2695 13628
rect 2631 13568 2695 13572
rect 2711 13628 2775 13632
rect 2711 13572 2715 13628
rect 2715 13572 2771 13628
rect 2771 13572 2775 13628
rect 2711 13568 2775 13572
rect 2791 13628 2855 13632
rect 2791 13572 2795 13628
rect 2795 13572 2851 13628
rect 2851 13572 2855 13628
rect 2791 13568 2855 13572
rect 2871 13628 2935 13632
rect 2871 13572 2875 13628
rect 2875 13572 2931 13628
rect 2931 13572 2935 13628
rect 2871 13568 2935 13572
rect 5989 13628 6053 13632
rect 5989 13572 5993 13628
rect 5993 13572 6049 13628
rect 6049 13572 6053 13628
rect 5989 13568 6053 13572
rect 6069 13628 6133 13632
rect 6069 13572 6073 13628
rect 6073 13572 6129 13628
rect 6129 13572 6133 13628
rect 6069 13568 6133 13572
rect 6149 13628 6213 13632
rect 6149 13572 6153 13628
rect 6153 13572 6209 13628
rect 6209 13572 6213 13628
rect 6149 13568 6213 13572
rect 6229 13628 6293 13632
rect 6229 13572 6233 13628
rect 6233 13572 6289 13628
rect 6289 13572 6293 13628
rect 6229 13568 6293 13572
rect 9347 13628 9411 13632
rect 9347 13572 9351 13628
rect 9351 13572 9407 13628
rect 9407 13572 9411 13628
rect 9347 13568 9411 13572
rect 9427 13628 9491 13632
rect 9427 13572 9431 13628
rect 9431 13572 9487 13628
rect 9487 13572 9491 13628
rect 9427 13568 9491 13572
rect 9507 13628 9571 13632
rect 9507 13572 9511 13628
rect 9511 13572 9567 13628
rect 9567 13572 9571 13628
rect 9507 13568 9571 13572
rect 9587 13628 9651 13632
rect 9587 13572 9591 13628
rect 9591 13572 9647 13628
rect 9647 13572 9651 13628
rect 9587 13568 9651 13572
rect 12705 13628 12769 13632
rect 12705 13572 12709 13628
rect 12709 13572 12765 13628
rect 12765 13572 12769 13628
rect 12705 13568 12769 13572
rect 12785 13628 12849 13632
rect 12785 13572 12789 13628
rect 12789 13572 12845 13628
rect 12845 13572 12849 13628
rect 12785 13568 12849 13572
rect 12865 13628 12929 13632
rect 12865 13572 12869 13628
rect 12869 13572 12925 13628
rect 12925 13572 12929 13628
rect 12865 13568 12929 13572
rect 12945 13628 13009 13632
rect 12945 13572 12949 13628
rect 12949 13572 13005 13628
rect 13005 13572 13009 13628
rect 12945 13568 13009 13572
rect 8892 13364 8956 13428
rect 11468 13228 11532 13292
rect 4310 13084 4374 13088
rect 4310 13028 4314 13084
rect 4314 13028 4370 13084
rect 4370 13028 4374 13084
rect 4310 13024 4374 13028
rect 4390 13084 4454 13088
rect 4390 13028 4394 13084
rect 4394 13028 4450 13084
rect 4450 13028 4454 13084
rect 4390 13024 4454 13028
rect 4470 13084 4534 13088
rect 4470 13028 4474 13084
rect 4474 13028 4530 13084
rect 4530 13028 4534 13084
rect 4470 13024 4534 13028
rect 4550 13084 4614 13088
rect 4550 13028 4554 13084
rect 4554 13028 4610 13084
rect 4610 13028 4614 13084
rect 4550 13024 4614 13028
rect 7668 13084 7732 13088
rect 7668 13028 7672 13084
rect 7672 13028 7728 13084
rect 7728 13028 7732 13084
rect 7668 13024 7732 13028
rect 7748 13084 7812 13088
rect 7748 13028 7752 13084
rect 7752 13028 7808 13084
rect 7808 13028 7812 13084
rect 7748 13024 7812 13028
rect 7828 13084 7892 13088
rect 7828 13028 7832 13084
rect 7832 13028 7888 13084
rect 7888 13028 7892 13084
rect 7828 13024 7892 13028
rect 7908 13084 7972 13088
rect 7908 13028 7912 13084
rect 7912 13028 7968 13084
rect 7968 13028 7972 13084
rect 7908 13024 7972 13028
rect 11026 13084 11090 13088
rect 11026 13028 11030 13084
rect 11030 13028 11086 13084
rect 11086 13028 11090 13084
rect 11026 13024 11090 13028
rect 11106 13084 11170 13088
rect 11106 13028 11110 13084
rect 11110 13028 11166 13084
rect 11166 13028 11170 13084
rect 11106 13024 11170 13028
rect 11186 13084 11250 13088
rect 11186 13028 11190 13084
rect 11190 13028 11246 13084
rect 11246 13028 11250 13084
rect 11186 13024 11250 13028
rect 11266 13084 11330 13088
rect 11266 13028 11270 13084
rect 11270 13028 11326 13084
rect 11326 13028 11330 13084
rect 11266 13024 11330 13028
rect 14384 13084 14448 13088
rect 14384 13028 14388 13084
rect 14388 13028 14444 13084
rect 14444 13028 14448 13084
rect 14384 13024 14448 13028
rect 14464 13084 14528 13088
rect 14464 13028 14468 13084
rect 14468 13028 14524 13084
rect 14524 13028 14528 13084
rect 14464 13024 14528 13028
rect 14544 13084 14608 13088
rect 14544 13028 14548 13084
rect 14548 13028 14604 13084
rect 14604 13028 14608 13084
rect 14544 13024 14608 13028
rect 14624 13084 14688 13088
rect 14624 13028 14628 13084
rect 14628 13028 14684 13084
rect 14684 13028 14688 13084
rect 14624 13024 14688 13028
rect 2631 12540 2695 12544
rect 2631 12484 2635 12540
rect 2635 12484 2691 12540
rect 2691 12484 2695 12540
rect 2631 12480 2695 12484
rect 2711 12540 2775 12544
rect 2711 12484 2715 12540
rect 2715 12484 2771 12540
rect 2771 12484 2775 12540
rect 2711 12480 2775 12484
rect 2791 12540 2855 12544
rect 2791 12484 2795 12540
rect 2795 12484 2851 12540
rect 2851 12484 2855 12540
rect 2791 12480 2855 12484
rect 2871 12540 2935 12544
rect 2871 12484 2875 12540
rect 2875 12484 2931 12540
rect 2931 12484 2935 12540
rect 2871 12480 2935 12484
rect 5989 12540 6053 12544
rect 5989 12484 5993 12540
rect 5993 12484 6049 12540
rect 6049 12484 6053 12540
rect 5989 12480 6053 12484
rect 6069 12540 6133 12544
rect 6069 12484 6073 12540
rect 6073 12484 6129 12540
rect 6129 12484 6133 12540
rect 6069 12480 6133 12484
rect 6149 12540 6213 12544
rect 6149 12484 6153 12540
rect 6153 12484 6209 12540
rect 6209 12484 6213 12540
rect 6149 12480 6213 12484
rect 6229 12540 6293 12544
rect 6229 12484 6233 12540
rect 6233 12484 6289 12540
rect 6289 12484 6293 12540
rect 6229 12480 6293 12484
rect 9347 12540 9411 12544
rect 9347 12484 9351 12540
rect 9351 12484 9407 12540
rect 9407 12484 9411 12540
rect 9347 12480 9411 12484
rect 9427 12540 9491 12544
rect 9427 12484 9431 12540
rect 9431 12484 9487 12540
rect 9487 12484 9491 12540
rect 9427 12480 9491 12484
rect 9507 12540 9571 12544
rect 9507 12484 9511 12540
rect 9511 12484 9567 12540
rect 9567 12484 9571 12540
rect 9507 12480 9571 12484
rect 9587 12540 9651 12544
rect 9587 12484 9591 12540
rect 9591 12484 9647 12540
rect 9647 12484 9651 12540
rect 9587 12480 9651 12484
rect 12705 12540 12769 12544
rect 12705 12484 12709 12540
rect 12709 12484 12765 12540
rect 12765 12484 12769 12540
rect 12705 12480 12769 12484
rect 12785 12540 12849 12544
rect 12785 12484 12789 12540
rect 12789 12484 12845 12540
rect 12845 12484 12849 12540
rect 12785 12480 12849 12484
rect 12865 12540 12929 12544
rect 12865 12484 12869 12540
rect 12869 12484 12925 12540
rect 12925 12484 12929 12540
rect 12865 12480 12929 12484
rect 12945 12540 13009 12544
rect 12945 12484 12949 12540
rect 12949 12484 13005 12540
rect 13005 12484 13009 12540
rect 12945 12480 13009 12484
rect 4310 11996 4374 12000
rect 4310 11940 4314 11996
rect 4314 11940 4370 11996
rect 4370 11940 4374 11996
rect 4310 11936 4374 11940
rect 4390 11996 4454 12000
rect 4390 11940 4394 11996
rect 4394 11940 4450 11996
rect 4450 11940 4454 11996
rect 4390 11936 4454 11940
rect 4470 11996 4534 12000
rect 4470 11940 4474 11996
rect 4474 11940 4530 11996
rect 4530 11940 4534 11996
rect 4470 11936 4534 11940
rect 4550 11996 4614 12000
rect 4550 11940 4554 11996
rect 4554 11940 4610 11996
rect 4610 11940 4614 11996
rect 4550 11936 4614 11940
rect 7668 11996 7732 12000
rect 7668 11940 7672 11996
rect 7672 11940 7728 11996
rect 7728 11940 7732 11996
rect 7668 11936 7732 11940
rect 7748 11996 7812 12000
rect 7748 11940 7752 11996
rect 7752 11940 7808 11996
rect 7808 11940 7812 11996
rect 7748 11936 7812 11940
rect 7828 11996 7892 12000
rect 7828 11940 7832 11996
rect 7832 11940 7888 11996
rect 7888 11940 7892 11996
rect 7828 11936 7892 11940
rect 7908 11996 7972 12000
rect 7908 11940 7912 11996
rect 7912 11940 7968 11996
rect 7968 11940 7972 11996
rect 7908 11936 7972 11940
rect 11026 11996 11090 12000
rect 11026 11940 11030 11996
rect 11030 11940 11086 11996
rect 11086 11940 11090 11996
rect 11026 11936 11090 11940
rect 11106 11996 11170 12000
rect 11106 11940 11110 11996
rect 11110 11940 11166 11996
rect 11166 11940 11170 11996
rect 11106 11936 11170 11940
rect 11186 11996 11250 12000
rect 11186 11940 11190 11996
rect 11190 11940 11246 11996
rect 11246 11940 11250 11996
rect 11186 11936 11250 11940
rect 11266 11996 11330 12000
rect 11266 11940 11270 11996
rect 11270 11940 11326 11996
rect 11326 11940 11330 11996
rect 11266 11936 11330 11940
rect 14384 11996 14448 12000
rect 14384 11940 14388 11996
rect 14388 11940 14444 11996
rect 14444 11940 14448 11996
rect 14384 11936 14448 11940
rect 14464 11996 14528 12000
rect 14464 11940 14468 11996
rect 14468 11940 14524 11996
rect 14524 11940 14528 11996
rect 14464 11936 14528 11940
rect 14544 11996 14608 12000
rect 14544 11940 14548 11996
rect 14548 11940 14604 11996
rect 14604 11940 14608 11996
rect 14544 11936 14608 11940
rect 14624 11996 14688 12000
rect 14624 11940 14628 11996
rect 14628 11940 14684 11996
rect 14684 11940 14688 11996
rect 14624 11936 14688 11940
rect 2631 11452 2695 11456
rect 2631 11396 2635 11452
rect 2635 11396 2691 11452
rect 2691 11396 2695 11452
rect 2631 11392 2695 11396
rect 2711 11452 2775 11456
rect 2711 11396 2715 11452
rect 2715 11396 2771 11452
rect 2771 11396 2775 11452
rect 2711 11392 2775 11396
rect 2791 11452 2855 11456
rect 2791 11396 2795 11452
rect 2795 11396 2851 11452
rect 2851 11396 2855 11452
rect 2791 11392 2855 11396
rect 2871 11452 2935 11456
rect 2871 11396 2875 11452
rect 2875 11396 2931 11452
rect 2931 11396 2935 11452
rect 2871 11392 2935 11396
rect 5989 11452 6053 11456
rect 5989 11396 5993 11452
rect 5993 11396 6049 11452
rect 6049 11396 6053 11452
rect 5989 11392 6053 11396
rect 6069 11452 6133 11456
rect 6069 11396 6073 11452
rect 6073 11396 6129 11452
rect 6129 11396 6133 11452
rect 6069 11392 6133 11396
rect 6149 11452 6213 11456
rect 6149 11396 6153 11452
rect 6153 11396 6209 11452
rect 6209 11396 6213 11452
rect 6149 11392 6213 11396
rect 6229 11452 6293 11456
rect 6229 11396 6233 11452
rect 6233 11396 6289 11452
rect 6289 11396 6293 11452
rect 6229 11392 6293 11396
rect 9347 11452 9411 11456
rect 9347 11396 9351 11452
rect 9351 11396 9407 11452
rect 9407 11396 9411 11452
rect 9347 11392 9411 11396
rect 9427 11452 9491 11456
rect 9427 11396 9431 11452
rect 9431 11396 9487 11452
rect 9487 11396 9491 11452
rect 9427 11392 9491 11396
rect 9507 11452 9571 11456
rect 9507 11396 9511 11452
rect 9511 11396 9567 11452
rect 9567 11396 9571 11452
rect 9507 11392 9571 11396
rect 9587 11452 9651 11456
rect 9587 11396 9591 11452
rect 9591 11396 9647 11452
rect 9647 11396 9651 11452
rect 9587 11392 9651 11396
rect 12705 11452 12769 11456
rect 12705 11396 12709 11452
rect 12709 11396 12765 11452
rect 12765 11396 12769 11452
rect 12705 11392 12769 11396
rect 12785 11452 12849 11456
rect 12785 11396 12789 11452
rect 12789 11396 12845 11452
rect 12845 11396 12849 11452
rect 12785 11392 12849 11396
rect 12865 11452 12929 11456
rect 12865 11396 12869 11452
rect 12869 11396 12925 11452
rect 12925 11396 12929 11452
rect 12865 11392 12929 11396
rect 12945 11452 13009 11456
rect 12945 11396 12949 11452
rect 12949 11396 13005 11452
rect 13005 11396 13009 11452
rect 12945 11392 13009 11396
rect 3740 11052 3804 11116
rect 4310 10908 4374 10912
rect 4310 10852 4314 10908
rect 4314 10852 4370 10908
rect 4370 10852 4374 10908
rect 4310 10848 4374 10852
rect 4390 10908 4454 10912
rect 4390 10852 4394 10908
rect 4394 10852 4450 10908
rect 4450 10852 4454 10908
rect 4390 10848 4454 10852
rect 4470 10908 4534 10912
rect 4470 10852 4474 10908
rect 4474 10852 4530 10908
rect 4530 10852 4534 10908
rect 4470 10848 4534 10852
rect 4550 10908 4614 10912
rect 4550 10852 4554 10908
rect 4554 10852 4610 10908
rect 4610 10852 4614 10908
rect 4550 10848 4614 10852
rect 7668 10908 7732 10912
rect 7668 10852 7672 10908
rect 7672 10852 7728 10908
rect 7728 10852 7732 10908
rect 7668 10848 7732 10852
rect 7748 10908 7812 10912
rect 7748 10852 7752 10908
rect 7752 10852 7808 10908
rect 7808 10852 7812 10908
rect 7748 10848 7812 10852
rect 7828 10908 7892 10912
rect 7828 10852 7832 10908
rect 7832 10852 7888 10908
rect 7888 10852 7892 10908
rect 7828 10848 7892 10852
rect 7908 10908 7972 10912
rect 7908 10852 7912 10908
rect 7912 10852 7968 10908
rect 7968 10852 7972 10908
rect 7908 10848 7972 10852
rect 11026 10908 11090 10912
rect 11026 10852 11030 10908
rect 11030 10852 11086 10908
rect 11086 10852 11090 10908
rect 11026 10848 11090 10852
rect 11106 10908 11170 10912
rect 11106 10852 11110 10908
rect 11110 10852 11166 10908
rect 11166 10852 11170 10908
rect 11106 10848 11170 10852
rect 11186 10908 11250 10912
rect 11186 10852 11190 10908
rect 11190 10852 11246 10908
rect 11246 10852 11250 10908
rect 11186 10848 11250 10852
rect 11266 10908 11330 10912
rect 11266 10852 11270 10908
rect 11270 10852 11326 10908
rect 11326 10852 11330 10908
rect 11266 10848 11330 10852
rect 14384 10908 14448 10912
rect 14384 10852 14388 10908
rect 14388 10852 14444 10908
rect 14444 10852 14448 10908
rect 14384 10848 14448 10852
rect 14464 10908 14528 10912
rect 14464 10852 14468 10908
rect 14468 10852 14524 10908
rect 14524 10852 14528 10908
rect 14464 10848 14528 10852
rect 14544 10908 14608 10912
rect 14544 10852 14548 10908
rect 14548 10852 14604 10908
rect 14604 10852 14608 10908
rect 14544 10848 14608 10852
rect 14624 10908 14688 10912
rect 14624 10852 14628 10908
rect 14628 10852 14684 10908
rect 14684 10852 14688 10908
rect 14624 10848 14688 10852
rect 11468 10644 11532 10708
rect 12572 10508 12636 10572
rect 2631 10364 2695 10368
rect 2631 10308 2635 10364
rect 2635 10308 2691 10364
rect 2691 10308 2695 10364
rect 2631 10304 2695 10308
rect 2711 10364 2775 10368
rect 2711 10308 2715 10364
rect 2715 10308 2771 10364
rect 2771 10308 2775 10364
rect 2711 10304 2775 10308
rect 2791 10364 2855 10368
rect 2791 10308 2795 10364
rect 2795 10308 2851 10364
rect 2851 10308 2855 10364
rect 2791 10304 2855 10308
rect 2871 10364 2935 10368
rect 2871 10308 2875 10364
rect 2875 10308 2931 10364
rect 2931 10308 2935 10364
rect 2871 10304 2935 10308
rect 5989 10364 6053 10368
rect 5989 10308 5993 10364
rect 5993 10308 6049 10364
rect 6049 10308 6053 10364
rect 5989 10304 6053 10308
rect 6069 10364 6133 10368
rect 6069 10308 6073 10364
rect 6073 10308 6129 10364
rect 6129 10308 6133 10364
rect 6069 10304 6133 10308
rect 6149 10364 6213 10368
rect 6149 10308 6153 10364
rect 6153 10308 6209 10364
rect 6209 10308 6213 10364
rect 6149 10304 6213 10308
rect 6229 10364 6293 10368
rect 6229 10308 6233 10364
rect 6233 10308 6289 10364
rect 6289 10308 6293 10364
rect 6229 10304 6293 10308
rect 9347 10364 9411 10368
rect 9347 10308 9351 10364
rect 9351 10308 9407 10364
rect 9407 10308 9411 10364
rect 9347 10304 9411 10308
rect 9427 10364 9491 10368
rect 9427 10308 9431 10364
rect 9431 10308 9487 10364
rect 9487 10308 9491 10364
rect 9427 10304 9491 10308
rect 9507 10364 9571 10368
rect 9507 10308 9511 10364
rect 9511 10308 9567 10364
rect 9567 10308 9571 10364
rect 9507 10304 9571 10308
rect 9587 10364 9651 10368
rect 9587 10308 9591 10364
rect 9591 10308 9647 10364
rect 9647 10308 9651 10364
rect 9587 10304 9651 10308
rect 12705 10364 12769 10368
rect 12705 10308 12709 10364
rect 12709 10308 12765 10364
rect 12765 10308 12769 10364
rect 12705 10304 12769 10308
rect 12785 10364 12849 10368
rect 12785 10308 12789 10364
rect 12789 10308 12845 10364
rect 12845 10308 12849 10364
rect 12785 10304 12849 10308
rect 12865 10364 12929 10368
rect 12865 10308 12869 10364
rect 12869 10308 12925 10364
rect 12925 10308 12929 10364
rect 12865 10304 12929 10308
rect 12945 10364 13009 10368
rect 12945 10308 12949 10364
rect 12949 10308 13005 10364
rect 13005 10308 13009 10364
rect 12945 10304 13009 10308
rect 4310 9820 4374 9824
rect 4310 9764 4314 9820
rect 4314 9764 4370 9820
rect 4370 9764 4374 9820
rect 4310 9760 4374 9764
rect 4390 9820 4454 9824
rect 4390 9764 4394 9820
rect 4394 9764 4450 9820
rect 4450 9764 4454 9820
rect 4390 9760 4454 9764
rect 4470 9820 4534 9824
rect 4470 9764 4474 9820
rect 4474 9764 4530 9820
rect 4530 9764 4534 9820
rect 4470 9760 4534 9764
rect 4550 9820 4614 9824
rect 4550 9764 4554 9820
rect 4554 9764 4610 9820
rect 4610 9764 4614 9820
rect 4550 9760 4614 9764
rect 7668 9820 7732 9824
rect 7668 9764 7672 9820
rect 7672 9764 7728 9820
rect 7728 9764 7732 9820
rect 7668 9760 7732 9764
rect 7748 9820 7812 9824
rect 7748 9764 7752 9820
rect 7752 9764 7808 9820
rect 7808 9764 7812 9820
rect 7748 9760 7812 9764
rect 7828 9820 7892 9824
rect 7828 9764 7832 9820
rect 7832 9764 7888 9820
rect 7888 9764 7892 9820
rect 7828 9760 7892 9764
rect 7908 9820 7972 9824
rect 7908 9764 7912 9820
rect 7912 9764 7968 9820
rect 7968 9764 7972 9820
rect 7908 9760 7972 9764
rect 11026 9820 11090 9824
rect 11026 9764 11030 9820
rect 11030 9764 11086 9820
rect 11086 9764 11090 9820
rect 11026 9760 11090 9764
rect 11106 9820 11170 9824
rect 11106 9764 11110 9820
rect 11110 9764 11166 9820
rect 11166 9764 11170 9820
rect 11106 9760 11170 9764
rect 11186 9820 11250 9824
rect 11186 9764 11190 9820
rect 11190 9764 11246 9820
rect 11246 9764 11250 9820
rect 11186 9760 11250 9764
rect 11266 9820 11330 9824
rect 11266 9764 11270 9820
rect 11270 9764 11326 9820
rect 11326 9764 11330 9820
rect 11266 9760 11330 9764
rect 14384 9820 14448 9824
rect 14384 9764 14388 9820
rect 14388 9764 14444 9820
rect 14444 9764 14448 9820
rect 14384 9760 14448 9764
rect 14464 9820 14528 9824
rect 14464 9764 14468 9820
rect 14468 9764 14524 9820
rect 14524 9764 14528 9820
rect 14464 9760 14528 9764
rect 14544 9820 14608 9824
rect 14544 9764 14548 9820
rect 14548 9764 14604 9820
rect 14604 9764 14608 9820
rect 14544 9760 14608 9764
rect 14624 9820 14688 9824
rect 14624 9764 14628 9820
rect 14628 9764 14684 9820
rect 14684 9764 14688 9820
rect 14624 9760 14688 9764
rect 13124 9692 13188 9756
rect 10732 9420 10796 9484
rect 10180 9344 10244 9348
rect 10180 9288 10194 9344
rect 10194 9288 10244 9344
rect 10180 9284 10244 9288
rect 2631 9276 2695 9280
rect 2631 9220 2635 9276
rect 2635 9220 2691 9276
rect 2691 9220 2695 9276
rect 2631 9216 2695 9220
rect 2711 9276 2775 9280
rect 2711 9220 2715 9276
rect 2715 9220 2771 9276
rect 2771 9220 2775 9276
rect 2711 9216 2775 9220
rect 2791 9276 2855 9280
rect 2791 9220 2795 9276
rect 2795 9220 2851 9276
rect 2851 9220 2855 9276
rect 2791 9216 2855 9220
rect 2871 9276 2935 9280
rect 2871 9220 2875 9276
rect 2875 9220 2931 9276
rect 2931 9220 2935 9276
rect 2871 9216 2935 9220
rect 5989 9276 6053 9280
rect 5989 9220 5993 9276
rect 5993 9220 6049 9276
rect 6049 9220 6053 9276
rect 5989 9216 6053 9220
rect 6069 9276 6133 9280
rect 6069 9220 6073 9276
rect 6073 9220 6129 9276
rect 6129 9220 6133 9276
rect 6069 9216 6133 9220
rect 6149 9276 6213 9280
rect 6149 9220 6153 9276
rect 6153 9220 6209 9276
rect 6209 9220 6213 9276
rect 6149 9216 6213 9220
rect 6229 9276 6293 9280
rect 6229 9220 6233 9276
rect 6233 9220 6289 9276
rect 6289 9220 6293 9276
rect 6229 9216 6293 9220
rect 9347 9276 9411 9280
rect 9347 9220 9351 9276
rect 9351 9220 9407 9276
rect 9407 9220 9411 9276
rect 9347 9216 9411 9220
rect 9427 9276 9491 9280
rect 9427 9220 9431 9276
rect 9431 9220 9487 9276
rect 9487 9220 9491 9276
rect 9427 9216 9491 9220
rect 9507 9276 9571 9280
rect 9507 9220 9511 9276
rect 9511 9220 9567 9276
rect 9567 9220 9571 9276
rect 9507 9216 9571 9220
rect 9587 9276 9651 9280
rect 9587 9220 9591 9276
rect 9591 9220 9647 9276
rect 9647 9220 9651 9276
rect 9587 9216 9651 9220
rect 12705 9276 12769 9280
rect 12705 9220 12709 9276
rect 12709 9220 12765 9276
rect 12765 9220 12769 9276
rect 12705 9216 12769 9220
rect 12785 9276 12849 9280
rect 12785 9220 12789 9276
rect 12789 9220 12845 9276
rect 12845 9220 12849 9276
rect 12785 9216 12849 9220
rect 12865 9276 12929 9280
rect 12865 9220 12869 9276
rect 12869 9220 12925 9276
rect 12925 9220 12929 9276
rect 12865 9216 12929 9220
rect 12945 9276 13009 9280
rect 12945 9220 12949 9276
rect 12949 9220 13005 9276
rect 13005 9220 13009 9276
rect 12945 9216 13009 9220
rect 8892 8740 8956 8804
rect 4310 8732 4374 8736
rect 4310 8676 4314 8732
rect 4314 8676 4370 8732
rect 4370 8676 4374 8732
rect 4310 8672 4374 8676
rect 4390 8732 4454 8736
rect 4390 8676 4394 8732
rect 4394 8676 4450 8732
rect 4450 8676 4454 8732
rect 4390 8672 4454 8676
rect 4470 8732 4534 8736
rect 4470 8676 4474 8732
rect 4474 8676 4530 8732
rect 4530 8676 4534 8732
rect 4470 8672 4534 8676
rect 4550 8732 4614 8736
rect 4550 8676 4554 8732
rect 4554 8676 4610 8732
rect 4610 8676 4614 8732
rect 4550 8672 4614 8676
rect 7668 8732 7732 8736
rect 7668 8676 7672 8732
rect 7672 8676 7728 8732
rect 7728 8676 7732 8732
rect 7668 8672 7732 8676
rect 7748 8732 7812 8736
rect 7748 8676 7752 8732
rect 7752 8676 7808 8732
rect 7808 8676 7812 8732
rect 7748 8672 7812 8676
rect 7828 8732 7892 8736
rect 7828 8676 7832 8732
rect 7832 8676 7888 8732
rect 7888 8676 7892 8732
rect 7828 8672 7892 8676
rect 7908 8732 7972 8736
rect 7908 8676 7912 8732
rect 7912 8676 7968 8732
rect 7968 8676 7972 8732
rect 7908 8672 7972 8676
rect 11026 8732 11090 8736
rect 11026 8676 11030 8732
rect 11030 8676 11086 8732
rect 11086 8676 11090 8732
rect 11026 8672 11090 8676
rect 11106 8732 11170 8736
rect 11106 8676 11110 8732
rect 11110 8676 11166 8732
rect 11166 8676 11170 8732
rect 11106 8672 11170 8676
rect 11186 8732 11250 8736
rect 11186 8676 11190 8732
rect 11190 8676 11246 8732
rect 11246 8676 11250 8732
rect 11186 8672 11250 8676
rect 11266 8732 11330 8736
rect 11266 8676 11270 8732
rect 11270 8676 11326 8732
rect 11326 8676 11330 8732
rect 11266 8672 11330 8676
rect 14384 8732 14448 8736
rect 14384 8676 14388 8732
rect 14388 8676 14444 8732
rect 14444 8676 14448 8732
rect 14384 8672 14448 8676
rect 14464 8732 14528 8736
rect 14464 8676 14468 8732
rect 14468 8676 14524 8732
rect 14524 8676 14528 8732
rect 14464 8672 14528 8676
rect 14544 8732 14608 8736
rect 14544 8676 14548 8732
rect 14548 8676 14604 8732
rect 14604 8676 14608 8732
rect 14544 8672 14608 8676
rect 14624 8732 14688 8736
rect 14624 8676 14628 8732
rect 14628 8676 14684 8732
rect 14684 8676 14688 8732
rect 14624 8672 14688 8676
rect 9812 8664 9876 8668
rect 9812 8608 9862 8664
rect 9862 8608 9876 8664
rect 9812 8604 9876 8608
rect 2631 8188 2695 8192
rect 2631 8132 2635 8188
rect 2635 8132 2691 8188
rect 2691 8132 2695 8188
rect 2631 8128 2695 8132
rect 2711 8188 2775 8192
rect 2711 8132 2715 8188
rect 2715 8132 2771 8188
rect 2771 8132 2775 8188
rect 2711 8128 2775 8132
rect 2791 8188 2855 8192
rect 2791 8132 2795 8188
rect 2795 8132 2851 8188
rect 2851 8132 2855 8188
rect 2791 8128 2855 8132
rect 2871 8188 2935 8192
rect 2871 8132 2875 8188
rect 2875 8132 2931 8188
rect 2931 8132 2935 8188
rect 2871 8128 2935 8132
rect 5989 8188 6053 8192
rect 5989 8132 5993 8188
rect 5993 8132 6049 8188
rect 6049 8132 6053 8188
rect 5989 8128 6053 8132
rect 6069 8188 6133 8192
rect 6069 8132 6073 8188
rect 6073 8132 6129 8188
rect 6129 8132 6133 8188
rect 6069 8128 6133 8132
rect 6149 8188 6213 8192
rect 6149 8132 6153 8188
rect 6153 8132 6209 8188
rect 6209 8132 6213 8188
rect 6149 8128 6213 8132
rect 6229 8188 6293 8192
rect 6229 8132 6233 8188
rect 6233 8132 6289 8188
rect 6289 8132 6293 8188
rect 6229 8128 6293 8132
rect 9347 8188 9411 8192
rect 9347 8132 9351 8188
rect 9351 8132 9407 8188
rect 9407 8132 9411 8188
rect 9347 8128 9411 8132
rect 9427 8188 9491 8192
rect 9427 8132 9431 8188
rect 9431 8132 9487 8188
rect 9487 8132 9491 8188
rect 9427 8128 9491 8132
rect 9507 8188 9571 8192
rect 9507 8132 9511 8188
rect 9511 8132 9567 8188
rect 9567 8132 9571 8188
rect 9507 8128 9571 8132
rect 9587 8188 9651 8192
rect 9587 8132 9591 8188
rect 9591 8132 9647 8188
rect 9647 8132 9651 8188
rect 9587 8128 9651 8132
rect 12705 8188 12769 8192
rect 12705 8132 12709 8188
rect 12709 8132 12765 8188
rect 12765 8132 12769 8188
rect 12705 8128 12769 8132
rect 12785 8188 12849 8192
rect 12785 8132 12789 8188
rect 12789 8132 12845 8188
rect 12845 8132 12849 8188
rect 12785 8128 12849 8132
rect 12865 8188 12929 8192
rect 12865 8132 12869 8188
rect 12869 8132 12925 8188
rect 12925 8132 12929 8188
rect 12865 8128 12929 8132
rect 12945 8188 13009 8192
rect 12945 8132 12949 8188
rect 12949 8132 13005 8188
rect 13005 8132 13009 8188
rect 12945 8128 13009 8132
rect 8156 8060 8220 8124
rect 8892 7652 8956 7716
rect 4310 7644 4374 7648
rect 4310 7588 4314 7644
rect 4314 7588 4370 7644
rect 4370 7588 4374 7644
rect 4310 7584 4374 7588
rect 4390 7644 4454 7648
rect 4390 7588 4394 7644
rect 4394 7588 4450 7644
rect 4450 7588 4454 7644
rect 4390 7584 4454 7588
rect 4470 7644 4534 7648
rect 4470 7588 4474 7644
rect 4474 7588 4530 7644
rect 4530 7588 4534 7644
rect 4470 7584 4534 7588
rect 4550 7644 4614 7648
rect 4550 7588 4554 7644
rect 4554 7588 4610 7644
rect 4610 7588 4614 7644
rect 4550 7584 4614 7588
rect 7668 7644 7732 7648
rect 7668 7588 7672 7644
rect 7672 7588 7728 7644
rect 7728 7588 7732 7644
rect 7668 7584 7732 7588
rect 7748 7644 7812 7648
rect 7748 7588 7752 7644
rect 7752 7588 7808 7644
rect 7808 7588 7812 7644
rect 7748 7584 7812 7588
rect 7828 7644 7892 7648
rect 7828 7588 7832 7644
rect 7832 7588 7888 7644
rect 7888 7588 7892 7644
rect 7828 7584 7892 7588
rect 7908 7644 7972 7648
rect 7908 7588 7912 7644
rect 7912 7588 7968 7644
rect 7968 7588 7972 7644
rect 7908 7584 7972 7588
rect 11026 7644 11090 7648
rect 11026 7588 11030 7644
rect 11030 7588 11086 7644
rect 11086 7588 11090 7644
rect 11026 7584 11090 7588
rect 11106 7644 11170 7648
rect 11106 7588 11110 7644
rect 11110 7588 11166 7644
rect 11166 7588 11170 7644
rect 11106 7584 11170 7588
rect 11186 7644 11250 7648
rect 11186 7588 11190 7644
rect 11190 7588 11246 7644
rect 11246 7588 11250 7644
rect 11186 7584 11250 7588
rect 11266 7644 11330 7648
rect 11266 7588 11270 7644
rect 11270 7588 11326 7644
rect 11326 7588 11330 7644
rect 11266 7584 11330 7588
rect 14384 7644 14448 7648
rect 14384 7588 14388 7644
rect 14388 7588 14444 7644
rect 14444 7588 14448 7644
rect 14384 7584 14448 7588
rect 14464 7644 14528 7648
rect 14464 7588 14468 7644
rect 14468 7588 14524 7644
rect 14524 7588 14528 7644
rect 14464 7584 14528 7588
rect 14544 7644 14608 7648
rect 14544 7588 14548 7644
rect 14548 7588 14604 7644
rect 14604 7588 14608 7644
rect 14544 7584 14608 7588
rect 14624 7644 14688 7648
rect 14624 7588 14628 7644
rect 14628 7588 14684 7644
rect 14684 7588 14688 7644
rect 14624 7584 14688 7588
rect 2631 7100 2695 7104
rect 2631 7044 2635 7100
rect 2635 7044 2691 7100
rect 2691 7044 2695 7100
rect 2631 7040 2695 7044
rect 2711 7100 2775 7104
rect 2711 7044 2715 7100
rect 2715 7044 2771 7100
rect 2771 7044 2775 7100
rect 2711 7040 2775 7044
rect 2791 7100 2855 7104
rect 2791 7044 2795 7100
rect 2795 7044 2851 7100
rect 2851 7044 2855 7100
rect 2791 7040 2855 7044
rect 2871 7100 2935 7104
rect 2871 7044 2875 7100
rect 2875 7044 2931 7100
rect 2931 7044 2935 7100
rect 2871 7040 2935 7044
rect 5989 7100 6053 7104
rect 5989 7044 5993 7100
rect 5993 7044 6049 7100
rect 6049 7044 6053 7100
rect 5989 7040 6053 7044
rect 6069 7100 6133 7104
rect 6069 7044 6073 7100
rect 6073 7044 6129 7100
rect 6129 7044 6133 7100
rect 6069 7040 6133 7044
rect 6149 7100 6213 7104
rect 6149 7044 6153 7100
rect 6153 7044 6209 7100
rect 6209 7044 6213 7100
rect 6149 7040 6213 7044
rect 6229 7100 6293 7104
rect 6229 7044 6233 7100
rect 6233 7044 6289 7100
rect 6289 7044 6293 7100
rect 6229 7040 6293 7044
rect 9347 7100 9411 7104
rect 9347 7044 9351 7100
rect 9351 7044 9407 7100
rect 9407 7044 9411 7100
rect 9347 7040 9411 7044
rect 9427 7100 9491 7104
rect 9427 7044 9431 7100
rect 9431 7044 9487 7100
rect 9487 7044 9491 7100
rect 9427 7040 9491 7044
rect 9507 7100 9571 7104
rect 9507 7044 9511 7100
rect 9511 7044 9567 7100
rect 9567 7044 9571 7100
rect 9507 7040 9571 7044
rect 9587 7100 9651 7104
rect 9587 7044 9591 7100
rect 9591 7044 9647 7100
rect 9647 7044 9651 7100
rect 9587 7040 9651 7044
rect 12705 7100 12769 7104
rect 12705 7044 12709 7100
rect 12709 7044 12765 7100
rect 12765 7044 12769 7100
rect 12705 7040 12769 7044
rect 12785 7100 12849 7104
rect 12785 7044 12789 7100
rect 12789 7044 12845 7100
rect 12845 7044 12849 7100
rect 12785 7040 12849 7044
rect 12865 7100 12929 7104
rect 12865 7044 12869 7100
rect 12869 7044 12925 7100
rect 12925 7044 12929 7100
rect 12865 7040 12929 7044
rect 12945 7100 13009 7104
rect 12945 7044 12949 7100
rect 12949 7044 13005 7100
rect 13005 7044 13009 7100
rect 12945 7040 13009 7044
rect 9812 6760 9876 6764
rect 9812 6704 9826 6760
rect 9826 6704 9876 6760
rect 9812 6700 9876 6704
rect 4310 6556 4374 6560
rect 4310 6500 4314 6556
rect 4314 6500 4370 6556
rect 4370 6500 4374 6556
rect 4310 6496 4374 6500
rect 4390 6556 4454 6560
rect 4390 6500 4394 6556
rect 4394 6500 4450 6556
rect 4450 6500 4454 6556
rect 4390 6496 4454 6500
rect 4470 6556 4534 6560
rect 4470 6500 4474 6556
rect 4474 6500 4530 6556
rect 4530 6500 4534 6556
rect 4470 6496 4534 6500
rect 4550 6556 4614 6560
rect 4550 6500 4554 6556
rect 4554 6500 4610 6556
rect 4610 6500 4614 6556
rect 4550 6496 4614 6500
rect 7668 6556 7732 6560
rect 7668 6500 7672 6556
rect 7672 6500 7728 6556
rect 7728 6500 7732 6556
rect 7668 6496 7732 6500
rect 7748 6556 7812 6560
rect 7748 6500 7752 6556
rect 7752 6500 7808 6556
rect 7808 6500 7812 6556
rect 7748 6496 7812 6500
rect 7828 6556 7892 6560
rect 7828 6500 7832 6556
rect 7832 6500 7888 6556
rect 7888 6500 7892 6556
rect 7828 6496 7892 6500
rect 7908 6556 7972 6560
rect 7908 6500 7912 6556
rect 7912 6500 7968 6556
rect 7968 6500 7972 6556
rect 7908 6496 7972 6500
rect 11026 6556 11090 6560
rect 11026 6500 11030 6556
rect 11030 6500 11086 6556
rect 11086 6500 11090 6556
rect 11026 6496 11090 6500
rect 11106 6556 11170 6560
rect 11106 6500 11110 6556
rect 11110 6500 11166 6556
rect 11166 6500 11170 6556
rect 11106 6496 11170 6500
rect 11186 6556 11250 6560
rect 11186 6500 11190 6556
rect 11190 6500 11246 6556
rect 11246 6500 11250 6556
rect 11186 6496 11250 6500
rect 11266 6556 11330 6560
rect 11266 6500 11270 6556
rect 11270 6500 11326 6556
rect 11326 6500 11330 6556
rect 11266 6496 11330 6500
rect 14384 6556 14448 6560
rect 14384 6500 14388 6556
rect 14388 6500 14444 6556
rect 14444 6500 14448 6556
rect 14384 6496 14448 6500
rect 14464 6556 14528 6560
rect 14464 6500 14468 6556
rect 14468 6500 14524 6556
rect 14524 6500 14528 6556
rect 14464 6496 14528 6500
rect 14544 6556 14608 6560
rect 14544 6500 14548 6556
rect 14548 6500 14604 6556
rect 14604 6500 14608 6556
rect 14544 6496 14608 6500
rect 14624 6556 14688 6560
rect 14624 6500 14628 6556
rect 14628 6500 14684 6556
rect 14684 6500 14688 6556
rect 14624 6496 14688 6500
rect 8156 6216 8220 6220
rect 8156 6160 8206 6216
rect 8206 6160 8220 6216
rect 8156 6156 8220 6160
rect 2631 6012 2695 6016
rect 2631 5956 2635 6012
rect 2635 5956 2691 6012
rect 2691 5956 2695 6012
rect 2631 5952 2695 5956
rect 2711 6012 2775 6016
rect 2711 5956 2715 6012
rect 2715 5956 2771 6012
rect 2771 5956 2775 6012
rect 2711 5952 2775 5956
rect 2791 6012 2855 6016
rect 2791 5956 2795 6012
rect 2795 5956 2851 6012
rect 2851 5956 2855 6012
rect 2791 5952 2855 5956
rect 2871 6012 2935 6016
rect 2871 5956 2875 6012
rect 2875 5956 2931 6012
rect 2931 5956 2935 6012
rect 2871 5952 2935 5956
rect 5989 6012 6053 6016
rect 5989 5956 5993 6012
rect 5993 5956 6049 6012
rect 6049 5956 6053 6012
rect 5989 5952 6053 5956
rect 6069 6012 6133 6016
rect 6069 5956 6073 6012
rect 6073 5956 6129 6012
rect 6129 5956 6133 6012
rect 6069 5952 6133 5956
rect 6149 6012 6213 6016
rect 6149 5956 6153 6012
rect 6153 5956 6209 6012
rect 6209 5956 6213 6012
rect 6149 5952 6213 5956
rect 6229 6012 6293 6016
rect 6229 5956 6233 6012
rect 6233 5956 6289 6012
rect 6289 5956 6293 6012
rect 6229 5952 6293 5956
rect 9347 6012 9411 6016
rect 9347 5956 9351 6012
rect 9351 5956 9407 6012
rect 9407 5956 9411 6012
rect 9347 5952 9411 5956
rect 9427 6012 9491 6016
rect 9427 5956 9431 6012
rect 9431 5956 9487 6012
rect 9487 5956 9491 6012
rect 9427 5952 9491 5956
rect 9507 6012 9571 6016
rect 9507 5956 9511 6012
rect 9511 5956 9567 6012
rect 9567 5956 9571 6012
rect 9507 5952 9571 5956
rect 9587 6012 9651 6016
rect 9587 5956 9591 6012
rect 9591 5956 9647 6012
rect 9647 5956 9651 6012
rect 9587 5952 9651 5956
rect 12705 6012 12769 6016
rect 12705 5956 12709 6012
rect 12709 5956 12765 6012
rect 12765 5956 12769 6012
rect 12705 5952 12769 5956
rect 12785 6012 12849 6016
rect 12785 5956 12789 6012
rect 12789 5956 12845 6012
rect 12845 5956 12849 6012
rect 12785 5952 12849 5956
rect 12865 6012 12929 6016
rect 12865 5956 12869 6012
rect 12869 5956 12925 6012
rect 12925 5956 12929 6012
rect 12865 5952 12929 5956
rect 12945 6012 13009 6016
rect 12945 5956 12949 6012
rect 12949 5956 13005 6012
rect 13005 5956 13009 6012
rect 12945 5952 13009 5956
rect 14964 5612 15028 5676
rect 4310 5468 4374 5472
rect 4310 5412 4314 5468
rect 4314 5412 4370 5468
rect 4370 5412 4374 5468
rect 4310 5408 4374 5412
rect 4390 5468 4454 5472
rect 4390 5412 4394 5468
rect 4394 5412 4450 5468
rect 4450 5412 4454 5468
rect 4390 5408 4454 5412
rect 4470 5468 4534 5472
rect 4470 5412 4474 5468
rect 4474 5412 4530 5468
rect 4530 5412 4534 5468
rect 4470 5408 4534 5412
rect 4550 5468 4614 5472
rect 4550 5412 4554 5468
rect 4554 5412 4610 5468
rect 4610 5412 4614 5468
rect 4550 5408 4614 5412
rect 7668 5468 7732 5472
rect 7668 5412 7672 5468
rect 7672 5412 7728 5468
rect 7728 5412 7732 5468
rect 7668 5408 7732 5412
rect 7748 5468 7812 5472
rect 7748 5412 7752 5468
rect 7752 5412 7808 5468
rect 7808 5412 7812 5468
rect 7748 5408 7812 5412
rect 7828 5468 7892 5472
rect 7828 5412 7832 5468
rect 7832 5412 7888 5468
rect 7888 5412 7892 5468
rect 7828 5408 7892 5412
rect 7908 5468 7972 5472
rect 7908 5412 7912 5468
rect 7912 5412 7968 5468
rect 7968 5412 7972 5468
rect 7908 5408 7972 5412
rect 11026 5468 11090 5472
rect 11026 5412 11030 5468
rect 11030 5412 11086 5468
rect 11086 5412 11090 5468
rect 11026 5408 11090 5412
rect 11106 5468 11170 5472
rect 11106 5412 11110 5468
rect 11110 5412 11166 5468
rect 11166 5412 11170 5468
rect 11106 5408 11170 5412
rect 11186 5468 11250 5472
rect 11186 5412 11190 5468
rect 11190 5412 11246 5468
rect 11246 5412 11250 5468
rect 11186 5408 11250 5412
rect 11266 5468 11330 5472
rect 11266 5412 11270 5468
rect 11270 5412 11326 5468
rect 11326 5412 11330 5468
rect 11266 5408 11330 5412
rect 14384 5468 14448 5472
rect 14384 5412 14388 5468
rect 14388 5412 14444 5468
rect 14444 5412 14448 5468
rect 14384 5408 14448 5412
rect 14464 5468 14528 5472
rect 14464 5412 14468 5468
rect 14468 5412 14524 5468
rect 14524 5412 14528 5468
rect 14464 5408 14528 5412
rect 14544 5468 14608 5472
rect 14544 5412 14548 5468
rect 14548 5412 14604 5468
rect 14604 5412 14608 5468
rect 14544 5408 14608 5412
rect 14624 5468 14688 5472
rect 14624 5412 14628 5468
rect 14628 5412 14684 5468
rect 14684 5412 14688 5468
rect 14624 5408 14688 5412
rect 2631 4924 2695 4928
rect 2631 4868 2635 4924
rect 2635 4868 2691 4924
rect 2691 4868 2695 4924
rect 2631 4864 2695 4868
rect 2711 4924 2775 4928
rect 2711 4868 2715 4924
rect 2715 4868 2771 4924
rect 2771 4868 2775 4924
rect 2711 4864 2775 4868
rect 2791 4924 2855 4928
rect 2791 4868 2795 4924
rect 2795 4868 2851 4924
rect 2851 4868 2855 4924
rect 2791 4864 2855 4868
rect 2871 4924 2935 4928
rect 2871 4868 2875 4924
rect 2875 4868 2931 4924
rect 2931 4868 2935 4924
rect 2871 4864 2935 4868
rect 5989 4924 6053 4928
rect 5989 4868 5993 4924
rect 5993 4868 6049 4924
rect 6049 4868 6053 4924
rect 5989 4864 6053 4868
rect 6069 4924 6133 4928
rect 6069 4868 6073 4924
rect 6073 4868 6129 4924
rect 6129 4868 6133 4924
rect 6069 4864 6133 4868
rect 6149 4924 6213 4928
rect 6149 4868 6153 4924
rect 6153 4868 6209 4924
rect 6209 4868 6213 4924
rect 6149 4864 6213 4868
rect 6229 4924 6293 4928
rect 6229 4868 6233 4924
rect 6233 4868 6289 4924
rect 6289 4868 6293 4924
rect 6229 4864 6293 4868
rect 9347 4924 9411 4928
rect 9347 4868 9351 4924
rect 9351 4868 9407 4924
rect 9407 4868 9411 4924
rect 9347 4864 9411 4868
rect 9427 4924 9491 4928
rect 9427 4868 9431 4924
rect 9431 4868 9487 4924
rect 9487 4868 9491 4924
rect 9427 4864 9491 4868
rect 9507 4924 9571 4928
rect 9507 4868 9511 4924
rect 9511 4868 9567 4924
rect 9567 4868 9571 4924
rect 9507 4864 9571 4868
rect 9587 4924 9651 4928
rect 9587 4868 9591 4924
rect 9591 4868 9647 4924
rect 9647 4868 9651 4924
rect 9587 4864 9651 4868
rect 12705 4924 12769 4928
rect 12705 4868 12709 4924
rect 12709 4868 12765 4924
rect 12765 4868 12769 4924
rect 12705 4864 12769 4868
rect 12785 4924 12849 4928
rect 12785 4868 12789 4924
rect 12789 4868 12845 4924
rect 12845 4868 12849 4924
rect 12785 4864 12849 4868
rect 12865 4924 12929 4928
rect 12865 4868 12869 4924
rect 12869 4868 12925 4924
rect 12925 4868 12929 4924
rect 12865 4864 12929 4868
rect 12945 4924 13009 4928
rect 12945 4868 12949 4924
rect 12949 4868 13005 4924
rect 13005 4868 13009 4924
rect 12945 4864 13009 4868
rect 4310 4380 4374 4384
rect 4310 4324 4314 4380
rect 4314 4324 4370 4380
rect 4370 4324 4374 4380
rect 4310 4320 4374 4324
rect 4390 4380 4454 4384
rect 4390 4324 4394 4380
rect 4394 4324 4450 4380
rect 4450 4324 4454 4380
rect 4390 4320 4454 4324
rect 4470 4380 4534 4384
rect 4470 4324 4474 4380
rect 4474 4324 4530 4380
rect 4530 4324 4534 4380
rect 4470 4320 4534 4324
rect 4550 4380 4614 4384
rect 4550 4324 4554 4380
rect 4554 4324 4610 4380
rect 4610 4324 4614 4380
rect 4550 4320 4614 4324
rect 7668 4380 7732 4384
rect 7668 4324 7672 4380
rect 7672 4324 7728 4380
rect 7728 4324 7732 4380
rect 7668 4320 7732 4324
rect 7748 4380 7812 4384
rect 7748 4324 7752 4380
rect 7752 4324 7808 4380
rect 7808 4324 7812 4380
rect 7748 4320 7812 4324
rect 7828 4380 7892 4384
rect 7828 4324 7832 4380
rect 7832 4324 7888 4380
rect 7888 4324 7892 4380
rect 7828 4320 7892 4324
rect 7908 4380 7972 4384
rect 7908 4324 7912 4380
rect 7912 4324 7968 4380
rect 7968 4324 7972 4380
rect 7908 4320 7972 4324
rect 11026 4380 11090 4384
rect 11026 4324 11030 4380
rect 11030 4324 11086 4380
rect 11086 4324 11090 4380
rect 11026 4320 11090 4324
rect 11106 4380 11170 4384
rect 11106 4324 11110 4380
rect 11110 4324 11166 4380
rect 11166 4324 11170 4380
rect 11106 4320 11170 4324
rect 11186 4380 11250 4384
rect 11186 4324 11190 4380
rect 11190 4324 11246 4380
rect 11246 4324 11250 4380
rect 11186 4320 11250 4324
rect 11266 4380 11330 4384
rect 11266 4324 11270 4380
rect 11270 4324 11326 4380
rect 11326 4324 11330 4380
rect 11266 4320 11330 4324
rect 14384 4380 14448 4384
rect 14384 4324 14388 4380
rect 14388 4324 14444 4380
rect 14444 4324 14448 4380
rect 14384 4320 14448 4324
rect 14464 4380 14528 4384
rect 14464 4324 14468 4380
rect 14468 4324 14524 4380
rect 14524 4324 14528 4380
rect 14464 4320 14528 4324
rect 14544 4380 14608 4384
rect 14544 4324 14548 4380
rect 14548 4324 14604 4380
rect 14604 4324 14608 4380
rect 14544 4320 14608 4324
rect 14624 4380 14688 4384
rect 14624 4324 14628 4380
rect 14628 4324 14684 4380
rect 14684 4324 14688 4380
rect 14624 4320 14688 4324
rect 2631 3836 2695 3840
rect 2631 3780 2635 3836
rect 2635 3780 2691 3836
rect 2691 3780 2695 3836
rect 2631 3776 2695 3780
rect 2711 3836 2775 3840
rect 2711 3780 2715 3836
rect 2715 3780 2771 3836
rect 2771 3780 2775 3836
rect 2711 3776 2775 3780
rect 2791 3836 2855 3840
rect 2791 3780 2795 3836
rect 2795 3780 2851 3836
rect 2851 3780 2855 3836
rect 2791 3776 2855 3780
rect 2871 3836 2935 3840
rect 2871 3780 2875 3836
rect 2875 3780 2931 3836
rect 2931 3780 2935 3836
rect 2871 3776 2935 3780
rect 5989 3836 6053 3840
rect 5989 3780 5993 3836
rect 5993 3780 6049 3836
rect 6049 3780 6053 3836
rect 5989 3776 6053 3780
rect 6069 3836 6133 3840
rect 6069 3780 6073 3836
rect 6073 3780 6129 3836
rect 6129 3780 6133 3836
rect 6069 3776 6133 3780
rect 6149 3836 6213 3840
rect 6149 3780 6153 3836
rect 6153 3780 6209 3836
rect 6209 3780 6213 3836
rect 6149 3776 6213 3780
rect 6229 3836 6293 3840
rect 6229 3780 6233 3836
rect 6233 3780 6289 3836
rect 6289 3780 6293 3836
rect 6229 3776 6293 3780
rect 9347 3836 9411 3840
rect 9347 3780 9351 3836
rect 9351 3780 9407 3836
rect 9407 3780 9411 3836
rect 9347 3776 9411 3780
rect 9427 3836 9491 3840
rect 9427 3780 9431 3836
rect 9431 3780 9487 3836
rect 9487 3780 9491 3836
rect 9427 3776 9491 3780
rect 9507 3836 9571 3840
rect 9507 3780 9511 3836
rect 9511 3780 9567 3836
rect 9567 3780 9571 3836
rect 9507 3776 9571 3780
rect 9587 3836 9651 3840
rect 9587 3780 9591 3836
rect 9591 3780 9647 3836
rect 9647 3780 9651 3836
rect 9587 3776 9651 3780
rect 12705 3836 12769 3840
rect 12705 3780 12709 3836
rect 12709 3780 12765 3836
rect 12765 3780 12769 3836
rect 12705 3776 12769 3780
rect 12785 3836 12849 3840
rect 12785 3780 12789 3836
rect 12789 3780 12845 3836
rect 12845 3780 12849 3836
rect 12785 3776 12849 3780
rect 12865 3836 12929 3840
rect 12865 3780 12869 3836
rect 12869 3780 12925 3836
rect 12925 3780 12929 3836
rect 12865 3776 12929 3780
rect 12945 3836 13009 3840
rect 12945 3780 12949 3836
rect 12949 3780 13005 3836
rect 13005 3780 13009 3836
rect 12945 3776 13009 3780
rect 4310 3292 4374 3296
rect 4310 3236 4314 3292
rect 4314 3236 4370 3292
rect 4370 3236 4374 3292
rect 4310 3232 4374 3236
rect 4390 3292 4454 3296
rect 4390 3236 4394 3292
rect 4394 3236 4450 3292
rect 4450 3236 4454 3292
rect 4390 3232 4454 3236
rect 4470 3292 4534 3296
rect 4470 3236 4474 3292
rect 4474 3236 4530 3292
rect 4530 3236 4534 3292
rect 4470 3232 4534 3236
rect 4550 3292 4614 3296
rect 4550 3236 4554 3292
rect 4554 3236 4610 3292
rect 4610 3236 4614 3292
rect 4550 3232 4614 3236
rect 7668 3292 7732 3296
rect 7668 3236 7672 3292
rect 7672 3236 7728 3292
rect 7728 3236 7732 3292
rect 7668 3232 7732 3236
rect 7748 3292 7812 3296
rect 7748 3236 7752 3292
rect 7752 3236 7808 3292
rect 7808 3236 7812 3292
rect 7748 3232 7812 3236
rect 7828 3292 7892 3296
rect 7828 3236 7832 3292
rect 7832 3236 7888 3292
rect 7888 3236 7892 3292
rect 7828 3232 7892 3236
rect 7908 3292 7972 3296
rect 7908 3236 7912 3292
rect 7912 3236 7968 3292
rect 7968 3236 7972 3292
rect 7908 3232 7972 3236
rect 11026 3292 11090 3296
rect 11026 3236 11030 3292
rect 11030 3236 11086 3292
rect 11086 3236 11090 3292
rect 11026 3232 11090 3236
rect 11106 3292 11170 3296
rect 11106 3236 11110 3292
rect 11110 3236 11166 3292
rect 11166 3236 11170 3292
rect 11106 3232 11170 3236
rect 11186 3292 11250 3296
rect 11186 3236 11190 3292
rect 11190 3236 11246 3292
rect 11246 3236 11250 3292
rect 11186 3232 11250 3236
rect 11266 3292 11330 3296
rect 11266 3236 11270 3292
rect 11270 3236 11326 3292
rect 11326 3236 11330 3292
rect 11266 3232 11330 3236
rect 14384 3292 14448 3296
rect 14384 3236 14388 3292
rect 14388 3236 14444 3292
rect 14444 3236 14448 3292
rect 14384 3232 14448 3236
rect 14464 3292 14528 3296
rect 14464 3236 14468 3292
rect 14468 3236 14524 3292
rect 14524 3236 14528 3292
rect 14464 3232 14528 3236
rect 14544 3292 14608 3296
rect 14544 3236 14548 3292
rect 14548 3236 14604 3292
rect 14604 3236 14608 3292
rect 14544 3232 14608 3236
rect 14624 3292 14688 3296
rect 14624 3236 14628 3292
rect 14628 3236 14684 3292
rect 14684 3236 14688 3292
rect 14624 3232 14688 3236
rect 2631 2748 2695 2752
rect 2631 2692 2635 2748
rect 2635 2692 2691 2748
rect 2691 2692 2695 2748
rect 2631 2688 2695 2692
rect 2711 2748 2775 2752
rect 2711 2692 2715 2748
rect 2715 2692 2771 2748
rect 2771 2692 2775 2748
rect 2711 2688 2775 2692
rect 2791 2748 2855 2752
rect 2791 2692 2795 2748
rect 2795 2692 2851 2748
rect 2851 2692 2855 2748
rect 2791 2688 2855 2692
rect 2871 2748 2935 2752
rect 2871 2692 2875 2748
rect 2875 2692 2931 2748
rect 2931 2692 2935 2748
rect 2871 2688 2935 2692
rect 5989 2748 6053 2752
rect 5989 2692 5993 2748
rect 5993 2692 6049 2748
rect 6049 2692 6053 2748
rect 5989 2688 6053 2692
rect 6069 2748 6133 2752
rect 6069 2692 6073 2748
rect 6073 2692 6129 2748
rect 6129 2692 6133 2748
rect 6069 2688 6133 2692
rect 6149 2748 6213 2752
rect 6149 2692 6153 2748
rect 6153 2692 6209 2748
rect 6209 2692 6213 2748
rect 6149 2688 6213 2692
rect 6229 2748 6293 2752
rect 6229 2692 6233 2748
rect 6233 2692 6289 2748
rect 6289 2692 6293 2748
rect 6229 2688 6293 2692
rect 9347 2748 9411 2752
rect 9347 2692 9351 2748
rect 9351 2692 9407 2748
rect 9407 2692 9411 2748
rect 9347 2688 9411 2692
rect 9427 2748 9491 2752
rect 9427 2692 9431 2748
rect 9431 2692 9487 2748
rect 9487 2692 9491 2748
rect 9427 2688 9491 2692
rect 9507 2748 9571 2752
rect 9507 2692 9511 2748
rect 9511 2692 9567 2748
rect 9567 2692 9571 2748
rect 9507 2688 9571 2692
rect 9587 2748 9651 2752
rect 9587 2692 9591 2748
rect 9591 2692 9647 2748
rect 9647 2692 9651 2748
rect 9587 2688 9651 2692
rect 12705 2748 12769 2752
rect 12705 2692 12709 2748
rect 12709 2692 12765 2748
rect 12765 2692 12769 2748
rect 12705 2688 12769 2692
rect 12785 2748 12849 2752
rect 12785 2692 12789 2748
rect 12789 2692 12845 2748
rect 12845 2692 12849 2748
rect 12785 2688 12849 2692
rect 12865 2748 12929 2752
rect 12865 2692 12869 2748
rect 12869 2692 12925 2748
rect 12925 2692 12929 2748
rect 12865 2688 12929 2692
rect 12945 2748 13009 2752
rect 12945 2692 12949 2748
rect 12949 2692 13005 2748
rect 13005 2692 13009 2748
rect 12945 2688 13009 2692
rect 6684 2680 6748 2684
rect 6684 2624 6698 2680
rect 6698 2624 6748 2680
rect 6684 2620 6748 2624
rect 10364 2620 10428 2684
rect 2084 2484 2148 2548
rect 9076 2484 9140 2548
rect 2268 2348 2332 2412
rect 4310 2204 4374 2208
rect 4310 2148 4314 2204
rect 4314 2148 4370 2204
rect 4370 2148 4374 2204
rect 4310 2144 4374 2148
rect 4390 2204 4454 2208
rect 4390 2148 4394 2204
rect 4394 2148 4450 2204
rect 4450 2148 4454 2204
rect 4390 2144 4454 2148
rect 4470 2204 4534 2208
rect 4470 2148 4474 2204
rect 4474 2148 4530 2204
rect 4530 2148 4534 2204
rect 4470 2144 4534 2148
rect 4550 2204 4614 2208
rect 4550 2148 4554 2204
rect 4554 2148 4610 2204
rect 4610 2148 4614 2204
rect 4550 2144 4614 2148
rect 7668 2204 7732 2208
rect 7668 2148 7672 2204
rect 7672 2148 7728 2204
rect 7728 2148 7732 2204
rect 7668 2144 7732 2148
rect 7748 2204 7812 2208
rect 7748 2148 7752 2204
rect 7752 2148 7808 2204
rect 7808 2148 7812 2204
rect 7748 2144 7812 2148
rect 7828 2204 7892 2208
rect 7828 2148 7832 2204
rect 7832 2148 7888 2204
rect 7888 2148 7892 2204
rect 7828 2144 7892 2148
rect 7908 2204 7972 2208
rect 7908 2148 7912 2204
rect 7912 2148 7968 2204
rect 7968 2148 7972 2204
rect 7908 2144 7972 2148
rect 11026 2204 11090 2208
rect 11026 2148 11030 2204
rect 11030 2148 11086 2204
rect 11086 2148 11090 2204
rect 11026 2144 11090 2148
rect 11106 2204 11170 2208
rect 11106 2148 11110 2204
rect 11110 2148 11166 2204
rect 11166 2148 11170 2204
rect 11106 2144 11170 2148
rect 11186 2204 11250 2208
rect 11186 2148 11190 2204
rect 11190 2148 11246 2204
rect 11246 2148 11250 2204
rect 11186 2144 11250 2148
rect 11266 2204 11330 2208
rect 11266 2148 11270 2204
rect 11270 2148 11326 2204
rect 11326 2148 11330 2204
rect 11266 2144 11330 2148
rect 14384 2204 14448 2208
rect 14384 2148 14388 2204
rect 14388 2148 14444 2204
rect 14444 2148 14448 2204
rect 14384 2144 14448 2148
rect 14464 2204 14528 2208
rect 14464 2148 14468 2204
rect 14468 2148 14524 2204
rect 14524 2148 14528 2204
rect 14464 2144 14528 2148
rect 14544 2204 14608 2208
rect 14544 2148 14548 2204
rect 14548 2148 14604 2204
rect 14604 2148 14608 2204
rect 14544 2144 14608 2148
rect 14624 2204 14688 2208
rect 14624 2148 14628 2204
rect 14628 2148 14684 2204
rect 14684 2148 14688 2204
rect 14624 2144 14688 2148
rect 3924 1940 3988 2004
rect 2631 1660 2695 1664
rect 2631 1604 2635 1660
rect 2635 1604 2691 1660
rect 2691 1604 2695 1660
rect 2631 1600 2695 1604
rect 2711 1660 2775 1664
rect 2711 1604 2715 1660
rect 2715 1604 2771 1660
rect 2771 1604 2775 1660
rect 2711 1600 2775 1604
rect 2791 1660 2855 1664
rect 2791 1604 2795 1660
rect 2795 1604 2851 1660
rect 2851 1604 2855 1660
rect 2791 1600 2855 1604
rect 2871 1660 2935 1664
rect 2871 1604 2875 1660
rect 2875 1604 2931 1660
rect 2931 1604 2935 1660
rect 2871 1600 2935 1604
rect 5989 1660 6053 1664
rect 5989 1604 5993 1660
rect 5993 1604 6049 1660
rect 6049 1604 6053 1660
rect 5989 1600 6053 1604
rect 6069 1660 6133 1664
rect 6069 1604 6073 1660
rect 6073 1604 6129 1660
rect 6129 1604 6133 1660
rect 6069 1600 6133 1604
rect 6149 1660 6213 1664
rect 6149 1604 6153 1660
rect 6153 1604 6209 1660
rect 6209 1604 6213 1660
rect 6149 1600 6213 1604
rect 6229 1660 6293 1664
rect 6229 1604 6233 1660
rect 6233 1604 6289 1660
rect 6289 1604 6293 1660
rect 6229 1600 6293 1604
rect 9347 1660 9411 1664
rect 9347 1604 9351 1660
rect 9351 1604 9407 1660
rect 9407 1604 9411 1660
rect 9347 1600 9411 1604
rect 9427 1660 9491 1664
rect 9427 1604 9431 1660
rect 9431 1604 9487 1660
rect 9487 1604 9491 1660
rect 9427 1600 9491 1604
rect 9507 1660 9571 1664
rect 9507 1604 9511 1660
rect 9511 1604 9567 1660
rect 9567 1604 9571 1660
rect 9507 1600 9571 1604
rect 9587 1660 9651 1664
rect 9587 1604 9591 1660
rect 9591 1604 9647 1660
rect 9647 1604 9651 1660
rect 9587 1600 9651 1604
rect 12705 1660 12769 1664
rect 12705 1604 12709 1660
rect 12709 1604 12765 1660
rect 12765 1604 12769 1660
rect 12705 1600 12769 1604
rect 12785 1660 12849 1664
rect 12785 1604 12789 1660
rect 12789 1604 12845 1660
rect 12845 1604 12849 1660
rect 12785 1600 12849 1604
rect 12865 1660 12929 1664
rect 12865 1604 12869 1660
rect 12869 1604 12925 1660
rect 12925 1604 12929 1660
rect 12865 1600 12929 1604
rect 12945 1660 13009 1664
rect 12945 1604 12949 1660
rect 12949 1604 13005 1660
rect 13005 1604 13009 1660
rect 12945 1600 13009 1604
rect 4844 1260 4908 1324
rect 5212 1320 5276 1324
rect 5212 1264 5226 1320
rect 5226 1264 5276 1320
rect 5212 1260 5276 1264
rect 6500 1260 6564 1324
rect 8708 1260 8772 1324
rect 4310 1116 4374 1120
rect 4310 1060 4314 1116
rect 4314 1060 4370 1116
rect 4370 1060 4374 1116
rect 4310 1056 4374 1060
rect 4390 1116 4454 1120
rect 4390 1060 4394 1116
rect 4394 1060 4450 1116
rect 4450 1060 4454 1116
rect 4390 1056 4454 1060
rect 4470 1116 4534 1120
rect 4470 1060 4474 1116
rect 4474 1060 4530 1116
rect 4530 1060 4534 1116
rect 4470 1056 4534 1060
rect 4550 1116 4614 1120
rect 4550 1060 4554 1116
rect 4554 1060 4610 1116
rect 4610 1060 4614 1116
rect 4550 1056 4614 1060
rect 7668 1116 7732 1120
rect 7668 1060 7672 1116
rect 7672 1060 7728 1116
rect 7728 1060 7732 1116
rect 7668 1056 7732 1060
rect 7748 1116 7812 1120
rect 7748 1060 7752 1116
rect 7752 1060 7808 1116
rect 7808 1060 7812 1116
rect 7748 1056 7812 1060
rect 7828 1116 7892 1120
rect 7828 1060 7832 1116
rect 7832 1060 7888 1116
rect 7888 1060 7892 1116
rect 7828 1056 7892 1060
rect 7908 1116 7972 1120
rect 7908 1060 7912 1116
rect 7912 1060 7968 1116
rect 7968 1060 7972 1116
rect 7908 1056 7972 1060
rect 11026 1116 11090 1120
rect 11026 1060 11030 1116
rect 11030 1060 11086 1116
rect 11086 1060 11090 1116
rect 11026 1056 11090 1060
rect 11106 1116 11170 1120
rect 11106 1060 11110 1116
rect 11110 1060 11166 1116
rect 11166 1060 11170 1116
rect 11106 1056 11170 1060
rect 11186 1116 11250 1120
rect 11186 1060 11190 1116
rect 11190 1060 11246 1116
rect 11246 1060 11250 1116
rect 11186 1056 11250 1060
rect 11266 1116 11330 1120
rect 11266 1060 11270 1116
rect 11270 1060 11326 1116
rect 11326 1060 11330 1116
rect 11266 1056 11330 1060
rect 14384 1116 14448 1120
rect 14384 1060 14388 1116
rect 14388 1060 14444 1116
rect 14444 1060 14448 1116
rect 14384 1056 14448 1060
rect 14464 1116 14528 1120
rect 14464 1060 14468 1116
rect 14468 1060 14524 1116
rect 14524 1060 14528 1116
rect 14464 1056 14528 1060
rect 14544 1116 14608 1120
rect 14544 1060 14548 1116
rect 14548 1060 14604 1116
rect 14604 1060 14608 1116
rect 14544 1056 14608 1060
rect 14624 1116 14688 1120
rect 14624 1060 14628 1116
rect 14628 1060 14684 1116
rect 14684 1060 14688 1116
rect 14624 1056 14688 1060
<< metal4 >>
rect 2623 43008 2943 43568
rect 2623 42944 2631 43008
rect 2695 42944 2711 43008
rect 2775 42944 2791 43008
rect 2855 42944 2871 43008
rect 2935 42944 2943 43008
rect 2267 42124 2333 42125
rect 2267 42060 2268 42124
rect 2332 42060 2333 42124
rect 2267 42059 2333 42060
rect 2083 41716 2149 41717
rect 2083 41652 2084 41716
rect 2148 41652 2149 41716
rect 2083 41651 2149 41652
rect 1531 41444 1597 41445
rect 1531 41380 1532 41444
rect 1596 41380 1597 41444
rect 1531 41379 1597 41380
rect 1534 20501 1594 41379
rect 1531 20500 1597 20501
rect 1531 20436 1532 20500
rect 1596 20436 1597 20500
rect 1531 20435 1597 20436
rect 2086 2549 2146 41651
rect 2083 2548 2149 2549
rect 2083 2484 2084 2548
rect 2148 2484 2149 2548
rect 2083 2483 2149 2484
rect 2270 2413 2330 42059
rect 2623 41920 2943 42944
rect 4302 43552 4622 43568
rect 4302 43488 4310 43552
rect 4374 43488 4390 43552
rect 4454 43488 4470 43552
rect 4534 43488 4550 43552
rect 4614 43488 4622 43552
rect 3923 42804 3989 42805
rect 3923 42740 3924 42804
rect 3988 42740 3989 42804
rect 3923 42739 3989 42740
rect 3739 42668 3805 42669
rect 3739 42604 3740 42668
rect 3804 42604 3805 42668
rect 3739 42603 3805 42604
rect 2623 41856 2631 41920
rect 2695 41856 2711 41920
rect 2775 41856 2791 41920
rect 2855 41856 2871 41920
rect 2935 41856 2943 41920
rect 2623 40832 2943 41856
rect 2623 40768 2631 40832
rect 2695 40768 2711 40832
rect 2775 40768 2791 40832
rect 2855 40768 2871 40832
rect 2935 40768 2943 40832
rect 2623 39744 2943 40768
rect 2623 39680 2631 39744
rect 2695 39680 2711 39744
rect 2775 39680 2791 39744
rect 2855 39680 2871 39744
rect 2935 39680 2943 39744
rect 2623 38656 2943 39680
rect 2623 38592 2631 38656
rect 2695 38592 2711 38656
rect 2775 38592 2791 38656
rect 2855 38592 2871 38656
rect 2935 38592 2943 38656
rect 2623 37568 2943 38592
rect 2623 37504 2631 37568
rect 2695 37504 2711 37568
rect 2775 37504 2791 37568
rect 2855 37504 2871 37568
rect 2935 37504 2943 37568
rect 2623 36480 2943 37504
rect 2623 36416 2631 36480
rect 2695 36416 2711 36480
rect 2775 36416 2791 36480
rect 2855 36416 2871 36480
rect 2935 36416 2943 36480
rect 2623 35392 2943 36416
rect 2623 35328 2631 35392
rect 2695 35328 2711 35392
rect 2775 35328 2791 35392
rect 2855 35328 2871 35392
rect 2935 35328 2943 35392
rect 2623 34304 2943 35328
rect 2623 34240 2631 34304
rect 2695 34240 2711 34304
rect 2775 34240 2791 34304
rect 2855 34240 2871 34304
rect 2935 34240 2943 34304
rect 2623 33216 2943 34240
rect 2623 33152 2631 33216
rect 2695 33152 2711 33216
rect 2775 33152 2791 33216
rect 2855 33152 2871 33216
rect 2935 33152 2943 33216
rect 2623 32128 2943 33152
rect 2623 32064 2631 32128
rect 2695 32064 2711 32128
rect 2775 32064 2791 32128
rect 2855 32064 2871 32128
rect 2935 32064 2943 32128
rect 2623 31040 2943 32064
rect 2623 30976 2631 31040
rect 2695 30976 2711 31040
rect 2775 30976 2791 31040
rect 2855 30976 2871 31040
rect 2935 30976 2943 31040
rect 2623 29952 2943 30976
rect 2623 29888 2631 29952
rect 2695 29888 2711 29952
rect 2775 29888 2791 29952
rect 2855 29888 2871 29952
rect 2935 29888 2943 29952
rect 2623 28864 2943 29888
rect 2623 28800 2631 28864
rect 2695 28800 2711 28864
rect 2775 28800 2791 28864
rect 2855 28800 2871 28864
rect 2935 28800 2943 28864
rect 2623 27776 2943 28800
rect 2623 27712 2631 27776
rect 2695 27712 2711 27776
rect 2775 27712 2791 27776
rect 2855 27712 2871 27776
rect 2935 27712 2943 27776
rect 2623 26688 2943 27712
rect 2623 26624 2631 26688
rect 2695 26624 2711 26688
rect 2775 26624 2791 26688
rect 2855 26624 2871 26688
rect 2935 26624 2943 26688
rect 2623 25600 2943 26624
rect 2623 25536 2631 25600
rect 2695 25536 2711 25600
rect 2775 25536 2791 25600
rect 2855 25536 2871 25600
rect 2935 25536 2943 25600
rect 2623 24512 2943 25536
rect 2623 24448 2631 24512
rect 2695 24448 2711 24512
rect 2775 24448 2791 24512
rect 2855 24448 2871 24512
rect 2935 24448 2943 24512
rect 2623 23424 2943 24448
rect 2623 23360 2631 23424
rect 2695 23360 2711 23424
rect 2775 23360 2791 23424
rect 2855 23360 2871 23424
rect 2935 23360 2943 23424
rect 2623 22336 2943 23360
rect 2623 22272 2631 22336
rect 2695 22272 2711 22336
rect 2775 22272 2791 22336
rect 2855 22272 2871 22336
rect 2935 22272 2943 22336
rect 2623 21248 2943 22272
rect 2623 21184 2631 21248
rect 2695 21184 2711 21248
rect 2775 21184 2791 21248
rect 2855 21184 2871 21248
rect 2935 21184 2943 21248
rect 2623 20160 2943 21184
rect 2623 20096 2631 20160
rect 2695 20096 2711 20160
rect 2775 20096 2791 20160
rect 2855 20096 2871 20160
rect 2935 20096 2943 20160
rect 2623 19072 2943 20096
rect 2623 19008 2631 19072
rect 2695 19008 2711 19072
rect 2775 19008 2791 19072
rect 2855 19008 2871 19072
rect 2935 19008 2943 19072
rect 2623 17984 2943 19008
rect 2623 17920 2631 17984
rect 2695 17920 2711 17984
rect 2775 17920 2791 17984
rect 2855 17920 2871 17984
rect 2935 17920 2943 17984
rect 2623 16896 2943 17920
rect 2623 16832 2631 16896
rect 2695 16832 2711 16896
rect 2775 16832 2791 16896
rect 2855 16832 2871 16896
rect 2935 16832 2943 16896
rect 2623 15808 2943 16832
rect 2623 15744 2631 15808
rect 2695 15744 2711 15808
rect 2775 15744 2791 15808
rect 2855 15744 2871 15808
rect 2935 15744 2943 15808
rect 2623 14720 2943 15744
rect 2623 14656 2631 14720
rect 2695 14656 2711 14720
rect 2775 14656 2791 14720
rect 2855 14656 2871 14720
rect 2935 14656 2943 14720
rect 2623 13632 2943 14656
rect 2623 13568 2631 13632
rect 2695 13568 2711 13632
rect 2775 13568 2791 13632
rect 2855 13568 2871 13632
rect 2935 13568 2943 13632
rect 2623 12544 2943 13568
rect 2623 12480 2631 12544
rect 2695 12480 2711 12544
rect 2775 12480 2791 12544
rect 2855 12480 2871 12544
rect 2935 12480 2943 12544
rect 2623 11456 2943 12480
rect 2623 11392 2631 11456
rect 2695 11392 2711 11456
rect 2775 11392 2791 11456
rect 2855 11392 2871 11456
rect 2935 11392 2943 11456
rect 2623 10368 2943 11392
rect 3742 11117 3802 42603
rect 3739 11116 3805 11117
rect 3739 11052 3740 11116
rect 3804 11052 3805 11116
rect 3739 11051 3805 11052
rect 2623 10304 2631 10368
rect 2695 10304 2711 10368
rect 2775 10304 2791 10368
rect 2855 10304 2871 10368
rect 2935 10304 2943 10368
rect 2623 9280 2943 10304
rect 2623 9216 2631 9280
rect 2695 9216 2711 9280
rect 2775 9216 2791 9280
rect 2855 9216 2871 9280
rect 2935 9216 2943 9280
rect 2623 8192 2943 9216
rect 2623 8128 2631 8192
rect 2695 8128 2711 8192
rect 2775 8128 2791 8192
rect 2855 8128 2871 8192
rect 2935 8128 2943 8192
rect 2623 7104 2943 8128
rect 2623 7040 2631 7104
rect 2695 7040 2711 7104
rect 2775 7040 2791 7104
rect 2855 7040 2871 7104
rect 2935 7040 2943 7104
rect 2623 6016 2943 7040
rect 2623 5952 2631 6016
rect 2695 5952 2711 6016
rect 2775 5952 2791 6016
rect 2855 5952 2871 6016
rect 2935 5952 2943 6016
rect 2623 4928 2943 5952
rect 2623 4864 2631 4928
rect 2695 4864 2711 4928
rect 2775 4864 2791 4928
rect 2855 4864 2871 4928
rect 2935 4864 2943 4928
rect 2623 3840 2943 4864
rect 2623 3776 2631 3840
rect 2695 3776 2711 3840
rect 2775 3776 2791 3840
rect 2855 3776 2871 3840
rect 2935 3776 2943 3840
rect 2623 2752 2943 3776
rect 2623 2688 2631 2752
rect 2695 2688 2711 2752
rect 2775 2688 2791 2752
rect 2855 2688 2871 2752
rect 2935 2688 2943 2752
rect 2267 2412 2333 2413
rect 2267 2348 2268 2412
rect 2332 2348 2333 2412
rect 2267 2347 2333 2348
rect 2623 1664 2943 2688
rect 3926 2005 3986 42739
rect 4302 42464 4622 43488
rect 4302 42400 4310 42464
rect 4374 42400 4390 42464
rect 4454 42400 4470 42464
rect 4534 42400 4550 42464
rect 4614 42400 4622 42464
rect 4302 41376 4622 42400
rect 5981 43008 6301 43568
rect 5981 42944 5989 43008
rect 6053 42944 6069 43008
rect 6133 42944 6149 43008
rect 6213 42944 6229 43008
rect 6293 42944 6301 43008
rect 5981 41920 6301 42944
rect 5981 41856 5989 41920
rect 6053 41856 6069 41920
rect 6133 41856 6149 41920
rect 6213 41856 6229 41920
rect 6293 41856 6301 41920
rect 4843 41580 4909 41581
rect 4843 41516 4844 41580
rect 4908 41516 4909 41580
rect 4843 41515 4909 41516
rect 4302 41312 4310 41376
rect 4374 41312 4390 41376
rect 4454 41312 4470 41376
rect 4534 41312 4550 41376
rect 4614 41312 4622 41376
rect 4302 40288 4622 41312
rect 4302 40224 4310 40288
rect 4374 40224 4390 40288
rect 4454 40224 4470 40288
rect 4534 40224 4550 40288
rect 4614 40224 4622 40288
rect 4302 39200 4622 40224
rect 4302 39136 4310 39200
rect 4374 39136 4390 39200
rect 4454 39136 4470 39200
rect 4534 39136 4550 39200
rect 4614 39136 4622 39200
rect 4302 38112 4622 39136
rect 4302 38048 4310 38112
rect 4374 38048 4390 38112
rect 4454 38048 4470 38112
rect 4534 38048 4550 38112
rect 4614 38048 4622 38112
rect 4302 37024 4622 38048
rect 4302 36960 4310 37024
rect 4374 36960 4390 37024
rect 4454 36960 4470 37024
rect 4534 36960 4550 37024
rect 4614 36960 4622 37024
rect 4302 35936 4622 36960
rect 4302 35872 4310 35936
rect 4374 35872 4390 35936
rect 4454 35872 4470 35936
rect 4534 35872 4550 35936
rect 4614 35872 4622 35936
rect 4302 34848 4622 35872
rect 4302 34784 4310 34848
rect 4374 34784 4390 34848
rect 4454 34784 4470 34848
rect 4534 34784 4550 34848
rect 4614 34784 4622 34848
rect 4302 33760 4622 34784
rect 4302 33696 4310 33760
rect 4374 33696 4390 33760
rect 4454 33696 4470 33760
rect 4534 33696 4550 33760
rect 4614 33696 4622 33760
rect 4302 32672 4622 33696
rect 4302 32608 4310 32672
rect 4374 32608 4390 32672
rect 4454 32608 4470 32672
rect 4534 32608 4550 32672
rect 4614 32608 4622 32672
rect 4302 31584 4622 32608
rect 4302 31520 4310 31584
rect 4374 31520 4390 31584
rect 4454 31520 4470 31584
rect 4534 31520 4550 31584
rect 4614 31520 4622 31584
rect 4302 30496 4622 31520
rect 4302 30432 4310 30496
rect 4374 30432 4390 30496
rect 4454 30432 4470 30496
rect 4534 30432 4550 30496
rect 4614 30432 4622 30496
rect 4302 29408 4622 30432
rect 4302 29344 4310 29408
rect 4374 29344 4390 29408
rect 4454 29344 4470 29408
rect 4534 29344 4550 29408
rect 4614 29344 4622 29408
rect 4302 28320 4622 29344
rect 4302 28256 4310 28320
rect 4374 28256 4390 28320
rect 4454 28256 4470 28320
rect 4534 28256 4550 28320
rect 4614 28256 4622 28320
rect 4302 27232 4622 28256
rect 4302 27168 4310 27232
rect 4374 27168 4390 27232
rect 4454 27168 4470 27232
rect 4534 27168 4550 27232
rect 4614 27168 4622 27232
rect 4302 26144 4622 27168
rect 4302 26080 4310 26144
rect 4374 26080 4390 26144
rect 4454 26080 4470 26144
rect 4534 26080 4550 26144
rect 4614 26080 4622 26144
rect 4302 25056 4622 26080
rect 4302 24992 4310 25056
rect 4374 24992 4390 25056
rect 4454 24992 4470 25056
rect 4534 24992 4550 25056
rect 4614 24992 4622 25056
rect 4302 23968 4622 24992
rect 4302 23904 4310 23968
rect 4374 23904 4390 23968
rect 4454 23904 4470 23968
rect 4534 23904 4550 23968
rect 4614 23904 4622 23968
rect 4302 22880 4622 23904
rect 4302 22816 4310 22880
rect 4374 22816 4390 22880
rect 4454 22816 4470 22880
rect 4534 22816 4550 22880
rect 4614 22816 4622 22880
rect 4302 21792 4622 22816
rect 4302 21728 4310 21792
rect 4374 21728 4390 21792
rect 4454 21728 4470 21792
rect 4534 21728 4550 21792
rect 4614 21728 4622 21792
rect 4302 20704 4622 21728
rect 4302 20640 4310 20704
rect 4374 20640 4390 20704
rect 4454 20640 4470 20704
rect 4534 20640 4550 20704
rect 4614 20640 4622 20704
rect 4302 19616 4622 20640
rect 4302 19552 4310 19616
rect 4374 19552 4390 19616
rect 4454 19552 4470 19616
rect 4534 19552 4550 19616
rect 4614 19552 4622 19616
rect 4302 18528 4622 19552
rect 4302 18464 4310 18528
rect 4374 18464 4390 18528
rect 4454 18464 4470 18528
rect 4534 18464 4550 18528
rect 4614 18464 4622 18528
rect 4302 17440 4622 18464
rect 4302 17376 4310 17440
rect 4374 17376 4390 17440
rect 4454 17376 4470 17440
rect 4534 17376 4550 17440
rect 4614 17376 4622 17440
rect 4302 16352 4622 17376
rect 4302 16288 4310 16352
rect 4374 16288 4390 16352
rect 4454 16288 4470 16352
rect 4534 16288 4550 16352
rect 4614 16288 4622 16352
rect 4302 15264 4622 16288
rect 4302 15200 4310 15264
rect 4374 15200 4390 15264
rect 4454 15200 4470 15264
rect 4534 15200 4550 15264
rect 4614 15200 4622 15264
rect 4302 14176 4622 15200
rect 4302 14112 4310 14176
rect 4374 14112 4390 14176
rect 4454 14112 4470 14176
rect 4534 14112 4550 14176
rect 4614 14112 4622 14176
rect 4302 13088 4622 14112
rect 4302 13024 4310 13088
rect 4374 13024 4390 13088
rect 4454 13024 4470 13088
rect 4534 13024 4550 13088
rect 4614 13024 4622 13088
rect 4302 12000 4622 13024
rect 4302 11936 4310 12000
rect 4374 11936 4390 12000
rect 4454 11936 4470 12000
rect 4534 11936 4550 12000
rect 4614 11936 4622 12000
rect 4302 10912 4622 11936
rect 4302 10848 4310 10912
rect 4374 10848 4390 10912
rect 4454 10848 4470 10912
rect 4534 10848 4550 10912
rect 4614 10848 4622 10912
rect 4302 9824 4622 10848
rect 4302 9760 4310 9824
rect 4374 9760 4390 9824
rect 4454 9760 4470 9824
rect 4534 9760 4550 9824
rect 4614 9760 4622 9824
rect 4302 8736 4622 9760
rect 4302 8672 4310 8736
rect 4374 8672 4390 8736
rect 4454 8672 4470 8736
rect 4534 8672 4550 8736
rect 4614 8672 4622 8736
rect 4302 7648 4622 8672
rect 4302 7584 4310 7648
rect 4374 7584 4390 7648
rect 4454 7584 4470 7648
rect 4534 7584 4550 7648
rect 4614 7584 4622 7648
rect 4302 6560 4622 7584
rect 4302 6496 4310 6560
rect 4374 6496 4390 6560
rect 4454 6496 4470 6560
rect 4534 6496 4550 6560
rect 4614 6496 4622 6560
rect 4302 5472 4622 6496
rect 4302 5408 4310 5472
rect 4374 5408 4390 5472
rect 4454 5408 4470 5472
rect 4534 5408 4550 5472
rect 4614 5408 4622 5472
rect 4302 4384 4622 5408
rect 4302 4320 4310 4384
rect 4374 4320 4390 4384
rect 4454 4320 4470 4384
rect 4534 4320 4550 4384
rect 4614 4320 4622 4384
rect 4302 3296 4622 4320
rect 4302 3232 4310 3296
rect 4374 3232 4390 3296
rect 4454 3232 4470 3296
rect 4534 3232 4550 3296
rect 4614 3232 4622 3296
rect 4302 2208 4622 3232
rect 4302 2144 4310 2208
rect 4374 2144 4390 2208
rect 4454 2144 4470 2208
rect 4534 2144 4550 2208
rect 4614 2144 4622 2208
rect 3923 2004 3989 2005
rect 3923 1940 3924 2004
rect 3988 1940 3989 2004
rect 3923 1939 3989 1940
rect 2623 1600 2631 1664
rect 2695 1600 2711 1664
rect 2775 1600 2791 1664
rect 2855 1600 2871 1664
rect 2935 1600 2943 1664
rect 2623 1040 2943 1600
rect 4302 1120 4622 2144
rect 4846 1325 4906 41515
rect 5211 41444 5277 41445
rect 5211 41380 5212 41444
rect 5276 41380 5277 41444
rect 5211 41379 5277 41380
rect 5214 1325 5274 41379
rect 5981 40832 6301 41856
rect 7660 43552 7980 43568
rect 7660 43488 7668 43552
rect 7732 43488 7748 43552
rect 7812 43488 7828 43552
rect 7892 43488 7908 43552
rect 7972 43488 7980 43552
rect 7660 42464 7980 43488
rect 7660 42400 7668 42464
rect 7732 42400 7748 42464
rect 7812 42400 7828 42464
rect 7892 42400 7908 42464
rect 7972 42400 7980 42464
rect 6683 41444 6749 41445
rect 6683 41380 6684 41444
rect 6748 41380 6749 41444
rect 6683 41379 6749 41380
rect 5981 40768 5989 40832
rect 6053 40768 6069 40832
rect 6133 40768 6149 40832
rect 6213 40768 6229 40832
rect 6293 40768 6301 40832
rect 5981 39744 6301 40768
rect 5981 39680 5989 39744
rect 6053 39680 6069 39744
rect 6133 39680 6149 39744
rect 6213 39680 6229 39744
rect 6293 39680 6301 39744
rect 5981 38656 6301 39680
rect 5981 38592 5989 38656
rect 6053 38592 6069 38656
rect 6133 38592 6149 38656
rect 6213 38592 6229 38656
rect 6293 38592 6301 38656
rect 5981 37568 6301 38592
rect 5981 37504 5989 37568
rect 6053 37504 6069 37568
rect 6133 37504 6149 37568
rect 6213 37504 6229 37568
rect 6293 37504 6301 37568
rect 5981 36480 6301 37504
rect 5981 36416 5989 36480
rect 6053 36416 6069 36480
rect 6133 36416 6149 36480
rect 6213 36416 6229 36480
rect 6293 36416 6301 36480
rect 5981 35392 6301 36416
rect 5981 35328 5989 35392
rect 6053 35328 6069 35392
rect 6133 35328 6149 35392
rect 6213 35328 6229 35392
rect 6293 35328 6301 35392
rect 5981 34304 6301 35328
rect 6499 34644 6565 34645
rect 6499 34580 6500 34644
rect 6564 34580 6565 34644
rect 6499 34579 6565 34580
rect 5981 34240 5989 34304
rect 6053 34240 6069 34304
rect 6133 34240 6149 34304
rect 6213 34240 6229 34304
rect 6293 34240 6301 34304
rect 5981 33216 6301 34240
rect 5981 33152 5989 33216
rect 6053 33152 6069 33216
rect 6133 33152 6149 33216
rect 6213 33152 6229 33216
rect 6293 33152 6301 33216
rect 5981 32128 6301 33152
rect 5981 32064 5989 32128
rect 6053 32064 6069 32128
rect 6133 32064 6149 32128
rect 6213 32064 6229 32128
rect 6293 32064 6301 32128
rect 5981 31040 6301 32064
rect 5981 30976 5989 31040
rect 6053 30976 6069 31040
rect 6133 30976 6149 31040
rect 6213 30976 6229 31040
rect 6293 30976 6301 31040
rect 5981 29952 6301 30976
rect 5981 29888 5989 29952
rect 6053 29888 6069 29952
rect 6133 29888 6149 29952
rect 6213 29888 6229 29952
rect 6293 29888 6301 29952
rect 5981 28864 6301 29888
rect 5981 28800 5989 28864
rect 6053 28800 6069 28864
rect 6133 28800 6149 28864
rect 6213 28800 6229 28864
rect 6293 28800 6301 28864
rect 5981 27776 6301 28800
rect 5981 27712 5989 27776
rect 6053 27712 6069 27776
rect 6133 27712 6149 27776
rect 6213 27712 6229 27776
rect 6293 27712 6301 27776
rect 5981 26688 6301 27712
rect 5981 26624 5989 26688
rect 6053 26624 6069 26688
rect 6133 26624 6149 26688
rect 6213 26624 6229 26688
rect 6293 26624 6301 26688
rect 5981 25600 6301 26624
rect 5981 25536 5989 25600
rect 6053 25536 6069 25600
rect 6133 25536 6149 25600
rect 6213 25536 6229 25600
rect 6293 25536 6301 25600
rect 5981 24512 6301 25536
rect 5981 24448 5989 24512
rect 6053 24448 6069 24512
rect 6133 24448 6149 24512
rect 6213 24448 6229 24512
rect 6293 24448 6301 24512
rect 5981 23424 6301 24448
rect 5981 23360 5989 23424
rect 6053 23360 6069 23424
rect 6133 23360 6149 23424
rect 6213 23360 6229 23424
rect 6293 23360 6301 23424
rect 5981 22336 6301 23360
rect 5981 22272 5989 22336
rect 6053 22272 6069 22336
rect 6133 22272 6149 22336
rect 6213 22272 6229 22336
rect 6293 22272 6301 22336
rect 5981 21248 6301 22272
rect 5981 21184 5989 21248
rect 6053 21184 6069 21248
rect 6133 21184 6149 21248
rect 6213 21184 6229 21248
rect 6293 21184 6301 21248
rect 5981 20160 6301 21184
rect 5981 20096 5989 20160
rect 6053 20096 6069 20160
rect 6133 20096 6149 20160
rect 6213 20096 6229 20160
rect 6293 20096 6301 20160
rect 5981 19072 6301 20096
rect 5981 19008 5989 19072
rect 6053 19008 6069 19072
rect 6133 19008 6149 19072
rect 6213 19008 6229 19072
rect 6293 19008 6301 19072
rect 5981 17984 6301 19008
rect 5981 17920 5989 17984
rect 6053 17920 6069 17984
rect 6133 17920 6149 17984
rect 6213 17920 6229 17984
rect 6293 17920 6301 17984
rect 5981 16896 6301 17920
rect 5981 16832 5989 16896
rect 6053 16832 6069 16896
rect 6133 16832 6149 16896
rect 6213 16832 6229 16896
rect 6293 16832 6301 16896
rect 5981 15808 6301 16832
rect 5981 15744 5989 15808
rect 6053 15744 6069 15808
rect 6133 15744 6149 15808
rect 6213 15744 6229 15808
rect 6293 15744 6301 15808
rect 5981 14720 6301 15744
rect 5981 14656 5989 14720
rect 6053 14656 6069 14720
rect 6133 14656 6149 14720
rect 6213 14656 6229 14720
rect 6293 14656 6301 14720
rect 5981 13632 6301 14656
rect 5981 13568 5989 13632
rect 6053 13568 6069 13632
rect 6133 13568 6149 13632
rect 6213 13568 6229 13632
rect 6293 13568 6301 13632
rect 5981 12544 6301 13568
rect 5981 12480 5989 12544
rect 6053 12480 6069 12544
rect 6133 12480 6149 12544
rect 6213 12480 6229 12544
rect 6293 12480 6301 12544
rect 5981 11456 6301 12480
rect 5981 11392 5989 11456
rect 6053 11392 6069 11456
rect 6133 11392 6149 11456
rect 6213 11392 6229 11456
rect 6293 11392 6301 11456
rect 5981 10368 6301 11392
rect 5981 10304 5989 10368
rect 6053 10304 6069 10368
rect 6133 10304 6149 10368
rect 6213 10304 6229 10368
rect 6293 10304 6301 10368
rect 5981 9280 6301 10304
rect 5981 9216 5989 9280
rect 6053 9216 6069 9280
rect 6133 9216 6149 9280
rect 6213 9216 6229 9280
rect 6293 9216 6301 9280
rect 5981 8192 6301 9216
rect 5981 8128 5989 8192
rect 6053 8128 6069 8192
rect 6133 8128 6149 8192
rect 6213 8128 6229 8192
rect 6293 8128 6301 8192
rect 5981 7104 6301 8128
rect 5981 7040 5989 7104
rect 6053 7040 6069 7104
rect 6133 7040 6149 7104
rect 6213 7040 6229 7104
rect 6293 7040 6301 7104
rect 5981 6016 6301 7040
rect 5981 5952 5989 6016
rect 6053 5952 6069 6016
rect 6133 5952 6149 6016
rect 6213 5952 6229 6016
rect 6293 5952 6301 6016
rect 5981 4928 6301 5952
rect 5981 4864 5989 4928
rect 6053 4864 6069 4928
rect 6133 4864 6149 4928
rect 6213 4864 6229 4928
rect 6293 4864 6301 4928
rect 5981 3840 6301 4864
rect 5981 3776 5989 3840
rect 6053 3776 6069 3840
rect 6133 3776 6149 3840
rect 6213 3776 6229 3840
rect 6293 3776 6301 3840
rect 5981 2752 6301 3776
rect 5981 2688 5989 2752
rect 6053 2688 6069 2752
rect 6133 2688 6149 2752
rect 6213 2688 6229 2752
rect 6293 2688 6301 2752
rect 5981 1664 6301 2688
rect 5981 1600 5989 1664
rect 6053 1600 6069 1664
rect 6133 1600 6149 1664
rect 6213 1600 6229 1664
rect 6293 1600 6301 1664
rect 4843 1324 4909 1325
rect 4843 1260 4844 1324
rect 4908 1260 4909 1324
rect 4843 1259 4909 1260
rect 5211 1324 5277 1325
rect 5211 1260 5212 1324
rect 5276 1260 5277 1324
rect 5211 1259 5277 1260
rect 4302 1056 4310 1120
rect 4374 1056 4390 1120
rect 4454 1056 4470 1120
rect 4534 1056 4550 1120
rect 4614 1056 4622 1120
rect 4302 1040 4622 1056
rect 5981 1040 6301 1600
rect 6502 1325 6562 34579
rect 6686 2685 6746 41379
rect 7660 41376 7980 42400
rect 7660 41312 7668 41376
rect 7732 41312 7748 41376
rect 7812 41312 7828 41376
rect 7892 41312 7908 41376
rect 7972 41312 7980 41376
rect 7660 40288 7980 41312
rect 7660 40224 7668 40288
rect 7732 40224 7748 40288
rect 7812 40224 7828 40288
rect 7892 40224 7908 40288
rect 7972 40224 7980 40288
rect 7660 39200 7980 40224
rect 7660 39136 7668 39200
rect 7732 39136 7748 39200
rect 7812 39136 7828 39200
rect 7892 39136 7908 39200
rect 7972 39136 7980 39200
rect 7660 38112 7980 39136
rect 7660 38048 7668 38112
rect 7732 38048 7748 38112
rect 7812 38048 7828 38112
rect 7892 38048 7908 38112
rect 7972 38048 7980 38112
rect 7660 37024 7980 38048
rect 7660 36960 7668 37024
rect 7732 36960 7748 37024
rect 7812 36960 7828 37024
rect 7892 36960 7908 37024
rect 7972 36960 7980 37024
rect 7660 35936 7980 36960
rect 7660 35872 7668 35936
rect 7732 35872 7748 35936
rect 7812 35872 7828 35936
rect 7892 35872 7908 35936
rect 7972 35872 7980 35936
rect 7660 34848 7980 35872
rect 7660 34784 7668 34848
rect 7732 34784 7748 34848
rect 7812 34784 7828 34848
rect 7892 34784 7908 34848
rect 7972 34784 7980 34848
rect 7660 33760 7980 34784
rect 7660 33696 7668 33760
rect 7732 33696 7748 33760
rect 7812 33696 7828 33760
rect 7892 33696 7908 33760
rect 7972 33696 7980 33760
rect 7660 32672 7980 33696
rect 7660 32608 7668 32672
rect 7732 32608 7748 32672
rect 7812 32608 7828 32672
rect 7892 32608 7908 32672
rect 7972 32608 7980 32672
rect 7660 31584 7980 32608
rect 7660 31520 7668 31584
rect 7732 31520 7748 31584
rect 7812 31520 7828 31584
rect 7892 31520 7908 31584
rect 7972 31520 7980 31584
rect 7660 30496 7980 31520
rect 7660 30432 7668 30496
rect 7732 30432 7748 30496
rect 7812 30432 7828 30496
rect 7892 30432 7908 30496
rect 7972 30432 7980 30496
rect 7660 29408 7980 30432
rect 7660 29344 7668 29408
rect 7732 29344 7748 29408
rect 7812 29344 7828 29408
rect 7892 29344 7908 29408
rect 7972 29344 7980 29408
rect 7660 28320 7980 29344
rect 9339 43008 9659 43568
rect 9339 42944 9347 43008
rect 9411 42944 9427 43008
rect 9491 42944 9507 43008
rect 9571 42944 9587 43008
rect 9651 42944 9659 43008
rect 9339 41920 9659 42944
rect 9339 41856 9347 41920
rect 9411 41856 9427 41920
rect 9491 41856 9507 41920
rect 9571 41856 9587 41920
rect 9651 41856 9659 41920
rect 9339 40832 9659 41856
rect 9339 40768 9347 40832
rect 9411 40768 9427 40832
rect 9491 40768 9507 40832
rect 9571 40768 9587 40832
rect 9651 40768 9659 40832
rect 9339 39744 9659 40768
rect 9339 39680 9347 39744
rect 9411 39680 9427 39744
rect 9491 39680 9507 39744
rect 9571 39680 9587 39744
rect 9651 39680 9659 39744
rect 9339 38656 9659 39680
rect 9339 38592 9347 38656
rect 9411 38592 9427 38656
rect 9491 38592 9507 38656
rect 9571 38592 9587 38656
rect 9651 38592 9659 38656
rect 9339 37568 9659 38592
rect 9339 37504 9347 37568
rect 9411 37504 9427 37568
rect 9491 37504 9507 37568
rect 9571 37504 9587 37568
rect 9651 37504 9659 37568
rect 9339 36480 9659 37504
rect 11018 43552 11338 43568
rect 11018 43488 11026 43552
rect 11090 43488 11106 43552
rect 11170 43488 11186 43552
rect 11250 43488 11266 43552
rect 11330 43488 11338 43552
rect 11018 42464 11338 43488
rect 11018 42400 11026 42464
rect 11090 42400 11106 42464
rect 11170 42400 11186 42464
rect 11250 42400 11266 42464
rect 11330 42400 11338 42464
rect 11018 41376 11338 42400
rect 11018 41312 11026 41376
rect 11090 41312 11106 41376
rect 11170 41312 11186 41376
rect 11250 41312 11266 41376
rect 11330 41312 11338 41376
rect 11018 40288 11338 41312
rect 11018 40224 11026 40288
rect 11090 40224 11106 40288
rect 11170 40224 11186 40288
rect 11250 40224 11266 40288
rect 11330 40224 11338 40288
rect 11018 39200 11338 40224
rect 11018 39136 11026 39200
rect 11090 39136 11106 39200
rect 11170 39136 11186 39200
rect 11250 39136 11266 39200
rect 11330 39136 11338 39200
rect 11018 38112 11338 39136
rect 11018 38048 11026 38112
rect 11090 38048 11106 38112
rect 11170 38048 11186 38112
rect 11250 38048 11266 38112
rect 11330 38048 11338 38112
rect 10363 37364 10429 37365
rect 10363 37300 10364 37364
rect 10428 37300 10429 37364
rect 10363 37299 10429 37300
rect 9339 36416 9347 36480
rect 9411 36416 9427 36480
rect 9491 36416 9507 36480
rect 9571 36416 9587 36480
rect 9651 36416 9659 36480
rect 9339 35392 9659 36416
rect 9339 35328 9347 35392
rect 9411 35328 9427 35392
rect 9491 35328 9507 35392
rect 9571 35328 9587 35392
rect 9651 35328 9659 35392
rect 9339 34304 9659 35328
rect 9339 34240 9347 34304
rect 9411 34240 9427 34304
rect 9491 34240 9507 34304
rect 9571 34240 9587 34304
rect 9651 34240 9659 34304
rect 9339 33216 9659 34240
rect 10179 33964 10245 33965
rect 10179 33900 10180 33964
rect 10244 33900 10245 33964
rect 10179 33899 10245 33900
rect 9339 33152 9347 33216
rect 9411 33152 9427 33216
rect 9491 33152 9507 33216
rect 9571 33152 9587 33216
rect 9651 33152 9659 33216
rect 9339 32128 9659 33152
rect 10182 32877 10242 33899
rect 10179 32876 10245 32877
rect 10179 32812 10180 32876
rect 10244 32812 10245 32876
rect 10179 32811 10245 32812
rect 9339 32064 9347 32128
rect 9411 32064 9427 32128
rect 9491 32064 9507 32128
rect 9571 32064 9587 32128
rect 9651 32064 9659 32128
rect 9339 31040 9659 32064
rect 9339 30976 9347 31040
rect 9411 30976 9427 31040
rect 9491 30976 9507 31040
rect 9571 30976 9587 31040
rect 9651 30976 9659 31040
rect 9339 29952 9659 30976
rect 10182 30837 10242 32811
rect 10179 30836 10245 30837
rect 10179 30772 10180 30836
rect 10244 30772 10245 30836
rect 10179 30771 10245 30772
rect 9339 29888 9347 29952
rect 9411 29888 9427 29952
rect 9491 29888 9507 29952
rect 9571 29888 9587 29952
rect 9651 29888 9659 29952
rect 9075 29068 9141 29069
rect 9075 29004 9076 29068
rect 9140 29004 9141 29068
rect 9075 29003 9141 29004
rect 7660 28256 7668 28320
rect 7732 28256 7748 28320
rect 7812 28256 7828 28320
rect 7892 28256 7908 28320
rect 7972 28256 7980 28320
rect 7660 27232 7980 28256
rect 8523 28116 8589 28117
rect 8523 28052 8524 28116
rect 8588 28052 8589 28116
rect 8523 28051 8589 28052
rect 7660 27168 7668 27232
rect 7732 27168 7748 27232
rect 7812 27168 7828 27232
rect 7892 27168 7908 27232
rect 7972 27168 7980 27232
rect 7419 26348 7485 26349
rect 7419 26284 7420 26348
rect 7484 26284 7485 26348
rect 7419 26283 7485 26284
rect 7422 21861 7482 26283
rect 7660 26144 7980 27168
rect 7660 26080 7668 26144
rect 7732 26080 7748 26144
rect 7812 26080 7828 26144
rect 7892 26080 7908 26144
rect 7972 26080 7980 26144
rect 7660 25056 7980 26080
rect 7660 24992 7668 25056
rect 7732 24992 7748 25056
rect 7812 24992 7828 25056
rect 7892 24992 7908 25056
rect 7972 24992 7980 25056
rect 7660 23968 7980 24992
rect 7660 23904 7668 23968
rect 7732 23904 7748 23968
rect 7812 23904 7828 23968
rect 7892 23904 7908 23968
rect 7972 23904 7980 23968
rect 7660 22880 7980 23904
rect 8526 23629 8586 28051
rect 8891 27708 8957 27709
rect 8891 27644 8892 27708
rect 8956 27644 8957 27708
rect 8891 27643 8957 27644
rect 8155 23628 8221 23629
rect 8155 23564 8156 23628
rect 8220 23564 8221 23628
rect 8155 23563 8221 23564
rect 8523 23628 8589 23629
rect 8523 23564 8524 23628
rect 8588 23564 8589 23628
rect 8523 23563 8589 23564
rect 7660 22816 7668 22880
rect 7732 22816 7748 22880
rect 7812 22816 7828 22880
rect 7892 22816 7908 22880
rect 7972 22816 7980 22880
rect 7419 21860 7485 21861
rect 7419 21796 7420 21860
rect 7484 21796 7485 21860
rect 7419 21795 7485 21796
rect 7660 21792 7980 22816
rect 7660 21728 7668 21792
rect 7732 21728 7748 21792
rect 7812 21728 7828 21792
rect 7892 21728 7908 21792
rect 7972 21728 7980 21792
rect 7051 20772 7117 20773
rect 7051 20708 7052 20772
rect 7116 20708 7117 20772
rect 7051 20707 7117 20708
rect 7054 17645 7114 20707
rect 7660 20704 7980 21728
rect 7660 20640 7668 20704
rect 7732 20640 7748 20704
rect 7812 20640 7828 20704
rect 7892 20640 7908 20704
rect 7972 20640 7980 20704
rect 7660 19616 7980 20640
rect 7660 19552 7668 19616
rect 7732 19552 7748 19616
rect 7812 19552 7828 19616
rect 7892 19552 7908 19616
rect 7972 19552 7980 19616
rect 7419 18868 7485 18869
rect 7419 18804 7420 18868
rect 7484 18804 7485 18868
rect 7419 18803 7485 18804
rect 7235 18732 7301 18733
rect 7235 18668 7236 18732
rect 7300 18668 7301 18732
rect 7235 18667 7301 18668
rect 7051 17644 7117 17645
rect 7051 17580 7052 17644
rect 7116 17580 7117 17644
rect 7051 17579 7117 17580
rect 7238 15877 7298 18667
rect 7235 15876 7301 15877
rect 7235 15812 7236 15876
rect 7300 15812 7301 15876
rect 7235 15811 7301 15812
rect 7422 13701 7482 18803
rect 7660 18528 7980 19552
rect 8158 18733 8218 23563
rect 8707 22540 8773 22541
rect 8707 22476 8708 22540
rect 8772 22476 8773 22540
rect 8707 22475 8773 22476
rect 8155 18732 8221 18733
rect 8155 18668 8156 18732
rect 8220 18668 8221 18732
rect 8155 18667 8221 18668
rect 7660 18464 7668 18528
rect 7732 18464 7748 18528
rect 7812 18464 7828 18528
rect 7892 18464 7908 18528
rect 7972 18464 7980 18528
rect 7660 17440 7980 18464
rect 7660 17376 7668 17440
rect 7732 17376 7748 17440
rect 7812 17376 7828 17440
rect 7892 17376 7908 17440
rect 7972 17376 7980 17440
rect 7660 16352 7980 17376
rect 7660 16288 7668 16352
rect 7732 16288 7748 16352
rect 7812 16288 7828 16352
rect 7892 16288 7908 16352
rect 7972 16288 7980 16352
rect 7660 15264 7980 16288
rect 7660 15200 7668 15264
rect 7732 15200 7748 15264
rect 7812 15200 7828 15264
rect 7892 15200 7908 15264
rect 7972 15200 7980 15264
rect 7660 14176 7980 15200
rect 7660 14112 7668 14176
rect 7732 14112 7748 14176
rect 7812 14112 7828 14176
rect 7892 14112 7908 14176
rect 7972 14112 7980 14176
rect 7419 13700 7485 13701
rect 7419 13636 7420 13700
rect 7484 13636 7485 13700
rect 7419 13635 7485 13636
rect 7660 13088 7980 14112
rect 7660 13024 7668 13088
rect 7732 13024 7748 13088
rect 7812 13024 7828 13088
rect 7892 13024 7908 13088
rect 7972 13024 7980 13088
rect 7660 12000 7980 13024
rect 7660 11936 7668 12000
rect 7732 11936 7748 12000
rect 7812 11936 7828 12000
rect 7892 11936 7908 12000
rect 7972 11936 7980 12000
rect 7660 10912 7980 11936
rect 7660 10848 7668 10912
rect 7732 10848 7748 10912
rect 7812 10848 7828 10912
rect 7892 10848 7908 10912
rect 7972 10848 7980 10912
rect 7660 9824 7980 10848
rect 7660 9760 7668 9824
rect 7732 9760 7748 9824
rect 7812 9760 7828 9824
rect 7892 9760 7908 9824
rect 7972 9760 7980 9824
rect 7660 8736 7980 9760
rect 7660 8672 7668 8736
rect 7732 8672 7748 8736
rect 7812 8672 7828 8736
rect 7892 8672 7908 8736
rect 7972 8672 7980 8736
rect 7660 7648 7980 8672
rect 8155 8124 8221 8125
rect 8155 8060 8156 8124
rect 8220 8060 8221 8124
rect 8155 8059 8221 8060
rect 7660 7584 7668 7648
rect 7732 7584 7748 7648
rect 7812 7584 7828 7648
rect 7892 7584 7908 7648
rect 7972 7584 7980 7648
rect 7660 6560 7980 7584
rect 7660 6496 7668 6560
rect 7732 6496 7748 6560
rect 7812 6496 7828 6560
rect 7892 6496 7908 6560
rect 7972 6496 7980 6560
rect 7660 5472 7980 6496
rect 8158 6221 8218 8059
rect 8155 6220 8221 6221
rect 8155 6156 8156 6220
rect 8220 6156 8221 6220
rect 8155 6155 8221 6156
rect 7660 5408 7668 5472
rect 7732 5408 7748 5472
rect 7812 5408 7828 5472
rect 7892 5408 7908 5472
rect 7972 5408 7980 5472
rect 7660 4384 7980 5408
rect 7660 4320 7668 4384
rect 7732 4320 7748 4384
rect 7812 4320 7828 4384
rect 7892 4320 7908 4384
rect 7972 4320 7980 4384
rect 7660 3296 7980 4320
rect 7660 3232 7668 3296
rect 7732 3232 7748 3296
rect 7812 3232 7828 3296
rect 7892 3232 7908 3296
rect 7972 3232 7980 3296
rect 6683 2684 6749 2685
rect 6683 2620 6684 2684
rect 6748 2620 6749 2684
rect 6683 2619 6749 2620
rect 7660 2208 7980 3232
rect 7660 2144 7668 2208
rect 7732 2144 7748 2208
rect 7812 2144 7828 2208
rect 7892 2144 7908 2208
rect 7972 2144 7980 2208
rect 6499 1324 6565 1325
rect 6499 1260 6500 1324
rect 6564 1260 6565 1324
rect 6499 1259 6565 1260
rect 7660 1120 7980 2144
rect 8710 1325 8770 22475
rect 8894 19277 8954 27643
rect 9078 19413 9138 29003
rect 9339 28864 9659 29888
rect 9339 28800 9347 28864
rect 9411 28800 9427 28864
rect 9491 28800 9507 28864
rect 9571 28800 9587 28864
rect 9651 28800 9659 28864
rect 9339 27776 9659 28800
rect 9339 27712 9347 27776
rect 9411 27712 9427 27776
rect 9491 27712 9507 27776
rect 9571 27712 9587 27776
rect 9651 27712 9659 27776
rect 9339 26688 9659 27712
rect 9339 26624 9347 26688
rect 9411 26624 9427 26688
rect 9491 26624 9507 26688
rect 9571 26624 9587 26688
rect 9651 26624 9659 26688
rect 9339 25600 9659 26624
rect 10366 25941 10426 37299
rect 11018 37024 11338 38048
rect 12697 43008 13017 43568
rect 12697 42944 12705 43008
rect 12769 42944 12785 43008
rect 12849 42944 12865 43008
rect 12929 42944 12945 43008
rect 13009 42944 13017 43008
rect 12697 41920 13017 42944
rect 12697 41856 12705 41920
rect 12769 41856 12785 41920
rect 12849 41856 12865 41920
rect 12929 41856 12945 41920
rect 13009 41856 13017 41920
rect 12697 40832 13017 41856
rect 12697 40768 12705 40832
rect 12769 40768 12785 40832
rect 12849 40768 12865 40832
rect 12929 40768 12945 40832
rect 13009 40768 13017 40832
rect 12697 39744 13017 40768
rect 12697 39680 12705 39744
rect 12769 39680 12785 39744
rect 12849 39680 12865 39744
rect 12929 39680 12945 39744
rect 13009 39680 13017 39744
rect 12697 38656 13017 39680
rect 12697 38592 12705 38656
rect 12769 38592 12785 38656
rect 12849 38592 12865 38656
rect 12929 38592 12945 38656
rect 13009 38592 13017 38656
rect 12697 37568 13017 38592
rect 12697 37504 12705 37568
rect 12769 37504 12785 37568
rect 12849 37504 12865 37568
rect 12929 37504 12945 37568
rect 13009 37504 13017 37568
rect 11835 37364 11901 37365
rect 11835 37300 11836 37364
rect 11900 37300 11901 37364
rect 11835 37299 11901 37300
rect 11018 36960 11026 37024
rect 11090 36960 11106 37024
rect 11170 36960 11186 37024
rect 11250 36960 11266 37024
rect 11330 36960 11338 37024
rect 11018 35936 11338 36960
rect 11018 35872 11026 35936
rect 11090 35872 11106 35936
rect 11170 35872 11186 35936
rect 11250 35872 11266 35936
rect 11330 35872 11338 35936
rect 11018 34848 11338 35872
rect 11018 34784 11026 34848
rect 11090 34784 11106 34848
rect 11170 34784 11186 34848
rect 11250 34784 11266 34848
rect 11330 34784 11338 34848
rect 10731 33964 10797 33965
rect 10731 33900 10732 33964
rect 10796 33900 10797 33964
rect 10731 33899 10797 33900
rect 10363 25940 10429 25941
rect 10363 25876 10364 25940
rect 10428 25876 10429 25940
rect 10363 25875 10429 25876
rect 9339 25536 9347 25600
rect 9411 25536 9427 25600
rect 9491 25536 9507 25600
rect 9571 25536 9587 25600
rect 9651 25536 9659 25600
rect 9339 24512 9659 25536
rect 10734 25397 10794 33899
rect 11018 33760 11338 34784
rect 11018 33696 11026 33760
rect 11090 33696 11106 33760
rect 11170 33696 11186 33760
rect 11250 33696 11266 33760
rect 11330 33696 11338 33760
rect 11018 32672 11338 33696
rect 11018 32608 11026 32672
rect 11090 32608 11106 32672
rect 11170 32608 11186 32672
rect 11250 32608 11266 32672
rect 11330 32608 11338 32672
rect 11018 31584 11338 32608
rect 11838 31770 11898 37299
rect 12697 36480 13017 37504
rect 12697 36416 12705 36480
rect 12769 36416 12785 36480
rect 12849 36416 12865 36480
rect 12929 36416 12945 36480
rect 13009 36416 13017 36480
rect 12697 35392 13017 36416
rect 12697 35328 12705 35392
rect 12769 35328 12785 35392
rect 12849 35328 12865 35392
rect 12929 35328 12945 35392
rect 13009 35328 13017 35392
rect 12571 34644 12637 34645
rect 12571 34580 12572 34644
rect 12636 34580 12637 34644
rect 12571 34579 12637 34580
rect 12574 33013 12634 34579
rect 12697 34304 13017 35328
rect 12697 34240 12705 34304
rect 12769 34240 12785 34304
rect 12849 34240 12865 34304
rect 12929 34240 12945 34304
rect 13009 34240 13017 34304
rect 12697 33216 13017 34240
rect 12697 33152 12705 33216
rect 12769 33152 12785 33216
rect 12849 33152 12865 33216
rect 12929 33152 12945 33216
rect 13009 33152 13017 33216
rect 12571 33012 12637 33013
rect 12571 32948 12572 33012
rect 12636 32948 12637 33012
rect 12571 32947 12637 32948
rect 11018 31520 11026 31584
rect 11090 31520 11106 31584
rect 11170 31520 11186 31584
rect 11250 31520 11266 31584
rect 11330 31520 11338 31584
rect 11018 30496 11338 31520
rect 11018 30432 11026 30496
rect 11090 30432 11106 30496
rect 11170 30432 11186 30496
rect 11250 30432 11266 30496
rect 11330 30432 11338 30496
rect 11018 29408 11338 30432
rect 11018 29344 11026 29408
rect 11090 29344 11106 29408
rect 11170 29344 11186 29408
rect 11250 29344 11266 29408
rect 11330 29344 11338 29408
rect 11018 28320 11338 29344
rect 11470 31710 11898 31770
rect 12697 32128 13017 33152
rect 12697 32064 12705 32128
rect 12769 32064 12785 32128
rect 12849 32064 12865 32128
rect 12929 32064 12945 32128
rect 13009 32064 13017 32128
rect 11470 29205 11530 31710
rect 12697 31040 13017 32064
rect 14376 43552 14696 43568
rect 14376 43488 14384 43552
rect 14448 43488 14464 43552
rect 14528 43488 14544 43552
rect 14608 43488 14624 43552
rect 14688 43488 14696 43552
rect 14376 42464 14696 43488
rect 14376 42400 14384 42464
rect 14448 42400 14464 42464
rect 14528 42400 14544 42464
rect 14608 42400 14624 42464
rect 14688 42400 14696 42464
rect 14376 41376 14696 42400
rect 14963 41580 15029 41581
rect 14963 41516 14964 41580
rect 15028 41516 15029 41580
rect 14963 41515 15029 41516
rect 14376 41312 14384 41376
rect 14448 41312 14464 41376
rect 14528 41312 14544 41376
rect 14608 41312 14624 41376
rect 14688 41312 14696 41376
rect 14376 40288 14696 41312
rect 14376 40224 14384 40288
rect 14448 40224 14464 40288
rect 14528 40224 14544 40288
rect 14608 40224 14624 40288
rect 14688 40224 14696 40288
rect 14376 39200 14696 40224
rect 14376 39136 14384 39200
rect 14448 39136 14464 39200
rect 14528 39136 14544 39200
rect 14608 39136 14624 39200
rect 14688 39136 14696 39200
rect 14376 38112 14696 39136
rect 14376 38048 14384 38112
rect 14448 38048 14464 38112
rect 14528 38048 14544 38112
rect 14608 38048 14624 38112
rect 14688 38048 14696 38112
rect 14376 37024 14696 38048
rect 14376 36960 14384 37024
rect 14448 36960 14464 37024
rect 14528 36960 14544 37024
rect 14608 36960 14624 37024
rect 14688 36960 14696 37024
rect 14376 35936 14696 36960
rect 14376 35872 14384 35936
rect 14448 35872 14464 35936
rect 14528 35872 14544 35936
rect 14608 35872 14624 35936
rect 14688 35872 14696 35936
rect 14376 34848 14696 35872
rect 14376 34784 14384 34848
rect 14448 34784 14464 34848
rect 14528 34784 14544 34848
rect 14608 34784 14624 34848
rect 14688 34784 14696 34848
rect 14376 33760 14696 34784
rect 14376 33696 14384 33760
rect 14448 33696 14464 33760
rect 14528 33696 14544 33760
rect 14608 33696 14624 33760
rect 14688 33696 14696 33760
rect 14376 32672 14696 33696
rect 14376 32608 14384 32672
rect 14448 32608 14464 32672
rect 14528 32608 14544 32672
rect 14608 32608 14624 32672
rect 14688 32608 14696 32672
rect 14227 32060 14293 32061
rect 14227 31996 14228 32060
rect 14292 31996 14293 32060
rect 14227 31995 14293 31996
rect 14230 31381 14290 31995
rect 14376 31584 14696 32608
rect 14376 31520 14384 31584
rect 14448 31520 14464 31584
rect 14528 31520 14544 31584
rect 14608 31520 14624 31584
rect 14688 31520 14696 31584
rect 14227 31380 14293 31381
rect 14227 31316 14228 31380
rect 14292 31316 14293 31380
rect 14227 31315 14293 31316
rect 12697 30976 12705 31040
rect 12769 30976 12785 31040
rect 12849 30976 12865 31040
rect 12929 30976 12945 31040
rect 13009 30976 13017 31040
rect 11835 30428 11901 30429
rect 11835 30364 11836 30428
rect 11900 30364 11901 30428
rect 11835 30363 11901 30364
rect 11467 29204 11533 29205
rect 11467 29140 11468 29204
rect 11532 29140 11533 29204
rect 11467 29139 11533 29140
rect 11018 28256 11026 28320
rect 11090 28256 11106 28320
rect 11170 28256 11186 28320
rect 11250 28256 11266 28320
rect 11330 28256 11338 28320
rect 11018 27232 11338 28256
rect 11018 27168 11026 27232
rect 11090 27168 11106 27232
rect 11170 27168 11186 27232
rect 11250 27168 11266 27232
rect 11330 27168 11338 27232
rect 11018 26144 11338 27168
rect 11838 26757 11898 30363
rect 12697 29952 13017 30976
rect 13491 30700 13557 30701
rect 13491 30636 13492 30700
rect 13556 30636 13557 30700
rect 13491 30635 13557 30636
rect 12697 29888 12705 29952
rect 12769 29888 12785 29952
rect 12849 29888 12865 29952
rect 12929 29888 12945 29952
rect 13009 29888 13017 29952
rect 12387 28932 12453 28933
rect 12387 28868 12388 28932
rect 12452 28868 12453 28932
rect 12387 28867 12453 28868
rect 12019 28796 12085 28797
rect 12019 28732 12020 28796
rect 12084 28732 12085 28796
rect 12019 28731 12085 28732
rect 12022 27845 12082 28731
rect 12019 27844 12085 27845
rect 12019 27780 12020 27844
rect 12084 27780 12085 27844
rect 12019 27779 12085 27780
rect 12019 27708 12085 27709
rect 12019 27644 12020 27708
rect 12084 27644 12085 27708
rect 12019 27643 12085 27644
rect 11835 26756 11901 26757
rect 11835 26692 11836 26756
rect 11900 26692 11901 26756
rect 11835 26691 11901 26692
rect 11018 26080 11026 26144
rect 11090 26080 11106 26144
rect 11170 26080 11186 26144
rect 11250 26080 11266 26144
rect 11330 26080 11338 26144
rect 10731 25396 10797 25397
rect 10731 25332 10732 25396
rect 10796 25332 10797 25396
rect 10731 25331 10797 25332
rect 9339 24448 9347 24512
rect 9411 24448 9427 24512
rect 9491 24448 9507 24512
rect 9571 24448 9587 24512
rect 9651 24448 9659 24512
rect 9339 23424 9659 24448
rect 11018 25056 11338 26080
rect 11018 24992 11026 25056
rect 11090 24992 11106 25056
rect 11170 24992 11186 25056
rect 11250 24992 11266 25056
rect 11330 24992 11338 25056
rect 10731 24172 10797 24173
rect 10731 24108 10732 24172
rect 10796 24108 10797 24172
rect 10731 24107 10797 24108
rect 9339 23360 9347 23424
rect 9411 23360 9427 23424
rect 9491 23360 9507 23424
rect 9571 23360 9587 23424
rect 9651 23360 9659 23424
rect 9339 22336 9659 23360
rect 9811 22540 9877 22541
rect 9811 22476 9812 22540
rect 9876 22476 9877 22540
rect 9811 22475 9877 22476
rect 9339 22272 9347 22336
rect 9411 22272 9427 22336
rect 9491 22272 9507 22336
rect 9571 22272 9587 22336
rect 9651 22272 9659 22336
rect 9339 21248 9659 22272
rect 9339 21184 9347 21248
rect 9411 21184 9427 21248
rect 9491 21184 9507 21248
rect 9571 21184 9587 21248
rect 9651 21184 9659 21248
rect 9339 20160 9659 21184
rect 9814 20909 9874 22475
rect 9811 20908 9877 20909
rect 9811 20844 9812 20908
rect 9876 20844 9877 20908
rect 9811 20843 9877 20844
rect 9339 20096 9347 20160
rect 9411 20096 9427 20160
rect 9491 20096 9507 20160
rect 9571 20096 9587 20160
rect 9651 20096 9659 20160
rect 9075 19412 9141 19413
rect 9075 19348 9076 19412
rect 9140 19348 9141 19412
rect 9075 19347 9141 19348
rect 8891 19276 8957 19277
rect 8891 19212 8892 19276
rect 8956 19212 8957 19276
rect 8891 19211 8957 19212
rect 8894 13429 8954 19211
rect 9339 19072 9659 20096
rect 9339 19008 9347 19072
rect 9411 19008 9427 19072
rect 9491 19008 9507 19072
rect 9571 19008 9587 19072
rect 9651 19008 9659 19072
rect 9075 18324 9141 18325
rect 9075 18260 9076 18324
rect 9140 18260 9141 18324
rect 9075 18259 9141 18260
rect 8891 13428 8957 13429
rect 8891 13364 8892 13428
rect 8956 13364 8957 13428
rect 8891 13363 8957 13364
rect 8891 8804 8957 8805
rect 8891 8740 8892 8804
rect 8956 8740 8957 8804
rect 8891 8739 8957 8740
rect 8894 7717 8954 8739
rect 8891 7716 8957 7717
rect 8891 7652 8892 7716
rect 8956 7652 8957 7716
rect 8891 7651 8957 7652
rect 9078 2549 9138 18259
rect 9339 17984 9659 19008
rect 9339 17920 9347 17984
rect 9411 17920 9427 17984
rect 9491 17920 9507 17984
rect 9571 17920 9587 17984
rect 9651 17920 9659 17984
rect 9339 16896 9659 17920
rect 9814 17917 9874 20843
rect 9995 19412 10061 19413
rect 9995 19348 9996 19412
rect 10060 19348 10061 19412
rect 9995 19347 10061 19348
rect 9811 17916 9877 17917
rect 9811 17852 9812 17916
rect 9876 17852 9877 17916
rect 9811 17851 9877 17852
rect 9339 16832 9347 16896
rect 9411 16832 9427 16896
rect 9491 16832 9507 16896
rect 9571 16832 9587 16896
rect 9651 16832 9659 16896
rect 9339 15808 9659 16832
rect 9339 15744 9347 15808
rect 9411 15744 9427 15808
rect 9491 15744 9507 15808
rect 9571 15744 9587 15808
rect 9651 15744 9659 15808
rect 9339 14720 9659 15744
rect 9998 15469 10058 19347
rect 10363 17100 10429 17101
rect 10363 17036 10364 17100
rect 10428 17036 10429 17100
rect 10363 17035 10429 17036
rect 9995 15468 10061 15469
rect 9995 15404 9996 15468
rect 10060 15404 10061 15468
rect 9995 15403 10061 15404
rect 9339 14656 9347 14720
rect 9411 14656 9427 14720
rect 9491 14656 9507 14720
rect 9571 14656 9587 14720
rect 9651 14656 9659 14720
rect 9339 13632 9659 14656
rect 10179 14652 10245 14653
rect 10179 14588 10180 14652
rect 10244 14588 10245 14652
rect 10179 14587 10245 14588
rect 9339 13568 9347 13632
rect 9411 13568 9427 13632
rect 9491 13568 9507 13632
rect 9571 13568 9587 13632
rect 9651 13568 9659 13632
rect 9339 12544 9659 13568
rect 9339 12480 9347 12544
rect 9411 12480 9427 12544
rect 9491 12480 9507 12544
rect 9571 12480 9587 12544
rect 9651 12480 9659 12544
rect 9339 11456 9659 12480
rect 9339 11392 9347 11456
rect 9411 11392 9427 11456
rect 9491 11392 9507 11456
rect 9571 11392 9587 11456
rect 9651 11392 9659 11456
rect 9339 10368 9659 11392
rect 9339 10304 9347 10368
rect 9411 10304 9427 10368
rect 9491 10304 9507 10368
rect 9571 10304 9587 10368
rect 9651 10304 9659 10368
rect 9339 9280 9659 10304
rect 10182 9349 10242 14587
rect 10179 9348 10245 9349
rect 10179 9284 10180 9348
rect 10244 9284 10245 9348
rect 10179 9283 10245 9284
rect 9339 9216 9347 9280
rect 9411 9216 9427 9280
rect 9491 9216 9507 9280
rect 9571 9216 9587 9280
rect 9651 9216 9659 9280
rect 9339 8192 9659 9216
rect 9811 8668 9877 8669
rect 9811 8604 9812 8668
rect 9876 8604 9877 8668
rect 9811 8603 9877 8604
rect 9339 8128 9347 8192
rect 9411 8128 9427 8192
rect 9491 8128 9507 8192
rect 9571 8128 9587 8192
rect 9651 8128 9659 8192
rect 9339 7104 9659 8128
rect 9339 7040 9347 7104
rect 9411 7040 9427 7104
rect 9491 7040 9507 7104
rect 9571 7040 9587 7104
rect 9651 7040 9659 7104
rect 9339 6016 9659 7040
rect 9814 6765 9874 8603
rect 9811 6764 9877 6765
rect 9811 6700 9812 6764
rect 9876 6700 9877 6764
rect 9811 6699 9877 6700
rect 9339 5952 9347 6016
rect 9411 5952 9427 6016
rect 9491 5952 9507 6016
rect 9571 5952 9587 6016
rect 9651 5952 9659 6016
rect 9339 4928 9659 5952
rect 9339 4864 9347 4928
rect 9411 4864 9427 4928
rect 9491 4864 9507 4928
rect 9571 4864 9587 4928
rect 9651 4864 9659 4928
rect 9339 3840 9659 4864
rect 9339 3776 9347 3840
rect 9411 3776 9427 3840
rect 9491 3776 9507 3840
rect 9571 3776 9587 3840
rect 9651 3776 9659 3840
rect 9339 2752 9659 3776
rect 9339 2688 9347 2752
rect 9411 2688 9427 2752
rect 9491 2688 9507 2752
rect 9571 2688 9587 2752
rect 9651 2688 9659 2752
rect 9075 2548 9141 2549
rect 9075 2484 9076 2548
rect 9140 2484 9141 2548
rect 9075 2483 9141 2484
rect 9339 1664 9659 2688
rect 10366 2685 10426 17035
rect 10734 16557 10794 24107
rect 11018 23968 11338 24992
rect 11018 23904 11026 23968
rect 11090 23904 11106 23968
rect 11170 23904 11186 23968
rect 11250 23904 11266 23968
rect 11330 23904 11338 23968
rect 11018 22880 11338 23904
rect 11018 22816 11026 22880
rect 11090 22816 11106 22880
rect 11170 22816 11186 22880
rect 11250 22816 11266 22880
rect 11330 22816 11338 22880
rect 11018 21792 11338 22816
rect 11018 21728 11026 21792
rect 11090 21728 11106 21792
rect 11170 21728 11186 21792
rect 11250 21728 11266 21792
rect 11330 21728 11338 21792
rect 11018 20704 11338 21728
rect 11018 20640 11026 20704
rect 11090 20640 11106 20704
rect 11170 20640 11186 20704
rect 11250 20640 11266 20704
rect 11330 20640 11338 20704
rect 11018 19616 11338 20640
rect 11018 19552 11026 19616
rect 11090 19552 11106 19616
rect 11170 19552 11186 19616
rect 11250 19552 11266 19616
rect 11330 19552 11338 19616
rect 11018 18528 11338 19552
rect 11018 18464 11026 18528
rect 11090 18464 11106 18528
rect 11170 18464 11186 18528
rect 11250 18464 11266 18528
rect 11330 18464 11338 18528
rect 11018 17440 11338 18464
rect 11467 18324 11533 18325
rect 11467 18260 11468 18324
rect 11532 18260 11533 18324
rect 11467 18259 11533 18260
rect 11018 17376 11026 17440
rect 11090 17376 11106 17440
rect 11170 17376 11186 17440
rect 11250 17376 11266 17440
rect 11330 17376 11338 17440
rect 10731 16556 10797 16557
rect 10731 16492 10732 16556
rect 10796 16492 10797 16556
rect 10731 16491 10797 16492
rect 11018 16352 11338 17376
rect 11018 16288 11026 16352
rect 11090 16288 11106 16352
rect 11170 16288 11186 16352
rect 11250 16288 11266 16352
rect 11330 16288 11338 16352
rect 10731 15604 10797 15605
rect 10731 15540 10732 15604
rect 10796 15540 10797 15604
rect 10731 15539 10797 15540
rect 10734 9485 10794 15539
rect 11018 15264 11338 16288
rect 11470 15605 11530 18259
rect 11467 15604 11533 15605
rect 11467 15540 11468 15604
rect 11532 15540 11533 15604
rect 11467 15539 11533 15540
rect 11018 15200 11026 15264
rect 11090 15200 11106 15264
rect 11170 15200 11186 15264
rect 11250 15200 11266 15264
rect 11330 15200 11338 15264
rect 11018 14176 11338 15200
rect 11018 14112 11026 14176
rect 11090 14112 11106 14176
rect 11170 14112 11186 14176
rect 11250 14112 11266 14176
rect 11330 14112 11338 14176
rect 11018 13088 11338 14112
rect 12022 13970 12082 27643
rect 12390 25941 12450 28867
rect 12697 28864 13017 29888
rect 12697 28800 12705 28864
rect 12769 28800 12785 28864
rect 12849 28800 12865 28864
rect 12929 28800 12945 28864
rect 13009 28800 13017 28864
rect 12697 27776 13017 28800
rect 12697 27712 12705 27776
rect 12769 27712 12785 27776
rect 12849 27712 12865 27776
rect 12929 27712 12945 27776
rect 13009 27712 13017 27776
rect 12571 27164 12637 27165
rect 12571 27100 12572 27164
rect 12636 27100 12637 27164
rect 12571 27099 12637 27100
rect 12387 25940 12453 25941
rect 12387 25876 12388 25940
rect 12452 25876 12453 25940
rect 12387 25875 12453 25876
rect 12574 22110 12634 27099
rect 12390 22050 12634 22110
rect 12697 26688 13017 27712
rect 12697 26624 12705 26688
rect 12769 26624 12785 26688
rect 12849 26624 12865 26688
rect 12929 26624 12945 26688
rect 13009 26624 13017 26688
rect 12697 25600 13017 26624
rect 12697 25536 12705 25600
rect 12769 25536 12785 25600
rect 12849 25536 12865 25600
rect 12929 25536 12945 25600
rect 13009 25536 13017 25600
rect 12697 24512 13017 25536
rect 12697 24448 12705 24512
rect 12769 24448 12785 24512
rect 12849 24448 12865 24512
rect 12929 24448 12945 24512
rect 13009 24448 13017 24512
rect 12697 23424 13017 24448
rect 12697 23360 12705 23424
rect 12769 23360 12785 23424
rect 12849 23360 12865 23424
rect 12929 23360 12945 23424
rect 13009 23360 13017 23424
rect 12697 22336 13017 23360
rect 12697 22272 12705 22336
rect 12769 22272 12785 22336
rect 12849 22272 12865 22336
rect 12929 22272 12945 22336
rect 13009 22272 13017 22336
rect 12390 21450 12450 22050
rect 12206 21390 12450 21450
rect 12206 20637 12266 21390
rect 12697 21248 13017 22272
rect 12697 21184 12705 21248
rect 12769 21184 12785 21248
rect 12849 21184 12865 21248
rect 12929 21184 12945 21248
rect 13009 21184 13017 21248
rect 12203 20636 12269 20637
rect 12203 20572 12204 20636
rect 12268 20572 12269 20636
rect 12203 20571 12269 20572
rect 12697 20160 13017 21184
rect 12697 20096 12705 20160
rect 12769 20096 12785 20160
rect 12849 20096 12865 20160
rect 12929 20096 12945 20160
rect 13009 20096 13017 20160
rect 12697 19072 13017 20096
rect 12697 19008 12705 19072
rect 12769 19008 12785 19072
rect 12849 19008 12865 19072
rect 12929 19008 12945 19072
rect 13009 19008 13017 19072
rect 12387 18324 12453 18325
rect 12387 18260 12388 18324
rect 12452 18260 12453 18324
rect 12387 18259 12453 18260
rect 12390 18050 12450 18259
rect 12390 17990 12634 18050
rect 12203 13972 12269 13973
rect 12203 13970 12204 13972
rect 12022 13910 12204 13970
rect 12203 13908 12204 13910
rect 12268 13908 12269 13972
rect 12203 13907 12269 13908
rect 11467 13292 11533 13293
rect 11467 13228 11468 13292
rect 11532 13228 11533 13292
rect 11467 13227 11533 13228
rect 11018 13024 11026 13088
rect 11090 13024 11106 13088
rect 11170 13024 11186 13088
rect 11250 13024 11266 13088
rect 11330 13024 11338 13088
rect 11018 12000 11338 13024
rect 11018 11936 11026 12000
rect 11090 11936 11106 12000
rect 11170 11936 11186 12000
rect 11250 11936 11266 12000
rect 11330 11936 11338 12000
rect 11018 10912 11338 11936
rect 11018 10848 11026 10912
rect 11090 10848 11106 10912
rect 11170 10848 11186 10912
rect 11250 10848 11266 10912
rect 11330 10848 11338 10912
rect 11018 9824 11338 10848
rect 11470 10709 11530 13227
rect 11467 10708 11533 10709
rect 11467 10644 11468 10708
rect 11532 10644 11533 10708
rect 11467 10643 11533 10644
rect 12574 10573 12634 17990
rect 12697 17984 13017 19008
rect 13307 18460 13373 18461
rect 13307 18396 13308 18460
rect 13372 18396 13373 18460
rect 13307 18395 13373 18396
rect 12697 17920 12705 17984
rect 12769 17920 12785 17984
rect 12849 17920 12865 17984
rect 12929 17920 12945 17984
rect 13009 17920 13017 17984
rect 12697 16896 13017 17920
rect 12697 16832 12705 16896
rect 12769 16832 12785 16896
rect 12849 16832 12865 16896
rect 12929 16832 12945 16896
rect 13009 16832 13017 16896
rect 12697 15808 13017 16832
rect 12697 15744 12705 15808
rect 12769 15744 12785 15808
rect 12849 15744 12865 15808
rect 12929 15744 12945 15808
rect 13009 15744 13017 15808
rect 12697 14720 13017 15744
rect 13123 15060 13189 15061
rect 13123 14996 13124 15060
rect 13188 14996 13189 15060
rect 13123 14995 13189 14996
rect 12697 14656 12705 14720
rect 12769 14656 12785 14720
rect 12849 14656 12865 14720
rect 12929 14656 12945 14720
rect 13009 14656 13017 14720
rect 12697 13632 13017 14656
rect 12697 13568 12705 13632
rect 12769 13568 12785 13632
rect 12849 13568 12865 13632
rect 12929 13568 12945 13632
rect 13009 13568 13017 13632
rect 12697 12544 13017 13568
rect 12697 12480 12705 12544
rect 12769 12480 12785 12544
rect 12849 12480 12865 12544
rect 12929 12480 12945 12544
rect 13009 12480 13017 12544
rect 12697 11456 13017 12480
rect 12697 11392 12705 11456
rect 12769 11392 12785 11456
rect 12849 11392 12865 11456
rect 12929 11392 12945 11456
rect 13009 11392 13017 11456
rect 12571 10572 12637 10573
rect 12571 10508 12572 10572
rect 12636 10508 12637 10572
rect 12571 10507 12637 10508
rect 11018 9760 11026 9824
rect 11090 9760 11106 9824
rect 11170 9760 11186 9824
rect 11250 9760 11266 9824
rect 11330 9760 11338 9824
rect 10731 9484 10797 9485
rect 10731 9420 10732 9484
rect 10796 9420 10797 9484
rect 10731 9419 10797 9420
rect 11018 8736 11338 9760
rect 11018 8672 11026 8736
rect 11090 8672 11106 8736
rect 11170 8672 11186 8736
rect 11250 8672 11266 8736
rect 11330 8672 11338 8736
rect 11018 7648 11338 8672
rect 11018 7584 11026 7648
rect 11090 7584 11106 7648
rect 11170 7584 11186 7648
rect 11250 7584 11266 7648
rect 11330 7584 11338 7648
rect 11018 6560 11338 7584
rect 11018 6496 11026 6560
rect 11090 6496 11106 6560
rect 11170 6496 11186 6560
rect 11250 6496 11266 6560
rect 11330 6496 11338 6560
rect 11018 5472 11338 6496
rect 11018 5408 11026 5472
rect 11090 5408 11106 5472
rect 11170 5408 11186 5472
rect 11250 5408 11266 5472
rect 11330 5408 11338 5472
rect 11018 4384 11338 5408
rect 11018 4320 11026 4384
rect 11090 4320 11106 4384
rect 11170 4320 11186 4384
rect 11250 4320 11266 4384
rect 11330 4320 11338 4384
rect 11018 3296 11338 4320
rect 11018 3232 11026 3296
rect 11090 3232 11106 3296
rect 11170 3232 11186 3296
rect 11250 3232 11266 3296
rect 11330 3232 11338 3296
rect 10363 2684 10429 2685
rect 10363 2620 10364 2684
rect 10428 2620 10429 2684
rect 10363 2619 10429 2620
rect 9339 1600 9347 1664
rect 9411 1600 9427 1664
rect 9491 1600 9507 1664
rect 9571 1600 9587 1664
rect 9651 1600 9659 1664
rect 8707 1324 8773 1325
rect 8707 1260 8708 1324
rect 8772 1260 8773 1324
rect 8707 1259 8773 1260
rect 7660 1056 7668 1120
rect 7732 1056 7748 1120
rect 7812 1056 7828 1120
rect 7892 1056 7908 1120
rect 7972 1056 7980 1120
rect 7660 1040 7980 1056
rect 9339 1040 9659 1600
rect 11018 2208 11338 3232
rect 11018 2144 11026 2208
rect 11090 2144 11106 2208
rect 11170 2144 11186 2208
rect 11250 2144 11266 2208
rect 11330 2144 11338 2208
rect 11018 1120 11338 2144
rect 11018 1056 11026 1120
rect 11090 1056 11106 1120
rect 11170 1056 11186 1120
rect 11250 1056 11266 1120
rect 11330 1056 11338 1120
rect 11018 1040 11338 1056
rect 12697 10368 13017 11392
rect 12697 10304 12705 10368
rect 12769 10304 12785 10368
rect 12849 10304 12865 10368
rect 12929 10304 12945 10368
rect 13009 10304 13017 10368
rect 12697 9280 13017 10304
rect 13126 9757 13186 14995
rect 13310 14517 13370 18395
rect 13494 18325 13554 30635
rect 14376 30496 14696 31520
rect 14376 30432 14384 30496
rect 14448 30432 14464 30496
rect 14528 30432 14544 30496
rect 14608 30432 14624 30496
rect 14688 30432 14696 30496
rect 14376 29408 14696 30432
rect 14376 29344 14384 29408
rect 14448 29344 14464 29408
rect 14528 29344 14544 29408
rect 14608 29344 14624 29408
rect 14688 29344 14696 29408
rect 14376 28320 14696 29344
rect 14376 28256 14384 28320
rect 14448 28256 14464 28320
rect 14528 28256 14544 28320
rect 14608 28256 14624 28320
rect 14688 28256 14696 28320
rect 14043 28252 14109 28253
rect 14043 28188 14044 28252
rect 14108 28188 14109 28252
rect 14043 28187 14109 28188
rect 13675 24988 13741 24989
rect 13675 24924 13676 24988
rect 13740 24924 13741 24988
rect 13675 24923 13741 24924
rect 13678 19277 13738 24923
rect 13859 20772 13925 20773
rect 13859 20708 13860 20772
rect 13924 20708 13925 20772
rect 13859 20707 13925 20708
rect 13675 19276 13741 19277
rect 13675 19212 13676 19276
rect 13740 19212 13741 19276
rect 13675 19211 13741 19212
rect 13491 18324 13557 18325
rect 13491 18260 13492 18324
rect 13556 18260 13557 18324
rect 13491 18259 13557 18260
rect 13494 16557 13554 18259
rect 13491 16556 13557 16557
rect 13491 16492 13492 16556
rect 13556 16492 13557 16556
rect 13491 16491 13557 16492
rect 13307 14516 13373 14517
rect 13307 14452 13308 14516
rect 13372 14452 13373 14516
rect 13307 14451 13373 14452
rect 13862 14381 13922 20707
rect 14046 17645 14106 28187
rect 14227 27708 14293 27709
rect 14227 27644 14228 27708
rect 14292 27644 14293 27708
rect 14227 27643 14293 27644
rect 14043 17644 14109 17645
rect 14043 17580 14044 17644
rect 14108 17580 14109 17644
rect 14043 17579 14109 17580
rect 14230 17373 14290 27643
rect 14376 27232 14696 28256
rect 14376 27168 14384 27232
rect 14448 27168 14464 27232
rect 14528 27168 14544 27232
rect 14608 27168 14624 27232
rect 14688 27168 14696 27232
rect 14376 26144 14696 27168
rect 14376 26080 14384 26144
rect 14448 26080 14464 26144
rect 14528 26080 14544 26144
rect 14608 26080 14624 26144
rect 14688 26080 14696 26144
rect 14376 25056 14696 26080
rect 14376 24992 14384 25056
rect 14448 24992 14464 25056
rect 14528 24992 14544 25056
rect 14608 24992 14624 25056
rect 14688 24992 14696 25056
rect 14376 23968 14696 24992
rect 14376 23904 14384 23968
rect 14448 23904 14464 23968
rect 14528 23904 14544 23968
rect 14608 23904 14624 23968
rect 14688 23904 14696 23968
rect 14376 22880 14696 23904
rect 14376 22816 14384 22880
rect 14448 22816 14464 22880
rect 14528 22816 14544 22880
rect 14608 22816 14624 22880
rect 14688 22816 14696 22880
rect 14376 21792 14696 22816
rect 14376 21728 14384 21792
rect 14448 21728 14464 21792
rect 14528 21728 14544 21792
rect 14608 21728 14624 21792
rect 14688 21728 14696 21792
rect 14376 20704 14696 21728
rect 14376 20640 14384 20704
rect 14448 20640 14464 20704
rect 14528 20640 14544 20704
rect 14608 20640 14624 20704
rect 14688 20640 14696 20704
rect 14376 19616 14696 20640
rect 14376 19552 14384 19616
rect 14448 19552 14464 19616
rect 14528 19552 14544 19616
rect 14608 19552 14624 19616
rect 14688 19552 14696 19616
rect 14376 18528 14696 19552
rect 14376 18464 14384 18528
rect 14448 18464 14464 18528
rect 14528 18464 14544 18528
rect 14608 18464 14624 18528
rect 14688 18464 14696 18528
rect 14376 17440 14696 18464
rect 14376 17376 14384 17440
rect 14448 17376 14464 17440
rect 14528 17376 14544 17440
rect 14608 17376 14624 17440
rect 14688 17376 14696 17440
rect 14227 17372 14293 17373
rect 14227 17308 14228 17372
rect 14292 17308 14293 17372
rect 14227 17307 14293 17308
rect 14230 14653 14290 17307
rect 14376 16352 14696 17376
rect 14376 16288 14384 16352
rect 14448 16288 14464 16352
rect 14528 16288 14544 16352
rect 14608 16288 14624 16352
rect 14688 16288 14696 16352
rect 14376 15264 14696 16288
rect 14376 15200 14384 15264
rect 14448 15200 14464 15264
rect 14528 15200 14544 15264
rect 14608 15200 14624 15264
rect 14688 15200 14696 15264
rect 14227 14652 14293 14653
rect 14227 14588 14228 14652
rect 14292 14588 14293 14652
rect 14227 14587 14293 14588
rect 13859 14380 13925 14381
rect 13859 14316 13860 14380
rect 13924 14316 13925 14380
rect 13859 14315 13925 14316
rect 14376 14176 14696 15200
rect 14376 14112 14384 14176
rect 14448 14112 14464 14176
rect 14528 14112 14544 14176
rect 14608 14112 14624 14176
rect 14688 14112 14696 14176
rect 14376 13088 14696 14112
rect 14376 13024 14384 13088
rect 14448 13024 14464 13088
rect 14528 13024 14544 13088
rect 14608 13024 14624 13088
rect 14688 13024 14696 13088
rect 14376 12000 14696 13024
rect 14376 11936 14384 12000
rect 14448 11936 14464 12000
rect 14528 11936 14544 12000
rect 14608 11936 14624 12000
rect 14688 11936 14696 12000
rect 14376 10912 14696 11936
rect 14376 10848 14384 10912
rect 14448 10848 14464 10912
rect 14528 10848 14544 10912
rect 14608 10848 14624 10912
rect 14688 10848 14696 10912
rect 14376 9824 14696 10848
rect 14376 9760 14384 9824
rect 14448 9760 14464 9824
rect 14528 9760 14544 9824
rect 14608 9760 14624 9824
rect 14688 9760 14696 9824
rect 13123 9756 13189 9757
rect 13123 9692 13124 9756
rect 13188 9692 13189 9756
rect 13123 9691 13189 9692
rect 12697 9216 12705 9280
rect 12769 9216 12785 9280
rect 12849 9216 12865 9280
rect 12929 9216 12945 9280
rect 13009 9216 13017 9280
rect 12697 8192 13017 9216
rect 12697 8128 12705 8192
rect 12769 8128 12785 8192
rect 12849 8128 12865 8192
rect 12929 8128 12945 8192
rect 13009 8128 13017 8192
rect 12697 7104 13017 8128
rect 12697 7040 12705 7104
rect 12769 7040 12785 7104
rect 12849 7040 12865 7104
rect 12929 7040 12945 7104
rect 13009 7040 13017 7104
rect 12697 6016 13017 7040
rect 12697 5952 12705 6016
rect 12769 5952 12785 6016
rect 12849 5952 12865 6016
rect 12929 5952 12945 6016
rect 13009 5952 13017 6016
rect 12697 4928 13017 5952
rect 12697 4864 12705 4928
rect 12769 4864 12785 4928
rect 12849 4864 12865 4928
rect 12929 4864 12945 4928
rect 13009 4864 13017 4928
rect 12697 3840 13017 4864
rect 12697 3776 12705 3840
rect 12769 3776 12785 3840
rect 12849 3776 12865 3840
rect 12929 3776 12945 3840
rect 13009 3776 13017 3840
rect 12697 2752 13017 3776
rect 12697 2688 12705 2752
rect 12769 2688 12785 2752
rect 12849 2688 12865 2752
rect 12929 2688 12945 2752
rect 13009 2688 13017 2752
rect 12697 1664 13017 2688
rect 12697 1600 12705 1664
rect 12769 1600 12785 1664
rect 12849 1600 12865 1664
rect 12929 1600 12945 1664
rect 13009 1600 13017 1664
rect 12697 1040 13017 1600
rect 14376 8736 14696 9760
rect 14376 8672 14384 8736
rect 14448 8672 14464 8736
rect 14528 8672 14544 8736
rect 14608 8672 14624 8736
rect 14688 8672 14696 8736
rect 14376 7648 14696 8672
rect 14376 7584 14384 7648
rect 14448 7584 14464 7648
rect 14528 7584 14544 7648
rect 14608 7584 14624 7648
rect 14688 7584 14696 7648
rect 14376 6560 14696 7584
rect 14376 6496 14384 6560
rect 14448 6496 14464 6560
rect 14528 6496 14544 6560
rect 14608 6496 14624 6560
rect 14688 6496 14696 6560
rect 14376 5472 14696 6496
rect 14966 5677 15026 41515
rect 15331 22540 15397 22541
rect 15331 22476 15332 22540
rect 15396 22476 15397 22540
rect 15331 22475 15397 22476
rect 15147 21452 15213 21453
rect 15147 21388 15148 21452
rect 15212 21388 15213 21452
rect 15147 21387 15213 21388
rect 15150 14925 15210 21387
rect 15334 16013 15394 22475
rect 15331 16012 15397 16013
rect 15331 15948 15332 16012
rect 15396 15948 15397 16012
rect 15331 15947 15397 15948
rect 15147 14924 15213 14925
rect 15147 14860 15148 14924
rect 15212 14860 15213 14924
rect 15147 14859 15213 14860
rect 14963 5676 15029 5677
rect 14963 5612 14964 5676
rect 15028 5612 15029 5676
rect 14963 5611 15029 5612
rect 14376 5408 14384 5472
rect 14448 5408 14464 5472
rect 14528 5408 14544 5472
rect 14608 5408 14624 5472
rect 14688 5408 14696 5472
rect 14376 4384 14696 5408
rect 14376 4320 14384 4384
rect 14448 4320 14464 4384
rect 14528 4320 14544 4384
rect 14608 4320 14624 4384
rect 14688 4320 14696 4384
rect 14376 3296 14696 4320
rect 14376 3232 14384 3296
rect 14448 3232 14464 3296
rect 14528 3232 14544 3296
rect 14608 3232 14624 3296
rect 14688 3232 14696 3296
rect 14376 2208 14696 3232
rect 14376 2144 14384 2208
rect 14448 2144 14464 2208
rect 14528 2144 14544 2208
rect 14608 2144 14624 2208
rect 14688 2144 14696 2208
rect 14376 1120 14696 2144
rect 14376 1056 14384 1120
rect 14448 1056 14464 1120
rect 14528 1056 14544 1120
rect 14608 1056 14624 1120
rect 14688 1056 14696 1120
rect 14376 1040 14696 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9660 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 10304 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 12972 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 10488 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0__0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1__0_
timestamp 1688980957
transform 1 0 13892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2__0_
timestamp 1688980957
transform 1 0 9936 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3__0_
timestamp 1688980957
transform 1 0 10488 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4__0_
timestamp 1688980957
transform 1 0 9936 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5__0_
timestamp 1688980957
transform 1 0 10212 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6__0_
timestamp 1688980957
transform 1 0 9476 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7__0_
timestamp 1688980957
transform 1 0 10672 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8__0_
timestamp 1688980957
transform 1 0 12880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9__0_
timestamp 1688980957
transform 1 0 9844 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10__0_
timestamp 1688980957
transform 1 0 11868 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11__0_
timestamp 1688980957
transform 1 0 10120 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12__0_
timestamp 1688980957
transform 1 0 10672 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13__0_
timestamp 1688980957
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14__0_
timestamp 1688980957
transform 1 0 10396 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15__0_
timestamp 1688980957
transform 1 0 10580 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16__0_
timestamp 1688980957
transform 1 0 10856 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17__0_
timestamp 1688980957
transform 1 0 11592 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18__0_
timestamp 1688980957
transform 1 0 9476 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19__0_
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20__0_
timestamp 1688980957
transform 1 0 11868 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21__0_
timestamp 1688980957
transform 1 0 11960 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22__0_
timestamp 1688980957
transform 1 0 12512 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23__0_
timestamp 1688980957
transform 1 0 11684 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24__0_
timestamp 1688980957
transform 1 0 12236 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25__0_
timestamp 1688980957
transform 1 0 12420 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26__0_
timestamp 1688980957
transform 1 0 10304 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27__0_
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28__0_
timestamp 1688980957
transform 1 0 12052 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29__0_
timestamp 1688980957
transform 1 0 13248 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30__0_
timestamp 1688980957
transform 1 0 7728 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31__0_
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0__0_
timestamp 1688980957
transform 1 0 10120 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1__0_
timestamp 1688980957
transform 1 0 13432 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2__0_
timestamp 1688980957
transform 1 0 10764 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3__0_
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4__0_
timestamp 1688980957
transform 1 0 10488 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5__0_
timestamp 1688980957
transform 1 0 11132 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6__0_
timestamp 1688980957
transform 1 0 10488 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7__0_
timestamp 1688980957
transform 1 0 10396 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8__0_
timestamp 1688980957
transform 1 0 11224 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9__0_
timestamp 1688980957
transform 1 0 10396 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10__0_
timestamp 1688980957
transform 1 0 10672 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11__0_
timestamp 1688980957
transform 1 0 10948 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12__0_
timestamp 1688980957
transform 1 0 11500 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13__0_
timestamp 1688980957
transform 1 0 10580 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14__0_
timestamp 1688980957
transform 1 0 11040 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15__0_
timestamp 1688980957
transform 1 0 10764 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16__0_
timestamp 1688980957
transform 1 0 11316 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17__0_
timestamp 1688980957
transform 1 0 11592 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18__0_
timestamp 1688980957
transform 1 0 10212 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19__0_
timestamp 1688980957
transform 1 0 9292 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20__0_
timestamp 1688980957
transform 1 0 12236 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21__0_
timestamp 1688980957
transform 1 0 11960 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22__0_
timestamp 1688980957
transform 1 0 11684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23__0_
timestamp 1688980957
transform 1 0 12604 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24__0_
timestamp 1688980957
transform 1 0 12696 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25__0_
timestamp 1688980957
transform 1 0 11868 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26__0_
timestamp 1688980957
transform 1 0 10948 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27__0_
timestamp 1688980957
transform 1 0 12144 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28__0_
timestamp 1688980957
transform 1 0 12328 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29__0_
timestamp 1688980957
transform 1 0 12420 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30__0_
timestamp 1688980957
transform 1 0 8372 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31__0_
timestamp 1688980957
transform 1 0 9476 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_15 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2484 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_39 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4692 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_52
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_70 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77
timestamp 1688980957
transform 1 0 8188 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_88 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_93
timestamp 1688980957
transform 1 0 9660 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10764 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_117
timestamp 1688980957
transform 1 0 11868 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 1688980957
transform 1 0 1932 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_34
timestamp 1688980957
transform 1 0 4232 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_46 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5336 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_54
timestamp 1688980957
transform 1 0 6072 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_61
timestamp 1688980957
transform 1 0 6716 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_68
timestamp 1688980957
transform 1 0 7360 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_76
timestamp 1688980957
transform 1 0 8096 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_84
timestamp 1688980957
transform 1 0 8832 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_92
timestamp 1688980957
transform 1 0 9568 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_100
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_108
timestamp 1688980957
transform 1 0 11040 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_117
timestamp 1688980957
transform 1 0 11868 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_124
timestamp 1688980957
transform 1 0 12512 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_131
timestamp 1688980957
transform 1 0 13156 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1688980957
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_18
timestamp 1688980957
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_30
timestamp 1688980957
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_42
timestamp 1688980957
transform 1 0 4968 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_54
timestamp 1688980957
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_101
timestamp 1688980957
transform 1 0 10396 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_133
timestamp 1688980957
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_115
timestamp 1688980957
transform 1 0 11684 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_12
timestamp 1688980957
transform 1 0 2208 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_24
timestamp 1688980957
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_36
timestamp 1688980957
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_48
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_104
timestamp 1688980957
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_9
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_16
timestamp 1688980957
transform 1 0 2576 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_82
timestamp 1688980957
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_18
timestamp 1688980957
transform 1 0 2760 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 1688980957
transform 1 0 3864 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_42
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_73
timestamp 1688980957
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 1688980957
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_61
timestamp 1688980957
transform 1 0 6716 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_106
timestamp 1688980957
transform 1 0 10856 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_12
timestamp 1688980957
transform 1 0 2208 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_24
timestamp 1688980957
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_36
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_48
timestamp 1688980957
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_65
timestamp 1688980957
transform 1 0 7084 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_87
timestamp 1688980957
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 1688980957
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 1688980957
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_91
timestamp 1688980957
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_113
timestamp 1688980957
transform 1 0 11500 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_67
timestamp 1688980957
transform 1 0 7268 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_75
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_84
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_92
timestamp 1688980957
transform 1 0 9568 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_123
timestamp 1688980957
transform 1 0 12420 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1688980957
transform 1 0 2852 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_18
timestamp 1688980957
transform 1 0 2760 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_30
timestamp 1688980957
transform 1 0 3864 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_42
timestamp 1688980957
transform 1 0 4968 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_54
timestamp 1688980957
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_87
timestamp 1688980957
transform 1 0 9108 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_109
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_117
timestamp 1688980957
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_21
timestamp 1688980957
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_137
timestamp 1688980957
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_12
timestamp 1688980957
transform 1 0 2208 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_24
timestamp 1688980957
transform 1 0 3312 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_36
timestamp 1688980957
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_48
timestamp 1688980957
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_63
timestamp 1688980957
transform 1 0 6900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_70
timestamp 1688980957
transform 1 0 7544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_92
timestamp 1688980957
transform 1 0 9568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_96
timestamp 1688980957
transform 1 0 9936 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_74
timestamp 1688980957
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_101
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_21
timestamp 1688980957
transform 1 0 3036 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_33
timestamp 1688980957
transform 1 0 4140 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_86
timestamp 1688980957
transform 1 0 9016 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_98
timestamp 1688980957
transform 1 0 10120 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_12
timestamp 1688980957
transform 1 0 2208 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_24
timestamp 1688980957
transform 1 0 3312 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_80
timestamp 1688980957
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_101
timestamp 1688980957
transform 1 0 10396 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_135
timestamp 1688980957
transform 1 0 13524 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_18
timestamp 1688980957
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_30
timestamp 1688980957
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_42
timestamp 1688980957
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_63
timestamp 1688980957
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_79
timestamp 1688980957
transform 1 0 8372 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_83
timestamp 1688980957
transform 1 0 8740 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_99
timestamp 1688980957
transform 1 0 10212 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_12
timestamp 1688980957
transform 1 0 2208 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_24
timestamp 1688980957
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_106
timestamp 1688980957
transform 1 0 10856 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_134
timestamp 1688980957
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_9
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_21
timestamp 1688980957
transform 1 0 3036 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_33
timestamp 1688980957
transform 1 0 4140 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_45
timestamp 1688980957
transform 1 0 5244 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_53
timestamp 1688980957
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_65
timestamp 1688980957
transform 1 0 7084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_87
timestamp 1688980957
transform 1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_106
timestamp 1688980957
transform 1 0 10856 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_142
timestamp 1688980957
transform 1 0 14168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_18
timestamp 1688980957
transform 1 0 2760 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_26
timestamp 1688980957
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_49
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_72
timestamp 1688980957
transform 1 0 7728 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_119
timestamp 1688980957
transform 1 0 12052 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_12
timestamp 1688980957
transform 1 0 2208 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_24
timestamp 1688980957
transform 1 0 3312 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_36
timestamp 1688980957
transform 1 0 4416 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_40
timestamp 1688980957
transform 1 0 4784 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_72
timestamp 1688980957
transform 1 0 7728 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_7
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_19
timestamp 1688980957
transform 1 0 2852 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_134
timestamp 1688980957
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_18
timestamp 1688980957
transform 1 0 2760 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_30
timestamp 1688980957
transform 1 0 3864 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_42
timestamp 1688980957
transform 1 0 4968 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_54
timestamp 1688980957
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_61
timestamp 1688980957
transform 1 0 6716 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_77
timestamp 1688980957
transform 1 0 8188 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_85
timestamp 1688980957
transform 1 0 8924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_101
timestamp 1688980957
transform 1 0 10396 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_109
timestamp 1688980957
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_131
timestamp 1688980957
transform 1 0 13156 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_7
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_53
timestamp 1688980957
transform 1 0 5980 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_76
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_10
timestamp 1688980957
transform 1 0 2024 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_22
timestamp 1688980957
transform 1 0 3128 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_34
timestamp 1688980957
transform 1 0 4232 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_46
timestamp 1688980957
transform 1 0 5336 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_54
timestamp 1688980957
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_61
timestamp 1688980957
transform 1 0 6716 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_98
timestamp 1688980957
transform 1 0 10120 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_117
timestamp 1688980957
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_18
timestamp 1688980957
transform 1 0 2760 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1688980957
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_73
timestamp 1688980957
transform 1 0 7820 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_101
timestamp 1688980957
transform 1 0 10396 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_108
timestamp 1688980957
transform 1 0 11040 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_7
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_19
timestamp 1688980957
transform 1 0 2852 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_31
timestamp 1688980957
transform 1 0 3956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_61
timestamp 1688980957
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_77
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_89
timestamp 1688980957
transform 1 0 9292 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_93
timestamp 1688980957
transform 1 0 9660 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_121
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_7
timestamp 1688980957
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_19
timestamp 1688980957
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_47
timestamp 1688980957
transform 1 0 5428 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_62
timestamp 1688980957
transform 1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 1688980957
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_115
timestamp 1688980957
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_122
timestamp 1688980957
transform 1 0 12328 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_138
timestamp 1688980957
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 1688980957
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 1688980957
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 1688980957
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 1688980957
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_75
timestamp 1688980957
transform 1 0 8004 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_102
timestamp 1688980957
transform 1 0 10488 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_121
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_19
timestamp 1688980957
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_37
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_58
timestamp 1688980957
transform 1 0 6440 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_65
timestamp 1688980957
transform 1 0 7084 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_100
timestamp 1688980957
transform 1 0 10304 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_117
timestamp 1688980957
transform 1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_13
timestamp 1688980957
transform 1 0 2300 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_25
timestamp 1688980957
transform 1 0 3404 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_37
timestamp 1688980957
transform 1 0 4508 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_49
timestamp 1688980957
transform 1 0 5612 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_63
timestamp 1688980957
transform 1 0 6900 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_79
timestamp 1688980957
transform 1 0 8372 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_91
timestamp 1688980957
transform 1 0 9476 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_116
timestamp 1688980957
transform 1 0 11776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_138
timestamp 1688980957
transform 1 0 13800 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_142
timestamp 1688980957
transform 1 0 14168 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_15
timestamp 1688980957
transform 1 0 2484 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_24
timestamp 1688980957
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_49
timestamp 1688980957
transform 1 0 5612 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_69
timestamp 1688980957
transform 1 0 7452 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_81
timestamp 1688980957
transform 1 0 8556 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_93
timestamp 1688980957
transform 1 0 9660 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_7
timestamp 1688980957
transform 1 0 1748 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_19
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_31
timestamp 1688980957
transform 1 0 3956 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_39
timestamp 1688980957
transform 1 0 4692 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_7
timestamp 1688980957
transform 1 0 1748 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_19
timestamp 1688980957
transform 1 0 2852 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_47
timestamp 1688980957
transform 1 0 5428 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_63
timestamp 1688980957
transform 1 0 6900 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_93
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_130
timestamp 1688980957
transform 1 0 13064 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_138
timestamp 1688980957
transform 1 0 13800 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_61
timestamp 1688980957
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_77
timestamp 1688980957
transform 1 0 8188 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_98
timestamp 1688980957
transform 1 0 10120 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_110
timestamp 1688980957
transform 1 0 11224 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_138
timestamp 1688980957
transform 1 0 13800 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_7
timestamp 1688980957
transform 1 0 1748 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_19
timestamp 1688980957
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_124
timestamp 1688980957
transform 1 0 12512 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_7
timestamp 1688980957
transform 1 0 1748 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_19
timestamp 1688980957
transform 1 0 2852 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_31
timestamp 1688980957
transform 1 0 3956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_43
timestamp 1688980957
transform 1 0 5060 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_65
timestamp 1688980957
transform 1 0 7084 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_89
timestamp 1688980957
transform 1 0 9292 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_110
timestamp 1688980957
transform 1 0 11224 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 1688980957
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_35
timestamp 1688980957
transform 1 0 4324 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_72
timestamp 1688980957
transform 1 0 7728 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_100
timestamp 1688980957
transform 1 0 10304 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 1688980957
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_7
timestamp 1688980957
transform 1 0 1748 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_19
timestamp 1688980957
transform 1 0 2852 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_31
timestamp 1688980957
transform 1 0 3956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_43
timestamp 1688980957
transform 1 0 5060 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_72
timestamp 1688980957
transform 1 0 7728 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_84
timestamp 1688980957
transform 1 0 8832 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_96
timestamp 1688980957
transform 1 0 9936 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_138
timestamp 1688980957
transform 1 0 13800 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_142
timestamp 1688980957
transform 1 0 14168 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_13
timestamp 1688980957
transform 1 0 2300 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_25
timestamp 1688980957
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_57
timestamp 1688980957
transform 1 0 6348 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_73
timestamp 1688980957
transform 1 0 7820 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_81
timestamp 1688980957
transform 1 0 8556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_106
timestamp 1688980957
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_110
timestamp 1688980957
transform 1 0 11224 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_132
timestamp 1688980957
transform 1 0 13248 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_108
timestamp 1688980957
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_119
timestamp 1688980957
transform 1 0 12052 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_7
timestamp 1688980957
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_19
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_78
timestamp 1688980957
transform 1 0 8280 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_97
timestamp 1688980957
transform 1 0 10028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_101
timestamp 1688980957
transform 1 0 10396 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_123
timestamp 1688980957
transform 1 0 12420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_7
timestamp 1688980957
transform 1 0 1748 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_21
timestamp 1688980957
transform 1 0 3036 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_33
timestamp 1688980957
transform 1 0 4140 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_78
timestamp 1688980957
transform 1 0 8280 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_90
timestamp 1688980957
transform 1 0 9384 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_94
timestamp 1688980957
transform 1 0 9752 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 1688980957
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_119
timestamp 1688980957
transform 1 0 12052 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_20
timestamp 1688980957
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_65
timestamp 1688980957
transform 1 0 7084 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_135
timestamp 1688980957
transform 1 0 13524 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_7
timestamp 1688980957
transform 1 0 1748 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_19
timestamp 1688980957
transform 1 0 2852 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_31
timestamp 1688980957
transform 1 0 3956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_43
timestamp 1688980957
transform 1 0 5060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_63
timestamp 1688980957
transform 1 0 6900 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_119
timestamp 1688980957
transform 1 0 12052 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_7
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_19
timestamp 1688980957
transform 1 0 2852 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 1688980957
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_80
timestamp 1688980957
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_97
timestamp 1688980957
transform 1 0 10028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_101
timestamp 1688980957
transform 1 0 10396 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_104
timestamp 1688980957
transform 1 0 10672 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 1688980957
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 1688980957
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_110
timestamp 1688980957
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_131
timestamp 1688980957
transform 1 0 13156 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_140
timestamp 1688980957
transform 1 0 13984 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_7
timestamp 1688980957
transform 1 0 1748 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_12
timestamp 1688980957
transform 1 0 2208 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_24
timestamp 1688980957
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_69
timestamp 1688980957
transform 1 0 7452 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_81
timestamp 1688980957
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_93
timestamp 1688980957
transform 1 0 9660 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_115
timestamp 1688980957
transform 1 0 11684 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_7
timestamp 1688980957
transform 1 0 1748 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_19
timestamp 1688980957
transform 1 0 2852 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_31
timestamp 1688980957
transform 1 0 3956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_43
timestamp 1688980957
transform 1 0 5060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_81
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_85
timestamp 1688980957
transform 1 0 8924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_107
timestamp 1688980957
transform 1 0 10948 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_117
timestamp 1688980957
transform 1 0 11868 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_142
timestamp 1688980957
transform 1 0 14168 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 1688980957
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_65
timestamp 1688980957
transform 1 0 7084 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_82
timestamp 1688980957
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_100
timestamp 1688980957
transform 1 0 10304 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_7
timestamp 1688980957
transform 1 0 1748 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_19
timestamp 1688980957
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_31
timestamp 1688980957
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_43
timestamp 1688980957
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_99
timestamp 1688980957
transform 1 0 10212 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_142
timestamp 1688980957
transform 1 0 14168 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_7
timestamp 1688980957
transform 1 0 1748 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_19
timestamp 1688980957
transform 1 0 2852 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 1688980957
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 1688980957
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_94
timestamp 1688980957
transform 1 0 9752 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_108
timestamp 1688980957
transform 1 0 11040 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_112
timestamp 1688980957
transform 1 0 11408 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_120
timestamp 1688980957
transform 1 0 12144 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_7
timestamp 1688980957
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_19
timestamp 1688980957
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 1688980957
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 1688980957
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 1688980957
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 1688980957
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_7
timestamp 1688980957
transform 1 0 1748 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_19
timestamp 1688980957
transform 1 0 2852 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_31
timestamp 1688980957
transform 1 0 3956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_43
timestamp 1688980957
transform 1 0 5060 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_107
timestamp 1688980957
transform 1 0 10948 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_128
timestamp 1688980957
transform 1 0 12880 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_142
timestamp 1688980957
transform 1 0 14168 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 1688980957
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_93
timestamp 1688980957
transform 1 0 9660 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_7
timestamp 1688980957
transform 1 0 1748 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_19
timestamp 1688980957
transform 1 0 2852 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_31
timestamp 1688980957
transform 1 0 3956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_43
timestamp 1688980957
transform 1 0 5060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_47
timestamp 1688980957
transform 1 0 5428 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_101
timestamp 1688980957
transform 1 0 10396 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_130
timestamp 1688980957
transform 1 0 13064 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_7
timestamp 1688980957
transform 1 0 1748 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_19
timestamp 1688980957
transform 1 0 2852 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_47
timestamp 1688980957
transform 1 0 5428 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_51
timestamp 1688980957
transform 1 0 5796 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_63
timestamp 1688980957
transform 1 0 6900 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_75
timestamp 1688980957
transform 1 0 8004 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_88
timestamp 1688980957
transform 1 0 9200 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_94
timestamp 1688980957
transform 1 0 9752 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_102
timestamp 1688980957
transform 1 0 10488 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_111
timestamp 1688980957
transform 1 0 11316 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_131
timestamp 1688980957
transform 1 0 13156 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_138
timestamp 1688980957
transform 1 0 13800 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_92
timestamp 1688980957
transform 1 0 9568 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_98
timestamp 1688980957
transform 1 0 10120 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_102
timestamp 1688980957
transform 1 0 10488 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_142
timestamp 1688980957
transform 1 0 14168 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_12
timestamp 1688980957
transform 1 0 2208 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_24
timestamp 1688980957
transform 1 0 3312 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_138
timestamp 1688980957
transform 1 0 13800 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_10
timestamp 1688980957
transform 1 0 2024 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_22
timestamp 1688980957
transform 1 0 3128 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_34
timestamp 1688980957
transform 1 0 4232 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_46
timestamp 1688980957
transform 1 0 5336 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_54
timestamp 1688980957
transform 1 0 6072 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_105
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_124
timestamp 1688980957
transform 1 0 12512 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_142
timestamp 1688980957
transform 1 0 14168 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_103
timestamp 1688980957
transform 1 0 10580 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_127
timestamp 1688980957
transform 1 0 12788 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_7
timestamp 1688980957
transform 1 0 1748 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_19
timestamp 1688980957
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_31
timestamp 1688980957
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_43
timestamp 1688980957
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_110
timestamp 1688980957
transform 1 0 11224 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_116
timestamp 1688980957
transform 1 0 11776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_142
timestamp 1688980957
transform 1 0 14168 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_7
timestamp 1688980957
transform 1 0 1748 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_19
timestamp 1688980957
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_65
timestamp 1688980957
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_77
timestamp 1688980957
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_117
timestamp 1688980957
transform 1 0 11868 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_138
timestamp 1688980957
transform 1 0 13800 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_39
timestamp 1688980957
transform 1 0 4692 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_51
timestamp 1688980957
transform 1 0 5796 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_121
timestamp 1688980957
transform 1 0 12236 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_141
timestamp 1688980957
transform 1 0 14076 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_9
timestamp 1688980957
transform 1 0 1932 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_21
timestamp 1688980957
transform 1 0 3036 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_27
timestamp 1688980957
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_71
timestamp 1688980957
transform 1 0 7636 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_75
timestamp 1688980957
transform 1 0 8004 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_82
timestamp 1688980957
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_88
timestamp 1688980957
transform 1 0 9200 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_94
timestamp 1688980957
transform 1 0 9752 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_106
timestamp 1688980957
transform 1 0 10856 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_118
timestamp 1688980957
transform 1 0 11960 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_126
timestamp 1688980957
transform 1 0 12696 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_138
timestamp 1688980957
transform 1 0 13800 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_7
timestamp 1688980957
transform 1 0 1748 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_19
timestamp 1688980957
transform 1 0 2852 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_31
timestamp 1688980957
transform 1 0 3956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_43
timestamp 1688980957
transform 1 0 5060 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_131
timestamp 1688980957
transform 1 0 13156 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_135
timestamp 1688980957
transform 1 0 13524 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_7
timestamp 1688980957
transform 1 0 1748 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_19
timestamp 1688980957
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_31
timestamp 1688980957
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_43
timestamp 1688980957
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_129
timestamp 1688980957
transform 1 0 12972 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_12
timestamp 1688980957
transform 1 0 2208 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_24
timestamp 1688980957
transform 1 0 3312 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_35
timestamp 1688980957
transform 1 0 4324 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_42
timestamp 1688980957
transform 1 0 4968 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_54
timestamp 1688980957
transform 1 0 6072 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_131
timestamp 1688980957
transform 1 0 13156 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_142
timestamp 1688980957
transform 1 0 14168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_26
timestamp 1688980957
transform 1 0 3496 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_35
timestamp 1688980957
transform 1 0 4324 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_39
timestamp 1688980957
transform 1 0 4692 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_43
timestamp 1688980957
transform 1 0 5060 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_55
timestamp 1688980957
transform 1 0 6164 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_59
timestamp 1688980957
transform 1 0 6532 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_63
timestamp 1688980957
transform 1 0 6900 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_67
timestamp 1688980957
transform 1 0 7268 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_71
timestamp 1688980957
transform 1 0 7636 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_75
timestamp 1688980957
transform 1 0 8004 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_79
timestamp 1688980957
transform 1 0 8372 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1688980957
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_91
timestamp 1688980957
transform 1 0 9476 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_98
timestamp 1688980957
transform 1 0 10120 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_102
timestamp 1688980957
transform 1 0 10488 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_107
timestamp 1688980957
transform 1 0 10948 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_111
timestamp 1688980957
transform 1 0 11316 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_115
timestamp 1688980957
transform 1 0 11684 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_119
timestamp 1688980957
transform 1 0 12052 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_123
timestamp 1688980957
transform 1 0 12420 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_129
timestamp 1688980957
transform 1 0 12972 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1688980957
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_9
timestamp 1688980957
transform 1 0 1932 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_14
timestamp 1688980957
transform 1 0 2392 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_25
timestamp 1688980957
transform 1 0 3404 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_33
timestamp 1688980957
transform 1 0 4140 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_40
timestamp 1688980957
transform 1 0 4784 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_46
timestamp 1688980957
transform 1 0 5336 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_54
timestamp 1688980957
transform 1 0 6072 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_62
timestamp 1688980957
transform 1 0 6808 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_70
timestamp 1688980957
transform 1 0 7544 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_78
timestamp 1688980957
transform 1 0 8280 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_89
timestamp 1688980957
transform 1 0 9292 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_94
timestamp 1688980957
transform 1 0 9752 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_102
timestamp 1688980957
transform 1 0 10488 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_118
timestamp 1688980957
transform 1 0 11960 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_128
timestamp 1688980957
transform 1 0 12880 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_141
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input10
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input16
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input18
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input19
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input20 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input21
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input22
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input24
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  input35 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 9384 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 11592 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 13064 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 13340 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 13984 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 12788 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input46
timestamp 1688980957
transform 1 0 2024 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input47
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  input48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1688980957
transform 1 0 4324 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1688980957
transform 1 0 4968 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 7268 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1688980957
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1688980957
transform 1 0 11868 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1688980957
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1688980957
transform 1 0 13524 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1688980957
transform 1 0 12788 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1688980957
transform 1 0 11960 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1688980957
transform 1 0 13892 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1688980957
transform 1 0 13892 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1688980957
transform 1 0 12236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1688980957
transform 1 0 10488 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform 1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1688980957
transform 1 0 11684 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1688980957
transform 1 0 11592 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1688980957
transform 1 0 9752 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1688980957
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input76
timestamp 1688980957
transform 1 0 11408 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input77
timestamp 1688980957
transform 1 0 10488 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1688980957
transform 1 0 13800 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1688980957
transform 1 0 11684 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1688980957
transform 1 0 13064 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1688980957
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1688980957
transform 1 0 13340 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1688980957
transform 1 0 13892 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1688980957
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1688980957
transform 1 0 11132 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input87
timestamp 1688980957
transform 1 0 12788 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1688980957
transform 1 0 12880 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input89
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1688980957
transform 1 0 13156 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input91
timestamp 1688980957
transform 1 0 13984 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input92
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input93
timestamp 1688980957
transform 1 0 11684 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input94
timestamp 1688980957
transform 1 0 13340 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp 1688980957
transform 1 0 11684 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input96
timestamp 1688980957
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input97
timestamp 1688980957
transform 1 0 12052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input98
timestamp 1688980957
transform 1 0 11684 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input99
timestamp 1688980957
transform 1 0 11868 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input100
timestamp 1688980957
transform 1 0 10488 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1688980957
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input102
timestamp 1688980957
transform 1 0 10488 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access__0_
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access__1_
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access__2_
timestamp 1688980957
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_config_Config_access__3_
timestamp 1688980957
transform 1 0 1748 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_A_IO_1_bidirectional_frame_config_pass__0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_A_IO_1_bidirectional_frame_config_pass__1_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  Inst_A_IO_1_bidirectional_frame_config_pass__2_
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_A_IO_1_bidirectional_frame_config_pass__3_
timestamp 1688980957
transform 1 0 5060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access__0_
timestamp 1688980957
transform 1 0 2300 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access__1_
timestamp 1688980957
transform 1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access__2_
timestamp 1688980957
transform 1 0 2300 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_config_Config_access__3_
timestamp 1688980957
transform 1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_B_IO_1_bidirectional_frame_config_pass__0_
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_B_IO_1_bidirectional_frame_config_pass__1_
timestamp 1688980957
transform 1 0 4600 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  Inst_B_IO_1_bidirectional_frame_config_pass__2_
timestamp 1688980957
transform 1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_B_IO_1_bidirectional_frame_config_pass__3_
timestamp 1688980957
transform 1 0 6072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8740 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit1
timestamp 1688980957
transform 1 0 9752 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit2
timestamp 1688980957
transform 1 0 6808 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit3
timestamp 1688980957
transform 1 0 7360 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit4
timestamp 1688980957
transform 1 0 9844 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit5
timestamp 1688980957
transform 1 0 10304 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit6
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit7
timestamp 1688980957
transform 1 0 9108 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit8
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit9
timestamp 1688980957
transform 1 0 11500 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit10
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit11
timestamp 1688980957
transform 1 0 5520 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit12
timestamp 1688980957
transform 1 0 10396 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit13
timestamp 1688980957
transform 1 0 11684 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit14
timestamp 1688980957
transform 1 0 7268 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit15
timestamp 1688980957
transform 1 0 7452 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit16
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit17
timestamp 1688980957
transform 1 0 11500 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit18
timestamp 1688980957
transform 1 0 7912 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit19
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit20
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit21
timestamp 1688980957
transform 1 0 11408 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit22
timestamp 1688980957
transform 1 0 6808 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit23
timestamp 1688980957
transform 1 0 7268 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit24
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit25
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit26
timestamp 1688980957
transform 1 0 9292 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit27
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit28
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit29
timestamp 1688980957
transform 1 0 4876 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit30
timestamp 1688980957
transform 1 0 5704 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame0_bit31
timestamp 1688980957
transform 1 0 4324 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit0
timestamp 1688980957
transform 1 0 7084 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit1
timestamp 1688980957
transform 1 0 8464 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit2
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit3
timestamp 1688980957
transform 1 0 7636 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit4
timestamp 1688980957
transform 1 0 12144 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit5
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit6
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit7
timestamp 1688980957
transform 1 0 10304 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit8
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit9
timestamp 1688980957
transform 1 0 12512 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit10
timestamp 1688980957
transform 1 0 11316 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit11
timestamp 1688980957
transform 1 0 12420 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit12
timestamp 1688980957
transform 1 0 4968 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit13
timestamp 1688980957
transform 1 0 6440 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit14
timestamp 1688980957
transform 1 0 9844 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit15
timestamp 1688980957
transform 1 0 10212 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit16
timestamp 1688980957
transform 1 0 11592 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit17
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit18
timestamp 1688980957
transform 1 0 4876 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit19
timestamp 1688980957
transform 1 0 6072 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit20
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit21
timestamp 1688980957
transform 1 0 7452 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit22
timestamp 1688980957
transform 1 0 12512 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit23
timestamp 1688980957
transform 1 0 12880 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit24
timestamp 1688980957
transform 1 0 10948 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit25
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit26
timestamp 1688980957
transform 1 0 6900 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit27
timestamp 1688980957
transform 1 0 8280 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit28
timestamp 1688980957
transform 1 0 11776 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit29
timestamp 1688980957
transform 1 0 12604 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit30
timestamp 1688980957
transform 1 0 6992 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame1_bit31
timestamp 1688980957
transform 1 0 7452 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit0
timestamp 1688980957
transform 1 0 11776 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit1
timestamp 1688980957
transform 1 0 12512 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit2
timestamp 1688980957
transform 1 0 9476 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit3
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit4
timestamp 1688980957
transform 1 0 10488 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit5
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit6
timestamp 1688980957
transform 1 0 7452 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit7
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit8
timestamp 1688980957
transform 1 0 11684 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit9
timestamp 1688980957
transform 1 0 12420 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit10
timestamp 1688980957
transform 1 0 11684 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit11
timestamp 1688980957
transform 1 0 12420 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit12
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit13
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit14
timestamp 1688980957
transform 1 0 4876 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit15
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit16
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit17
timestamp 1688980957
transform 1 0 12512 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit18
timestamp 1688980957
transform 1 0 6072 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit19
timestamp 1688980957
transform 1 0 6992 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit20
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit21
timestamp 1688980957
transform 1 0 12512 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit22
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit23
timestamp 1688980957
transform 1 0 8832 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit24
timestamp 1688980957
transform 1 0 11960 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit25
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit26
timestamp 1688980957
transform 1 0 9844 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit27
timestamp 1688980957
transform 1 0 10488 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit28
timestamp 1688980957
transform 1 0 11868 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit29
timestamp 1688980957
transform 1 0 12604 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit30
timestamp 1688980957
transform 1 0 4416 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame2_bit31
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit14
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit15
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit16
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit17
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit18
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit19
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit20
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit21
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit22
timestamp 1688980957
transform 1 0 9752 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit23
timestamp 1688980957
transform 1 0 5060 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit24
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit25
timestamp 1688980957
transform 1 0 9752 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit26
timestamp 1688980957
transform 1 0 6440 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit27
timestamp 1688980957
transform 1 0 6716 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit28
timestamp 1688980957
transform 1 0 8740 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit29
timestamp 1688980957
transform 1 0 9016 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit30
timestamp 1688980957
transform 1 0 6808 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_W_IO_ConfigMem_Inst_frame3_bit31
timestamp 1688980957
transform 1 0 7452 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__2_
timestamp 1688980957
transform 1 0 10764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10488 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 11040 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__2_
timestamp 1688980957
transform 1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__3_
timestamp 1688980957
transform 1 0 6440 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__4_
timestamp 1688980957
transform 1 0 6440 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 7912 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 6164 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__2_
timestamp 1688980957
transform 1 0 7360 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__3_
timestamp 1688980957
transform 1 0 7728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__4_
timestamp 1688980957
transform 1 0 6992 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 7636 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 6808 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__2_
timestamp 1688980957
transform 1 0 10672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__3_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__4_
timestamp 1688980957
transform 1 0 10948 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6808 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG1
timestamp 1688980957
transform 1 0 9200 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG2
timestamp 1688980957
transform 1 0 8096 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG3
timestamp 1688980957
transform 1 0 12052 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG4
timestamp 1688980957
transform 1 0 10120 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG5
timestamp 1688980957
transform 1 0 11224 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG6
timestamp 1688980957
transform 1 0 8556 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG7
timestamp 1688980957
transform 1 0 12328 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb0
timestamp 1688980957
transform 1 0 12328 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb1
timestamp 1688980957
transform 1 0 9476 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb2
timestamp 1688980957
transform 1 0 5796 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb3
timestamp 1688980957
transform 1 0 12052 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb4
timestamp 1688980957
transform 1 0 7176 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb5
timestamp 1688980957
transform 1 0 12328 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb6
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb7
timestamp 1688980957
transform 1 0 12328 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG0
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG1
timestamp 1688980957
transform 1 0 12328 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG2
timestamp 1688980957
transform 1 0 7544 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG3
timestamp 1688980957
transform 1 0 9752 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG4
timestamp 1688980957
transform 1 0 7360 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG5
timestamp 1688980957
transform 1 0 10856 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG6
timestamp 1688980957
transform 1 0 9016 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG7
timestamp 1688980957
transform 1 0 11776 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5796 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG9
timestamp 1688980957
transform 1 0 11960 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG10
timestamp 1688980957
transform 1 0 8004 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG11
timestamp 1688980957
transform 1 0 11684 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG0
timestamp 1688980957
transform 1 0 10580 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG1
timestamp 1688980957
transform 1 0 12328 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG2
timestamp 1688980957
transform 1 0 5796 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG3
timestamp 1688980957
transform 1 0 8924 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG4
timestamp 1688980957
transform 1 0 7912 0 -1 10880
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG5
timestamp 1688980957
transform 1 0 12328 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG6
timestamp 1688980957
transform 1 0 10120 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG7
timestamp 1688980957
transform 1 0 12328 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG8
timestamp 1688980957
transform 1 0 12328 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG9
timestamp 1688980957
transform 1 0 6348 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG10
timestamp 1688980957
transform 1 0 10488 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG11
timestamp 1688980957
transform 1 0 12328 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG12
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG13
timestamp 1688980957
transform 1 0 6992 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG14
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG15
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 6992 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6900 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1_216 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8280 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1_218
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 6624 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 5612 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 6072 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 6348 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6624 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1_217
timestamp 1688980957
transform 1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1_219
timestamp 1688980957
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9200 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst2
timestamp 1688980957
transform 1 0 10856 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst3
timestamp 1688980957
transform 1 0 9476 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst4
timestamp 1688980957
transform 1 0 10488 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst2
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst3
timestamp 1688980957
transform 1 0 9568 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst4
timestamp 1688980957
transform 1 0 10580 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 11960 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 11684 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 11132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output119
timestamp 1688980957
transform 1 0 11776 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 11684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform 1 0 11316 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1688980957
transform 1 0 13892 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform 1 0 12328 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 12880 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform 1 0 11776 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform 1 0 11224 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 13248 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 11776 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 11868 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 13248 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1688980957
transform 1 0 13892 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output134
timestamp 1688980957
transform 1 0 13248 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 12052 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 12880 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 13616 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 12788 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform 1 0 9752 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 10856 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 11592 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 13616 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 13432 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output147
timestamp 1688980957
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output148
timestamp 1688980957
transform 1 0 12788 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output149
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output150
timestamp 1688980957
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output151
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output152
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output153
timestamp 1688980957
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output154
timestamp 1688980957
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output155
timestamp 1688980957
transform 1 0 10304 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output156
timestamp 1688980957
transform 1 0 11776 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output157
timestamp 1688980957
transform 1 0 12972 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output158
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output159
timestamp 1688980957
transform 1 0 12696 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output160
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output161
timestamp 1688980957
transform 1 0 13432 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output162
timestamp 1688980957
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output163
timestamp 1688980957
transform 1 0 12880 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output164
timestamp 1688980957
transform 1 0 12512 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output165
timestamp 1688980957
transform 1 0 10856 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output166
timestamp 1688980957
transform 1 0 13064 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output167
timestamp 1688980957
transform 1 0 13616 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output168
timestamp 1688980957
transform 1 0 13248 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1688980957
transform 1 0 12144 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output170
timestamp 1688980957
transform 1 0 12696 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output171
timestamp 1688980957
transform 1 0 12144 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output172
timestamp 1688980957
transform 1 0 13064 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1688980957
transform 1 0 12696 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output174
timestamp 1688980957
transform 1 0 13064 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output175
timestamp 1688980957
transform 1 0 13432 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output176
timestamp 1688980957
transform 1 0 13616 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output177
timestamp 1688980957
transform 1 0 12880 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1688980957
transform 1 0 12696 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output179
timestamp 1688980957
transform 1 0 13064 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1688980957
transform 1 0 12880 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output181
timestamp 1688980957
transform 1 0 13248 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output182
timestamp 1688980957
transform 1 0 12972 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output183
timestamp 1688980957
transform 1 0 13524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1688980957
transform 1 0 12880 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output185
timestamp 1688980957
transform 1 0 10948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output186
timestamp 1688980957
transform 1 0 13248 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output187
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output188
timestamp 1688980957
transform 1 0 13432 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output189
timestamp 1688980957
transform 1 0 11776 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output190
timestamp 1688980957
transform 1 0 12328 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output191
timestamp 1688980957
transform 1 0 12880 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 13156 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output193
timestamp 1688980957
transform 1 0 13616 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output194
timestamp 1688980957
transform 1 0 13248 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output195
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1688980957
transform 1 0 9384 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1688980957
transform 1 0 10120 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output199
timestamp 1688980957
transform 1 0 10856 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1688980957
transform 1 0 11592 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output201
timestamp 1688980957
transform 1 0 12328 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1688980957
transform 1 0 13064 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output203
timestamp 1688980957
transform 1 0 13616 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output204
timestamp 1688980957
transform 1 0 13064 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 13432 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1688980957
transform 1 0 2024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output207
timestamp 1688980957
transform 1 0 2576 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output209
timestamp 1688980957
transform 1 0 4232 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1688980957
transform 1 0 4968 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1688980957
transform 1 0 5704 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1688980957
transform 1 0 6440 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1688980957
transform 1 0 7176 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1688980957
transform 1 0 7912 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  output215
timestamp 1688980957
transform 1 0 3128 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 14536 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 14536 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 14536 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 14536 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 14536 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 14536 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 14536 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 14536 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 14536 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 14536 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 14536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 14536 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 14536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 14536 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 14536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 14536 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 14536 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 14536 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 14536 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 14536 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 14536 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 14536 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 14536 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 14536 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 14536 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 14536 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 14536 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 14536 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 14536 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 14536 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 14536 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 14536 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 14536 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 14536 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 14536 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 14536 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 14536 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 14536 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 14536 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 14536 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 14536 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 14536 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 14536 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 14536 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 14536 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 14536 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 14536 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 14536 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 14536 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 14536 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 14536 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 14536 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 14536 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 14536 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 14536 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 14536 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 14536 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 14536 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 14536 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 14536 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 14536 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 14536 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 14536 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 14536 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 14536 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 14536 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 14536 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 14536 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 14536 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 14536 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 14536 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 14536 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 1932 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 1932 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 2760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 4048 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 4692 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 5520 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 6992 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 7728 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 8464 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 9936 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 10672 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 12144 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 12788 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 13248 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 13616 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 1748 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 2668 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 3220 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 4048 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 4784 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 5520 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 6256 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 6992 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 7728 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 8464 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 9200 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 9844 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 10672 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 11408 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 12144 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 13616 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 13616 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 13064 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 13340 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s -300 11160 160 11280 0 FreeSans 480 0 0 0 A_I_top
port 0 nsew signal tristate
flabel metal3 s -300 9528 160 9648 0 FreeSans 480 0 0 0 A_O_top
port 1 nsew signal input
flabel metal3 s -300 10344 160 10464 0 FreeSans 480 0 0 0 A_T_top
port 2 nsew signal tristate
flabel metal3 s -300 11976 160 12096 0 FreeSans 480 0 0 0 A_config_C_bit0
port 3 nsew signal tristate
flabel metal3 s -300 12792 160 12912 0 FreeSans 480 0 0 0 A_config_C_bit1
port 4 nsew signal tristate
flabel metal3 s -300 13608 160 13728 0 FreeSans 480 0 0 0 A_config_C_bit2
port 5 nsew signal tristate
flabel metal3 s -300 14424 160 14544 0 FreeSans 480 0 0 0 A_config_C_bit3
port 6 nsew signal tristate
flabel metal3 s -300 5448 160 5568 0 FreeSans 480 0 0 0 B_I_top
port 7 nsew signal tristate
flabel metal3 s -300 3816 160 3936 0 FreeSans 480 0 0 0 B_O_top
port 8 nsew signal input
flabel metal3 s -300 4632 160 4752 0 FreeSans 480 0 0 0 B_T_top
port 9 nsew signal tristate
flabel metal3 s -300 6264 160 6384 0 FreeSans 480 0 0 0 B_config_C_bit0
port 10 nsew signal tristate
flabel metal3 s -300 7080 160 7200 0 FreeSans 480 0 0 0 B_config_C_bit1
port 11 nsew signal tristate
flabel metal3 s -300 7896 160 8016 0 FreeSans 480 0 0 0 B_config_C_bit2
port 12 nsew signal tristate
flabel metal3 s -300 8712 160 8832 0 FreeSans 480 0 0 0 B_config_C_bit3
port 13 nsew signal tristate
flabel metal3 s 15540 17960 16000 18080 0 FreeSans 480 0 0 0 E1BEG[0]
port 14 nsew signal tristate
flabel metal3 s 15540 18232 16000 18352 0 FreeSans 480 0 0 0 E1BEG[1]
port 15 nsew signal tristate
flabel metal3 s 15540 18504 16000 18624 0 FreeSans 480 0 0 0 E1BEG[2]
port 16 nsew signal tristate
flabel metal3 s 15540 18776 16000 18896 0 FreeSans 480 0 0 0 E1BEG[3]
port 17 nsew signal tristate
flabel metal3 s 15540 19048 16000 19168 0 FreeSans 480 0 0 0 E2BEG[0]
port 18 nsew signal tristate
flabel metal3 s 15540 19320 16000 19440 0 FreeSans 480 0 0 0 E2BEG[1]
port 19 nsew signal tristate
flabel metal3 s 15540 19592 16000 19712 0 FreeSans 480 0 0 0 E2BEG[2]
port 20 nsew signal tristate
flabel metal3 s 15540 19864 16000 19984 0 FreeSans 480 0 0 0 E2BEG[3]
port 21 nsew signal tristate
flabel metal3 s 15540 20136 16000 20256 0 FreeSans 480 0 0 0 E2BEG[4]
port 22 nsew signal tristate
flabel metal3 s 15540 20408 16000 20528 0 FreeSans 480 0 0 0 E2BEG[5]
port 23 nsew signal tristate
flabel metal3 s 15540 20680 16000 20800 0 FreeSans 480 0 0 0 E2BEG[6]
port 24 nsew signal tristate
flabel metal3 s 15540 20952 16000 21072 0 FreeSans 480 0 0 0 E2BEG[7]
port 25 nsew signal tristate
flabel metal3 s 15540 21224 16000 21344 0 FreeSans 480 0 0 0 E2BEGb[0]
port 26 nsew signal tristate
flabel metal3 s 15540 21496 16000 21616 0 FreeSans 480 0 0 0 E2BEGb[1]
port 27 nsew signal tristate
flabel metal3 s 15540 21768 16000 21888 0 FreeSans 480 0 0 0 E2BEGb[2]
port 28 nsew signal tristate
flabel metal3 s 15540 22040 16000 22160 0 FreeSans 480 0 0 0 E2BEGb[3]
port 29 nsew signal tristate
flabel metal3 s 15540 22312 16000 22432 0 FreeSans 480 0 0 0 E2BEGb[4]
port 30 nsew signal tristate
flabel metal3 s 15540 22584 16000 22704 0 FreeSans 480 0 0 0 E2BEGb[5]
port 31 nsew signal tristate
flabel metal3 s 15540 22856 16000 22976 0 FreeSans 480 0 0 0 E2BEGb[6]
port 32 nsew signal tristate
flabel metal3 s 15540 23128 16000 23248 0 FreeSans 480 0 0 0 E2BEGb[7]
port 33 nsew signal tristate
flabel metal3 s 15540 27752 16000 27872 0 FreeSans 480 0 0 0 E6BEG[0]
port 34 nsew signal tristate
flabel metal3 s 15540 30472 16000 30592 0 FreeSans 480 0 0 0 E6BEG[10]
port 35 nsew signal tristate
flabel metal3 s 15540 30744 16000 30864 0 FreeSans 480 0 0 0 E6BEG[11]
port 36 nsew signal tristate
flabel metal3 s 15540 28024 16000 28144 0 FreeSans 480 0 0 0 E6BEG[1]
port 37 nsew signal tristate
flabel metal3 s 15540 28296 16000 28416 0 FreeSans 480 0 0 0 E6BEG[2]
port 38 nsew signal tristate
flabel metal3 s 15540 28568 16000 28688 0 FreeSans 480 0 0 0 E6BEG[3]
port 39 nsew signal tristate
flabel metal3 s 15540 28840 16000 28960 0 FreeSans 480 0 0 0 E6BEG[4]
port 40 nsew signal tristate
flabel metal3 s 15540 29112 16000 29232 0 FreeSans 480 0 0 0 E6BEG[5]
port 41 nsew signal tristate
flabel metal3 s 15540 29384 16000 29504 0 FreeSans 480 0 0 0 E6BEG[6]
port 42 nsew signal tristate
flabel metal3 s 15540 29656 16000 29776 0 FreeSans 480 0 0 0 E6BEG[7]
port 43 nsew signal tristate
flabel metal3 s 15540 29928 16000 30048 0 FreeSans 480 0 0 0 E6BEG[8]
port 44 nsew signal tristate
flabel metal3 s 15540 30200 16000 30320 0 FreeSans 480 0 0 0 E6BEG[9]
port 45 nsew signal tristate
flabel metal3 s 15540 23400 16000 23520 0 FreeSans 480 0 0 0 EE4BEG[0]
port 46 nsew signal tristate
flabel metal3 s 15540 26120 16000 26240 0 FreeSans 480 0 0 0 EE4BEG[10]
port 47 nsew signal tristate
flabel metal3 s 15540 26392 16000 26512 0 FreeSans 480 0 0 0 EE4BEG[11]
port 48 nsew signal tristate
flabel metal3 s 15540 26664 16000 26784 0 FreeSans 480 0 0 0 EE4BEG[12]
port 49 nsew signal tristate
flabel metal3 s 15540 26936 16000 27056 0 FreeSans 480 0 0 0 EE4BEG[13]
port 50 nsew signal tristate
flabel metal3 s 15540 27208 16000 27328 0 FreeSans 480 0 0 0 EE4BEG[14]
port 51 nsew signal tristate
flabel metal3 s 15540 27480 16000 27600 0 FreeSans 480 0 0 0 EE4BEG[15]
port 52 nsew signal tristate
flabel metal3 s 15540 23672 16000 23792 0 FreeSans 480 0 0 0 EE4BEG[1]
port 53 nsew signal tristate
flabel metal3 s 15540 23944 16000 24064 0 FreeSans 480 0 0 0 EE4BEG[2]
port 54 nsew signal tristate
flabel metal3 s 15540 24216 16000 24336 0 FreeSans 480 0 0 0 EE4BEG[3]
port 55 nsew signal tristate
flabel metal3 s 15540 24488 16000 24608 0 FreeSans 480 0 0 0 EE4BEG[4]
port 56 nsew signal tristate
flabel metal3 s 15540 24760 16000 24880 0 FreeSans 480 0 0 0 EE4BEG[5]
port 57 nsew signal tristate
flabel metal3 s 15540 25032 16000 25152 0 FreeSans 480 0 0 0 EE4BEG[6]
port 58 nsew signal tristate
flabel metal3 s 15540 25304 16000 25424 0 FreeSans 480 0 0 0 EE4BEG[7]
port 59 nsew signal tristate
flabel metal3 s 15540 25576 16000 25696 0 FreeSans 480 0 0 0 EE4BEG[8]
port 60 nsew signal tristate
flabel metal3 s 15540 25848 16000 25968 0 FreeSans 480 0 0 0 EE4BEG[9]
port 61 nsew signal tristate
flabel metal3 s -300 15240 160 15360 0 FreeSans 480 0 0 0 FrameData[0]
port 62 nsew signal input
flabel metal3 s -300 23400 160 23520 0 FreeSans 480 0 0 0 FrameData[10]
port 63 nsew signal input
flabel metal3 s -300 24216 160 24336 0 FreeSans 480 0 0 0 FrameData[11]
port 64 nsew signal input
flabel metal3 s -300 25032 160 25152 0 FreeSans 480 0 0 0 FrameData[12]
port 65 nsew signal input
flabel metal3 s -300 25848 160 25968 0 FreeSans 480 0 0 0 FrameData[13]
port 66 nsew signal input
flabel metal3 s -300 26664 160 26784 0 FreeSans 480 0 0 0 FrameData[14]
port 67 nsew signal input
flabel metal3 s -300 27480 160 27600 0 FreeSans 480 0 0 0 FrameData[15]
port 68 nsew signal input
flabel metal3 s -300 28296 160 28416 0 FreeSans 480 0 0 0 FrameData[16]
port 69 nsew signal input
flabel metal3 s -300 29112 160 29232 0 FreeSans 480 0 0 0 FrameData[17]
port 70 nsew signal input
flabel metal3 s -300 29928 160 30048 0 FreeSans 480 0 0 0 FrameData[18]
port 71 nsew signal input
flabel metal3 s -300 30744 160 30864 0 FreeSans 480 0 0 0 FrameData[19]
port 72 nsew signal input
flabel metal3 s -300 16056 160 16176 0 FreeSans 480 0 0 0 FrameData[1]
port 73 nsew signal input
flabel metal3 s -300 31560 160 31680 0 FreeSans 480 0 0 0 FrameData[20]
port 74 nsew signal input
flabel metal3 s -300 32376 160 32496 0 FreeSans 480 0 0 0 FrameData[21]
port 75 nsew signal input
flabel metal3 s -300 33192 160 33312 0 FreeSans 480 0 0 0 FrameData[22]
port 76 nsew signal input
flabel metal3 s -300 34008 160 34128 0 FreeSans 480 0 0 0 FrameData[23]
port 77 nsew signal input
flabel metal3 s -300 34824 160 34944 0 FreeSans 480 0 0 0 FrameData[24]
port 78 nsew signal input
flabel metal3 s -300 35640 160 35760 0 FreeSans 480 0 0 0 FrameData[25]
port 79 nsew signal input
flabel metal3 s -300 36456 160 36576 0 FreeSans 480 0 0 0 FrameData[26]
port 80 nsew signal input
flabel metal3 s -300 37272 160 37392 0 FreeSans 480 0 0 0 FrameData[27]
port 81 nsew signal input
flabel metal3 s -300 38088 160 38208 0 FreeSans 480 0 0 0 FrameData[28]
port 82 nsew signal input
flabel metal3 s -300 38904 160 39024 0 FreeSans 480 0 0 0 FrameData[29]
port 83 nsew signal input
flabel metal3 s -300 16872 160 16992 0 FreeSans 480 0 0 0 FrameData[2]
port 84 nsew signal input
flabel metal3 s -300 39720 160 39840 0 FreeSans 480 0 0 0 FrameData[30]
port 85 nsew signal input
flabel metal3 s -300 40536 160 40656 0 FreeSans 480 0 0 0 FrameData[31]
port 86 nsew signal input
flabel metal3 s -300 17688 160 17808 0 FreeSans 480 0 0 0 FrameData[3]
port 87 nsew signal input
flabel metal3 s -300 18504 160 18624 0 FreeSans 480 0 0 0 FrameData[4]
port 88 nsew signal input
flabel metal3 s -300 19320 160 19440 0 FreeSans 480 0 0 0 FrameData[5]
port 89 nsew signal input
flabel metal3 s -300 20136 160 20256 0 FreeSans 480 0 0 0 FrameData[6]
port 90 nsew signal input
flabel metal3 s -300 20952 160 21072 0 FreeSans 480 0 0 0 FrameData[7]
port 91 nsew signal input
flabel metal3 s -300 21768 160 21888 0 FreeSans 480 0 0 0 FrameData[8]
port 92 nsew signal input
flabel metal3 s -300 22584 160 22704 0 FreeSans 480 0 0 0 FrameData[9]
port 93 nsew signal input
flabel metal3 s 15540 31016 16000 31136 0 FreeSans 480 0 0 0 FrameData_O[0]
port 94 nsew signal tristate
flabel metal3 s 15540 33736 16000 33856 0 FreeSans 480 0 0 0 FrameData_O[10]
port 95 nsew signal tristate
flabel metal3 s 15540 34008 16000 34128 0 FreeSans 480 0 0 0 FrameData_O[11]
port 96 nsew signal tristate
flabel metal3 s 15540 34280 16000 34400 0 FreeSans 480 0 0 0 FrameData_O[12]
port 97 nsew signal tristate
flabel metal3 s 15540 34552 16000 34672 0 FreeSans 480 0 0 0 FrameData_O[13]
port 98 nsew signal tristate
flabel metal3 s 15540 34824 16000 34944 0 FreeSans 480 0 0 0 FrameData_O[14]
port 99 nsew signal tristate
flabel metal3 s 15540 35096 16000 35216 0 FreeSans 480 0 0 0 FrameData_O[15]
port 100 nsew signal tristate
flabel metal3 s 15540 35368 16000 35488 0 FreeSans 480 0 0 0 FrameData_O[16]
port 101 nsew signal tristate
flabel metal3 s 15540 35640 16000 35760 0 FreeSans 480 0 0 0 FrameData_O[17]
port 102 nsew signal tristate
flabel metal3 s 15540 35912 16000 36032 0 FreeSans 480 0 0 0 FrameData_O[18]
port 103 nsew signal tristate
flabel metal3 s 15540 36184 16000 36304 0 FreeSans 480 0 0 0 FrameData_O[19]
port 104 nsew signal tristate
flabel metal3 s 15540 31288 16000 31408 0 FreeSans 480 0 0 0 FrameData_O[1]
port 105 nsew signal tristate
flabel metal3 s 15540 36456 16000 36576 0 FreeSans 480 0 0 0 FrameData_O[20]
port 106 nsew signal tristate
flabel metal3 s 15540 36728 16000 36848 0 FreeSans 480 0 0 0 FrameData_O[21]
port 107 nsew signal tristate
flabel metal3 s 15540 37000 16000 37120 0 FreeSans 480 0 0 0 FrameData_O[22]
port 108 nsew signal tristate
flabel metal3 s 15540 37272 16000 37392 0 FreeSans 480 0 0 0 FrameData_O[23]
port 109 nsew signal tristate
flabel metal3 s 15540 37544 16000 37664 0 FreeSans 480 0 0 0 FrameData_O[24]
port 110 nsew signal tristate
flabel metal3 s 15540 37816 16000 37936 0 FreeSans 480 0 0 0 FrameData_O[25]
port 111 nsew signal tristate
flabel metal3 s 15540 38088 16000 38208 0 FreeSans 480 0 0 0 FrameData_O[26]
port 112 nsew signal tristate
flabel metal3 s 15540 38360 16000 38480 0 FreeSans 480 0 0 0 FrameData_O[27]
port 113 nsew signal tristate
flabel metal3 s 15540 38632 16000 38752 0 FreeSans 480 0 0 0 FrameData_O[28]
port 114 nsew signal tristate
flabel metal3 s 15540 38904 16000 39024 0 FreeSans 480 0 0 0 FrameData_O[29]
port 115 nsew signal tristate
flabel metal3 s 15540 31560 16000 31680 0 FreeSans 480 0 0 0 FrameData_O[2]
port 116 nsew signal tristate
flabel metal3 s 15540 39176 16000 39296 0 FreeSans 480 0 0 0 FrameData_O[30]
port 117 nsew signal tristate
flabel metal3 s 15540 39448 16000 39568 0 FreeSans 480 0 0 0 FrameData_O[31]
port 118 nsew signal tristate
flabel metal3 s 15540 31832 16000 31952 0 FreeSans 480 0 0 0 FrameData_O[3]
port 119 nsew signal tristate
flabel metal3 s 15540 32104 16000 32224 0 FreeSans 480 0 0 0 FrameData_O[4]
port 120 nsew signal tristate
flabel metal3 s 15540 32376 16000 32496 0 FreeSans 480 0 0 0 FrameData_O[5]
port 121 nsew signal tristate
flabel metal3 s 15540 32648 16000 32768 0 FreeSans 480 0 0 0 FrameData_O[6]
port 122 nsew signal tristate
flabel metal3 s 15540 32920 16000 33040 0 FreeSans 480 0 0 0 FrameData_O[7]
port 123 nsew signal tristate
flabel metal3 s 15540 33192 16000 33312 0 FreeSans 480 0 0 0 FrameData_O[8]
port 124 nsew signal tristate
flabel metal3 s 15540 33464 16000 33584 0 FreeSans 480 0 0 0 FrameData_O[9]
port 125 nsew signal tristate
flabel metal2 s 1214 -300 1270 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 126 nsew signal input
flabel metal2 s 8574 -300 8630 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 127 nsew signal input
flabel metal2 s 9310 -300 9366 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 128 nsew signal input
flabel metal2 s 10046 -300 10102 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 129 nsew signal input
flabel metal2 s 10782 -300 10838 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 130 nsew signal input
flabel metal2 s 11518 -300 11574 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 131 nsew signal input
flabel metal2 s 12254 -300 12310 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 132 nsew signal input
flabel metal2 s 12990 -300 13046 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 133 nsew signal input
flabel metal2 s 13726 -300 13782 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 134 nsew signal input
flabel metal2 s 14462 -300 14518 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 135 nsew signal input
flabel metal2 s 15198 -300 15254 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 136 nsew signal input
flabel metal2 s 1950 -300 2006 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 137 nsew signal input
flabel metal2 s 2686 -300 2742 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 138 nsew signal input
flabel metal2 s 3422 -300 3478 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 139 nsew signal input
flabel metal2 s 4158 -300 4214 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 140 nsew signal input
flabel metal2 s 4894 -300 4950 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 141 nsew signal input
flabel metal2 s 5630 -300 5686 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 142 nsew signal input
flabel metal2 s 6366 -300 6422 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 143 nsew signal input
flabel metal2 s 7102 -300 7158 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 144 nsew signal input
flabel metal2 s 7838 -300 7894 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 145 nsew signal input
flabel metal2 s 1214 44540 1270 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 146 nsew signal tristate
flabel metal2 s 8574 44540 8630 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 147 nsew signal tristate
flabel metal2 s 9310 44540 9366 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 148 nsew signal tristate
flabel metal2 s 10046 44540 10102 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 149 nsew signal tristate
flabel metal2 s 10782 44540 10838 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 150 nsew signal tristate
flabel metal2 s 11518 44540 11574 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 151 nsew signal tristate
flabel metal2 s 12254 44540 12310 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 152 nsew signal tristate
flabel metal2 s 12990 44540 13046 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 153 nsew signal tristate
flabel metal2 s 13726 44540 13782 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 154 nsew signal tristate
flabel metal2 s 14462 44540 14518 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 155 nsew signal tristate
flabel metal2 s 15198 44540 15254 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 156 nsew signal tristate
flabel metal2 s 1950 44540 2006 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 157 nsew signal tristate
flabel metal2 s 2686 44540 2742 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 158 nsew signal tristate
flabel metal2 s 3422 44540 3478 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 159 nsew signal tristate
flabel metal2 s 4158 44540 4214 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 160 nsew signal tristate
flabel metal2 s 4894 44540 4950 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 161 nsew signal tristate
flabel metal2 s 5630 44540 5686 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 162 nsew signal tristate
flabel metal2 s 6366 44540 6422 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 163 nsew signal tristate
flabel metal2 s 7102 44540 7158 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 164 nsew signal tristate
flabel metal2 s 7838 44540 7894 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 165 nsew signal tristate
flabel metal2 s 478 -300 534 160 0 FreeSans 224 90 0 0 UserCLK
port 166 nsew signal input
flabel metal2 s 478 44540 534 45000 0 FreeSans 224 90 0 0 UserCLKo
port 167 nsew signal tristate
flabel metal4 s 4302 1040 4622 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 7660 1040 7980 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 11018 1040 11338 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 14376 1040 14696 43568 0 FreeSans 1920 90 0 0 VGND
port 168 nsew ground bidirectional
flabel metal4 s 2623 1040 2943 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 5981 1040 6301 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 9339 1040 9659 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal4 s 12697 1040 13017 43568 0 FreeSans 1920 90 0 0 VPWR
port 169 nsew power bidirectional
flabel metal3 s 15540 4904 16000 5024 0 FreeSans 480 0 0 0 W1END[0]
port 170 nsew signal input
flabel metal3 s 15540 5176 16000 5296 0 FreeSans 480 0 0 0 W1END[1]
port 171 nsew signal input
flabel metal3 s 15540 5448 16000 5568 0 FreeSans 480 0 0 0 W1END[2]
port 172 nsew signal input
flabel metal3 s 15540 5720 16000 5840 0 FreeSans 480 0 0 0 W1END[3]
port 173 nsew signal input
flabel metal3 s 15540 8168 16000 8288 0 FreeSans 480 0 0 0 W2END[0]
port 174 nsew signal input
flabel metal3 s 15540 8440 16000 8560 0 FreeSans 480 0 0 0 W2END[1]
port 175 nsew signal input
flabel metal3 s 15540 8712 16000 8832 0 FreeSans 480 0 0 0 W2END[2]
port 176 nsew signal input
flabel metal3 s 15540 8984 16000 9104 0 FreeSans 480 0 0 0 W2END[3]
port 177 nsew signal input
flabel metal3 s 15540 9256 16000 9376 0 FreeSans 480 0 0 0 W2END[4]
port 178 nsew signal input
flabel metal3 s 15540 9528 16000 9648 0 FreeSans 480 0 0 0 W2END[5]
port 179 nsew signal input
flabel metal3 s 15540 9800 16000 9920 0 FreeSans 480 0 0 0 W2END[6]
port 180 nsew signal input
flabel metal3 s 15540 10072 16000 10192 0 FreeSans 480 0 0 0 W2END[7]
port 181 nsew signal input
flabel metal3 s 15540 5992 16000 6112 0 FreeSans 480 0 0 0 W2MID[0]
port 182 nsew signal input
flabel metal3 s 15540 6264 16000 6384 0 FreeSans 480 0 0 0 W2MID[1]
port 183 nsew signal input
flabel metal3 s 15540 6536 16000 6656 0 FreeSans 480 0 0 0 W2MID[2]
port 184 nsew signal input
flabel metal3 s 15540 6808 16000 6928 0 FreeSans 480 0 0 0 W2MID[3]
port 185 nsew signal input
flabel metal3 s 15540 7080 16000 7200 0 FreeSans 480 0 0 0 W2MID[4]
port 186 nsew signal input
flabel metal3 s 15540 7352 16000 7472 0 FreeSans 480 0 0 0 W2MID[5]
port 187 nsew signal input
flabel metal3 s 15540 7624 16000 7744 0 FreeSans 480 0 0 0 W2MID[6]
port 188 nsew signal input
flabel metal3 s 15540 7896 16000 8016 0 FreeSans 480 0 0 0 W2MID[7]
port 189 nsew signal input
flabel metal3 s 15540 14696 16000 14816 0 FreeSans 480 0 0 0 W6END[0]
port 190 nsew signal input
flabel metal3 s 15540 17416 16000 17536 0 FreeSans 480 0 0 0 W6END[10]
port 191 nsew signal input
flabel metal3 s 15540 17688 16000 17808 0 FreeSans 480 0 0 0 W6END[11]
port 192 nsew signal input
flabel metal3 s 15540 14968 16000 15088 0 FreeSans 480 0 0 0 W6END[1]
port 193 nsew signal input
flabel metal3 s 15540 15240 16000 15360 0 FreeSans 480 0 0 0 W6END[2]
port 194 nsew signal input
flabel metal3 s 15540 15512 16000 15632 0 FreeSans 480 0 0 0 W6END[3]
port 195 nsew signal input
flabel metal3 s 15540 15784 16000 15904 0 FreeSans 480 0 0 0 W6END[4]
port 196 nsew signal input
flabel metal3 s 15540 16056 16000 16176 0 FreeSans 480 0 0 0 W6END[5]
port 197 nsew signal input
flabel metal3 s 15540 16328 16000 16448 0 FreeSans 480 0 0 0 W6END[6]
port 198 nsew signal input
flabel metal3 s 15540 16600 16000 16720 0 FreeSans 480 0 0 0 W6END[7]
port 199 nsew signal input
flabel metal3 s 15540 16872 16000 16992 0 FreeSans 480 0 0 0 W6END[8]
port 200 nsew signal input
flabel metal3 s 15540 17144 16000 17264 0 FreeSans 480 0 0 0 W6END[9]
port 201 nsew signal input
flabel metal3 s 15540 10344 16000 10464 0 FreeSans 480 0 0 0 WW4END[0]
port 202 nsew signal input
flabel metal3 s 15540 13064 16000 13184 0 FreeSans 480 0 0 0 WW4END[10]
port 203 nsew signal input
flabel metal3 s 15540 13336 16000 13456 0 FreeSans 480 0 0 0 WW4END[11]
port 204 nsew signal input
flabel metal3 s 15540 13608 16000 13728 0 FreeSans 480 0 0 0 WW4END[12]
port 205 nsew signal input
flabel metal3 s 15540 13880 16000 14000 0 FreeSans 480 0 0 0 WW4END[13]
port 206 nsew signal input
flabel metal3 s 15540 14152 16000 14272 0 FreeSans 480 0 0 0 WW4END[14]
port 207 nsew signal input
flabel metal3 s 15540 14424 16000 14544 0 FreeSans 480 0 0 0 WW4END[15]
port 208 nsew signal input
flabel metal3 s 15540 10616 16000 10736 0 FreeSans 480 0 0 0 WW4END[1]
port 209 nsew signal input
flabel metal3 s 15540 10888 16000 11008 0 FreeSans 480 0 0 0 WW4END[2]
port 210 nsew signal input
flabel metal3 s 15540 11160 16000 11280 0 FreeSans 480 0 0 0 WW4END[3]
port 211 nsew signal input
flabel metal3 s 15540 11432 16000 11552 0 FreeSans 480 0 0 0 WW4END[4]
port 212 nsew signal input
flabel metal3 s 15540 11704 16000 11824 0 FreeSans 480 0 0 0 WW4END[5]
port 213 nsew signal input
flabel metal3 s 15540 11976 16000 12096 0 FreeSans 480 0 0 0 WW4END[6]
port 214 nsew signal input
flabel metal3 s 15540 12248 16000 12368 0 FreeSans 480 0 0 0 WW4END[7]
port 215 nsew signal input
flabel metal3 s 15540 12520 16000 12640 0 FreeSans 480 0 0 0 WW4END[8]
port 216 nsew signal input
flabel metal3 s 15540 12792 16000 12912 0 FreeSans 480 0 0 0 WW4END[9]
port 217 nsew signal input
rlabel via1 7900 43520 7900 43520 0 VGND
rlabel metal1 7820 42976 7820 42976 0 VPWR
rlabel metal2 2162 10812 2162 10812 0 A_I
rlabel metal3 498 11220 498 11220 0 A_I_top
rlabel metal1 8740 21114 8740 21114 0 A_O
rlabel metal2 2806 9809 2806 9809 0 A_O_top
rlabel metal1 6394 20842 6394 20842 0 A_Q
rlabel metal2 2622 8772 2622 8772 0 A_T
rlabel metal3 498 10404 498 10404 0 A_T_top
rlabel metal3 498 12036 498 12036 0 A_config_C_bit0
rlabel metal3 498 12852 498 12852 0 A_config_C_bit1
rlabel metal3 866 13668 866 13668 0 A_config_C_bit2
rlabel metal3 498 14484 498 14484 0 A_config_C_bit3
rlabel metal1 2254 5644 2254 5644 0 B_I
rlabel metal3 866 5508 866 5508 0 B_I_top
rlabel metal1 7038 19924 7038 19924 0 B_O
rlabel metal3 452 3876 452 3876 0 B_O_top
rlabel metal2 8326 19958 8326 19958 0 B_Q
rlabel metal2 4738 7548 4738 7548 0 B_T
rlabel metal3 498 4692 498 4692 0 B_T_top
rlabel metal3 498 6324 498 6324 0 B_config_C_bit0
rlabel metal3 498 7140 498 7140 0 B_config_C_bit1
rlabel metal3 475 7956 475 7956 0 B_config_C_bit2
rlabel metal3 498 8772 498 8772 0 B_config_C_bit3
rlabel metal1 2300 12206 2300 12206 0 ConfigBits\[0\]
rlabel metal2 9614 10030 9614 10030 0 ConfigBits\[100\]
rlabel metal1 10500 9010 10500 9010 0 ConfigBits\[101\]
rlabel metal1 10902 10778 10902 10778 0 ConfigBits\[102\]
rlabel metal2 11730 10132 11730 10132 0 ConfigBits\[103\]
rlabel metal1 7728 7310 7728 7310 0 ConfigBits\[104\]
rlabel metal2 8418 6596 8418 6596 0 ConfigBits\[105\]
rlabel metal1 6164 8466 6164 8466 0 ConfigBits\[106\]
rlabel metal2 9614 6511 9614 6511 0 ConfigBits\[107\]
rlabel metal2 10534 5814 10534 5814 0 ConfigBits\[108\]
rlabel metal1 11408 4794 11408 4794 0 ConfigBits\[109\]
rlabel metal1 7636 19346 7636 19346 0 ConfigBits\[10\]
rlabel metal2 11822 5508 11822 5508 0 ConfigBits\[110\]
rlabel metal1 6394 11186 6394 11186 0 ConfigBits\[111\]
rlabel metal2 7222 11594 7222 11594 0 ConfigBits\[112\]
rlabel metal2 5658 11050 5658 11050 0 ConfigBits\[113\]
rlabel metal1 11178 20298 11178 20298 0 ConfigBits\[11\]
rlabel metal2 7498 17306 7498 17306 0 ConfigBits\[12\]
rlabel metal1 7912 16762 7912 16762 0 ConfigBits\[13\]
rlabel metal1 9890 16728 9890 16728 0 ConfigBits\[14\]
rlabel metal1 10258 16218 10258 16218 0 ConfigBits\[15\]
rlabel metal1 8602 14926 8602 14926 0 ConfigBits\[16\]
rlabel metal2 9338 15164 9338 15164 0 ConfigBits\[17\]
rlabel metal1 12788 16218 12788 16218 0 ConfigBits\[18\]
rlabel metal1 13386 16626 13386 16626 0 ConfigBits\[19\]
rlabel metal1 2300 13294 2300 13294 0 ConfigBits\[1\]
rlabel metal1 10672 14042 10672 14042 0 ConfigBits\[20\]
rlabel metal2 11362 14586 11362 14586 0 ConfigBits\[21\]
rlabel metal1 11730 12410 11730 12410 0 ConfigBits\[22\]
rlabel metal2 12466 13532 12466 13532 0 ConfigBits\[23\]
rlabel metal1 9062 19278 9062 19278 0 ConfigBits\[24\]
rlabel metal1 9890 18938 9890 18938 0 ConfigBits\[25\]
rlabel metal1 12696 17850 12696 17850 0 ConfigBits\[26\]
rlabel metal2 13570 18428 13570 18428 0 ConfigBits\[27\]
rlabel metal2 13018 21658 13018 21658 0 ConfigBits\[28\]
rlabel metal2 13524 22236 13524 22236 0 ConfigBits\[29\]
rlabel metal1 2300 14994 2300 14994 0 ConfigBits\[2\]
rlabel metal2 10120 21454 10120 21454 0 ConfigBits\[30\]
rlabel metal2 10718 23596 10718 23596 0 ConfigBits\[31\]
rlabel metal1 6210 14518 6210 14518 0 ConfigBits\[32\]
rlabel metal1 7222 14450 7222 14450 0 ConfigBits\[33\]
rlabel metal2 12742 19958 12742 19958 0 ConfigBits\[34\]
rlabel metal1 13432 19482 13432 19482 0 ConfigBits\[35\]
rlabel metal1 7498 13498 7498 13498 0 ConfigBits\[36\]
rlabel metal1 8234 12954 8234 12954 0 ConfigBits\[37\]
rlabel metal1 12972 10574 12972 10574 0 ConfigBits\[38\]
rlabel metal2 13570 9588 13570 9588 0 ConfigBits\[39\]
rlabel metal1 2208 17170 2208 17170 0 ConfigBits\[3\]
rlabel metal1 9062 13430 9062 13430 0 ConfigBits\[40\]
rlabel metal1 10028 12954 10028 12954 0 ConfigBits\[41\]
rlabel metal1 13064 7514 13064 7514 0 ConfigBits\[42\]
rlabel metal1 13708 8058 13708 8058 0 ConfigBits\[43\]
rlabel metal1 11178 23222 11178 23222 0 ConfigBits\[44\]
rlabel metal2 11822 23562 11822 23562 0 ConfigBits\[45\]
rlabel metal1 12972 23630 12972 23630 0 ConfigBits\[46\]
rlabel metal1 13616 23290 13616 23290 0 ConfigBits\[47\]
rlabel metal1 5980 24310 5980 24310 0 ConfigBits\[48\]
rlabel metal1 7222 24242 7222 24242 0 ConfigBits\[49\]
rlabel metal1 2484 5678 2484 5678 0 ConfigBits\[4\]
rlabel metal1 9246 27914 9246 27914 0 ConfigBits\[50\]
rlabel metal2 10166 28492 10166 28492 0 ConfigBits\[51\]
rlabel metal2 8142 11254 8142 11254 0 ConfigBits\[52\]
rlabel metal1 8602 10710 8602 10710 0 ConfigBits\[53\]
rlabel metal2 13064 12682 13064 12682 0 ConfigBits\[54\]
rlabel metal1 13616 11866 13616 11866 0 ConfigBits\[55\]
rlabel metal1 10396 15606 10396 15606 0 ConfigBits\[56\]
rlabel metal1 11454 15538 11454 15538 0 ConfigBits\[57\]
rlabel metal2 13018 15130 13018 15130 0 ConfigBits\[58\]
rlabel metal2 13570 14756 13570 14756 0 ConfigBits\[59\]
rlabel metal1 2300 7378 2300 7378 0 ConfigBits\[5\]
rlabel metal1 12512 25466 12512 25466 0 ConfigBits\[60\]
rlabel metal1 13524 24922 13524 24922 0 ConfigBits\[61\]
rlabel metal1 6532 26486 6532 26486 0 ConfigBits\[62\]
rlabel metal1 7544 25466 7544 25466 0 ConfigBits\[63\]
rlabel metal1 11040 26486 11040 26486 0 ConfigBits\[64\]
rlabel metal2 11730 26826 11730 26826 0 ConfigBits\[65\]
rlabel metal1 12880 26894 12880 26894 0 ConfigBits\[66\]
rlabel metal1 13616 26554 13616 26554 0 ConfigBits\[67\]
rlabel metal1 6486 26826 6486 26826 0 ConfigBits\[68\]
rlabel metal2 7590 27404 7590 27404 0 ConfigBits\[69\]
rlabel metal2 2530 9418 2530 9418 0 ConfigBits\[6\]
rlabel metal1 7636 27982 7636 27982 0 ConfigBits\[70\]
rlabel metal1 8372 27574 8372 27574 0 ConfigBits\[71\]
rlabel metal1 13662 5542 13662 5542 0 ConfigBits\[72\]
rlabel metal1 13570 5338 13570 5338 0 ConfigBits\[73\]
rlabel metal1 12183 6834 12183 6834 0 ConfigBits\[74\]
rlabel metal1 13524 4794 13524 4794 0 ConfigBits\[75\]
rlabel metal1 8786 25398 8786 25398 0 ConfigBits\[76\]
rlabel metal2 9706 25449 9706 25449 0 ConfigBits\[77\]
rlabel metal1 12880 27982 12880 27982 0 ConfigBits\[78\]
rlabel metal2 13570 28764 13570 28764 0 ConfigBits\[79\]
rlabel metal1 2346 8942 2346 8942 0 ConfigBits\[7\]
rlabel metal1 8142 20570 8142 20570 0 ConfigBits\[80\]
rlabel metal1 8648 21862 8648 21862 0 ConfigBits\[81\]
rlabel metal1 10120 22134 10120 22134 0 ConfigBits\[82\]
rlabel metal1 10856 21114 10856 21114 0 ConfigBits\[83\]
rlabel metal1 7958 22746 7958 22746 0 ConfigBits\[84\]
rlabel metal1 8602 23222 8602 23222 0 ConfigBits\[85\]
rlabel metal1 11224 28662 11224 28662 0 ConfigBits\[86\]
rlabel metal2 12098 29002 12098 29002 0 ConfigBits\[87\]
rlabel metal1 9660 30158 9660 30158 0 ConfigBits\[88\]
rlabel metal2 10212 32198 10212 32198 0 ConfigBits\[89\]
rlabel metal1 10534 17612 10534 17612 0 ConfigBits\[8\]
rlabel metal2 12466 31110 12466 31110 0 ConfigBits\[90\]
rlabel metal2 12972 32198 12972 32198 0 ConfigBits\[91\]
rlabel metal2 5934 21148 5934 21148 0 ConfigBits\[92\]
rlabel metal1 6486 21862 6486 21862 0 ConfigBits\[93\]
rlabel metal2 12282 30362 12282 30362 0 ConfigBits\[94\]
rlabel metal2 13110 32436 13110 32436 0 ConfigBits\[95\]
rlabel metal1 8510 30906 8510 30906 0 ConfigBits\[96\]
rlabel metal1 8878 31654 8878 31654 0 ConfigBits\[97\]
rlabel metal2 12512 32810 12512 32810 0 ConfigBits\[98\]
rlabel metal2 12558 33932 12558 33932 0 ConfigBits\[99\]
rlabel metal1 6486 18700 6486 18700 0 ConfigBits\[9\]
rlabel metal3 14797 18020 14797 18020 0 E1BEG[0]
rlabel metal1 14720 16218 14720 16218 0 E1BEG[1]
rlabel metal3 15280 18564 15280 18564 0 E1BEG[2]
rlabel metal1 11822 17850 11822 17850 0 E1BEG[3]
rlabel metal3 14774 19108 14774 19108 0 E2BEG[0]
rlabel metal2 11270 19329 11270 19329 0 E2BEG[1]
rlabel metal3 15165 19652 15165 19652 0 E2BEG[2]
rlabel metal3 14084 19924 14084 19924 0 E2BEG[3]
rlabel metal2 14122 19839 14122 19839 0 E2BEG[4]
rlabel metal3 14797 20468 14797 20468 0 E2BEG[5]
rlabel metal3 15280 20740 15280 20740 0 E2BEG[6]
rlabel metal3 14820 21012 14820 21012 0 E2BEG[7]
rlabel metal3 14774 21284 14774 21284 0 E2BEGb[0]
rlabel metal1 13708 20570 13708 20570 0 E2BEGb[1]
rlabel metal3 15418 21828 15418 21828 0 E2BEGb[2]
rlabel metal3 14682 22100 14682 22100 0 E2BEGb[3]
rlabel metal1 13708 22066 13708 22066 0 E2BEGb[4]
rlabel metal1 14122 20910 14122 20910 0 E2BEGb[5]
rlabel metal1 14536 22746 14536 22746 0 E2BEGb[6]
rlabel metal3 14636 23188 14636 23188 0 E2BEGb[7]
rlabel metal3 15165 27812 15165 27812 0 E6BEG[0]
rlabel metal3 15165 30532 15165 30532 0 E6BEG[10]
rlabel metal1 13432 32946 13432 32946 0 E6BEG[11]
rlabel metal3 14912 28084 14912 28084 0 E6BEG[1]
rlabel metal1 13478 31790 13478 31790 0 E6BEG[2]
rlabel metal1 14030 31994 14030 31994 0 E6BEG[3]
rlabel metal3 14728 28900 14728 28900 0 E6BEG[4]
rlabel metal2 11638 30141 11638 30141 0 E6BEG[5]
rlabel metal3 15165 29444 15165 29444 0 E6BEG[6]
rlabel metal1 14536 33286 14536 33286 0 E6BEG[7]
rlabel metal1 14122 32810 14122 32810 0 E6BEG[8]
rlabel metal1 14582 34578 14582 34578 0 E6BEG[9]
rlabel metal3 14682 23460 14682 23460 0 EE4BEG[0]
rlabel metal3 15280 26180 15280 26180 0 EE4BEG[10]
rlabel metal3 14774 26452 14774 26452 0 EE4BEG[11]
rlabel metal3 14728 26724 14728 26724 0 EE4BEG[12]
rlabel metal2 12098 27421 12098 27421 0 EE4BEG[13]
rlabel metal1 14674 32198 14674 32198 0 EE4BEG[14]
rlabel metal3 15464 27540 15464 27540 0 EE4BEG[15]
rlabel metal3 14912 23732 14912 23732 0 EE4BEG[1]
rlabel metal3 15165 24004 15165 24004 0 EE4BEG[2]
rlabel metal3 14774 24276 14774 24276 0 EE4BEG[3]
rlabel metal3 14498 24548 14498 24548 0 EE4BEG[4]
rlabel metal3 14774 24820 14774 24820 0 EE4BEG[5]
rlabel metal3 15165 25092 15165 25092 0 EE4BEG[6]
rlabel metal3 13716 25364 13716 25364 0 EE4BEG[7]
rlabel metal3 14682 25636 14682 25636 0 EE4BEG[8]
rlabel metal3 14636 25908 14636 25908 0 EE4BEG[9]
rlabel metal3 452 15300 452 15300 0 FrameData[0]
rlabel metal3 452 23460 452 23460 0 FrameData[10]
rlabel metal3 452 24276 452 24276 0 FrameData[11]
rlabel metal3 452 25092 452 25092 0 FrameData[12]
rlabel metal3 475 25908 475 25908 0 FrameData[13]
rlabel metal3 452 26724 452 26724 0 FrameData[14]
rlabel metal3 774 27540 774 27540 0 FrameData[15]
rlabel metal3 452 28356 452 28356 0 FrameData[16]
rlabel metal3 452 29172 452 29172 0 FrameData[17]
rlabel metal3 452 29988 452 29988 0 FrameData[18]
rlabel metal3 452 30804 452 30804 0 FrameData[19]
rlabel metal3 452 16116 452 16116 0 FrameData[1]
rlabel metal3 774 31620 774 31620 0 FrameData[20]
rlabel metal3 452 32436 452 32436 0 FrameData[21]
rlabel metal3 452 33252 452 33252 0 FrameData[22]
rlabel metal3 475 34068 475 34068 0 FrameData[23]
rlabel metal3 452 34884 452 34884 0 FrameData[24]
rlabel metal3 820 35700 820 35700 0 FrameData[25]
rlabel metal3 452 36516 452 36516 0 FrameData[26]
rlabel metal3 452 37332 452 37332 0 FrameData[27]
rlabel metal3 452 38148 452 38148 0 FrameData[28]
rlabel metal3 452 38964 452 38964 0 FrameData[29]
rlabel metal3 452 16932 452 16932 0 FrameData[2]
rlabel metal3 820 39780 820 39780 0 FrameData[30]
rlabel metal3 452 40596 452 40596 0 FrameData[31]
rlabel metal3 475 17748 475 17748 0 FrameData[3]
rlabel metal3 452 18564 452 18564 0 FrameData[4]
rlabel metal3 452 19380 452 19380 0 FrameData[5]
rlabel metal3 452 20196 452 20196 0 FrameData[6]
rlabel metal3 452 21012 452 21012 0 FrameData[7]
rlabel metal3 452 21828 452 21828 0 FrameData[8]
rlabel metal3 452 22644 452 22644 0 FrameData[9]
rlabel metal3 14429 31076 14429 31076 0 FrameData_O[0]
rlabel metal3 15165 33796 15165 33796 0 FrameData_O[10]
rlabel metal2 11362 34323 11362 34323 0 FrameData_O[11]
rlabel metal3 14498 34340 14498 34340 0 FrameData_O[12]
rlabel metal3 14544 34612 14544 34612 0 FrameData_O[13]
rlabel metal3 15165 34884 15165 34884 0 FrameData_O[14]
rlabel metal3 14774 35156 14774 35156 0 FrameData_O[15]
rlabel metal3 14360 35428 14360 35428 0 FrameData_O[16]
rlabel metal3 14084 35700 14084 35700 0 FrameData_O[17]
rlabel metal3 15280 35972 15280 35972 0 FrameData_O[18]
rlabel metal3 14866 36244 14866 36244 0 FrameData_O[19]
rlabel metal3 14889 31348 14889 31348 0 FrameData_O[1]
rlabel metal3 14590 36516 14590 36516 0 FrameData_O[20]
rlabel metal3 14636 36788 14636 36788 0 FrameData_O[21]
rlabel metal3 15165 37060 15165 37060 0 FrameData_O[22]
rlabel metal3 14866 37332 14866 37332 0 FrameData_O[23]
rlabel metal3 14958 37604 14958 37604 0 FrameData_O[24]
rlabel metal3 14912 37876 14912 37876 0 FrameData_O[25]
rlabel metal3 15188 38148 15188 38148 0 FrameData_O[26]
rlabel metal3 14452 38420 14452 38420 0 FrameData_O[27]
rlabel metal3 14728 38692 14728 38692 0 FrameData_O[28]
rlabel metal3 14912 38964 14912 38964 0 FrameData_O[29]
rlabel metal3 15165 31620 15165 31620 0 FrameData_O[2]
rlabel metal3 15188 39236 15188 39236 0 FrameData_O[30]
rlabel metal3 14820 39508 14820 39508 0 FrameData_O[31]
rlabel metal3 14590 31892 14590 31892 0 FrameData_O[3]
rlabel metal3 14797 32164 14797 32164 0 FrameData_O[4]
rlabel metal3 14222 32436 14222 32436 0 FrameData_O[5]
rlabel metal3 15165 32708 15165 32708 0 FrameData_O[6]
rlabel metal3 14981 32980 14981 32980 0 FrameData_O[7]
rlabel metal3 14820 33252 14820 33252 0 FrameData_O[8]
rlabel metal3 14590 33524 14590 33524 0 FrameData_O[9]
rlabel metal1 13754 30668 13754 30668 0 FrameData_O_i\[0\]
rlabel via1 10902 33964 10902 33964 0 FrameData_O_i\[10\]
rlabel metal1 11178 33898 11178 33898 0 FrameData_O_i\[11\]
rlabel metal1 11086 33286 11086 33286 0 FrameData_O_i\[12\]
rlabel metal1 10810 35700 10810 35700 0 FrameData_O_i\[13\]
rlabel metal2 10442 34578 10442 34578 0 FrameData_O_i\[14\]
rlabel metal2 10626 34884 10626 34884 0 FrameData_O_i\[15\]
rlabel metal2 10902 35972 10902 35972 0 FrameData_O_i\[16\]
rlabel metal2 11822 35836 11822 35836 0 FrameData_O_i\[17\]
rlabel metal1 9982 35258 9982 35258 0 FrameData_O_i\[18\]
rlabel metal2 8970 35462 8970 35462 0 FrameData_O_i\[19\]
rlabel metal1 13800 32334 13800 32334 0 FrameData_O_i\[1\]
rlabel metal2 12466 36550 12466 36550 0 FrameData_O_i\[20\]
rlabel metal1 12098 36754 12098 36754 0 FrameData_O_i\[21\]
rlabel via1 11914 37213 11914 37213 0 FrameData_O_i\[22\]
rlabel metal2 12834 36975 12834 36975 0 FrameData_O_i\[23\]
rlabel metal1 12926 38896 12926 38896 0 FrameData_O_i\[24\]
rlabel metal1 12466 37944 12466 37944 0 FrameData_O_i\[25\]
rlabel metal2 10350 37638 10350 37638 0 FrameData_O_i\[26\]
rlabel metal1 12374 37808 12374 37808 0 FrameData_O_i\[27\]
rlabel metal1 12489 38318 12489 38318 0 FrameData_O_i\[28\]
rlabel metal1 12650 38964 12650 38964 0 FrameData_O_i\[29\]
rlabel metal1 10902 31790 10902 31790 0 FrameData_O_i\[2\]
rlabel metal1 8602 39440 8602 39440 0 FrameData_O_i\[30\]
rlabel metal1 9706 39440 9706 39440 0 FrameData_O_i\[31\]
rlabel metal2 11408 31756 11408 31756 0 FrameData_O_i\[3\]
rlabel metal1 10718 31824 10718 31824 0 FrameData_O_i\[4\]
rlabel metal1 10764 31926 10764 31926 0 FrameData_O_i\[5\]
rlabel metal1 10120 31994 10120 31994 0 FrameData_O_i\[6\]
rlabel metal1 10626 32810 10626 32810 0 FrameData_O_i\[7\]
rlabel metal2 12650 34476 12650 34476 0 FrameData_O_i\[8\]
rlabel metal1 10258 33490 10258 33490 0 FrameData_O_i\[9\]
rlabel metal2 1242 704 1242 704 0 FrameStrobe[0]
rlabel metal2 8602 704 8602 704 0 FrameStrobe[10]
rlabel metal2 9338 704 9338 704 0 FrameStrobe[11]
rlabel metal2 10074 704 10074 704 0 FrameStrobe[12]
rlabel metal2 10810 704 10810 704 0 FrameStrobe[13]
rlabel metal2 11546 704 11546 704 0 FrameStrobe[14]
rlabel metal2 12282 704 12282 704 0 FrameStrobe[15]
rlabel metal2 13018 143 13018 143 0 FrameStrobe[16]
rlabel metal2 13754 704 13754 704 0 FrameStrobe[17]
rlabel metal2 14345 68 14345 68 0 FrameStrobe[18]
rlabel metal2 15226 704 15226 704 0 FrameStrobe[19]
rlabel metal2 1978 1010 1978 1010 0 FrameStrobe[1]
rlabel metal2 2714 704 2714 704 0 FrameStrobe[2]
rlabel metal2 3641 68 3641 68 0 FrameStrobe[3]
rlabel metal2 4186 670 4186 670 0 FrameStrobe[4]
rlabel metal2 5021 68 5021 68 0 FrameStrobe[5]
rlabel metal2 5658 670 5658 670 0 FrameStrobe[6]
rlabel metal2 6295 68 6295 68 0 FrameStrobe[7]
rlabel metal2 7130 704 7130 704 0 FrameStrobe[8]
rlabel metal2 7866 143 7866 143 0 FrameStrobe[9]
rlabel metal2 1242 43785 1242 43785 0 FrameStrobe_O[0]
rlabel metal1 8878 43418 8878 43418 0 FrameStrobe_O[10]
rlabel metal1 9476 43418 9476 43418 0 FrameStrobe_O[11]
rlabel metal1 10212 43418 10212 43418 0 FrameStrobe_O[12]
rlabel metal2 10810 43972 10810 43972 0 FrameStrobe_O[13]
rlabel metal1 11684 43418 11684 43418 0 FrameStrobe_O[14]
rlabel metal2 12282 43972 12282 43972 0 FrameStrobe_O[15]
rlabel metal1 13156 43418 13156 43418 0 FrameStrobe_O[16]
rlabel metal2 13754 43428 13754 43428 0 FrameStrobe_O[17]
rlabel metal1 13892 42738 13892 42738 0 FrameStrobe_O[18]
rlabel metal1 14536 43418 14536 43418 0 FrameStrobe_O[19]
rlabel metal1 2116 43146 2116 43146 0 FrameStrobe_O[1]
rlabel metal2 2714 44193 2714 44193 0 FrameStrobe_O[2]
rlabel metal1 3726 43418 3726 43418 0 FrameStrobe_O[3]
rlabel metal2 4186 43972 4186 43972 0 FrameStrobe_O[4]
rlabel metal1 5060 43418 5060 43418 0 FrameStrobe_O[5]
rlabel metal1 5796 43418 5796 43418 0 FrameStrobe_O[6]
rlabel metal1 6532 43418 6532 43418 0 FrameStrobe_O[7]
rlabel metal1 7268 43418 7268 43418 0 FrameStrobe_O[8]
rlabel metal1 8096 43418 8096 43418 0 FrameStrobe_O[9]
rlabel metal2 1978 36550 1978 36550 0 FrameStrobe_O_i\[0\]
rlabel metal2 8694 2227 8694 2227 0 FrameStrobe_O_i\[10\]
rlabel metal3 9269 2516 9269 2516 0 FrameStrobe_O_i\[11\]
rlabel metal2 10166 2023 10166 2023 0 FrameStrobe_O_i\[12\]
rlabel metal3 10649 2652 10649 2652 0 FrameStrobe_O_i\[13\]
rlabel metal1 12742 1870 12742 1870 0 FrameStrobe_O_i\[14\]
rlabel metal1 12374 1768 12374 1768 0 FrameStrobe_O_i\[15\]
rlabel metal3 14421 41548 14421 41548 0 FrameStrobe_O_i\[16\]
rlabel metal1 14352 1870 14352 1870 0 FrameStrobe_O_i\[17\]
rlabel metal2 13432 2074 13432 2074 0 FrameStrobe_O_i\[18\]
rlabel metal3 11293 1292 11293 1292 0 FrameStrobe_O_i\[19\]
rlabel metal2 2162 36006 2162 36006 0 FrameStrobe_O_i\[1\]
rlabel metal2 2714 27268 2714 27268 0 FrameStrobe_O_i\[2\]
rlabel metal2 3266 21597 3266 21597 0 FrameStrobe_O_i\[3\]
rlabel metal2 4094 42500 4094 42500 0 FrameStrobe_O_i\[4\]
rlabel metal1 4876 42330 4876 42330 0 FrameStrobe_O_i\[5\]
rlabel metal1 5658 34714 5658 34714 0 FrameStrobe_O_i\[6\]
rlabel metal1 6624 2074 6624 2074 0 FrameStrobe_O_i\[7\]
rlabel metal2 7222 2295 7222 2295 0 FrameStrobe_O_i\[8\]
rlabel metal1 7728 2074 7728 2074 0 FrameStrobe_O_i\[9\]
rlabel metal1 10994 9418 10994 9418 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out0
rlabel metal1 10672 10234 10672 10234 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out1
rlabel metal1 12190 10234 12190 10234 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out2
rlabel metal1 11454 9146 11454 9146 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_A_I/cus_mux41_buf_out3
rlabel metal1 10994 5746 10994 5746 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out0
rlabel metal1 10672 5746 10672 5746 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out1
rlabel via1 11650 5746 11650 5746 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out2
rlabel metal2 11546 6800 11546 6800 0 Inst_W_IO_switch_matrix/inst_cus_mux161_buf_B_I/cus_mux41_buf_out3
rlabel metal2 10948 16966 10948 16966 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN\[0\]
rlabel metal1 10718 17714 10718 17714 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/AIN\[1\]
rlabel metal1 11316 17102 11316 17102 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_0_
rlabel metal1 11822 17068 11822 17068 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG0/_1_
rlabel metal1 7176 18258 7176 18258 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN\[0\]
rlabel metal1 6624 18258 6624 18258 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/AIN\[1\]
rlabel metal2 6946 18564 6946 18564 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_0_
rlabel metal1 6716 18394 6716 18394 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG1/_1_
rlabel metal1 7544 18734 7544 18734 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN\[0\]
rlabel metal1 7958 19380 7958 19380 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/AIN\[1\]
rlabel metal1 7314 18666 7314 18666 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_0_
rlabel metal1 7314 18870 7314 18870 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG2/_1_
rlabel metal2 10718 20570 10718 20570 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN\[0\]
rlabel metal1 11730 20468 11730 20468 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/AIN\[1\]
rlabel metal1 10948 19890 10948 19890 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_0_
rlabel metal1 11454 19890 11454 19890 0 Inst_W_IO_switch_matrix/inst_cus_mux21_E1BEG3/_1_
rlabel metal1 6578 8058 6578 8058 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN\[0\]
rlabel metal1 6946 7990 6946 7990 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/AIN\[1\]
rlabel metal1 6670 8330 6670 8330 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_0_
rlabel metal1 6900 8398 6900 8398 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux21_inst/_1_
rlabel metal1 6670 7854 6670 7854 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out0
rlabel metal1 7958 7514 7958 7514 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_A_T/cus_mux41_buf_out1
rlabel metal1 6256 9894 6256 9894 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN\[0\]
rlabel metal1 6486 10166 6486 10166 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/AIN\[1\]
rlabel metal2 5750 10336 5750 10336 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_0_
rlabel metal1 6348 10098 6348 10098 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux21_inst/_1_
rlabel metal1 6394 10030 6394 10030 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out0
rlabel metal2 6578 10081 6578 10081 0 Inst_W_IO_switch_matrix/inst_cus_mux81_buf_B_T/cus_mux41_buf_out1
rlabel metal3 1495 41412 1495 41412 0 UserCLK
rlabel metal1 1932 43418 1932 43418 0 UserCLKo
rlabel metal3 14728 4964 14728 4964 0 W1END[0]
rlabel metal3 15234 5236 15234 5236 0 W1END[1]
rlabel metal3 15165 5508 15165 5508 0 W1END[2]
rlabel metal3 15073 5780 15073 5780 0 W1END[3]
rlabel metal3 14797 8228 14797 8228 0 W2END[0]
rlabel metal3 14866 8500 14866 8500 0 W2END[1]
rlabel metal3 15188 8772 15188 8772 0 W2END[2]
rlabel metal1 10994 8466 10994 8466 0 W2END[3]
rlabel metal3 14774 9316 14774 9316 0 W2END[4]
rlabel metal3 15418 9588 15418 9588 0 W2END[5]
rlabel metal3 15165 9860 15165 9860 0 W2END[6]
rlabel metal3 14774 10132 14774 10132 0 W2END[7]
rlabel metal3 14797 6052 14797 6052 0 W2MID[0]
rlabel metal2 12282 5372 12282 5372 0 W2MID[1]
rlabel metal3 15165 6596 15165 6596 0 W2MID[2]
rlabel metal2 9476 7242 9476 7242 0 W2MID[3]
rlabel metal3 14797 7140 14797 7140 0 W2MID[4]
rlabel metal2 11730 7973 11730 7973 0 W2MID[5]
rlabel metal3 15188 7684 15188 7684 0 W2MID[6]
rlabel metal3 14889 7956 14889 7956 0 W2MID[7]
rlabel metal3 14958 14756 14958 14756 0 W6END[0]
rlabel metal3 15165 17476 15165 17476 0 W6END[10]
rlabel metal2 10534 17459 10534 17459 0 W6END[11]
rlabel metal3 14728 15028 14728 15028 0 W6END[1]
rlabel metal3 15165 15300 15165 15300 0 W6END[2]
rlabel metal3 14682 15572 14682 15572 0 W6END[3]
rlabel metal3 14314 15844 14314 15844 0 W6END[4]
rlabel metal3 15096 16116 15096 16116 0 W6END[5]
rlabel metal3 15280 16388 15280 16388 0 W6END[6]
rlabel metal3 14774 16660 14774 16660 0 W6END[7]
rlabel metal3 14797 16932 14797 16932 0 W6END[8]
rlabel metal3 15280 17204 15280 17204 0 W6END[9]
rlabel metal1 13478 10098 13478 10098 0 WW4END[0]
rlabel metal3 15165 13124 15165 13124 0 WW4END[10]
rlabel metal3 14774 13396 14774 13396 0 WW4END[11]
rlabel metal3 14958 13668 14958 13668 0 WW4END[12]
rlabel metal3 14820 13940 14820 13940 0 WW4END[13]
rlabel metal3 15280 14212 15280 14212 0 WW4END[14]
rlabel metal3 14774 14484 14774 14484 0 WW4END[15]
rlabel metal1 13386 7242 13386 7242 0 WW4END[1]
rlabel metal3 15165 10948 15165 10948 0 WW4END[2]
rlabel metal2 11822 10931 11822 10931 0 WW4END[3]
rlabel metal3 14797 11492 14797 11492 0 WW4END[4]
rlabel metal1 11730 11764 11730 11764 0 WW4END[5]
rlabel metal3 15165 12036 15165 12036 0 WW4END[6]
rlabel metal1 11362 12682 11362 12682 0 WW4END[7]
rlabel metal3 14636 12580 14636 12580 0 WW4END[8]
rlabel metal3 13946 12852 13946 12852 0 WW4END[9]
rlabel metal1 3900 18258 3900 18258 0 net1
rlabel metal2 2024 17476 2024 17476 0 net10
rlabel metal2 9706 16813 9706 16813 0 net100
rlabel via1 13455 18258 13455 18258 0 net101
rlabel metal1 9856 13362 9856 13362 0 net102
rlabel metal1 1748 10778 1748 10778 0 net103
rlabel metal1 2438 8874 2438 8874 0 net104
rlabel metal1 1748 12138 1748 12138 0 net105
rlabel metal1 1748 13226 1748 13226 0 net106
rlabel metal1 1518 14008 1518 14008 0 net107
rlabel metal2 1518 16014 1518 16014 0 net108
rlabel metal1 1794 5610 1794 5610 0 net109
rlabel metal1 1885 17646 1885 17646 0 net11
rlabel metal1 1794 5270 1794 5270 0 net110
rlabel metal1 1932 5882 1932 5882 0 net111
rlabel metal1 1748 7446 1748 7446 0 net112
rlabel metal1 1932 8534 1932 8534 0 net113
rlabel metal1 1794 8874 1794 8874 0 net114
rlabel metal1 11960 17238 11960 17238 0 net115
rlabel metal1 8142 18360 8142 18360 0 net116
rlabel metal1 10028 18326 10028 18326 0 net117
rlabel metal1 11362 17646 11362 17646 0 net118
rlabel metal2 8694 17952 8694 17952 0 net119
rlabel viali 6385 13264 6385 13264 0 net12
rlabel metal1 11362 16762 11362 16762 0 net120
rlabel metal1 10166 15130 10166 15130 0 net121
rlabel metal1 13892 16762 13892 16762 0 net122
rlabel metal1 14030 19346 14030 19346 0 net123
rlabel metal1 13294 13498 13294 13498 0 net124
rlabel metal2 12558 19992 12558 19992 0 net125
rlabel metal1 14076 18190 14076 18190 0 net126
rlabel metal1 14582 21182 14582 21182 0 net127
rlabel metal1 12282 20502 12282 20502 0 net128
rlabel metal1 7866 14586 7866 14586 0 net129
rlabel metal1 8648 35054 8648 35054 0 net13
rlabel metal2 13938 20723 13938 20723 0 net130
rlabel via3 13869 20740 13869 20740 0 net131
rlabel metal2 14168 20332 14168 20332 0 net132
rlabel metal4 15180 18156 15180 18156 0 net133
rlabel metal1 14214 20332 14214 20332 0 net134
rlabel metal1 11132 25466 11132 25466 0 net135
rlabel metal1 10442 32334 10442 32334 0 net136
rlabel metal1 13202 32810 13202 32810 0 net137
rlabel metal2 14214 29750 14214 29750 0 net138
rlabel metal2 13984 26860 13984 26860 0 net139
rlabel metal1 12742 30056 12742 30056 0 net14
rlabel metal2 11638 22559 11638 22559 0 net140
rlabel metal2 9246 26180 9246 26180 0 net141
rlabel metal1 13018 28662 13018 28662 0 net142
rlabel metal1 11316 30294 11316 30294 0 net143
rlabel metal1 13708 30838 13708 30838 0 net144
rlabel metal2 7268 26180 7268 26180 0 net145
rlabel metal2 13846 32436 13846 32436 0 net146
rlabel metal1 12788 23290 12788 23290 0 net147
rlabel metal2 12650 27200 12650 27200 0 net148
rlabel metal1 13317 27098 13317 27098 0 net149
rlabel via2 12742 11101 12742 11101 0 net15
rlabel metal2 8234 27268 8234 27268 0 net150
rlabel metal1 11638 28152 11638 28152 0 net151
rlabel metal1 14490 32402 14490 32402 0 net152
rlabel metal1 14444 6630 14444 6630 0 net153
rlabel metal2 14214 23936 14214 23936 0 net154
rlabel metal1 9062 24378 9062 24378 0 net155
rlabel metal1 11362 23766 11362 23766 0 net156
rlabel metal1 5704 27574 5704 27574 0 net157
rlabel metal1 15502 21556 15502 21556 0 net158
rlabel metal1 12972 15674 12972 15674 0 net159
rlabel viali 1693 9584 1693 9584 0 net16
rlabel metal1 14720 15130 14720 15130 0 net160
rlabel metal1 13938 26010 13938 26010 0 net161
rlabel metal2 10074 27200 10074 27200 0 net162
rlabel metal1 10166 32504 10166 32504 0 net163
rlabel metal2 12558 34884 12558 34884 0 net164
rlabel metal2 10994 34374 10994 34374 0 net165
rlabel metal1 11960 34170 11960 34170 0 net166
rlabel metal2 10626 36312 10626 36312 0 net167
rlabel metal2 13386 35666 13386 35666 0 net168
rlabel metal1 10902 35258 10902 35258 0 net169
rlabel metal2 12742 37077 12742 37077 0 net17
rlabel metal1 12627 36142 12627 36142 0 net170
rlabel metal1 11960 35530 11960 35530 0 net171
rlabel metal1 13202 36720 13202 36720 0 net172
rlabel metal2 12466 35751 12466 35751 0 net173
rlabel metal1 13340 32538 13340 32538 0 net174
rlabel metal2 13570 37026 13570 37026 0 net175
rlabel metal1 13616 37910 13616 37910 0 net176
rlabel metal1 13018 37264 13018 37264 0 net177
rlabel metal1 12742 37876 12742 37876 0 net178
rlabel metal1 13156 37910 13156 37910 0 net179
rlabel metal1 1610 34680 1610 34680 0 net18
rlabel metal1 12926 38284 12926 38284 0 net180
rlabel metal1 12834 37706 12834 37706 0 net181
rlabel metal2 12466 38403 12466 38403 0 net182
rlabel metal2 13662 38726 13662 38726 0 net183
rlabel metal1 12696 39066 12696 39066 0 net184
rlabel metal2 10810 32402 10810 32402 0 net185
rlabel metal1 8418 39304 8418 39304 0 net186
rlabel metal2 13846 39814 13846 39814 0 net187
rlabel metal2 13570 33626 13570 33626 0 net188
rlabel metal1 11454 31858 11454 31858 0 net189
rlabel metal2 12742 35904 12742 35904 0 net19
rlabel metal1 12466 33864 12466 33864 0 net190
rlabel metal1 13110 32504 13110 32504 0 net191
rlabel via1 13570 33099 13570 33099 0 net192
rlabel metal2 11270 34408 11270 34408 0 net193
rlabel metal1 13202 33592 13202 33592 0 net194
rlabel metal2 1794 39950 1794 39950 0 net195
rlabel metal1 8740 42874 8740 42874 0 net196
rlabel metal2 9246 43078 9246 43078 0 net197
rlabel metal1 10028 42874 10028 42874 0 net198
rlabel metal1 10856 42874 10856 42874 0 net199
rlabel via1 4917 19754 4917 19754 0 net2
rlabel metal2 12650 37638 12650 37638 0 net20
rlabel metal1 11546 42874 11546 42874 0 net200
rlabel metal1 12328 42874 12328 42874 0 net201
rlabel metal1 13386 42874 13386 42874 0 net202
rlabel metal1 13708 41786 13708 41786 0 net203
rlabel metal1 13156 41786 13156 41786 0 net204
rlabel metal1 13478 42330 13478 42330 0 net205
rlabel metal1 2024 42330 2024 42330 0 net206
rlabel metal1 2898 43282 2898 43282 0 net207
rlabel metal1 3542 42874 3542 42874 0 net208
rlabel metal1 4232 42874 4232 42874 0 net209
rlabel metal3 7015 20740 7015 20740 0 net21
rlabel metal1 4922 42874 4922 42874 0 net210
rlabel metal2 5658 43282 5658 43282 0 net211
rlabel metal1 6394 42874 6394 42874 0 net212
rlabel metal1 7130 42874 7130 42874 0 net213
rlabel metal1 7866 42874 7866 42874 0 net214
rlabel metal1 3036 42874 3036 42874 0 net215
rlabel viali 8269 7378 8269 7378 0 net216
rlabel metal1 7176 10642 7176 10642 0 net217
rlabel metal1 8050 7310 8050 7310 0 net218
rlabel metal1 7130 10778 7130 10778 0 net219
rlabel metal1 8325 16558 8325 16558 0 net22
rlabel metal1 8861 17170 8861 17170 0 net23
rlabel metal2 2530 19584 2530 19584 0 net24
rlabel metal1 8372 31450 8372 31450 0 net25
rlabel metal1 7083 16082 7083 16082 0 net26
rlabel metal1 8924 39406 8924 39406 0 net27
rlabel metal1 9476 30362 9476 30362 0 net28
rlabel metal2 5888 21420 5888 21420 0 net29
rlabel metal1 11299 16082 11299 16082 0 net3
rlabel metal1 1656 20026 1656 20026 0 net30
rlabel metal1 9199 19822 9199 19822 0 net31
rlabel metal1 8907 18734 8907 18734 0 net32
rlabel metal2 2346 19465 2346 19465 0 net33
rlabel metal1 13109 18734 13109 18734 0 net34
rlabel metal2 2576 5678 2576 5678 0 net35
rlabel metal1 8786 1530 8786 1530 0 net36
rlabel metal1 9338 1530 9338 1530 0 net37
rlabel metal1 10120 1530 10120 1530 0 net38
rlabel metal1 10856 1530 10856 1530 0 net39
rlabel metal3 11431 33932 11431 33932 0 net4
rlabel metal2 11638 1734 11638 1734 0 net40
rlabel metal1 12328 1530 12328 1530 0 net41
rlabel metal2 13110 1734 13110 1734 0 net42
rlabel metal1 13570 1530 13570 1530 0 net43
rlabel metal1 13708 2006 13708 2006 0 net44
rlabel metal1 13294 1258 13294 1258 0 net45
rlabel metal1 5980 2006 5980 2006 0 net46
rlabel metal2 7498 19652 7498 19652 0 net47
rlabel metal1 1426 6154 1426 6154 0 net48
rlabel via2 4646 1309 4646 1309 0 net49
rlabel via1 12741 24786 12741 24786 0 net5
rlabel metal1 5244 1326 5244 1326 0 net50
rlabel metal3 6601 1292 6601 1292 0 net51
rlabel metal1 6256 1530 6256 1530 0 net52
rlabel metal1 7222 1530 7222 1530 0 net53
rlabel metal1 7912 1530 7912 1530 0 net54
rlabel metal1 13202 3944 13202 3944 0 net55
rlabel metal1 7866 18768 7866 18768 0 net56
rlabel metal1 8188 18734 8188 18734 0 net57
rlabel metal1 14628 4046 14628 4046 0 net58
rlabel via1 7694 10030 7694 10030 0 net59
rlabel metal1 9199 24174 9199 24174 0 net6
rlabel metal1 12834 9010 12834 9010 0 net60
rlabel metal1 13892 9146 13892 9146 0 net61
rlabel metal1 9596 7344 9596 7344 0 net62
rlabel metal1 13202 19448 13202 19448 0 net63
rlabel via1 13455 12750 13455 12750 0 net64
rlabel metal1 13294 8568 13294 8568 0 net65
rlabel metal2 13018 19924 13018 19924 0 net66
rlabel metal1 13202 5848 13202 5848 0 net67
rlabel via2 12558 15011 12558 15011 0 net68
rlabel via1 10362 6290 10362 6290 0 net69
rlabel metal1 10211 25874 10211 25874 0 net7
rlabel metal2 9614 7854 9614 7854 0 net70
rlabel metal1 9200 10098 9200 10098 0 net71
rlabel metal2 13386 14484 13386 14484 0 net72
rlabel metal2 6854 9894 6854 9894 0 net73
rlabel metal2 7130 7905 7130 7905 0 net74
rlabel metal1 12972 9486 12972 9486 0 net75
rlabel metal2 13340 25874 13340 25874 0 net76
rlabel metal1 10396 16966 10396 16966 0 net77
rlabel metal1 7452 31314 7452 31314 0 net78
rlabel metal1 14582 13498 14582 13498 0 net79
rlabel metal1 1656 27098 1656 27098 0 net8
rlabel metal2 10580 21522 10580 21522 0 net80
rlabel metal1 13294 17646 13294 17646 0 net81
rlabel metal2 9062 14722 9062 14722 0 net82
rlabel metal2 12558 26656 12558 26656 0 net83
rlabel metal1 13938 17306 13938 17306 0 net84
rlabel metal1 12650 30362 12650 30362 0 net85
rlabel metal2 12558 16830 12558 16830 0 net86
rlabel metal1 13110 9962 13110 9962 0 net87
rlabel metal1 13202 13804 13202 13804 0 net88
rlabel metal1 8832 21318 8832 21318 0 net89
rlabel metal2 1610 26860 1610 26860 0 net9
rlabel metal1 12984 19890 12984 19890 0 net90
rlabel metal1 13294 11560 13294 11560 0 net91
rlabel metal1 10833 21454 10833 21454 0 net92
rlabel via2 13386 21437 13386 21437 0 net93
rlabel metal2 13662 7582 13662 7582 0 net94
rlabel metal1 11040 13294 11040 13294 0 net95
rlabel metal1 6164 13906 6164 13906 0 net96
rlabel metal1 12144 16626 12144 16626 0 net97
rlabel metal2 8142 17884 8142 17884 0 net98
rlabel metal1 9430 21454 9430 21454 0 net99
<< properties >>
string FIXED_BBOX 0 0 15700 44700
<< end >>
