magic
tech sky130A
magscale 1 2
timestamp 1733615472
<< obsli1 >>
rect 1104 1071 43516 89233
<< obsm1 >>
rect 14 76 44698 90024
<< metal2 >>
rect 5170 90540 5226 91000
rect 5446 90540 5502 91000
rect 5722 90540 5778 91000
rect 5998 90540 6054 91000
rect 6274 90540 6330 91000
rect 6550 90540 6606 91000
rect 6826 90540 6882 91000
rect 7102 90540 7158 91000
rect 7378 90540 7434 91000
rect 7654 90540 7710 91000
rect 7930 90540 7986 91000
rect 8206 90540 8262 91000
rect 8482 90540 8538 91000
rect 8758 90540 8814 91000
rect 9034 90540 9090 91000
rect 9310 90540 9366 91000
rect 9586 90540 9642 91000
rect 9862 90540 9918 91000
rect 10138 90540 10194 91000
rect 10414 90540 10470 91000
rect 10690 90540 10746 91000
rect 10966 90540 11022 91000
rect 11242 90540 11298 91000
rect 11518 90540 11574 91000
rect 11794 90540 11850 91000
rect 12070 90540 12126 91000
rect 12346 90540 12402 91000
rect 12622 90540 12678 91000
rect 12898 90540 12954 91000
rect 13174 90540 13230 91000
rect 13450 90540 13506 91000
rect 13726 90540 13782 91000
rect 14002 90540 14058 91000
rect 14278 90540 14334 91000
rect 14554 90540 14610 91000
rect 14830 90540 14886 91000
rect 15106 90540 15162 91000
rect 15382 90540 15438 91000
rect 15658 90540 15714 91000
rect 15934 90540 15990 91000
rect 16210 90540 16266 91000
rect 16486 90540 16542 91000
rect 16762 90540 16818 91000
rect 17038 90540 17094 91000
rect 17314 90540 17370 91000
rect 17590 90540 17646 91000
rect 17866 90540 17922 91000
rect 18142 90540 18198 91000
rect 18418 90540 18474 91000
rect 18694 90540 18750 91000
rect 18970 90540 19026 91000
rect 19246 90540 19302 91000
rect 19522 90540 19578 91000
rect 19798 90540 19854 91000
rect 20074 90540 20130 91000
rect 20350 90540 20406 91000
rect 20626 90540 20682 91000
rect 20902 90540 20958 91000
rect 21178 90540 21234 91000
rect 21454 90540 21510 91000
rect 21730 90540 21786 91000
rect 22006 90540 22062 91000
rect 22282 90540 22338 91000
rect 22558 90540 22614 91000
rect 22834 90540 22890 91000
rect 23110 90540 23166 91000
rect 23386 90540 23442 91000
rect 23662 90540 23718 91000
rect 23938 90540 23994 91000
rect 24214 90540 24270 91000
rect 24490 90540 24546 91000
rect 24766 90540 24822 91000
rect 25042 90540 25098 91000
rect 25318 90540 25374 91000
rect 25594 90540 25650 91000
rect 25870 90540 25926 91000
rect 26146 90540 26202 91000
rect 26422 90540 26478 91000
rect 26698 90540 26754 91000
rect 26974 90540 27030 91000
rect 27250 90540 27306 91000
rect 27526 90540 27582 91000
rect 27802 90540 27858 91000
rect 28078 90540 28134 91000
rect 28354 90540 28410 91000
rect 28630 90540 28686 91000
rect 28906 90540 28962 91000
rect 29182 90540 29238 91000
rect 29458 90540 29514 91000
rect 29734 90540 29790 91000
rect 30010 90540 30066 91000
rect 30286 90540 30342 91000
rect 30562 90540 30618 91000
rect 30838 90540 30894 91000
rect 31114 90540 31170 91000
rect 31390 90540 31446 91000
rect 31666 90540 31722 91000
rect 31942 90540 31998 91000
rect 32218 90540 32274 91000
rect 32494 90540 32550 91000
rect 32770 90540 32826 91000
rect 33046 90540 33102 91000
rect 33322 90540 33378 91000
rect 33598 90540 33654 91000
rect 33874 90540 33930 91000
rect 34150 90540 34206 91000
rect 34426 90540 34482 91000
rect 34702 90540 34758 91000
rect 34978 90540 35034 91000
rect 35254 90540 35310 91000
rect 35530 90540 35586 91000
rect 35806 90540 35862 91000
rect 36082 90540 36138 91000
rect 36358 90540 36414 91000
rect 36634 90540 36690 91000
rect 36910 90540 36966 91000
rect 37186 90540 37242 91000
rect 37462 90540 37518 91000
rect 37738 90540 37794 91000
rect 38014 90540 38070 91000
rect 38290 90540 38346 91000
rect 38566 90540 38622 91000
rect 38842 90540 38898 91000
rect 39118 90540 39174 91000
rect 39394 90540 39450 91000
rect 5170 -300 5226 160
rect 5446 -300 5502 160
rect 5722 -300 5778 160
rect 5998 -300 6054 160
rect 6274 -300 6330 160
rect 6550 -300 6606 160
rect 6826 -300 6882 160
rect 7102 -300 7158 160
rect 7378 -300 7434 160
rect 7654 -300 7710 160
rect 7930 -300 7986 160
rect 8206 -300 8262 160
rect 8482 -300 8538 160
rect 8758 -300 8814 160
rect 9034 -300 9090 160
rect 9310 -300 9366 160
rect 9586 -300 9642 160
rect 9862 -300 9918 160
rect 10138 -300 10194 160
rect 10414 -300 10470 160
rect 10690 -300 10746 160
rect 10966 -300 11022 160
rect 11242 -300 11298 160
rect 11518 -300 11574 160
rect 11794 -300 11850 160
rect 12070 -300 12126 160
rect 12346 -300 12402 160
rect 12622 -300 12678 160
rect 12898 -300 12954 160
rect 13174 -300 13230 160
rect 13450 -300 13506 160
rect 13726 -300 13782 160
rect 14002 -300 14058 160
rect 14278 -300 14334 160
rect 14554 -300 14610 160
rect 14830 -300 14886 160
rect 15106 -300 15162 160
rect 15382 -300 15438 160
rect 15658 -300 15714 160
rect 15934 -300 15990 160
rect 16210 -300 16266 160
rect 16486 -300 16542 160
rect 16762 -300 16818 160
rect 17038 -300 17094 160
rect 17314 -300 17370 160
rect 17590 -300 17646 160
rect 17866 -300 17922 160
rect 18142 -300 18198 160
rect 18418 -300 18474 160
rect 18694 -300 18750 160
rect 18970 -300 19026 160
rect 19246 -300 19302 160
rect 19522 -300 19578 160
rect 19798 -300 19854 160
rect 20074 -300 20130 160
rect 20350 -300 20406 160
rect 20626 -300 20682 160
rect 20902 -300 20958 160
rect 21178 -300 21234 160
rect 21454 -300 21510 160
rect 21730 -300 21786 160
rect 22006 -300 22062 160
rect 22282 -300 22338 160
rect 22558 -300 22614 160
rect 22834 -300 22890 160
rect 23110 -300 23166 160
rect 23386 -300 23442 160
rect 23662 -300 23718 160
rect 23938 -300 23994 160
rect 24214 -300 24270 160
rect 24490 -300 24546 160
rect 24766 -300 24822 160
rect 25042 -300 25098 160
rect 25318 -300 25374 160
rect 25594 -300 25650 160
rect 25870 -300 25926 160
rect 26146 -300 26202 160
rect 26422 -300 26478 160
rect 26698 -300 26754 160
rect 26974 -300 27030 160
rect 27250 -300 27306 160
rect 27526 -300 27582 160
rect 27802 -300 27858 160
rect 28078 -300 28134 160
rect 28354 -300 28410 160
rect 28630 -300 28686 160
rect 28906 -300 28962 160
rect 29182 -300 29238 160
rect 29458 -300 29514 160
rect 29734 -300 29790 160
rect 30010 -300 30066 160
rect 30286 -300 30342 160
rect 30562 -300 30618 160
rect 30838 -300 30894 160
rect 31114 -300 31170 160
rect 31390 -300 31446 160
rect 31666 -300 31722 160
rect 31942 -300 31998 160
rect 32218 -300 32274 160
rect 32494 -300 32550 160
rect 32770 -300 32826 160
rect 33046 -300 33102 160
rect 33322 -300 33378 160
rect 33598 -300 33654 160
rect 33874 -300 33930 160
rect 34150 -300 34206 160
rect 34426 -300 34482 160
rect 34702 -300 34758 160
rect 34978 -300 35034 160
rect 35254 -300 35310 160
rect 35530 -300 35586 160
rect 35806 -300 35862 160
rect 36082 -300 36138 160
rect 36358 -300 36414 160
rect 36634 -300 36690 160
rect 36910 -300 36966 160
rect 37186 -300 37242 160
rect 37462 -300 37518 160
rect 37738 -300 37794 160
rect 38014 -300 38070 160
rect 38290 -300 38346 160
rect 38566 -300 38622 160
rect 38842 -300 38898 160
rect 39118 -300 39174 160
rect 39394 -300 39450 160
<< obsm2 >>
rect 20 90484 5114 90658
rect 5282 90484 5390 90658
rect 5558 90484 5666 90658
rect 5834 90484 5942 90658
rect 6110 90484 6218 90658
rect 6386 90484 6494 90658
rect 6662 90484 6770 90658
rect 6938 90484 7046 90658
rect 7214 90484 7322 90658
rect 7490 90484 7598 90658
rect 7766 90484 7874 90658
rect 8042 90484 8150 90658
rect 8318 90484 8426 90658
rect 8594 90484 8702 90658
rect 8870 90484 8978 90658
rect 9146 90484 9254 90658
rect 9422 90484 9530 90658
rect 9698 90484 9806 90658
rect 9974 90484 10082 90658
rect 10250 90484 10358 90658
rect 10526 90484 10634 90658
rect 10802 90484 10910 90658
rect 11078 90484 11186 90658
rect 11354 90484 11462 90658
rect 11630 90484 11738 90658
rect 11906 90484 12014 90658
rect 12182 90484 12290 90658
rect 12458 90484 12566 90658
rect 12734 90484 12842 90658
rect 13010 90484 13118 90658
rect 13286 90484 13394 90658
rect 13562 90484 13670 90658
rect 13838 90484 13946 90658
rect 14114 90484 14222 90658
rect 14390 90484 14498 90658
rect 14666 90484 14774 90658
rect 14942 90484 15050 90658
rect 15218 90484 15326 90658
rect 15494 90484 15602 90658
rect 15770 90484 15878 90658
rect 16046 90484 16154 90658
rect 16322 90484 16430 90658
rect 16598 90484 16706 90658
rect 16874 90484 16982 90658
rect 17150 90484 17258 90658
rect 17426 90484 17534 90658
rect 17702 90484 17810 90658
rect 17978 90484 18086 90658
rect 18254 90484 18362 90658
rect 18530 90484 18638 90658
rect 18806 90484 18914 90658
rect 19082 90484 19190 90658
rect 19358 90484 19466 90658
rect 19634 90484 19742 90658
rect 19910 90484 20018 90658
rect 20186 90484 20294 90658
rect 20462 90484 20570 90658
rect 20738 90484 20846 90658
rect 21014 90484 21122 90658
rect 21290 90484 21398 90658
rect 21566 90484 21674 90658
rect 21842 90484 21950 90658
rect 22118 90484 22226 90658
rect 22394 90484 22502 90658
rect 22670 90484 22778 90658
rect 22946 90484 23054 90658
rect 23222 90484 23330 90658
rect 23498 90484 23606 90658
rect 23774 90484 23882 90658
rect 24050 90484 24158 90658
rect 24326 90484 24434 90658
rect 24602 90484 24710 90658
rect 24878 90484 24986 90658
rect 25154 90484 25262 90658
rect 25430 90484 25538 90658
rect 25706 90484 25814 90658
rect 25982 90484 26090 90658
rect 26258 90484 26366 90658
rect 26534 90484 26642 90658
rect 26810 90484 26918 90658
rect 27086 90484 27194 90658
rect 27362 90484 27470 90658
rect 27638 90484 27746 90658
rect 27914 90484 28022 90658
rect 28190 90484 28298 90658
rect 28466 90484 28574 90658
rect 28742 90484 28850 90658
rect 29018 90484 29126 90658
rect 29294 90484 29402 90658
rect 29570 90484 29678 90658
rect 29846 90484 29954 90658
rect 30122 90484 30230 90658
rect 30398 90484 30506 90658
rect 30674 90484 30782 90658
rect 30950 90484 31058 90658
rect 31226 90484 31334 90658
rect 31502 90484 31610 90658
rect 31778 90484 31886 90658
rect 32054 90484 32162 90658
rect 32330 90484 32438 90658
rect 32606 90484 32714 90658
rect 32882 90484 32990 90658
rect 33158 90484 33266 90658
rect 33434 90484 33542 90658
rect 33710 90484 33818 90658
rect 33986 90484 34094 90658
rect 34262 90484 34370 90658
rect 34538 90484 34646 90658
rect 34814 90484 34922 90658
rect 35090 90484 35198 90658
rect 35366 90484 35474 90658
rect 35642 90484 35750 90658
rect 35918 90484 36026 90658
rect 36194 90484 36302 90658
rect 36470 90484 36578 90658
rect 36746 90484 36854 90658
rect 37022 90484 37130 90658
rect 37298 90484 37406 90658
rect 37574 90484 37682 90658
rect 37850 90484 37958 90658
rect 38126 90484 38234 90658
rect 38402 90484 38510 90658
rect 38678 90484 38786 90658
rect 38954 90484 39062 90658
rect 39230 90484 39338 90658
rect 39506 90484 44692 90658
rect 20 216 44692 90484
rect 20 54 5114 216
rect 5282 54 5390 216
rect 5558 54 5666 216
rect 5834 54 5942 216
rect 6110 54 6218 216
rect 6386 54 6494 216
rect 6662 54 6770 216
rect 6938 54 7046 216
rect 7214 54 7322 216
rect 7490 54 7598 216
rect 7766 54 7874 216
rect 8042 54 8150 216
rect 8318 54 8426 216
rect 8594 54 8702 216
rect 8870 54 8978 216
rect 9146 54 9254 216
rect 9422 54 9530 216
rect 9698 54 9806 216
rect 9974 54 10082 216
rect 10250 54 10358 216
rect 10526 54 10634 216
rect 10802 54 10910 216
rect 11078 54 11186 216
rect 11354 54 11462 216
rect 11630 54 11738 216
rect 11906 54 12014 216
rect 12182 54 12290 216
rect 12458 54 12566 216
rect 12734 54 12842 216
rect 13010 54 13118 216
rect 13286 54 13394 216
rect 13562 54 13670 216
rect 13838 54 13946 216
rect 14114 54 14222 216
rect 14390 54 14498 216
rect 14666 54 14774 216
rect 14942 54 15050 216
rect 15218 54 15326 216
rect 15494 54 15602 216
rect 15770 54 15878 216
rect 16046 54 16154 216
rect 16322 54 16430 216
rect 16598 54 16706 216
rect 16874 54 16982 216
rect 17150 54 17258 216
rect 17426 54 17534 216
rect 17702 54 17810 216
rect 17978 54 18086 216
rect 18254 54 18362 216
rect 18530 54 18638 216
rect 18806 54 18914 216
rect 19082 54 19190 216
rect 19358 54 19466 216
rect 19634 54 19742 216
rect 19910 54 20018 216
rect 20186 54 20294 216
rect 20462 54 20570 216
rect 20738 54 20846 216
rect 21014 54 21122 216
rect 21290 54 21398 216
rect 21566 54 21674 216
rect 21842 54 21950 216
rect 22118 54 22226 216
rect 22394 54 22502 216
rect 22670 54 22778 216
rect 22946 54 23054 216
rect 23222 54 23330 216
rect 23498 54 23606 216
rect 23774 54 23882 216
rect 24050 54 24158 216
rect 24326 54 24434 216
rect 24602 54 24710 216
rect 24878 54 24986 216
rect 25154 54 25262 216
rect 25430 54 25538 216
rect 25706 54 25814 216
rect 25982 54 26090 216
rect 26258 54 26366 216
rect 26534 54 26642 216
rect 26810 54 26918 216
rect 27086 54 27194 216
rect 27362 54 27470 216
rect 27638 54 27746 216
rect 27914 54 28022 216
rect 28190 54 28298 216
rect 28466 54 28574 216
rect 28742 54 28850 216
rect 29018 54 29126 216
rect 29294 54 29402 216
rect 29570 54 29678 216
rect 29846 54 29954 216
rect 30122 54 30230 216
rect 30398 54 30506 216
rect 30674 54 30782 216
rect 30950 54 31058 216
rect 31226 54 31334 216
rect 31502 54 31610 216
rect 31778 54 31886 216
rect 32054 54 32162 216
rect 32330 54 32438 216
rect 32606 54 32714 216
rect 32882 54 32990 216
rect 33158 54 33266 216
rect 33434 54 33542 216
rect 33710 54 33818 216
rect 33986 54 34094 216
rect 34262 54 34370 216
rect 34538 54 34646 216
rect 34814 54 34922 216
rect 35090 54 35198 216
rect 35366 54 35474 216
rect 35642 54 35750 216
rect 35918 54 36026 216
rect 36194 54 36302 216
rect 36470 54 36578 216
rect 36746 54 36854 216
rect 37022 54 37130 216
rect 37298 54 37406 216
rect 37574 54 37682 216
rect 37850 54 37958 216
rect 38126 54 38234 216
rect 38402 54 38510 216
rect 38678 54 38786 216
rect 38954 54 39062 216
rect 39230 54 39338 216
rect 39506 54 44692 216
<< metal3 >>
rect -300 85688 160 85808
rect -300 85416 160 85536
rect -300 85144 160 85264
rect -300 84872 160 84992
rect -300 84600 160 84720
rect -300 84328 160 84448
rect -300 84056 160 84176
rect -300 83784 160 83904
rect -300 83512 160 83632
rect -300 83240 160 83360
rect -300 82968 160 83088
rect -300 82696 160 82816
rect -300 82424 160 82544
rect -300 82152 160 82272
rect -300 81880 160 82000
rect -300 81608 160 81728
rect -300 81336 160 81456
rect -300 81064 160 81184
rect -300 80792 160 80912
rect -300 80520 160 80640
rect -300 80248 160 80368
rect -300 79976 160 80096
rect -300 79704 160 79824
rect -300 79432 160 79552
rect -300 79160 160 79280
rect -300 78888 160 79008
rect -300 78616 160 78736
rect -300 78344 160 78464
rect -300 78072 160 78192
rect -300 77800 160 77920
rect -300 77528 160 77648
rect -300 77256 160 77376
rect -300 76984 160 77104
rect -300 76712 160 76832
rect -300 76440 160 76560
rect -300 76168 160 76288
rect -300 75896 160 76016
rect -300 75624 160 75744
rect -300 75352 160 75472
rect -300 75080 160 75200
rect -300 74808 160 74928
rect -300 74536 160 74656
rect -300 74264 160 74384
rect -300 73992 160 74112
rect -300 73720 160 73840
rect -300 73448 160 73568
rect -300 73176 160 73296
rect -300 72904 160 73024
rect -300 72632 160 72752
rect -300 72360 160 72480
rect -300 72088 160 72208
rect -300 71816 160 71936
rect -300 71544 160 71664
rect -300 71272 160 71392
rect -300 71000 160 71120
rect -300 70728 160 70848
rect -300 70456 160 70576
rect -300 70184 160 70304
rect -300 69912 160 70032
rect -300 69640 160 69760
rect -300 69368 160 69488
rect -300 69096 160 69216
rect -300 68824 160 68944
rect -300 68552 160 68672
rect -300 68280 160 68400
rect -300 68008 160 68128
rect -300 67736 160 67856
rect -300 67464 160 67584
rect -300 67192 160 67312
rect -300 66920 160 67040
rect -300 66648 160 66768
rect -300 66376 160 66496
rect -300 66104 160 66224
rect -300 65832 160 65952
rect -300 65560 160 65680
rect -300 65288 160 65408
rect -300 65016 160 65136
rect -300 64744 160 64864
rect -300 64472 160 64592
rect -300 64200 160 64320
rect -300 63928 160 64048
rect -300 63656 160 63776
rect -300 63384 160 63504
rect -300 63112 160 63232
rect -300 62840 160 62960
rect -300 62568 160 62688
rect -300 62296 160 62416
rect -300 62024 160 62144
rect -300 61752 160 61872
rect -300 61480 160 61600
rect -300 61208 160 61328
rect -300 60936 160 61056
rect -300 60664 160 60784
rect -300 60392 160 60512
rect -300 60120 160 60240
rect -300 59848 160 59968
rect -300 59576 160 59696
rect -300 59304 160 59424
rect -300 59032 160 59152
rect -300 58760 160 58880
rect -300 58488 160 58608
rect -300 58216 160 58336
rect -300 57944 160 58064
rect -300 57672 160 57792
rect -300 57400 160 57520
rect -300 57128 160 57248
rect -300 56856 160 56976
rect -300 56584 160 56704
rect -300 56312 160 56432
rect -300 56040 160 56160
rect -300 55768 160 55888
rect -300 55496 160 55616
rect -300 55224 160 55344
rect -300 54952 160 55072
rect -300 54680 160 54800
rect -300 54408 160 54528
rect -300 54136 160 54256
rect -300 53864 160 53984
rect -300 53592 160 53712
rect -300 53320 160 53440
rect -300 53048 160 53168
rect -300 52776 160 52896
rect -300 52504 160 52624
rect -300 52232 160 52352
rect -300 51960 160 52080
rect -300 51688 160 51808
rect -300 51416 160 51536
rect -300 51144 160 51264
rect 44540 85688 45000 85808
rect 44540 85416 45000 85536
rect 44540 85144 45000 85264
rect 44540 84872 45000 84992
rect 44540 84600 45000 84720
rect 44540 84328 45000 84448
rect 44540 84056 45000 84176
rect 44540 83784 45000 83904
rect 44540 83512 45000 83632
rect 44540 83240 45000 83360
rect 44540 82968 45000 83088
rect 44540 82696 45000 82816
rect 44540 82424 45000 82544
rect 44540 82152 45000 82272
rect 44540 81880 45000 82000
rect 44540 81608 45000 81728
rect 44540 81336 45000 81456
rect 44540 81064 45000 81184
rect 44540 80792 45000 80912
rect 44540 80520 45000 80640
rect 44540 80248 45000 80368
rect 44540 79976 45000 80096
rect 44540 79704 45000 79824
rect 44540 79432 45000 79552
rect 44540 79160 45000 79280
rect 44540 78888 45000 79008
rect 44540 78616 45000 78736
rect 44540 78344 45000 78464
rect 44540 78072 45000 78192
rect 44540 77800 45000 77920
rect 44540 77528 45000 77648
rect 44540 77256 45000 77376
rect 44540 76984 45000 77104
rect 44540 76712 45000 76832
rect 44540 76440 45000 76560
rect 44540 76168 45000 76288
rect 44540 75896 45000 76016
rect 44540 75624 45000 75744
rect 44540 75352 45000 75472
rect 44540 75080 45000 75200
rect 44540 74808 45000 74928
rect 44540 74536 45000 74656
rect 44540 74264 45000 74384
rect 44540 73992 45000 74112
rect 44540 73720 45000 73840
rect 44540 73448 45000 73568
rect 44540 73176 45000 73296
rect 44540 72904 45000 73024
rect 44540 72632 45000 72752
rect 44540 72360 45000 72480
rect 44540 72088 45000 72208
rect 44540 71816 45000 71936
rect 44540 71544 45000 71664
rect 44540 71272 45000 71392
rect 44540 71000 45000 71120
rect 44540 70728 45000 70848
rect 44540 70456 45000 70576
rect 44540 70184 45000 70304
rect 44540 69912 45000 70032
rect 44540 69640 45000 69760
rect 44540 69368 45000 69488
rect 44540 69096 45000 69216
rect 44540 68824 45000 68944
rect 44540 68552 45000 68672
rect 44540 68280 45000 68400
rect 44540 68008 45000 68128
rect 44540 67736 45000 67856
rect 44540 67464 45000 67584
rect 44540 67192 45000 67312
rect 44540 66920 45000 67040
rect 44540 66648 45000 66768
rect 44540 66376 45000 66496
rect 44540 66104 45000 66224
rect 44540 65832 45000 65952
rect 44540 65560 45000 65680
rect 44540 65288 45000 65408
rect 44540 65016 45000 65136
rect 44540 64744 45000 64864
rect 44540 64472 45000 64592
rect 44540 64200 45000 64320
rect 44540 63928 45000 64048
rect 44540 63656 45000 63776
rect 44540 63384 45000 63504
rect 44540 63112 45000 63232
rect 44540 62840 45000 62960
rect 44540 62568 45000 62688
rect 44540 62296 45000 62416
rect 44540 62024 45000 62144
rect 44540 61752 45000 61872
rect 44540 61480 45000 61600
rect 44540 61208 45000 61328
rect 44540 60936 45000 61056
rect 44540 60664 45000 60784
rect 44540 60392 45000 60512
rect 44540 60120 45000 60240
rect 44540 59848 45000 59968
rect 44540 59576 45000 59696
rect 44540 59304 45000 59424
rect 44540 59032 45000 59152
rect 44540 58760 45000 58880
rect 44540 58488 45000 58608
rect 44540 58216 45000 58336
rect 44540 57944 45000 58064
rect 44540 57672 45000 57792
rect 44540 57400 45000 57520
rect 44540 57128 45000 57248
rect 44540 56856 45000 56976
rect 44540 56584 45000 56704
rect 44540 56312 45000 56432
rect 44540 56040 45000 56160
rect 44540 55768 45000 55888
rect 44540 55496 45000 55616
rect 44540 55224 45000 55344
rect 44540 54952 45000 55072
rect 44540 54680 45000 54800
rect 44540 54408 45000 54528
rect 44540 54136 45000 54256
rect 44540 53864 45000 53984
rect 44540 53592 45000 53712
rect 44540 53320 45000 53440
rect 44540 53048 45000 53168
rect 44540 52776 45000 52896
rect 44540 52504 45000 52624
rect 44540 52232 45000 52352
rect 44540 51960 45000 52080
rect 44540 51688 45000 51808
rect 44540 51416 45000 51536
rect 44540 51144 45000 51264
rect -300 39720 160 39840
rect -300 39448 160 39568
rect -300 39176 160 39296
rect -300 38904 160 39024
rect -300 38632 160 38752
rect -300 38360 160 38480
rect -300 38088 160 38208
rect -300 37816 160 37936
rect -300 37544 160 37664
rect -300 37272 160 37392
rect -300 37000 160 37120
rect -300 36728 160 36848
rect -300 36456 160 36576
rect -300 36184 160 36304
rect -300 35912 160 36032
rect -300 35640 160 35760
rect -300 35368 160 35488
rect -300 35096 160 35216
rect -300 34824 160 34944
rect -300 34552 160 34672
rect -300 34280 160 34400
rect -300 34008 160 34128
rect -300 33736 160 33856
rect -300 33464 160 33584
rect -300 33192 160 33312
rect -300 32920 160 33040
rect -300 32648 160 32768
rect -300 32376 160 32496
rect -300 32104 160 32224
rect -300 31832 160 31952
rect -300 31560 160 31680
rect -300 31288 160 31408
rect -300 31016 160 31136
rect -300 30744 160 30864
rect -300 30472 160 30592
rect -300 30200 160 30320
rect -300 29928 160 30048
rect -300 29656 160 29776
rect -300 29384 160 29504
rect -300 29112 160 29232
rect -300 28840 160 28960
rect -300 28568 160 28688
rect -300 28296 160 28416
rect -300 28024 160 28144
rect -300 27752 160 27872
rect -300 27480 160 27600
rect -300 27208 160 27328
rect -300 26936 160 27056
rect -300 26664 160 26784
rect -300 26392 160 26512
rect -300 26120 160 26240
rect -300 25848 160 25968
rect -300 25576 160 25696
rect -300 25304 160 25424
rect -300 25032 160 25152
rect -300 24760 160 24880
rect -300 24488 160 24608
rect -300 24216 160 24336
rect -300 23944 160 24064
rect -300 23672 160 23792
rect -300 23400 160 23520
rect -300 23128 160 23248
rect -300 22856 160 22976
rect -300 22584 160 22704
rect -300 22312 160 22432
rect -300 22040 160 22160
rect -300 21768 160 21888
rect -300 21496 160 21616
rect -300 21224 160 21344
rect -300 20952 160 21072
rect -300 20680 160 20800
rect -300 20408 160 20528
rect -300 20136 160 20256
rect -300 19864 160 19984
rect -300 19592 160 19712
rect -300 19320 160 19440
rect -300 19048 160 19168
rect -300 18776 160 18896
rect -300 18504 160 18624
rect -300 18232 160 18352
rect -300 17960 160 18080
rect -300 17688 160 17808
rect -300 17416 160 17536
rect -300 17144 160 17264
rect -300 16872 160 16992
rect -300 16600 160 16720
rect -300 16328 160 16448
rect -300 16056 160 16176
rect -300 15784 160 15904
rect -300 15512 160 15632
rect -300 15240 160 15360
rect -300 14968 160 15088
rect -300 14696 160 14816
rect -300 14424 160 14544
rect -300 14152 160 14272
rect -300 13880 160 14000
rect -300 13608 160 13728
rect -300 13336 160 13456
rect -300 13064 160 13184
rect -300 12792 160 12912
rect -300 12520 160 12640
rect -300 12248 160 12368
rect -300 11976 160 12096
rect -300 11704 160 11824
rect -300 11432 160 11552
rect -300 11160 160 11280
rect -300 10888 160 11008
rect -300 10616 160 10736
rect -300 10344 160 10464
rect -300 10072 160 10192
rect -300 9800 160 9920
rect -300 9528 160 9648
rect -300 9256 160 9376
rect -300 8984 160 9104
rect -300 8712 160 8832
rect -300 8440 160 8560
rect -300 8168 160 8288
rect -300 7896 160 8016
rect -300 7624 160 7744
rect -300 7352 160 7472
rect -300 7080 160 7200
rect -300 6808 160 6928
rect -300 6536 160 6656
rect -300 6264 160 6384
rect -300 5992 160 6112
rect -300 5720 160 5840
rect -300 5448 160 5568
rect -300 5176 160 5296
rect 44540 39720 45000 39840
rect 44540 39448 45000 39568
rect 44540 39176 45000 39296
rect 44540 38904 45000 39024
rect 44540 38632 45000 38752
rect 44540 38360 45000 38480
rect 44540 38088 45000 38208
rect 44540 37816 45000 37936
rect 44540 37544 45000 37664
rect 44540 37272 45000 37392
rect 44540 37000 45000 37120
rect 44540 36728 45000 36848
rect 44540 36456 45000 36576
rect 44540 36184 45000 36304
rect 44540 35912 45000 36032
rect 44540 35640 45000 35760
rect 44540 35368 45000 35488
rect 44540 35096 45000 35216
rect 44540 34824 45000 34944
rect 44540 34552 45000 34672
rect 44540 34280 45000 34400
rect 44540 34008 45000 34128
rect 44540 33736 45000 33856
rect 44540 33464 45000 33584
rect 44540 33192 45000 33312
rect 44540 32920 45000 33040
rect 44540 32648 45000 32768
rect 44540 32376 45000 32496
rect 44540 32104 45000 32224
rect 44540 31832 45000 31952
rect 44540 31560 45000 31680
rect 44540 31288 45000 31408
rect 44540 31016 45000 31136
rect 44540 30744 45000 30864
rect 44540 30472 45000 30592
rect 44540 30200 45000 30320
rect 44540 29928 45000 30048
rect 44540 29656 45000 29776
rect 44540 29384 45000 29504
rect 44540 29112 45000 29232
rect 44540 28840 45000 28960
rect 44540 28568 45000 28688
rect 44540 28296 45000 28416
rect 44540 28024 45000 28144
rect 44540 27752 45000 27872
rect 44540 27480 45000 27600
rect 44540 27208 45000 27328
rect 44540 26936 45000 27056
rect 44540 26664 45000 26784
rect 44540 26392 45000 26512
rect 44540 26120 45000 26240
rect 44540 25848 45000 25968
rect 44540 25576 45000 25696
rect 44540 25304 45000 25424
rect 44540 25032 45000 25152
rect 44540 24760 45000 24880
rect 44540 24488 45000 24608
rect 44540 24216 45000 24336
rect 44540 23944 45000 24064
rect 44540 23672 45000 23792
rect 44540 23400 45000 23520
rect 44540 23128 45000 23248
rect 44540 22856 45000 22976
rect 44540 22584 45000 22704
rect 44540 22312 45000 22432
rect 44540 22040 45000 22160
rect 44540 21768 45000 21888
rect 44540 21496 45000 21616
rect 44540 21224 45000 21344
rect 44540 20952 45000 21072
rect 44540 20680 45000 20800
rect 44540 20408 45000 20528
rect 44540 20136 45000 20256
rect 44540 19864 45000 19984
rect 44540 19592 45000 19712
rect 44540 19320 45000 19440
rect 44540 19048 45000 19168
rect 44540 18776 45000 18896
rect 44540 18504 45000 18624
rect 44540 18232 45000 18352
rect 44540 17960 45000 18080
rect 44540 17688 45000 17808
rect 44540 17416 45000 17536
rect 44540 17144 45000 17264
rect 44540 16872 45000 16992
rect 44540 16600 45000 16720
rect 44540 16328 45000 16448
rect 44540 16056 45000 16176
rect 44540 15784 45000 15904
rect 44540 15512 45000 15632
rect 44540 15240 45000 15360
rect 44540 14968 45000 15088
rect 44540 14696 45000 14816
rect 44540 14424 45000 14544
rect 44540 14152 45000 14272
rect 44540 13880 45000 14000
rect 44540 13608 45000 13728
rect 44540 13336 45000 13456
rect 44540 13064 45000 13184
rect 44540 12792 45000 12912
rect 44540 12520 45000 12640
rect 44540 12248 45000 12368
rect 44540 11976 45000 12096
rect 44540 11704 45000 11824
rect 44540 11432 45000 11552
rect 44540 11160 45000 11280
rect 44540 10888 45000 11008
rect 44540 10616 45000 10736
rect 44540 10344 45000 10464
rect 44540 10072 45000 10192
rect 44540 9800 45000 9920
rect 44540 9528 45000 9648
rect 44540 9256 45000 9376
rect 44540 8984 45000 9104
rect 44540 8712 45000 8832
rect 44540 8440 45000 8560
rect 44540 8168 45000 8288
rect 44540 7896 45000 8016
rect 44540 7624 45000 7744
rect 44540 7352 45000 7472
rect 44540 7080 45000 7200
rect 44540 6808 45000 6928
rect 44540 6536 45000 6656
rect 44540 6264 45000 6384
rect 44540 5992 45000 6112
rect 44540 5720 45000 5840
rect 44540 5448 45000 5568
rect 44540 5176 45000 5296
<< obsm3 >>
rect 160 85888 44540 89453
rect 240 51064 44460 85888
rect 160 39920 44540 51064
rect 240 5096 44460 39920
rect 160 715 44540 5096
<< metal4 >>
rect 4208 1040 4528 89264
rect 19568 1040 19888 89264
rect 34928 1040 35248 89264
<< obsm4 >>
rect 795 89344 42261 89453
rect 795 960 4128 89344
rect 4608 960 19488 89344
rect 19968 960 34848 89344
rect 35328 960 42261 89344
rect 795 715 42261 960
<< labels >>
rlabel metal3 s 44540 64200 45000 64320 6 Tile_X0Y0_E1BEG[0]
port 1 nsew signal output
rlabel metal3 s 44540 64472 45000 64592 6 Tile_X0Y0_E1BEG[1]
port 2 nsew signal output
rlabel metal3 s 44540 64744 45000 64864 6 Tile_X0Y0_E1BEG[2]
port 3 nsew signal output
rlabel metal3 s 44540 65016 45000 65136 6 Tile_X0Y0_E1BEG[3]
port 4 nsew signal output
rlabel metal3 s -300 64200 160 64320 4 Tile_X0Y0_E1END[0]
port 5 nsew signal input
rlabel metal3 s -300 64472 160 64592 4 Tile_X0Y0_E1END[1]
port 6 nsew signal input
rlabel metal3 s -300 64744 160 64864 4 Tile_X0Y0_E1END[2]
port 7 nsew signal input
rlabel metal3 s -300 65016 160 65136 4 Tile_X0Y0_E1END[3]
port 8 nsew signal input
rlabel metal3 s 44540 65288 45000 65408 6 Tile_X0Y0_E2BEG[0]
port 9 nsew signal output
rlabel metal3 s 44540 65560 45000 65680 6 Tile_X0Y0_E2BEG[1]
port 10 nsew signal output
rlabel metal3 s 44540 65832 45000 65952 6 Tile_X0Y0_E2BEG[2]
port 11 nsew signal output
rlabel metal3 s 44540 66104 45000 66224 6 Tile_X0Y0_E2BEG[3]
port 12 nsew signal output
rlabel metal3 s 44540 66376 45000 66496 6 Tile_X0Y0_E2BEG[4]
port 13 nsew signal output
rlabel metal3 s 44540 66648 45000 66768 6 Tile_X0Y0_E2BEG[5]
port 14 nsew signal output
rlabel metal3 s 44540 66920 45000 67040 6 Tile_X0Y0_E2BEG[6]
port 15 nsew signal output
rlabel metal3 s 44540 67192 45000 67312 6 Tile_X0Y0_E2BEG[7]
port 16 nsew signal output
rlabel metal3 s 44540 67464 45000 67584 6 Tile_X0Y0_E2BEGb[0]
port 17 nsew signal output
rlabel metal3 s 44540 67736 45000 67856 6 Tile_X0Y0_E2BEGb[1]
port 18 nsew signal output
rlabel metal3 s 44540 68008 45000 68128 6 Tile_X0Y0_E2BEGb[2]
port 19 nsew signal output
rlabel metal3 s 44540 68280 45000 68400 6 Tile_X0Y0_E2BEGb[3]
port 20 nsew signal output
rlabel metal3 s 44540 68552 45000 68672 6 Tile_X0Y0_E2BEGb[4]
port 21 nsew signal output
rlabel metal3 s 44540 68824 45000 68944 6 Tile_X0Y0_E2BEGb[5]
port 22 nsew signal output
rlabel metal3 s 44540 69096 45000 69216 6 Tile_X0Y0_E2BEGb[6]
port 23 nsew signal output
rlabel metal3 s 44540 69368 45000 69488 6 Tile_X0Y0_E2BEGb[7]
port 24 nsew signal output
rlabel metal3 s -300 67464 160 67584 4 Tile_X0Y0_E2END[0]
port 25 nsew signal input
rlabel metal3 s -300 67736 160 67856 4 Tile_X0Y0_E2END[1]
port 26 nsew signal input
rlabel metal3 s -300 68008 160 68128 4 Tile_X0Y0_E2END[2]
port 27 nsew signal input
rlabel metal3 s -300 68280 160 68400 4 Tile_X0Y0_E2END[3]
port 28 nsew signal input
rlabel metal3 s -300 68552 160 68672 4 Tile_X0Y0_E2END[4]
port 29 nsew signal input
rlabel metal3 s -300 68824 160 68944 4 Tile_X0Y0_E2END[5]
port 30 nsew signal input
rlabel metal3 s -300 69096 160 69216 4 Tile_X0Y0_E2END[6]
port 31 nsew signal input
rlabel metal3 s -300 69368 160 69488 4 Tile_X0Y0_E2END[7]
port 32 nsew signal input
rlabel metal3 s -300 65288 160 65408 4 Tile_X0Y0_E2MID[0]
port 33 nsew signal input
rlabel metal3 s -300 65560 160 65680 4 Tile_X0Y0_E2MID[1]
port 34 nsew signal input
rlabel metal3 s -300 65832 160 65952 4 Tile_X0Y0_E2MID[2]
port 35 nsew signal input
rlabel metal3 s -300 66104 160 66224 4 Tile_X0Y0_E2MID[3]
port 36 nsew signal input
rlabel metal3 s -300 66376 160 66496 4 Tile_X0Y0_E2MID[4]
port 37 nsew signal input
rlabel metal3 s -300 66648 160 66768 4 Tile_X0Y0_E2MID[5]
port 38 nsew signal input
rlabel metal3 s -300 66920 160 67040 4 Tile_X0Y0_E2MID[6]
port 39 nsew signal input
rlabel metal3 s -300 67192 160 67312 4 Tile_X0Y0_E2MID[7]
port 40 nsew signal input
rlabel metal3 s 44540 73992 45000 74112 6 Tile_X0Y0_E6BEG[0]
port 41 nsew signal output
rlabel metal3 s 44540 76712 45000 76832 6 Tile_X0Y0_E6BEG[10]
port 42 nsew signal output
rlabel metal3 s 44540 76984 45000 77104 6 Tile_X0Y0_E6BEG[11]
port 43 nsew signal output
rlabel metal3 s 44540 74264 45000 74384 6 Tile_X0Y0_E6BEG[1]
port 44 nsew signal output
rlabel metal3 s 44540 74536 45000 74656 6 Tile_X0Y0_E6BEG[2]
port 45 nsew signal output
rlabel metal3 s 44540 74808 45000 74928 6 Tile_X0Y0_E6BEG[3]
port 46 nsew signal output
rlabel metal3 s 44540 75080 45000 75200 6 Tile_X0Y0_E6BEG[4]
port 47 nsew signal output
rlabel metal3 s 44540 75352 45000 75472 6 Tile_X0Y0_E6BEG[5]
port 48 nsew signal output
rlabel metal3 s 44540 75624 45000 75744 6 Tile_X0Y0_E6BEG[6]
port 49 nsew signal output
rlabel metal3 s 44540 75896 45000 76016 6 Tile_X0Y0_E6BEG[7]
port 50 nsew signal output
rlabel metal3 s 44540 76168 45000 76288 6 Tile_X0Y0_E6BEG[8]
port 51 nsew signal output
rlabel metal3 s 44540 76440 45000 76560 6 Tile_X0Y0_E6BEG[9]
port 52 nsew signal output
rlabel metal3 s -300 73992 160 74112 4 Tile_X0Y0_E6END[0]
port 53 nsew signal input
rlabel metal3 s -300 76712 160 76832 4 Tile_X0Y0_E6END[10]
port 54 nsew signal input
rlabel metal3 s -300 76984 160 77104 4 Tile_X0Y0_E6END[11]
port 55 nsew signal input
rlabel metal3 s -300 74264 160 74384 4 Tile_X0Y0_E6END[1]
port 56 nsew signal input
rlabel metal3 s -300 74536 160 74656 4 Tile_X0Y0_E6END[2]
port 57 nsew signal input
rlabel metal3 s -300 74808 160 74928 4 Tile_X0Y0_E6END[3]
port 58 nsew signal input
rlabel metal3 s -300 75080 160 75200 4 Tile_X0Y0_E6END[4]
port 59 nsew signal input
rlabel metal3 s -300 75352 160 75472 4 Tile_X0Y0_E6END[5]
port 60 nsew signal input
rlabel metal3 s -300 75624 160 75744 4 Tile_X0Y0_E6END[6]
port 61 nsew signal input
rlabel metal3 s -300 75896 160 76016 4 Tile_X0Y0_E6END[7]
port 62 nsew signal input
rlabel metal3 s -300 76168 160 76288 4 Tile_X0Y0_E6END[8]
port 63 nsew signal input
rlabel metal3 s -300 76440 160 76560 4 Tile_X0Y0_E6END[9]
port 64 nsew signal input
rlabel metal3 s 44540 69640 45000 69760 6 Tile_X0Y0_EE4BEG[0]
port 65 nsew signal output
rlabel metal3 s 44540 72360 45000 72480 6 Tile_X0Y0_EE4BEG[10]
port 66 nsew signal output
rlabel metal3 s 44540 72632 45000 72752 6 Tile_X0Y0_EE4BEG[11]
port 67 nsew signal output
rlabel metal3 s 44540 72904 45000 73024 6 Tile_X0Y0_EE4BEG[12]
port 68 nsew signal output
rlabel metal3 s 44540 73176 45000 73296 6 Tile_X0Y0_EE4BEG[13]
port 69 nsew signal output
rlabel metal3 s 44540 73448 45000 73568 6 Tile_X0Y0_EE4BEG[14]
port 70 nsew signal output
rlabel metal3 s 44540 73720 45000 73840 6 Tile_X0Y0_EE4BEG[15]
port 71 nsew signal output
rlabel metal3 s 44540 69912 45000 70032 6 Tile_X0Y0_EE4BEG[1]
port 72 nsew signal output
rlabel metal3 s 44540 70184 45000 70304 6 Tile_X0Y0_EE4BEG[2]
port 73 nsew signal output
rlabel metal3 s 44540 70456 45000 70576 6 Tile_X0Y0_EE4BEG[3]
port 74 nsew signal output
rlabel metal3 s 44540 70728 45000 70848 6 Tile_X0Y0_EE4BEG[4]
port 75 nsew signal output
rlabel metal3 s 44540 71000 45000 71120 6 Tile_X0Y0_EE4BEG[5]
port 76 nsew signal output
rlabel metal3 s 44540 71272 45000 71392 6 Tile_X0Y0_EE4BEG[6]
port 77 nsew signal output
rlabel metal3 s 44540 71544 45000 71664 6 Tile_X0Y0_EE4BEG[7]
port 78 nsew signal output
rlabel metal3 s 44540 71816 45000 71936 6 Tile_X0Y0_EE4BEG[8]
port 79 nsew signal output
rlabel metal3 s 44540 72088 45000 72208 6 Tile_X0Y0_EE4BEG[9]
port 80 nsew signal output
rlabel metal3 s -300 69640 160 69760 4 Tile_X0Y0_EE4END[0]
port 81 nsew signal input
rlabel metal3 s -300 72360 160 72480 4 Tile_X0Y0_EE4END[10]
port 82 nsew signal input
rlabel metal3 s -300 72632 160 72752 4 Tile_X0Y0_EE4END[11]
port 83 nsew signal input
rlabel metal3 s -300 72904 160 73024 4 Tile_X0Y0_EE4END[12]
port 84 nsew signal input
rlabel metal3 s -300 73176 160 73296 4 Tile_X0Y0_EE4END[13]
port 85 nsew signal input
rlabel metal3 s -300 73448 160 73568 4 Tile_X0Y0_EE4END[14]
port 86 nsew signal input
rlabel metal3 s -300 73720 160 73840 4 Tile_X0Y0_EE4END[15]
port 87 nsew signal input
rlabel metal3 s -300 69912 160 70032 4 Tile_X0Y0_EE4END[1]
port 88 nsew signal input
rlabel metal3 s -300 70184 160 70304 4 Tile_X0Y0_EE4END[2]
port 89 nsew signal input
rlabel metal3 s -300 70456 160 70576 4 Tile_X0Y0_EE4END[3]
port 90 nsew signal input
rlabel metal3 s -300 70728 160 70848 4 Tile_X0Y0_EE4END[4]
port 91 nsew signal input
rlabel metal3 s -300 71000 160 71120 4 Tile_X0Y0_EE4END[5]
port 92 nsew signal input
rlabel metal3 s -300 71272 160 71392 4 Tile_X0Y0_EE4END[6]
port 93 nsew signal input
rlabel metal3 s -300 71544 160 71664 4 Tile_X0Y0_EE4END[7]
port 94 nsew signal input
rlabel metal3 s -300 71816 160 71936 4 Tile_X0Y0_EE4END[8]
port 95 nsew signal input
rlabel metal3 s -300 72088 160 72208 4 Tile_X0Y0_EE4END[9]
port 96 nsew signal input
rlabel metal3 s -300 77256 160 77376 4 Tile_X0Y0_FrameData[0]
port 97 nsew signal input
rlabel metal3 s -300 79976 160 80096 4 Tile_X0Y0_FrameData[10]
port 98 nsew signal input
rlabel metal3 s -300 80248 160 80368 4 Tile_X0Y0_FrameData[11]
port 99 nsew signal input
rlabel metal3 s -300 80520 160 80640 4 Tile_X0Y0_FrameData[12]
port 100 nsew signal input
rlabel metal3 s -300 80792 160 80912 4 Tile_X0Y0_FrameData[13]
port 101 nsew signal input
rlabel metal3 s -300 81064 160 81184 4 Tile_X0Y0_FrameData[14]
port 102 nsew signal input
rlabel metal3 s -300 81336 160 81456 4 Tile_X0Y0_FrameData[15]
port 103 nsew signal input
rlabel metal3 s -300 81608 160 81728 4 Tile_X0Y0_FrameData[16]
port 104 nsew signal input
rlabel metal3 s -300 81880 160 82000 4 Tile_X0Y0_FrameData[17]
port 105 nsew signal input
rlabel metal3 s -300 82152 160 82272 4 Tile_X0Y0_FrameData[18]
port 106 nsew signal input
rlabel metal3 s -300 82424 160 82544 4 Tile_X0Y0_FrameData[19]
port 107 nsew signal input
rlabel metal3 s -300 77528 160 77648 4 Tile_X0Y0_FrameData[1]
port 108 nsew signal input
rlabel metal3 s -300 82696 160 82816 4 Tile_X0Y0_FrameData[20]
port 109 nsew signal input
rlabel metal3 s -300 82968 160 83088 4 Tile_X0Y0_FrameData[21]
port 110 nsew signal input
rlabel metal3 s -300 83240 160 83360 4 Tile_X0Y0_FrameData[22]
port 111 nsew signal input
rlabel metal3 s -300 83512 160 83632 4 Tile_X0Y0_FrameData[23]
port 112 nsew signal input
rlabel metal3 s -300 83784 160 83904 4 Tile_X0Y0_FrameData[24]
port 113 nsew signal input
rlabel metal3 s -300 84056 160 84176 4 Tile_X0Y0_FrameData[25]
port 114 nsew signal input
rlabel metal3 s -300 84328 160 84448 4 Tile_X0Y0_FrameData[26]
port 115 nsew signal input
rlabel metal3 s -300 84600 160 84720 4 Tile_X0Y0_FrameData[27]
port 116 nsew signal input
rlabel metal3 s -300 84872 160 84992 4 Tile_X0Y0_FrameData[28]
port 117 nsew signal input
rlabel metal3 s -300 85144 160 85264 4 Tile_X0Y0_FrameData[29]
port 118 nsew signal input
rlabel metal3 s -300 77800 160 77920 4 Tile_X0Y0_FrameData[2]
port 119 nsew signal input
rlabel metal3 s -300 85416 160 85536 4 Tile_X0Y0_FrameData[30]
port 120 nsew signal input
rlabel metal3 s -300 85688 160 85808 4 Tile_X0Y0_FrameData[31]
port 121 nsew signal input
rlabel metal3 s -300 78072 160 78192 4 Tile_X0Y0_FrameData[3]
port 122 nsew signal input
rlabel metal3 s -300 78344 160 78464 4 Tile_X0Y0_FrameData[4]
port 123 nsew signal input
rlabel metal3 s -300 78616 160 78736 4 Tile_X0Y0_FrameData[5]
port 124 nsew signal input
rlabel metal3 s -300 78888 160 79008 4 Tile_X0Y0_FrameData[6]
port 125 nsew signal input
rlabel metal3 s -300 79160 160 79280 4 Tile_X0Y0_FrameData[7]
port 126 nsew signal input
rlabel metal3 s -300 79432 160 79552 4 Tile_X0Y0_FrameData[8]
port 127 nsew signal input
rlabel metal3 s -300 79704 160 79824 4 Tile_X0Y0_FrameData[9]
port 128 nsew signal input
rlabel metal3 s 44540 77256 45000 77376 6 Tile_X0Y0_FrameData_O[0]
port 129 nsew signal output
rlabel metal3 s 44540 79976 45000 80096 6 Tile_X0Y0_FrameData_O[10]
port 130 nsew signal output
rlabel metal3 s 44540 80248 45000 80368 6 Tile_X0Y0_FrameData_O[11]
port 131 nsew signal output
rlabel metal3 s 44540 80520 45000 80640 6 Tile_X0Y0_FrameData_O[12]
port 132 nsew signal output
rlabel metal3 s 44540 80792 45000 80912 6 Tile_X0Y0_FrameData_O[13]
port 133 nsew signal output
rlabel metal3 s 44540 81064 45000 81184 6 Tile_X0Y0_FrameData_O[14]
port 134 nsew signal output
rlabel metal3 s 44540 81336 45000 81456 6 Tile_X0Y0_FrameData_O[15]
port 135 nsew signal output
rlabel metal3 s 44540 81608 45000 81728 6 Tile_X0Y0_FrameData_O[16]
port 136 nsew signal output
rlabel metal3 s 44540 81880 45000 82000 6 Tile_X0Y0_FrameData_O[17]
port 137 nsew signal output
rlabel metal3 s 44540 82152 45000 82272 6 Tile_X0Y0_FrameData_O[18]
port 138 nsew signal output
rlabel metal3 s 44540 82424 45000 82544 6 Tile_X0Y0_FrameData_O[19]
port 139 nsew signal output
rlabel metal3 s 44540 77528 45000 77648 6 Tile_X0Y0_FrameData_O[1]
port 140 nsew signal output
rlabel metal3 s 44540 82696 45000 82816 6 Tile_X0Y0_FrameData_O[20]
port 141 nsew signal output
rlabel metal3 s 44540 82968 45000 83088 6 Tile_X0Y0_FrameData_O[21]
port 142 nsew signal output
rlabel metal3 s 44540 83240 45000 83360 6 Tile_X0Y0_FrameData_O[22]
port 143 nsew signal output
rlabel metal3 s 44540 83512 45000 83632 6 Tile_X0Y0_FrameData_O[23]
port 144 nsew signal output
rlabel metal3 s 44540 83784 45000 83904 6 Tile_X0Y0_FrameData_O[24]
port 145 nsew signal output
rlabel metal3 s 44540 84056 45000 84176 6 Tile_X0Y0_FrameData_O[25]
port 146 nsew signal output
rlabel metal3 s 44540 84328 45000 84448 6 Tile_X0Y0_FrameData_O[26]
port 147 nsew signal output
rlabel metal3 s 44540 84600 45000 84720 6 Tile_X0Y0_FrameData_O[27]
port 148 nsew signal output
rlabel metal3 s 44540 84872 45000 84992 6 Tile_X0Y0_FrameData_O[28]
port 149 nsew signal output
rlabel metal3 s 44540 85144 45000 85264 6 Tile_X0Y0_FrameData_O[29]
port 150 nsew signal output
rlabel metal3 s 44540 77800 45000 77920 6 Tile_X0Y0_FrameData_O[2]
port 151 nsew signal output
rlabel metal3 s 44540 85416 45000 85536 6 Tile_X0Y0_FrameData_O[30]
port 152 nsew signal output
rlabel metal3 s 44540 85688 45000 85808 6 Tile_X0Y0_FrameData_O[31]
port 153 nsew signal output
rlabel metal3 s 44540 78072 45000 78192 6 Tile_X0Y0_FrameData_O[3]
port 154 nsew signal output
rlabel metal3 s 44540 78344 45000 78464 6 Tile_X0Y0_FrameData_O[4]
port 155 nsew signal output
rlabel metal3 s 44540 78616 45000 78736 6 Tile_X0Y0_FrameData_O[5]
port 156 nsew signal output
rlabel metal3 s 44540 78888 45000 79008 6 Tile_X0Y0_FrameData_O[6]
port 157 nsew signal output
rlabel metal3 s 44540 79160 45000 79280 6 Tile_X0Y0_FrameData_O[7]
port 158 nsew signal output
rlabel metal3 s 44540 79432 45000 79552 6 Tile_X0Y0_FrameData_O[8]
port 159 nsew signal output
rlabel metal3 s 44540 79704 45000 79824 6 Tile_X0Y0_FrameData_O[9]
port 160 nsew signal output
rlabel metal2 s 34150 90540 34206 91000 6 Tile_X0Y0_FrameStrobe_O[0]
port 161 nsew signal output
rlabel metal2 s 36910 90540 36966 91000 6 Tile_X0Y0_FrameStrobe_O[10]
port 162 nsew signal output
rlabel metal2 s 37186 90540 37242 91000 6 Tile_X0Y0_FrameStrobe_O[11]
port 163 nsew signal output
rlabel metal2 s 37462 90540 37518 91000 6 Tile_X0Y0_FrameStrobe_O[12]
port 164 nsew signal output
rlabel metal2 s 37738 90540 37794 91000 6 Tile_X0Y0_FrameStrobe_O[13]
port 165 nsew signal output
rlabel metal2 s 38014 90540 38070 91000 6 Tile_X0Y0_FrameStrobe_O[14]
port 166 nsew signal output
rlabel metal2 s 38290 90540 38346 91000 6 Tile_X0Y0_FrameStrobe_O[15]
port 167 nsew signal output
rlabel metal2 s 38566 90540 38622 91000 6 Tile_X0Y0_FrameStrobe_O[16]
port 168 nsew signal output
rlabel metal2 s 38842 90540 38898 91000 6 Tile_X0Y0_FrameStrobe_O[17]
port 169 nsew signal output
rlabel metal2 s 39118 90540 39174 91000 6 Tile_X0Y0_FrameStrobe_O[18]
port 170 nsew signal output
rlabel metal2 s 39394 90540 39450 91000 6 Tile_X0Y0_FrameStrobe_O[19]
port 171 nsew signal output
rlabel metal2 s 34426 90540 34482 91000 6 Tile_X0Y0_FrameStrobe_O[1]
port 172 nsew signal output
rlabel metal2 s 34702 90540 34758 91000 6 Tile_X0Y0_FrameStrobe_O[2]
port 173 nsew signal output
rlabel metal2 s 34978 90540 35034 91000 6 Tile_X0Y0_FrameStrobe_O[3]
port 174 nsew signal output
rlabel metal2 s 35254 90540 35310 91000 6 Tile_X0Y0_FrameStrobe_O[4]
port 175 nsew signal output
rlabel metal2 s 35530 90540 35586 91000 6 Tile_X0Y0_FrameStrobe_O[5]
port 176 nsew signal output
rlabel metal2 s 35806 90540 35862 91000 6 Tile_X0Y0_FrameStrobe_O[6]
port 177 nsew signal output
rlabel metal2 s 36082 90540 36138 91000 6 Tile_X0Y0_FrameStrobe_O[7]
port 178 nsew signal output
rlabel metal2 s 36358 90540 36414 91000 6 Tile_X0Y0_FrameStrobe_O[8]
port 179 nsew signal output
rlabel metal2 s 36634 90540 36690 91000 6 Tile_X0Y0_FrameStrobe_O[9]
port 180 nsew signal output
rlabel metal2 s 5170 90540 5226 91000 6 Tile_X0Y0_N1BEG[0]
port 181 nsew signal output
rlabel metal2 s 5446 90540 5502 91000 6 Tile_X0Y0_N1BEG[1]
port 182 nsew signal output
rlabel metal2 s 5722 90540 5778 91000 6 Tile_X0Y0_N1BEG[2]
port 183 nsew signal output
rlabel metal2 s 5998 90540 6054 91000 6 Tile_X0Y0_N1BEG[3]
port 184 nsew signal output
rlabel metal2 s 6274 90540 6330 91000 6 Tile_X0Y0_N2BEG[0]
port 185 nsew signal output
rlabel metal2 s 6550 90540 6606 91000 6 Tile_X0Y0_N2BEG[1]
port 186 nsew signal output
rlabel metal2 s 6826 90540 6882 91000 6 Tile_X0Y0_N2BEG[2]
port 187 nsew signal output
rlabel metal2 s 7102 90540 7158 91000 6 Tile_X0Y0_N2BEG[3]
port 188 nsew signal output
rlabel metal2 s 7378 90540 7434 91000 6 Tile_X0Y0_N2BEG[4]
port 189 nsew signal output
rlabel metal2 s 7654 90540 7710 91000 6 Tile_X0Y0_N2BEG[5]
port 190 nsew signal output
rlabel metal2 s 7930 90540 7986 91000 6 Tile_X0Y0_N2BEG[6]
port 191 nsew signal output
rlabel metal2 s 8206 90540 8262 91000 6 Tile_X0Y0_N2BEG[7]
port 192 nsew signal output
rlabel metal2 s 8482 90540 8538 91000 6 Tile_X0Y0_N2BEGb[0]
port 193 nsew signal output
rlabel metal2 s 8758 90540 8814 91000 6 Tile_X0Y0_N2BEGb[1]
port 194 nsew signal output
rlabel metal2 s 9034 90540 9090 91000 6 Tile_X0Y0_N2BEGb[2]
port 195 nsew signal output
rlabel metal2 s 9310 90540 9366 91000 6 Tile_X0Y0_N2BEGb[3]
port 196 nsew signal output
rlabel metal2 s 9586 90540 9642 91000 6 Tile_X0Y0_N2BEGb[4]
port 197 nsew signal output
rlabel metal2 s 9862 90540 9918 91000 6 Tile_X0Y0_N2BEGb[5]
port 198 nsew signal output
rlabel metal2 s 10138 90540 10194 91000 6 Tile_X0Y0_N2BEGb[6]
port 199 nsew signal output
rlabel metal2 s 10414 90540 10470 91000 6 Tile_X0Y0_N2BEGb[7]
port 200 nsew signal output
rlabel metal2 s 10690 90540 10746 91000 6 Tile_X0Y0_N4BEG[0]
port 201 nsew signal output
rlabel metal2 s 13450 90540 13506 91000 6 Tile_X0Y0_N4BEG[10]
port 202 nsew signal output
rlabel metal2 s 13726 90540 13782 91000 6 Tile_X0Y0_N4BEG[11]
port 203 nsew signal output
rlabel metal2 s 14002 90540 14058 91000 6 Tile_X0Y0_N4BEG[12]
port 204 nsew signal output
rlabel metal2 s 14278 90540 14334 91000 6 Tile_X0Y0_N4BEG[13]
port 205 nsew signal output
rlabel metal2 s 14554 90540 14610 91000 6 Tile_X0Y0_N4BEG[14]
port 206 nsew signal output
rlabel metal2 s 14830 90540 14886 91000 6 Tile_X0Y0_N4BEG[15]
port 207 nsew signal output
rlabel metal2 s 10966 90540 11022 91000 6 Tile_X0Y0_N4BEG[1]
port 208 nsew signal output
rlabel metal2 s 11242 90540 11298 91000 6 Tile_X0Y0_N4BEG[2]
port 209 nsew signal output
rlabel metal2 s 11518 90540 11574 91000 6 Tile_X0Y0_N4BEG[3]
port 210 nsew signal output
rlabel metal2 s 11794 90540 11850 91000 6 Tile_X0Y0_N4BEG[4]
port 211 nsew signal output
rlabel metal2 s 12070 90540 12126 91000 6 Tile_X0Y0_N4BEG[5]
port 212 nsew signal output
rlabel metal2 s 12346 90540 12402 91000 6 Tile_X0Y0_N4BEG[6]
port 213 nsew signal output
rlabel metal2 s 12622 90540 12678 91000 6 Tile_X0Y0_N4BEG[7]
port 214 nsew signal output
rlabel metal2 s 12898 90540 12954 91000 6 Tile_X0Y0_N4BEG[8]
port 215 nsew signal output
rlabel metal2 s 13174 90540 13230 91000 6 Tile_X0Y0_N4BEG[9]
port 216 nsew signal output
rlabel metal2 s 15106 90540 15162 91000 6 Tile_X0Y0_NN4BEG[0]
port 217 nsew signal output
rlabel metal2 s 17866 90540 17922 91000 6 Tile_X0Y0_NN4BEG[10]
port 218 nsew signal output
rlabel metal2 s 18142 90540 18198 91000 6 Tile_X0Y0_NN4BEG[11]
port 219 nsew signal output
rlabel metal2 s 18418 90540 18474 91000 6 Tile_X0Y0_NN4BEG[12]
port 220 nsew signal output
rlabel metal2 s 18694 90540 18750 91000 6 Tile_X0Y0_NN4BEG[13]
port 221 nsew signal output
rlabel metal2 s 18970 90540 19026 91000 6 Tile_X0Y0_NN4BEG[14]
port 222 nsew signal output
rlabel metal2 s 19246 90540 19302 91000 6 Tile_X0Y0_NN4BEG[15]
port 223 nsew signal output
rlabel metal2 s 15382 90540 15438 91000 6 Tile_X0Y0_NN4BEG[1]
port 224 nsew signal output
rlabel metal2 s 15658 90540 15714 91000 6 Tile_X0Y0_NN4BEG[2]
port 225 nsew signal output
rlabel metal2 s 15934 90540 15990 91000 6 Tile_X0Y0_NN4BEG[3]
port 226 nsew signal output
rlabel metal2 s 16210 90540 16266 91000 6 Tile_X0Y0_NN4BEG[4]
port 227 nsew signal output
rlabel metal2 s 16486 90540 16542 91000 6 Tile_X0Y0_NN4BEG[5]
port 228 nsew signal output
rlabel metal2 s 16762 90540 16818 91000 6 Tile_X0Y0_NN4BEG[6]
port 229 nsew signal output
rlabel metal2 s 17038 90540 17094 91000 6 Tile_X0Y0_NN4BEG[7]
port 230 nsew signal output
rlabel metal2 s 17314 90540 17370 91000 6 Tile_X0Y0_NN4BEG[8]
port 231 nsew signal output
rlabel metal2 s 17590 90540 17646 91000 6 Tile_X0Y0_NN4BEG[9]
port 232 nsew signal output
rlabel metal2 s 19522 90540 19578 91000 6 Tile_X0Y0_S1END[0]
port 233 nsew signal input
rlabel metal2 s 19798 90540 19854 91000 6 Tile_X0Y0_S1END[1]
port 234 nsew signal input
rlabel metal2 s 20074 90540 20130 91000 6 Tile_X0Y0_S1END[2]
port 235 nsew signal input
rlabel metal2 s 20350 90540 20406 91000 6 Tile_X0Y0_S1END[3]
port 236 nsew signal input
rlabel metal2 s 20626 90540 20682 91000 6 Tile_X0Y0_S2END[0]
port 237 nsew signal input
rlabel metal2 s 20902 90540 20958 91000 6 Tile_X0Y0_S2END[1]
port 238 nsew signal input
rlabel metal2 s 21178 90540 21234 91000 6 Tile_X0Y0_S2END[2]
port 239 nsew signal input
rlabel metal2 s 21454 90540 21510 91000 6 Tile_X0Y0_S2END[3]
port 240 nsew signal input
rlabel metal2 s 21730 90540 21786 91000 6 Tile_X0Y0_S2END[4]
port 241 nsew signal input
rlabel metal2 s 22006 90540 22062 91000 6 Tile_X0Y0_S2END[5]
port 242 nsew signal input
rlabel metal2 s 22282 90540 22338 91000 6 Tile_X0Y0_S2END[6]
port 243 nsew signal input
rlabel metal2 s 22558 90540 22614 91000 6 Tile_X0Y0_S2END[7]
port 244 nsew signal input
rlabel metal2 s 22834 90540 22890 91000 6 Tile_X0Y0_S2MID[0]
port 245 nsew signal input
rlabel metal2 s 23110 90540 23166 91000 6 Tile_X0Y0_S2MID[1]
port 246 nsew signal input
rlabel metal2 s 23386 90540 23442 91000 6 Tile_X0Y0_S2MID[2]
port 247 nsew signal input
rlabel metal2 s 23662 90540 23718 91000 6 Tile_X0Y0_S2MID[3]
port 248 nsew signal input
rlabel metal2 s 23938 90540 23994 91000 6 Tile_X0Y0_S2MID[4]
port 249 nsew signal input
rlabel metal2 s 24214 90540 24270 91000 6 Tile_X0Y0_S2MID[5]
port 250 nsew signal input
rlabel metal2 s 24490 90540 24546 91000 6 Tile_X0Y0_S2MID[6]
port 251 nsew signal input
rlabel metal2 s 24766 90540 24822 91000 6 Tile_X0Y0_S2MID[7]
port 252 nsew signal input
rlabel metal2 s 25042 90540 25098 91000 6 Tile_X0Y0_S4END[0]
port 253 nsew signal input
rlabel metal2 s 27802 90540 27858 91000 6 Tile_X0Y0_S4END[10]
port 254 nsew signal input
rlabel metal2 s 28078 90540 28134 91000 6 Tile_X0Y0_S4END[11]
port 255 nsew signal input
rlabel metal2 s 28354 90540 28410 91000 6 Tile_X0Y0_S4END[12]
port 256 nsew signal input
rlabel metal2 s 28630 90540 28686 91000 6 Tile_X0Y0_S4END[13]
port 257 nsew signal input
rlabel metal2 s 28906 90540 28962 91000 6 Tile_X0Y0_S4END[14]
port 258 nsew signal input
rlabel metal2 s 29182 90540 29238 91000 6 Tile_X0Y0_S4END[15]
port 259 nsew signal input
rlabel metal2 s 25318 90540 25374 91000 6 Tile_X0Y0_S4END[1]
port 260 nsew signal input
rlabel metal2 s 25594 90540 25650 91000 6 Tile_X0Y0_S4END[2]
port 261 nsew signal input
rlabel metal2 s 25870 90540 25926 91000 6 Tile_X0Y0_S4END[3]
port 262 nsew signal input
rlabel metal2 s 26146 90540 26202 91000 6 Tile_X0Y0_S4END[4]
port 263 nsew signal input
rlabel metal2 s 26422 90540 26478 91000 6 Tile_X0Y0_S4END[5]
port 264 nsew signal input
rlabel metal2 s 26698 90540 26754 91000 6 Tile_X0Y0_S4END[6]
port 265 nsew signal input
rlabel metal2 s 26974 90540 27030 91000 6 Tile_X0Y0_S4END[7]
port 266 nsew signal input
rlabel metal2 s 27250 90540 27306 91000 6 Tile_X0Y0_S4END[8]
port 267 nsew signal input
rlabel metal2 s 27526 90540 27582 91000 6 Tile_X0Y0_S4END[9]
port 268 nsew signal input
rlabel metal2 s 29458 90540 29514 91000 6 Tile_X0Y0_SS4END[0]
port 269 nsew signal input
rlabel metal2 s 32218 90540 32274 91000 6 Tile_X0Y0_SS4END[10]
port 270 nsew signal input
rlabel metal2 s 32494 90540 32550 91000 6 Tile_X0Y0_SS4END[11]
port 271 nsew signal input
rlabel metal2 s 32770 90540 32826 91000 6 Tile_X0Y0_SS4END[12]
port 272 nsew signal input
rlabel metal2 s 33046 90540 33102 91000 6 Tile_X0Y0_SS4END[13]
port 273 nsew signal input
rlabel metal2 s 33322 90540 33378 91000 6 Tile_X0Y0_SS4END[14]
port 274 nsew signal input
rlabel metal2 s 33598 90540 33654 91000 6 Tile_X0Y0_SS4END[15]
port 275 nsew signal input
rlabel metal2 s 29734 90540 29790 91000 6 Tile_X0Y0_SS4END[1]
port 276 nsew signal input
rlabel metal2 s 30010 90540 30066 91000 6 Tile_X0Y0_SS4END[2]
port 277 nsew signal input
rlabel metal2 s 30286 90540 30342 91000 6 Tile_X0Y0_SS4END[3]
port 278 nsew signal input
rlabel metal2 s 30562 90540 30618 91000 6 Tile_X0Y0_SS4END[4]
port 279 nsew signal input
rlabel metal2 s 30838 90540 30894 91000 6 Tile_X0Y0_SS4END[5]
port 280 nsew signal input
rlabel metal2 s 31114 90540 31170 91000 6 Tile_X0Y0_SS4END[6]
port 281 nsew signal input
rlabel metal2 s 31390 90540 31446 91000 6 Tile_X0Y0_SS4END[7]
port 282 nsew signal input
rlabel metal2 s 31666 90540 31722 91000 6 Tile_X0Y0_SS4END[8]
port 283 nsew signal input
rlabel metal2 s 31942 90540 31998 91000 6 Tile_X0Y0_SS4END[9]
port 284 nsew signal input
rlabel metal2 s 33874 90540 33930 91000 6 Tile_X0Y0_UserCLKo
port 285 nsew signal output
rlabel metal3 s -300 51144 160 51264 4 Tile_X0Y0_W1BEG[0]
port 286 nsew signal output
rlabel metal3 s -300 51416 160 51536 4 Tile_X0Y0_W1BEG[1]
port 287 nsew signal output
rlabel metal3 s -300 51688 160 51808 4 Tile_X0Y0_W1BEG[2]
port 288 nsew signal output
rlabel metal3 s -300 51960 160 52080 4 Tile_X0Y0_W1BEG[3]
port 289 nsew signal output
rlabel metal3 s 44540 51144 45000 51264 6 Tile_X0Y0_W1END[0]
port 290 nsew signal input
rlabel metal3 s 44540 51416 45000 51536 6 Tile_X0Y0_W1END[1]
port 291 nsew signal input
rlabel metal3 s 44540 51688 45000 51808 6 Tile_X0Y0_W1END[2]
port 292 nsew signal input
rlabel metal3 s 44540 51960 45000 52080 6 Tile_X0Y0_W1END[3]
port 293 nsew signal input
rlabel metal3 s -300 52232 160 52352 4 Tile_X0Y0_W2BEG[0]
port 294 nsew signal output
rlabel metal3 s -300 52504 160 52624 4 Tile_X0Y0_W2BEG[1]
port 295 nsew signal output
rlabel metal3 s -300 52776 160 52896 4 Tile_X0Y0_W2BEG[2]
port 296 nsew signal output
rlabel metal3 s -300 53048 160 53168 4 Tile_X0Y0_W2BEG[3]
port 297 nsew signal output
rlabel metal3 s -300 53320 160 53440 4 Tile_X0Y0_W2BEG[4]
port 298 nsew signal output
rlabel metal3 s -300 53592 160 53712 4 Tile_X0Y0_W2BEG[5]
port 299 nsew signal output
rlabel metal3 s -300 53864 160 53984 4 Tile_X0Y0_W2BEG[6]
port 300 nsew signal output
rlabel metal3 s -300 54136 160 54256 4 Tile_X0Y0_W2BEG[7]
port 301 nsew signal output
rlabel metal3 s -300 54408 160 54528 4 Tile_X0Y0_W2BEGb[0]
port 302 nsew signal output
rlabel metal3 s -300 54680 160 54800 4 Tile_X0Y0_W2BEGb[1]
port 303 nsew signal output
rlabel metal3 s -300 54952 160 55072 4 Tile_X0Y0_W2BEGb[2]
port 304 nsew signal output
rlabel metal3 s -300 55224 160 55344 4 Tile_X0Y0_W2BEGb[3]
port 305 nsew signal output
rlabel metal3 s -300 55496 160 55616 4 Tile_X0Y0_W2BEGb[4]
port 306 nsew signal output
rlabel metal3 s -300 55768 160 55888 4 Tile_X0Y0_W2BEGb[5]
port 307 nsew signal output
rlabel metal3 s -300 56040 160 56160 4 Tile_X0Y0_W2BEGb[6]
port 308 nsew signal output
rlabel metal3 s -300 56312 160 56432 4 Tile_X0Y0_W2BEGb[7]
port 309 nsew signal output
rlabel metal3 s 44540 54408 45000 54528 6 Tile_X0Y0_W2END[0]
port 310 nsew signal input
rlabel metal3 s 44540 54680 45000 54800 6 Tile_X0Y0_W2END[1]
port 311 nsew signal input
rlabel metal3 s 44540 54952 45000 55072 6 Tile_X0Y0_W2END[2]
port 312 nsew signal input
rlabel metal3 s 44540 55224 45000 55344 6 Tile_X0Y0_W2END[3]
port 313 nsew signal input
rlabel metal3 s 44540 55496 45000 55616 6 Tile_X0Y0_W2END[4]
port 314 nsew signal input
rlabel metal3 s 44540 55768 45000 55888 6 Tile_X0Y0_W2END[5]
port 315 nsew signal input
rlabel metal3 s 44540 56040 45000 56160 6 Tile_X0Y0_W2END[6]
port 316 nsew signal input
rlabel metal3 s 44540 56312 45000 56432 6 Tile_X0Y0_W2END[7]
port 317 nsew signal input
rlabel metal3 s 44540 52232 45000 52352 6 Tile_X0Y0_W2MID[0]
port 318 nsew signal input
rlabel metal3 s 44540 52504 45000 52624 6 Tile_X0Y0_W2MID[1]
port 319 nsew signal input
rlabel metal3 s 44540 52776 45000 52896 6 Tile_X0Y0_W2MID[2]
port 320 nsew signal input
rlabel metal3 s 44540 53048 45000 53168 6 Tile_X0Y0_W2MID[3]
port 321 nsew signal input
rlabel metal3 s 44540 53320 45000 53440 6 Tile_X0Y0_W2MID[4]
port 322 nsew signal input
rlabel metal3 s 44540 53592 45000 53712 6 Tile_X0Y0_W2MID[5]
port 323 nsew signal input
rlabel metal3 s 44540 53864 45000 53984 6 Tile_X0Y0_W2MID[6]
port 324 nsew signal input
rlabel metal3 s 44540 54136 45000 54256 6 Tile_X0Y0_W2MID[7]
port 325 nsew signal input
rlabel metal3 s -300 60936 160 61056 4 Tile_X0Y0_W6BEG[0]
port 326 nsew signal output
rlabel metal3 s -300 63656 160 63776 4 Tile_X0Y0_W6BEG[10]
port 327 nsew signal output
rlabel metal3 s -300 63928 160 64048 4 Tile_X0Y0_W6BEG[11]
port 328 nsew signal output
rlabel metal3 s -300 61208 160 61328 4 Tile_X0Y0_W6BEG[1]
port 329 nsew signal output
rlabel metal3 s -300 61480 160 61600 4 Tile_X0Y0_W6BEG[2]
port 330 nsew signal output
rlabel metal3 s -300 61752 160 61872 4 Tile_X0Y0_W6BEG[3]
port 331 nsew signal output
rlabel metal3 s -300 62024 160 62144 4 Tile_X0Y0_W6BEG[4]
port 332 nsew signal output
rlabel metal3 s -300 62296 160 62416 4 Tile_X0Y0_W6BEG[5]
port 333 nsew signal output
rlabel metal3 s -300 62568 160 62688 4 Tile_X0Y0_W6BEG[6]
port 334 nsew signal output
rlabel metal3 s -300 62840 160 62960 4 Tile_X0Y0_W6BEG[7]
port 335 nsew signal output
rlabel metal3 s -300 63112 160 63232 4 Tile_X0Y0_W6BEG[8]
port 336 nsew signal output
rlabel metal3 s -300 63384 160 63504 4 Tile_X0Y0_W6BEG[9]
port 337 nsew signal output
rlabel metal3 s 44540 60936 45000 61056 6 Tile_X0Y0_W6END[0]
port 338 nsew signal input
rlabel metal3 s 44540 63656 45000 63776 6 Tile_X0Y0_W6END[10]
port 339 nsew signal input
rlabel metal3 s 44540 63928 45000 64048 6 Tile_X0Y0_W6END[11]
port 340 nsew signal input
rlabel metal3 s 44540 61208 45000 61328 6 Tile_X0Y0_W6END[1]
port 341 nsew signal input
rlabel metal3 s 44540 61480 45000 61600 6 Tile_X0Y0_W6END[2]
port 342 nsew signal input
rlabel metal3 s 44540 61752 45000 61872 6 Tile_X0Y0_W6END[3]
port 343 nsew signal input
rlabel metal3 s 44540 62024 45000 62144 6 Tile_X0Y0_W6END[4]
port 344 nsew signal input
rlabel metal3 s 44540 62296 45000 62416 6 Tile_X0Y0_W6END[5]
port 345 nsew signal input
rlabel metal3 s 44540 62568 45000 62688 6 Tile_X0Y0_W6END[6]
port 346 nsew signal input
rlabel metal3 s 44540 62840 45000 62960 6 Tile_X0Y0_W6END[7]
port 347 nsew signal input
rlabel metal3 s 44540 63112 45000 63232 6 Tile_X0Y0_W6END[8]
port 348 nsew signal input
rlabel metal3 s 44540 63384 45000 63504 6 Tile_X0Y0_W6END[9]
port 349 nsew signal input
rlabel metal3 s -300 56584 160 56704 4 Tile_X0Y0_WW4BEG[0]
port 350 nsew signal output
rlabel metal3 s -300 59304 160 59424 4 Tile_X0Y0_WW4BEG[10]
port 351 nsew signal output
rlabel metal3 s -300 59576 160 59696 4 Tile_X0Y0_WW4BEG[11]
port 352 nsew signal output
rlabel metal3 s -300 59848 160 59968 4 Tile_X0Y0_WW4BEG[12]
port 353 nsew signal output
rlabel metal3 s -300 60120 160 60240 4 Tile_X0Y0_WW4BEG[13]
port 354 nsew signal output
rlabel metal3 s -300 60392 160 60512 4 Tile_X0Y0_WW4BEG[14]
port 355 nsew signal output
rlabel metal3 s -300 60664 160 60784 4 Tile_X0Y0_WW4BEG[15]
port 356 nsew signal output
rlabel metal3 s -300 56856 160 56976 4 Tile_X0Y0_WW4BEG[1]
port 357 nsew signal output
rlabel metal3 s -300 57128 160 57248 4 Tile_X0Y0_WW4BEG[2]
port 358 nsew signal output
rlabel metal3 s -300 57400 160 57520 4 Tile_X0Y0_WW4BEG[3]
port 359 nsew signal output
rlabel metal3 s -300 57672 160 57792 4 Tile_X0Y0_WW4BEG[4]
port 360 nsew signal output
rlabel metal3 s -300 57944 160 58064 4 Tile_X0Y0_WW4BEG[5]
port 361 nsew signal output
rlabel metal3 s -300 58216 160 58336 4 Tile_X0Y0_WW4BEG[6]
port 362 nsew signal output
rlabel metal3 s -300 58488 160 58608 4 Tile_X0Y0_WW4BEG[7]
port 363 nsew signal output
rlabel metal3 s -300 58760 160 58880 4 Tile_X0Y0_WW4BEG[8]
port 364 nsew signal output
rlabel metal3 s -300 59032 160 59152 4 Tile_X0Y0_WW4BEG[9]
port 365 nsew signal output
rlabel metal3 s 44540 56584 45000 56704 6 Tile_X0Y0_WW4END[0]
port 366 nsew signal input
rlabel metal3 s 44540 59304 45000 59424 6 Tile_X0Y0_WW4END[10]
port 367 nsew signal input
rlabel metal3 s 44540 59576 45000 59696 6 Tile_X0Y0_WW4END[11]
port 368 nsew signal input
rlabel metal3 s 44540 59848 45000 59968 6 Tile_X0Y0_WW4END[12]
port 369 nsew signal input
rlabel metal3 s 44540 60120 45000 60240 6 Tile_X0Y0_WW4END[13]
port 370 nsew signal input
rlabel metal3 s 44540 60392 45000 60512 6 Tile_X0Y0_WW4END[14]
port 371 nsew signal input
rlabel metal3 s 44540 60664 45000 60784 6 Tile_X0Y0_WW4END[15]
port 372 nsew signal input
rlabel metal3 s 44540 56856 45000 56976 6 Tile_X0Y0_WW4END[1]
port 373 nsew signal input
rlabel metal3 s 44540 57128 45000 57248 6 Tile_X0Y0_WW4END[2]
port 374 nsew signal input
rlabel metal3 s 44540 57400 45000 57520 6 Tile_X0Y0_WW4END[3]
port 375 nsew signal input
rlabel metal3 s 44540 57672 45000 57792 6 Tile_X0Y0_WW4END[4]
port 376 nsew signal input
rlabel metal3 s 44540 57944 45000 58064 6 Tile_X0Y0_WW4END[5]
port 377 nsew signal input
rlabel metal3 s 44540 58216 45000 58336 6 Tile_X0Y0_WW4END[6]
port 378 nsew signal input
rlabel metal3 s 44540 58488 45000 58608 6 Tile_X0Y0_WW4END[7]
port 379 nsew signal input
rlabel metal3 s 44540 58760 45000 58880 6 Tile_X0Y0_WW4END[8]
port 380 nsew signal input
rlabel metal3 s 44540 59032 45000 59152 6 Tile_X0Y0_WW4END[9]
port 381 nsew signal input
rlabel metal3 s 44540 18232 45000 18352 6 Tile_X0Y1_E1BEG[0]
port 382 nsew signal output
rlabel metal3 s 44540 18504 45000 18624 6 Tile_X0Y1_E1BEG[1]
port 383 nsew signal output
rlabel metal3 s 44540 18776 45000 18896 6 Tile_X0Y1_E1BEG[2]
port 384 nsew signal output
rlabel metal3 s 44540 19048 45000 19168 6 Tile_X0Y1_E1BEG[3]
port 385 nsew signal output
rlabel metal3 s -300 18232 160 18352 4 Tile_X0Y1_E1END[0]
port 386 nsew signal input
rlabel metal3 s -300 18504 160 18624 4 Tile_X0Y1_E1END[1]
port 387 nsew signal input
rlabel metal3 s -300 18776 160 18896 4 Tile_X0Y1_E1END[2]
port 388 nsew signal input
rlabel metal3 s -300 19048 160 19168 4 Tile_X0Y1_E1END[3]
port 389 nsew signal input
rlabel metal3 s 44540 19320 45000 19440 6 Tile_X0Y1_E2BEG[0]
port 390 nsew signal output
rlabel metal3 s 44540 19592 45000 19712 6 Tile_X0Y1_E2BEG[1]
port 391 nsew signal output
rlabel metal3 s 44540 19864 45000 19984 6 Tile_X0Y1_E2BEG[2]
port 392 nsew signal output
rlabel metal3 s 44540 20136 45000 20256 6 Tile_X0Y1_E2BEG[3]
port 393 nsew signal output
rlabel metal3 s 44540 20408 45000 20528 6 Tile_X0Y1_E2BEG[4]
port 394 nsew signal output
rlabel metal3 s 44540 20680 45000 20800 6 Tile_X0Y1_E2BEG[5]
port 395 nsew signal output
rlabel metal3 s 44540 20952 45000 21072 6 Tile_X0Y1_E2BEG[6]
port 396 nsew signal output
rlabel metal3 s 44540 21224 45000 21344 6 Tile_X0Y1_E2BEG[7]
port 397 nsew signal output
rlabel metal3 s 44540 21496 45000 21616 6 Tile_X0Y1_E2BEGb[0]
port 398 nsew signal output
rlabel metal3 s 44540 21768 45000 21888 6 Tile_X0Y1_E2BEGb[1]
port 399 nsew signal output
rlabel metal3 s 44540 22040 45000 22160 6 Tile_X0Y1_E2BEGb[2]
port 400 nsew signal output
rlabel metal3 s 44540 22312 45000 22432 6 Tile_X0Y1_E2BEGb[3]
port 401 nsew signal output
rlabel metal3 s 44540 22584 45000 22704 6 Tile_X0Y1_E2BEGb[4]
port 402 nsew signal output
rlabel metal3 s 44540 22856 45000 22976 6 Tile_X0Y1_E2BEGb[5]
port 403 nsew signal output
rlabel metal3 s 44540 23128 45000 23248 6 Tile_X0Y1_E2BEGb[6]
port 404 nsew signal output
rlabel metal3 s 44540 23400 45000 23520 6 Tile_X0Y1_E2BEGb[7]
port 405 nsew signal output
rlabel metal3 s -300 21496 160 21616 4 Tile_X0Y1_E2END[0]
port 406 nsew signal input
rlabel metal3 s -300 21768 160 21888 4 Tile_X0Y1_E2END[1]
port 407 nsew signal input
rlabel metal3 s -300 22040 160 22160 4 Tile_X0Y1_E2END[2]
port 408 nsew signal input
rlabel metal3 s -300 22312 160 22432 4 Tile_X0Y1_E2END[3]
port 409 nsew signal input
rlabel metal3 s -300 22584 160 22704 4 Tile_X0Y1_E2END[4]
port 410 nsew signal input
rlabel metal3 s -300 22856 160 22976 4 Tile_X0Y1_E2END[5]
port 411 nsew signal input
rlabel metal3 s -300 23128 160 23248 4 Tile_X0Y1_E2END[6]
port 412 nsew signal input
rlabel metal3 s -300 23400 160 23520 4 Tile_X0Y1_E2END[7]
port 413 nsew signal input
rlabel metal3 s -300 19320 160 19440 4 Tile_X0Y1_E2MID[0]
port 414 nsew signal input
rlabel metal3 s -300 19592 160 19712 4 Tile_X0Y1_E2MID[1]
port 415 nsew signal input
rlabel metal3 s -300 19864 160 19984 4 Tile_X0Y1_E2MID[2]
port 416 nsew signal input
rlabel metal3 s -300 20136 160 20256 4 Tile_X0Y1_E2MID[3]
port 417 nsew signal input
rlabel metal3 s -300 20408 160 20528 4 Tile_X0Y1_E2MID[4]
port 418 nsew signal input
rlabel metal3 s -300 20680 160 20800 4 Tile_X0Y1_E2MID[5]
port 419 nsew signal input
rlabel metal3 s -300 20952 160 21072 4 Tile_X0Y1_E2MID[6]
port 420 nsew signal input
rlabel metal3 s -300 21224 160 21344 4 Tile_X0Y1_E2MID[7]
port 421 nsew signal input
rlabel metal3 s 44540 28024 45000 28144 6 Tile_X0Y1_E6BEG[0]
port 422 nsew signal output
rlabel metal3 s 44540 30744 45000 30864 6 Tile_X0Y1_E6BEG[10]
port 423 nsew signal output
rlabel metal3 s 44540 31016 45000 31136 6 Tile_X0Y1_E6BEG[11]
port 424 nsew signal output
rlabel metal3 s 44540 28296 45000 28416 6 Tile_X0Y1_E6BEG[1]
port 425 nsew signal output
rlabel metal3 s 44540 28568 45000 28688 6 Tile_X0Y1_E6BEG[2]
port 426 nsew signal output
rlabel metal3 s 44540 28840 45000 28960 6 Tile_X0Y1_E6BEG[3]
port 427 nsew signal output
rlabel metal3 s 44540 29112 45000 29232 6 Tile_X0Y1_E6BEG[4]
port 428 nsew signal output
rlabel metal3 s 44540 29384 45000 29504 6 Tile_X0Y1_E6BEG[5]
port 429 nsew signal output
rlabel metal3 s 44540 29656 45000 29776 6 Tile_X0Y1_E6BEG[6]
port 430 nsew signal output
rlabel metal3 s 44540 29928 45000 30048 6 Tile_X0Y1_E6BEG[7]
port 431 nsew signal output
rlabel metal3 s 44540 30200 45000 30320 6 Tile_X0Y1_E6BEG[8]
port 432 nsew signal output
rlabel metal3 s 44540 30472 45000 30592 6 Tile_X0Y1_E6BEG[9]
port 433 nsew signal output
rlabel metal3 s -300 28024 160 28144 4 Tile_X0Y1_E6END[0]
port 434 nsew signal input
rlabel metal3 s -300 30744 160 30864 4 Tile_X0Y1_E6END[10]
port 435 nsew signal input
rlabel metal3 s -300 31016 160 31136 4 Tile_X0Y1_E6END[11]
port 436 nsew signal input
rlabel metal3 s -300 28296 160 28416 4 Tile_X0Y1_E6END[1]
port 437 nsew signal input
rlabel metal3 s -300 28568 160 28688 4 Tile_X0Y1_E6END[2]
port 438 nsew signal input
rlabel metal3 s -300 28840 160 28960 4 Tile_X0Y1_E6END[3]
port 439 nsew signal input
rlabel metal3 s -300 29112 160 29232 4 Tile_X0Y1_E6END[4]
port 440 nsew signal input
rlabel metal3 s -300 29384 160 29504 4 Tile_X0Y1_E6END[5]
port 441 nsew signal input
rlabel metal3 s -300 29656 160 29776 4 Tile_X0Y1_E6END[6]
port 442 nsew signal input
rlabel metal3 s -300 29928 160 30048 4 Tile_X0Y1_E6END[7]
port 443 nsew signal input
rlabel metal3 s -300 30200 160 30320 4 Tile_X0Y1_E6END[8]
port 444 nsew signal input
rlabel metal3 s -300 30472 160 30592 4 Tile_X0Y1_E6END[9]
port 445 nsew signal input
rlabel metal3 s 44540 23672 45000 23792 6 Tile_X0Y1_EE4BEG[0]
port 446 nsew signal output
rlabel metal3 s 44540 26392 45000 26512 6 Tile_X0Y1_EE4BEG[10]
port 447 nsew signal output
rlabel metal3 s 44540 26664 45000 26784 6 Tile_X0Y1_EE4BEG[11]
port 448 nsew signal output
rlabel metal3 s 44540 26936 45000 27056 6 Tile_X0Y1_EE4BEG[12]
port 449 nsew signal output
rlabel metal3 s 44540 27208 45000 27328 6 Tile_X0Y1_EE4BEG[13]
port 450 nsew signal output
rlabel metal3 s 44540 27480 45000 27600 6 Tile_X0Y1_EE4BEG[14]
port 451 nsew signal output
rlabel metal3 s 44540 27752 45000 27872 6 Tile_X0Y1_EE4BEG[15]
port 452 nsew signal output
rlabel metal3 s 44540 23944 45000 24064 6 Tile_X0Y1_EE4BEG[1]
port 453 nsew signal output
rlabel metal3 s 44540 24216 45000 24336 6 Tile_X0Y1_EE4BEG[2]
port 454 nsew signal output
rlabel metal3 s 44540 24488 45000 24608 6 Tile_X0Y1_EE4BEG[3]
port 455 nsew signal output
rlabel metal3 s 44540 24760 45000 24880 6 Tile_X0Y1_EE4BEG[4]
port 456 nsew signal output
rlabel metal3 s 44540 25032 45000 25152 6 Tile_X0Y1_EE4BEG[5]
port 457 nsew signal output
rlabel metal3 s 44540 25304 45000 25424 6 Tile_X0Y1_EE4BEG[6]
port 458 nsew signal output
rlabel metal3 s 44540 25576 45000 25696 6 Tile_X0Y1_EE4BEG[7]
port 459 nsew signal output
rlabel metal3 s 44540 25848 45000 25968 6 Tile_X0Y1_EE4BEG[8]
port 460 nsew signal output
rlabel metal3 s 44540 26120 45000 26240 6 Tile_X0Y1_EE4BEG[9]
port 461 nsew signal output
rlabel metal3 s -300 23672 160 23792 4 Tile_X0Y1_EE4END[0]
port 462 nsew signal input
rlabel metal3 s -300 26392 160 26512 4 Tile_X0Y1_EE4END[10]
port 463 nsew signal input
rlabel metal3 s -300 26664 160 26784 4 Tile_X0Y1_EE4END[11]
port 464 nsew signal input
rlabel metal3 s -300 26936 160 27056 4 Tile_X0Y1_EE4END[12]
port 465 nsew signal input
rlabel metal3 s -300 27208 160 27328 4 Tile_X0Y1_EE4END[13]
port 466 nsew signal input
rlabel metal3 s -300 27480 160 27600 4 Tile_X0Y1_EE4END[14]
port 467 nsew signal input
rlabel metal3 s -300 27752 160 27872 4 Tile_X0Y1_EE4END[15]
port 468 nsew signal input
rlabel metal3 s -300 23944 160 24064 4 Tile_X0Y1_EE4END[1]
port 469 nsew signal input
rlabel metal3 s -300 24216 160 24336 4 Tile_X0Y1_EE4END[2]
port 470 nsew signal input
rlabel metal3 s -300 24488 160 24608 4 Tile_X0Y1_EE4END[3]
port 471 nsew signal input
rlabel metal3 s -300 24760 160 24880 4 Tile_X0Y1_EE4END[4]
port 472 nsew signal input
rlabel metal3 s -300 25032 160 25152 4 Tile_X0Y1_EE4END[5]
port 473 nsew signal input
rlabel metal3 s -300 25304 160 25424 4 Tile_X0Y1_EE4END[6]
port 474 nsew signal input
rlabel metal3 s -300 25576 160 25696 4 Tile_X0Y1_EE4END[7]
port 475 nsew signal input
rlabel metal3 s -300 25848 160 25968 4 Tile_X0Y1_EE4END[8]
port 476 nsew signal input
rlabel metal3 s -300 26120 160 26240 4 Tile_X0Y1_EE4END[9]
port 477 nsew signal input
rlabel metal3 s -300 31288 160 31408 4 Tile_X0Y1_FrameData[0]
port 478 nsew signal input
rlabel metal3 s -300 34008 160 34128 4 Tile_X0Y1_FrameData[10]
port 479 nsew signal input
rlabel metal3 s -300 34280 160 34400 4 Tile_X0Y1_FrameData[11]
port 480 nsew signal input
rlabel metal3 s -300 34552 160 34672 4 Tile_X0Y1_FrameData[12]
port 481 nsew signal input
rlabel metal3 s -300 34824 160 34944 4 Tile_X0Y1_FrameData[13]
port 482 nsew signal input
rlabel metal3 s -300 35096 160 35216 4 Tile_X0Y1_FrameData[14]
port 483 nsew signal input
rlabel metal3 s -300 35368 160 35488 4 Tile_X0Y1_FrameData[15]
port 484 nsew signal input
rlabel metal3 s -300 35640 160 35760 4 Tile_X0Y1_FrameData[16]
port 485 nsew signal input
rlabel metal3 s -300 35912 160 36032 4 Tile_X0Y1_FrameData[17]
port 486 nsew signal input
rlabel metal3 s -300 36184 160 36304 4 Tile_X0Y1_FrameData[18]
port 487 nsew signal input
rlabel metal3 s -300 36456 160 36576 4 Tile_X0Y1_FrameData[19]
port 488 nsew signal input
rlabel metal3 s -300 31560 160 31680 4 Tile_X0Y1_FrameData[1]
port 489 nsew signal input
rlabel metal3 s -300 36728 160 36848 4 Tile_X0Y1_FrameData[20]
port 490 nsew signal input
rlabel metal3 s -300 37000 160 37120 4 Tile_X0Y1_FrameData[21]
port 491 nsew signal input
rlabel metal3 s -300 37272 160 37392 4 Tile_X0Y1_FrameData[22]
port 492 nsew signal input
rlabel metal3 s -300 37544 160 37664 4 Tile_X0Y1_FrameData[23]
port 493 nsew signal input
rlabel metal3 s -300 37816 160 37936 4 Tile_X0Y1_FrameData[24]
port 494 nsew signal input
rlabel metal3 s -300 38088 160 38208 4 Tile_X0Y1_FrameData[25]
port 495 nsew signal input
rlabel metal3 s -300 38360 160 38480 4 Tile_X0Y1_FrameData[26]
port 496 nsew signal input
rlabel metal3 s -300 38632 160 38752 4 Tile_X0Y1_FrameData[27]
port 497 nsew signal input
rlabel metal3 s -300 38904 160 39024 4 Tile_X0Y1_FrameData[28]
port 498 nsew signal input
rlabel metal3 s -300 39176 160 39296 4 Tile_X0Y1_FrameData[29]
port 499 nsew signal input
rlabel metal3 s -300 31832 160 31952 4 Tile_X0Y1_FrameData[2]
port 500 nsew signal input
rlabel metal3 s -300 39448 160 39568 4 Tile_X0Y1_FrameData[30]
port 501 nsew signal input
rlabel metal3 s -300 39720 160 39840 4 Tile_X0Y1_FrameData[31]
port 502 nsew signal input
rlabel metal3 s -300 32104 160 32224 4 Tile_X0Y1_FrameData[3]
port 503 nsew signal input
rlabel metal3 s -300 32376 160 32496 4 Tile_X0Y1_FrameData[4]
port 504 nsew signal input
rlabel metal3 s -300 32648 160 32768 4 Tile_X0Y1_FrameData[5]
port 505 nsew signal input
rlabel metal3 s -300 32920 160 33040 4 Tile_X0Y1_FrameData[6]
port 506 nsew signal input
rlabel metal3 s -300 33192 160 33312 4 Tile_X0Y1_FrameData[7]
port 507 nsew signal input
rlabel metal3 s -300 33464 160 33584 4 Tile_X0Y1_FrameData[8]
port 508 nsew signal input
rlabel metal3 s -300 33736 160 33856 4 Tile_X0Y1_FrameData[9]
port 509 nsew signal input
rlabel metal3 s 44540 31288 45000 31408 6 Tile_X0Y1_FrameData_O[0]
port 510 nsew signal output
rlabel metal3 s 44540 34008 45000 34128 6 Tile_X0Y1_FrameData_O[10]
port 511 nsew signal output
rlabel metal3 s 44540 34280 45000 34400 6 Tile_X0Y1_FrameData_O[11]
port 512 nsew signal output
rlabel metal3 s 44540 34552 45000 34672 6 Tile_X0Y1_FrameData_O[12]
port 513 nsew signal output
rlabel metal3 s 44540 34824 45000 34944 6 Tile_X0Y1_FrameData_O[13]
port 514 nsew signal output
rlabel metal3 s 44540 35096 45000 35216 6 Tile_X0Y1_FrameData_O[14]
port 515 nsew signal output
rlabel metal3 s 44540 35368 45000 35488 6 Tile_X0Y1_FrameData_O[15]
port 516 nsew signal output
rlabel metal3 s 44540 35640 45000 35760 6 Tile_X0Y1_FrameData_O[16]
port 517 nsew signal output
rlabel metal3 s 44540 35912 45000 36032 6 Tile_X0Y1_FrameData_O[17]
port 518 nsew signal output
rlabel metal3 s 44540 36184 45000 36304 6 Tile_X0Y1_FrameData_O[18]
port 519 nsew signal output
rlabel metal3 s 44540 36456 45000 36576 6 Tile_X0Y1_FrameData_O[19]
port 520 nsew signal output
rlabel metal3 s 44540 31560 45000 31680 6 Tile_X0Y1_FrameData_O[1]
port 521 nsew signal output
rlabel metal3 s 44540 36728 45000 36848 6 Tile_X0Y1_FrameData_O[20]
port 522 nsew signal output
rlabel metal3 s 44540 37000 45000 37120 6 Tile_X0Y1_FrameData_O[21]
port 523 nsew signal output
rlabel metal3 s 44540 37272 45000 37392 6 Tile_X0Y1_FrameData_O[22]
port 524 nsew signal output
rlabel metal3 s 44540 37544 45000 37664 6 Tile_X0Y1_FrameData_O[23]
port 525 nsew signal output
rlabel metal3 s 44540 37816 45000 37936 6 Tile_X0Y1_FrameData_O[24]
port 526 nsew signal output
rlabel metal3 s 44540 38088 45000 38208 6 Tile_X0Y1_FrameData_O[25]
port 527 nsew signal output
rlabel metal3 s 44540 38360 45000 38480 6 Tile_X0Y1_FrameData_O[26]
port 528 nsew signal output
rlabel metal3 s 44540 38632 45000 38752 6 Tile_X0Y1_FrameData_O[27]
port 529 nsew signal output
rlabel metal3 s 44540 38904 45000 39024 6 Tile_X0Y1_FrameData_O[28]
port 530 nsew signal output
rlabel metal3 s 44540 39176 45000 39296 6 Tile_X0Y1_FrameData_O[29]
port 531 nsew signal output
rlabel metal3 s 44540 31832 45000 31952 6 Tile_X0Y1_FrameData_O[2]
port 532 nsew signal output
rlabel metal3 s 44540 39448 45000 39568 6 Tile_X0Y1_FrameData_O[30]
port 533 nsew signal output
rlabel metal3 s 44540 39720 45000 39840 6 Tile_X0Y1_FrameData_O[31]
port 534 nsew signal output
rlabel metal3 s 44540 32104 45000 32224 6 Tile_X0Y1_FrameData_O[3]
port 535 nsew signal output
rlabel metal3 s 44540 32376 45000 32496 6 Tile_X0Y1_FrameData_O[4]
port 536 nsew signal output
rlabel metal3 s 44540 32648 45000 32768 6 Tile_X0Y1_FrameData_O[5]
port 537 nsew signal output
rlabel metal3 s 44540 32920 45000 33040 6 Tile_X0Y1_FrameData_O[6]
port 538 nsew signal output
rlabel metal3 s 44540 33192 45000 33312 6 Tile_X0Y1_FrameData_O[7]
port 539 nsew signal output
rlabel metal3 s 44540 33464 45000 33584 6 Tile_X0Y1_FrameData_O[8]
port 540 nsew signal output
rlabel metal3 s 44540 33736 45000 33856 6 Tile_X0Y1_FrameData_O[9]
port 541 nsew signal output
rlabel metal2 s 34150 -300 34206 160 8 Tile_X0Y1_FrameStrobe[0]
port 542 nsew signal input
rlabel metal2 s 36910 -300 36966 160 8 Tile_X0Y1_FrameStrobe[10]
port 543 nsew signal input
rlabel metal2 s 37186 -300 37242 160 8 Tile_X0Y1_FrameStrobe[11]
port 544 nsew signal input
rlabel metal2 s 37462 -300 37518 160 8 Tile_X0Y1_FrameStrobe[12]
port 545 nsew signal input
rlabel metal2 s 37738 -300 37794 160 8 Tile_X0Y1_FrameStrobe[13]
port 546 nsew signal input
rlabel metal2 s 38014 -300 38070 160 8 Tile_X0Y1_FrameStrobe[14]
port 547 nsew signal input
rlabel metal2 s 38290 -300 38346 160 8 Tile_X0Y1_FrameStrobe[15]
port 548 nsew signal input
rlabel metal2 s 38566 -300 38622 160 8 Tile_X0Y1_FrameStrobe[16]
port 549 nsew signal input
rlabel metal2 s 38842 -300 38898 160 8 Tile_X0Y1_FrameStrobe[17]
port 550 nsew signal input
rlabel metal2 s 39118 -300 39174 160 8 Tile_X0Y1_FrameStrobe[18]
port 551 nsew signal input
rlabel metal2 s 39394 -300 39450 160 8 Tile_X0Y1_FrameStrobe[19]
port 552 nsew signal input
rlabel metal2 s 34426 -300 34482 160 8 Tile_X0Y1_FrameStrobe[1]
port 553 nsew signal input
rlabel metal2 s 34702 -300 34758 160 8 Tile_X0Y1_FrameStrobe[2]
port 554 nsew signal input
rlabel metal2 s 34978 -300 35034 160 8 Tile_X0Y1_FrameStrobe[3]
port 555 nsew signal input
rlabel metal2 s 35254 -300 35310 160 8 Tile_X0Y1_FrameStrobe[4]
port 556 nsew signal input
rlabel metal2 s 35530 -300 35586 160 8 Tile_X0Y1_FrameStrobe[5]
port 557 nsew signal input
rlabel metal2 s 35806 -300 35862 160 8 Tile_X0Y1_FrameStrobe[6]
port 558 nsew signal input
rlabel metal2 s 36082 -300 36138 160 8 Tile_X0Y1_FrameStrobe[7]
port 559 nsew signal input
rlabel metal2 s 36358 -300 36414 160 8 Tile_X0Y1_FrameStrobe[8]
port 560 nsew signal input
rlabel metal2 s 36634 -300 36690 160 8 Tile_X0Y1_FrameStrobe[9]
port 561 nsew signal input
rlabel metal2 s 5170 -300 5226 160 8 Tile_X0Y1_N1END[0]
port 562 nsew signal input
rlabel metal2 s 5446 -300 5502 160 8 Tile_X0Y1_N1END[1]
port 563 nsew signal input
rlabel metal2 s 5722 -300 5778 160 8 Tile_X0Y1_N1END[2]
port 564 nsew signal input
rlabel metal2 s 5998 -300 6054 160 8 Tile_X0Y1_N1END[3]
port 565 nsew signal input
rlabel metal2 s 8482 -300 8538 160 8 Tile_X0Y1_N2END[0]
port 566 nsew signal input
rlabel metal2 s 8758 -300 8814 160 8 Tile_X0Y1_N2END[1]
port 567 nsew signal input
rlabel metal2 s 9034 -300 9090 160 8 Tile_X0Y1_N2END[2]
port 568 nsew signal input
rlabel metal2 s 9310 -300 9366 160 8 Tile_X0Y1_N2END[3]
port 569 nsew signal input
rlabel metal2 s 9586 -300 9642 160 8 Tile_X0Y1_N2END[4]
port 570 nsew signal input
rlabel metal2 s 9862 -300 9918 160 8 Tile_X0Y1_N2END[5]
port 571 nsew signal input
rlabel metal2 s 10138 -300 10194 160 8 Tile_X0Y1_N2END[6]
port 572 nsew signal input
rlabel metal2 s 10414 -300 10470 160 8 Tile_X0Y1_N2END[7]
port 573 nsew signal input
rlabel metal2 s 6274 -300 6330 160 8 Tile_X0Y1_N2MID[0]
port 574 nsew signal input
rlabel metal2 s 6550 -300 6606 160 8 Tile_X0Y1_N2MID[1]
port 575 nsew signal input
rlabel metal2 s 6826 -300 6882 160 8 Tile_X0Y1_N2MID[2]
port 576 nsew signal input
rlabel metal2 s 7102 -300 7158 160 8 Tile_X0Y1_N2MID[3]
port 577 nsew signal input
rlabel metal2 s 7378 -300 7434 160 8 Tile_X0Y1_N2MID[4]
port 578 nsew signal input
rlabel metal2 s 7654 -300 7710 160 8 Tile_X0Y1_N2MID[5]
port 579 nsew signal input
rlabel metal2 s 7930 -300 7986 160 8 Tile_X0Y1_N2MID[6]
port 580 nsew signal input
rlabel metal2 s 8206 -300 8262 160 8 Tile_X0Y1_N2MID[7]
port 581 nsew signal input
rlabel metal2 s 10690 -300 10746 160 8 Tile_X0Y1_N4END[0]
port 582 nsew signal input
rlabel metal2 s 13450 -300 13506 160 8 Tile_X0Y1_N4END[10]
port 583 nsew signal input
rlabel metal2 s 13726 -300 13782 160 8 Tile_X0Y1_N4END[11]
port 584 nsew signal input
rlabel metal2 s 14002 -300 14058 160 8 Tile_X0Y1_N4END[12]
port 585 nsew signal input
rlabel metal2 s 14278 -300 14334 160 8 Tile_X0Y1_N4END[13]
port 586 nsew signal input
rlabel metal2 s 14554 -300 14610 160 8 Tile_X0Y1_N4END[14]
port 587 nsew signal input
rlabel metal2 s 14830 -300 14886 160 8 Tile_X0Y1_N4END[15]
port 588 nsew signal input
rlabel metal2 s 10966 -300 11022 160 8 Tile_X0Y1_N4END[1]
port 589 nsew signal input
rlabel metal2 s 11242 -300 11298 160 8 Tile_X0Y1_N4END[2]
port 590 nsew signal input
rlabel metal2 s 11518 -300 11574 160 8 Tile_X0Y1_N4END[3]
port 591 nsew signal input
rlabel metal2 s 11794 -300 11850 160 8 Tile_X0Y1_N4END[4]
port 592 nsew signal input
rlabel metal2 s 12070 -300 12126 160 8 Tile_X0Y1_N4END[5]
port 593 nsew signal input
rlabel metal2 s 12346 -300 12402 160 8 Tile_X0Y1_N4END[6]
port 594 nsew signal input
rlabel metal2 s 12622 -300 12678 160 8 Tile_X0Y1_N4END[7]
port 595 nsew signal input
rlabel metal2 s 12898 -300 12954 160 8 Tile_X0Y1_N4END[8]
port 596 nsew signal input
rlabel metal2 s 13174 -300 13230 160 8 Tile_X0Y1_N4END[9]
port 597 nsew signal input
rlabel metal2 s 15106 -300 15162 160 8 Tile_X0Y1_NN4END[0]
port 598 nsew signal input
rlabel metal2 s 17866 -300 17922 160 8 Tile_X0Y1_NN4END[10]
port 599 nsew signal input
rlabel metal2 s 18142 -300 18198 160 8 Tile_X0Y1_NN4END[11]
port 600 nsew signal input
rlabel metal2 s 18418 -300 18474 160 8 Tile_X0Y1_NN4END[12]
port 601 nsew signal input
rlabel metal2 s 18694 -300 18750 160 8 Tile_X0Y1_NN4END[13]
port 602 nsew signal input
rlabel metal2 s 18970 -300 19026 160 8 Tile_X0Y1_NN4END[14]
port 603 nsew signal input
rlabel metal2 s 19246 -300 19302 160 8 Tile_X0Y1_NN4END[15]
port 604 nsew signal input
rlabel metal2 s 15382 -300 15438 160 8 Tile_X0Y1_NN4END[1]
port 605 nsew signal input
rlabel metal2 s 15658 -300 15714 160 8 Tile_X0Y1_NN4END[2]
port 606 nsew signal input
rlabel metal2 s 15934 -300 15990 160 8 Tile_X0Y1_NN4END[3]
port 607 nsew signal input
rlabel metal2 s 16210 -300 16266 160 8 Tile_X0Y1_NN4END[4]
port 608 nsew signal input
rlabel metal2 s 16486 -300 16542 160 8 Tile_X0Y1_NN4END[5]
port 609 nsew signal input
rlabel metal2 s 16762 -300 16818 160 8 Tile_X0Y1_NN4END[6]
port 610 nsew signal input
rlabel metal2 s 17038 -300 17094 160 8 Tile_X0Y1_NN4END[7]
port 611 nsew signal input
rlabel metal2 s 17314 -300 17370 160 8 Tile_X0Y1_NN4END[8]
port 612 nsew signal input
rlabel metal2 s 17590 -300 17646 160 8 Tile_X0Y1_NN4END[9]
port 613 nsew signal input
rlabel metal2 s 19522 -300 19578 160 8 Tile_X0Y1_S1BEG[0]
port 614 nsew signal output
rlabel metal2 s 19798 -300 19854 160 8 Tile_X0Y1_S1BEG[1]
port 615 nsew signal output
rlabel metal2 s 20074 -300 20130 160 8 Tile_X0Y1_S1BEG[2]
port 616 nsew signal output
rlabel metal2 s 20350 -300 20406 160 8 Tile_X0Y1_S1BEG[3]
port 617 nsew signal output
rlabel metal2 s 22834 -300 22890 160 8 Tile_X0Y1_S2BEG[0]
port 618 nsew signal output
rlabel metal2 s 23110 -300 23166 160 8 Tile_X0Y1_S2BEG[1]
port 619 nsew signal output
rlabel metal2 s 23386 -300 23442 160 8 Tile_X0Y1_S2BEG[2]
port 620 nsew signal output
rlabel metal2 s 23662 -300 23718 160 8 Tile_X0Y1_S2BEG[3]
port 621 nsew signal output
rlabel metal2 s 23938 -300 23994 160 8 Tile_X0Y1_S2BEG[4]
port 622 nsew signal output
rlabel metal2 s 24214 -300 24270 160 8 Tile_X0Y1_S2BEG[5]
port 623 nsew signal output
rlabel metal2 s 24490 -300 24546 160 8 Tile_X0Y1_S2BEG[6]
port 624 nsew signal output
rlabel metal2 s 24766 -300 24822 160 8 Tile_X0Y1_S2BEG[7]
port 625 nsew signal output
rlabel metal2 s 20626 -300 20682 160 8 Tile_X0Y1_S2BEGb[0]
port 626 nsew signal output
rlabel metal2 s 20902 -300 20958 160 8 Tile_X0Y1_S2BEGb[1]
port 627 nsew signal output
rlabel metal2 s 21178 -300 21234 160 8 Tile_X0Y1_S2BEGb[2]
port 628 nsew signal output
rlabel metal2 s 21454 -300 21510 160 8 Tile_X0Y1_S2BEGb[3]
port 629 nsew signal output
rlabel metal2 s 21730 -300 21786 160 8 Tile_X0Y1_S2BEGb[4]
port 630 nsew signal output
rlabel metal2 s 22006 -300 22062 160 8 Tile_X0Y1_S2BEGb[5]
port 631 nsew signal output
rlabel metal2 s 22282 -300 22338 160 8 Tile_X0Y1_S2BEGb[6]
port 632 nsew signal output
rlabel metal2 s 22558 -300 22614 160 8 Tile_X0Y1_S2BEGb[7]
port 633 nsew signal output
rlabel metal2 s 25042 -300 25098 160 8 Tile_X0Y1_S4BEG[0]
port 634 nsew signal output
rlabel metal2 s 27802 -300 27858 160 8 Tile_X0Y1_S4BEG[10]
port 635 nsew signal output
rlabel metal2 s 28078 -300 28134 160 8 Tile_X0Y1_S4BEG[11]
port 636 nsew signal output
rlabel metal2 s 28354 -300 28410 160 8 Tile_X0Y1_S4BEG[12]
port 637 nsew signal output
rlabel metal2 s 28630 -300 28686 160 8 Tile_X0Y1_S4BEG[13]
port 638 nsew signal output
rlabel metal2 s 28906 -300 28962 160 8 Tile_X0Y1_S4BEG[14]
port 639 nsew signal output
rlabel metal2 s 29182 -300 29238 160 8 Tile_X0Y1_S4BEG[15]
port 640 nsew signal output
rlabel metal2 s 25318 -300 25374 160 8 Tile_X0Y1_S4BEG[1]
port 641 nsew signal output
rlabel metal2 s 25594 -300 25650 160 8 Tile_X0Y1_S4BEG[2]
port 642 nsew signal output
rlabel metal2 s 25870 -300 25926 160 8 Tile_X0Y1_S4BEG[3]
port 643 nsew signal output
rlabel metal2 s 26146 -300 26202 160 8 Tile_X0Y1_S4BEG[4]
port 644 nsew signal output
rlabel metal2 s 26422 -300 26478 160 8 Tile_X0Y1_S4BEG[5]
port 645 nsew signal output
rlabel metal2 s 26698 -300 26754 160 8 Tile_X0Y1_S4BEG[6]
port 646 nsew signal output
rlabel metal2 s 26974 -300 27030 160 8 Tile_X0Y1_S4BEG[7]
port 647 nsew signal output
rlabel metal2 s 27250 -300 27306 160 8 Tile_X0Y1_S4BEG[8]
port 648 nsew signal output
rlabel metal2 s 27526 -300 27582 160 8 Tile_X0Y1_S4BEG[9]
port 649 nsew signal output
rlabel metal2 s 29458 -300 29514 160 8 Tile_X0Y1_SS4BEG[0]
port 650 nsew signal output
rlabel metal2 s 32218 -300 32274 160 8 Tile_X0Y1_SS4BEG[10]
port 651 nsew signal output
rlabel metal2 s 32494 -300 32550 160 8 Tile_X0Y1_SS4BEG[11]
port 652 nsew signal output
rlabel metal2 s 32770 -300 32826 160 8 Tile_X0Y1_SS4BEG[12]
port 653 nsew signal output
rlabel metal2 s 33046 -300 33102 160 8 Tile_X0Y1_SS4BEG[13]
port 654 nsew signal output
rlabel metal2 s 33322 -300 33378 160 8 Tile_X0Y1_SS4BEG[14]
port 655 nsew signal output
rlabel metal2 s 33598 -300 33654 160 8 Tile_X0Y1_SS4BEG[15]
port 656 nsew signal output
rlabel metal2 s 29734 -300 29790 160 8 Tile_X0Y1_SS4BEG[1]
port 657 nsew signal output
rlabel metal2 s 30010 -300 30066 160 8 Tile_X0Y1_SS4BEG[2]
port 658 nsew signal output
rlabel metal2 s 30286 -300 30342 160 8 Tile_X0Y1_SS4BEG[3]
port 659 nsew signal output
rlabel metal2 s 30562 -300 30618 160 8 Tile_X0Y1_SS4BEG[4]
port 660 nsew signal output
rlabel metal2 s 30838 -300 30894 160 8 Tile_X0Y1_SS4BEG[5]
port 661 nsew signal output
rlabel metal2 s 31114 -300 31170 160 8 Tile_X0Y1_SS4BEG[6]
port 662 nsew signal output
rlabel metal2 s 31390 -300 31446 160 8 Tile_X0Y1_SS4BEG[7]
port 663 nsew signal output
rlabel metal2 s 31666 -300 31722 160 8 Tile_X0Y1_SS4BEG[8]
port 664 nsew signal output
rlabel metal2 s 31942 -300 31998 160 8 Tile_X0Y1_SS4BEG[9]
port 665 nsew signal output
rlabel metal2 s 33874 -300 33930 160 8 Tile_X0Y1_UserCLK
port 666 nsew signal input
rlabel metal3 s -300 5176 160 5296 4 Tile_X0Y1_W1BEG[0]
port 667 nsew signal output
rlabel metal3 s -300 5448 160 5568 4 Tile_X0Y1_W1BEG[1]
port 668 nsew signal output
rlabel metal3 s -300 5720 160 5840 4 Tile_X0Y1_W1BEG[2]
port 669 nsew signal output
rlabel metal3 s -300 5992 160 6112 4 Tile_X0Y1_W1BEG[3]
port 670 nsew signal output
rlabel metal3 s 44540 5176 45000 5296 6 Tile_X0Y1_W1END[0]
port 671 nsew signal input
rlabel metal3 s 44540 5448 45000 5568 6 Tile_X0Y1_W1END[1]
port 672 nsew signal input
rlabel metal3 s 44540 5720 45000 5840 6 Tile_X0Y1_W1END[2]
port 673 nsew signal input
rlabel metal3 s 44540 5992 45000 6112 6 Tile_X0Y1_W1END[3]
port 674 nsew signal input
rlabel metal3 s -300 6264 160 6384 4 Tile_X0Y1_W2BEG[0]
port 675 nsew signal output
rlabel metal3 s -300 6536 160 6656 4 Tile_X0Y1_W2BEG[1]
port 676 nsew signal output
rlabel metal3 s -300 6808 160 6928 4 Tile_X0Y1_W2BEG[2]
port 677 nsew signal output
rlabel metal3 s -300 7080 160 7200 4 Tile_X0Y1_W2BEG[3]
port 678 nsew signal output
rlabel metal3 s -300 7352 160 7472 4 Tile_X0Y1_W2BEG[4]
port 679 nsew signal output
rlabel metal3 s -300 7624 160 7744 4 Tile_X0Y1_W2BEG[5]
port 680 nsew signal output
rlabel metal3 s -300 7896 160 8016 4 Tile_X0Y1_W2BEG[6]
port 681 nsew signal output
rlabel metal3 s -300 8168 160 8288 4 Tile_X0Y1_W2BEG[7]
port 682 nsew signal output
rlabel metal3 s -300 8440 160 8560 4 Tile_X0Y1_W2BEGb[0]
port 683 nsew signal output
rlabel metal3 s -300 8712 160 8832 4 Tile_X0Y1_W2BEGb[1]
port 684 nsew signal output
rlabel metal3 s -300 8984 160 9104 4 Tile_X0Y1_W2BEGb[2]
port 685 nsew signal output
rlabel metal3 s -300 9256 160 9376 4 Tile_X0Y1_W2BEGb[3]
port 686 nsew signal output
rlabel metal3 s -300 9528 160 9648 4 Tile_X0Y1_W2BEGb[4]
port 687 nsew signal output
rlabel metal3 s -300 9800 160 9920 4 Tile_X0Y1_W2BEGb[5]
port 688 nsew signal output
rlabel metal3 s -300 10072 160 10192 4 Tile_X0Y1_W2BEGb[6]
port 689 nsew signal output
rlabel metal3 s -300 10344 160 10464 4 Tile_X0Y1_W2BEGb[7]
port 690 nsew signal output
rlabel metal3 s 44540 8440 45000 8560 6 Tile_X0Y1_W2END[0]
port 691 nsew signal input
rlabel metal3 s 44540 8712 45000 8832 6 Tile_X0Y1_W2END[1]
port 692 nsew signal input
rlabel metal3 s 44540 8984 45000 9104 6 Tile_X0Y1_W2END[2]
port 693 nsew signal input
rlabel metal3 s 44540 9256 45000 9376 6 Tile_X0Y1_W2END[3]
port 694 nsew signal input
rlabel metal3 s 44540 9528 45000 9648 6 Tile_X0Y1_W2END[4]
port 695 nsew signal input
rlabel metal3 s 44540 9800 45000 9920 6 Tile_X0Y1_W2END[5]
port 696 nsew signal input
rlabel metal3 s 44540 10072 45000 10192 6 Tile_X0Y1_W2END[6]
port 697 nsew signal input
rlabel metal3 s 44540 10344 45000 10464 6 Tile_X0Y1_W2END[7]
port 698 nsew signal input
rlabel metal3 s 44540 6264 45000 6384 6 Tile_X0Y1_W2MID[0]
port 699 nsew signal input
rlabel metal3 s 44540 6536 45000 6656 6 Tile_X0Y1_W2MID[1]
port 700 nsew signal input
rlabel metal3 s 44540 6808 45000 6928 6 Tile_X0Y1_W2MID[2]
port 701 nsew signal input
rlabel metal3 s 44540 7080 45000 7200 6 Tile_X0Y1_W2MID[3]
port 702 nsew signal input
rlabel metal3 s 44540 7352 45000 7472 6 Tile_X0Y1_W2MID[4]
port 703 nsew signal input
rlabel metal3 s 44540 7624 45000 7744 6 Tile_X0Y1_W2MID[5]
port 704 nsew signal input
rlabel metal3 s 44540 7896 45000 8016 6 Tile_X0Y1_W2MID[6]
port 705 nsew signal input
rlabel metal3 s 44540 8168 45000 8288 6 Tile_X0Y1_W2MID[7]
port 706 nsew signal input
rlabel metal3 s -300 14968 160 15088 4 Tile_X0Y1_W6BEG[0]
port 707 nsew signal output
rlabel metal3 s -300 17688 160 17808 4 Tile_X0Y1_W6BEG[10]
port 708 nsew signal output
rlabel metal3 s -300 17960 160 18080 4 Tile_X0Y1_W6BEG[11]
port 709 nsew signal output
rlabel metal3 s -300 15240 160 15360 4 Tile_X0Y1_W6BEG[1]
port 710 nsew signal output
rlabel metal3 s -300 15512 160 15632 4 Tile_X0Y1_W6BEG[2]
port 711 nsew signal output
rlabel metal3 s -300 15784 160 15904 4 Tile_X0Y1_W6BEG[3]
port 712 nsew signal output
rlabel metal3 s -300 16056 160 16176 4 Tile_X0Y1_W6BEG[4]
port 713 nsew signal output
rlabel metal3 s -300 16328 160 16448 4 Tile_X0Y1_W6BEG[5]
port 714 nsew signal output
rlabel metal3 s -300 16600 160 16720 4 Tile_X0Y1_W6BEG[6]
port 715 nsew signal output
rlabel metal3 s -300 16872 160 16992 4 Tile_X0Y1_W6BEG[7]
port 716 nsew signal output
rlabel metal3 s -300 17144 160 17264 4 Tile_X0Y1_W6BEG[8]
port 717 nsew signal output
rlabel metal3 s -300 17416 160 17536 4 Tile_X0Y1_W6BEG[9]
port 718 nsew signal output
rlabel metal3 s 44540 14968 45000 15088 6 Tile_X0Y1_W6END[0]
port 719 nsew signal input
rlabel metal3 s 44540 17688 45000 17808 6 Tile_X0Y1_W6END[10]
port 720 nsew signal input
rlabel metal3 s 44540 17960 45000 18080 6 Tile_X0Y1_W6END[11]
port 721 nsew signal input
rlabel metal3 s 44540 15240 45000 15360 6 Tile_X0Y1_W6END[1]
port 722 nsew signal input
rlabel metal3 s 44540 15512 45000 15632 6 Tile_X0Y1_W6END[2]
port 723 nsew signal input
rlabel metal3 s 44540 15784 45000 15904 6 Tile_X0Y1_W6END[3]
port 724 nsew signal input
rlabel metal3 s 44540 16056 45000 16176 6 Tile_X0Y1_W6END[4]
port 725 nsew signal input
rlabel metal3 s 44540 16328 45000 16448 6 Tile_X0Y1_W6END[5]
port 726 nsew signal input
rlabel metal3 s 44540 16600 45000 16720 6 Tile_X0Y1_W6END[6]
port 727 nsew signal input
rlabel metal3 s 44540 16872 45000 16992 6 Tile_X0Y1_W6END[7]
port 728 nsew signal input
rlabel metal3 s 44540 17144 45000 17264 6 Tile_X0Y1_W6END[8]
port 729 nsew signal input
rlabel metal3 s 44540 17416 45000 17536 6 Tile_X0Y1_W6END[9]
port 730 nsew signal input
rlabel metal3 s -300 10616 160 10736 4 Tile_X0Y1_WW4BEG[0]
port 731 nsew signal output
rlabel metal3 s -300 13336 160 13456 4 Tile_X0Y1_WW4BEG[10]
port 732 nsew signal output
rlabel metal3 s -300 13608 160 13728 4 Tile_X0Y1_WW4BEG[11]
port 733 nsew signal output
rlabel metal3 s -300 13880 160 14000 4 Tile_X0Y1_WW4BEG[12]
port 734 nsew signal output
rlabel metal3 s -300 14152 160 14272 4 Tile_X0Y1_WW4BEG[13]
port 735 nsew signal output
rlabel metal3 s -300 14424 160 14544 4 Tile_X0Y1_WW4BEG[14]
port 736 nsew signal output
rlabel metal3 s -300 14696 160 14816 4 Tile_X0Y1_WW4BEG[15]
port 737 nsew signal output
rlabel metal3 s -300 10888 160 11008 4 Tile_X0Y1_WW4BEG[1]
port 738 nsew signal output
rlabel metal3 s -300 11160 160 11280 4 Tile_X0Y1_WW4BEG[2]
port 739 nsew signal output
rlabel metal3 s -300 11432 160 11552 4 Tile_X0Y1_WW4BEG[3]
port 740 nsew signal output
rlabel metal3 s -300 11704 160 11824 4 Tile_X0Y1_WW4BEG[4]
port 741 nsew signal output
rlabel metal3 s -300 11976 160 12096 4 Tile_X0Y1_WW4BEG[5]
port 742 nsew signal output
rlabel metal3 s -300 12248 160 12368 4 Tile_X0Y1_WW4BEG[6]
port 743 nsew signal output
rlabel metal3 s -300 12520 160 12640 4 Tile_X0Y1_WW4BEG[7]
port 744 nsew signal output
rlabel metal3 s -300 12792 160 12912 4 Tile_X0Y1_WW4BEG[8]
port 745 nsew signal output
rlabel metal3 s -300 13064 160 13184 4 Tile_X0Y1_WW4BEG[9]
port 746 nsew signal output
rlabel metal3 s 44540 10616 45000 10736 6 Tile_X0Y1_WW4END[0]
port 747 nsew signal input
rlabel metal3 s 44540 13336 45000 13456 6 Tile_X0Y1_WW4END[10]
port 748 nsew signal input
rlabel metal3 s 44540 13608 45000 13728 6 Tile_X0Y1_WW4END[11]
port 749 nsew signal input
rlabel metal3 s 44540 13880 45000 14000 6 Tile_X0Y1_WW4END[12]
port 750 nsew signal input
rlabel metal3 s 44540 14152 45000 14272 6 Tile_X0Y1_WW4END[13]
port 751 nsew signal input
rlabel metal3 s 44540 14424 45000 14544 6 Tile_X0Y1_WW4END[14]
port 752 nsew signal input
rlabel metal3 s 44540 14696 45000 14816 6 Tile_X0Y1_WW4END[15]
port 753 nsew signal input
rlabel metal3 s 44540 10888 45000 11008 6 Tile_X0Y1_WW4END[1]
port 754 nsew signal input
rlabel metal3 s 44540 11160 45000 11280 6 Tile_X0Y1_WW4END[2]
port 755 nsew signal input
rlabel metal3 s 44540 11432 45000 11552 6 Tile_X0Y1_WW4END[3]
port 756 nsew signal input
rlabel metal3 s 44540 11704 45000 11824 6 Tile_X0Y1_WW4END[4]
port 757 nsew signal input
rlabel metal3 s 44540 11976 45000 12096 6 Tile_X0Y1_WW4END[5]
port 758 nsew signal input
rlabel metal3 s 44540 12248 45000 12368 6 Tile_X0Y1_WW4END[6]
port 759 nsew signal input
rlabel metal3 s 44540 12520 45000 12640 6 Tile_X0Y1_WW4END[7]
port 760 nsew signal input
rlabel metal3 s 44540 12792 45000 12912 6 Tile_X0Y1_WW4END[8]
port 761 nsew signal input
rlabel metal3 s 44540 13064 45000 13184 6 Tile_X0Y1_WW4END[9]
port 762 nsew signal input
rlabel metal4 s 19568 1040 19888 89264 6 VGND
port 763 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 89264 6 VPWR
port 764 nsew power bidirectional
rlabel metal4 s 34928 1040 35248 89264 6 VPWR
port 764 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 44700 90700
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13987304
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/DSP/runs/24_12_07_23_46/results/signoff/DSP.magic.gds
string GDS_START 1107074
<< end >>

