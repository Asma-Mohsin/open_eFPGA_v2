* NGSPICE file created from LUT4AB.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxbp_1 abstract view
.subckt sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_8 abstract view
.subckt sky130_fd_sc_hd__mux2_8 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo W1BEG[0] W1BEG[1]
+ W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1] W2BEG[2]
+ W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2] W2BEGb[3]
+ W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3] W2END[4]
+ W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5]
+ W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3] W6BEG[4]
+ W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11] W6END[1]
+ W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9] WW4BEG[0]
+ WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1] WW4BEG[2]
+ WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9] WW4END[0]
+ WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1] WW4END[2]
+ WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9] vccd1 vssd1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit11 input52/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XW6END_inbuf_0__0_ input230/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_0__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit22 input64/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit28_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit19_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_394 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0_A3
+ input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_data_inbuf_11__0__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit19 input60/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__081__A Inst_LUT4AB_switch_matrix__081_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_26__0__A input68/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit3_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3 Inst_LUT4AB_ConfigMem_Inst_Frame18_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit21/Q Inst_LE_LUT4c_frame_config_dffesr__07_/A
+ Inst_LE_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XWW4END_inbuf_10__0_ input243/X vssd1 vssd1 vccd1 vccd1 WW4END_inbuf_10__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit15 input56/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit26 input68/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit4_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput401 output401/A vssd1 vssd1 vccd1 vccd1 NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput423 output423/A vssd1 vssd1 vccd1 vccd1 S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput412 output412/A vssd1 vssd1 vccd1 vccd1 S2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput434 output434/A vssd1 vssd1 vccd1 vccd1 S4BEG[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput467 output467/A vssd1 vssd1 vccd1 vccd1 W2BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput456 output456/A vssd1 vssd1 vccd1 vccd1 SS4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput445 output445/A vssd1 vssd1 vccd1 vccd1 SS4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput478 output478/A vssd1 vssd1 vccd1 vccd1 W2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput489 output489/A vssd1 vssd1 vccd1 vccd1 W6BEG[7] sky130_fd_sc_hd__clkbuf_4
XN4BEG_outbuf_11__0_ N4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 output377/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG1_A2 input22/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit2 input72/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I1_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__076__A input117/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit21 input63/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit10 input51/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XS4END_inbuf_9__0_ input178/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix__051_ input19/X vssd1 vssd1 vccd1 vccd1 output272/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit19 input60/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG3_A2 input158/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0_A0
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit14_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit23_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput286 output286/A vssd1 vssd1 vccd1 vccd1 E6BEG[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput264 output264/A vssd1 vssd1 vccd1 vccd1 E2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput275 output275/A vssd1 vssd1 vccd1 vccd1 E6BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput297 output297/A vssd1 vssd1 vccd1 vccd1 EE4BEG[4] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit18 input59/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S0_A0 Inst_LUT4AB_switch_matrix__069_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG2_A0 input158/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit29 input71/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG3_A2 input218/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0_A3
+ input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit14 input55/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit25 input67/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit19_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit7_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit28_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1 input22/X
+ input160/X input212/X input226/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit2_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__103_ ANTENNA_4/DIODE vssd1 vssd1 vccd1 vccd1 output470/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit8_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__034_ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__034_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit11_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit3_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0_A1
+ input108/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit5 input77/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG2_A2 input214/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit20 input62/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit18 input59/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit6 input78/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit29 input71/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit16_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit25_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0 input104/X
+ input110/X input122/X input10/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_W6BEG_outbuf_8__0__A W6END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG0_A3 input216/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_inbuf_20__0_ input62/X vssd1 vssd1 vccd1 vccd1 data_inbuf_20__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit17 input58/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit28 input70/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LG_LUT4c_frame_config_dffesr__12__A1 Inst_LG_LUT4c_frame_config_dffesr__09_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG1_A3 input221/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LH_LUT4c_frame_config_dffesr__08_ Inst_LH_LUT4c_frame_config_dffesr__08_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__08_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG0_A3 Inst_LUT4AB_switch_matrix__069_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_11__0_ input52/X vssd1 vssd1 vccd1 vccd1 data_inbuf_11__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit13 input54/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG1_A0 input117/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit24 input66/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG0_A0 input120/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__084__A Inst_LUT4AB_switch_matrix__084_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S3 Inst_LUT4AB_switch_matrix__072_/A
+ Inst_LUT4AB_switch_matrix__045_/A Inst_LUT4AB_switch_matrix__088_/A Inst_LUT4AB_switch_matrix__104_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit2/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_AH__0_/S sky130_fd_sc_hd__mux4_2
XFILLER_0_53_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_5 ANTENNA_5/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I1_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_SS4BEG_outbuf_4__0__A SS4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit28 input70/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit17 input58/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit0 input50/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit15/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit14/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit14/Q Inst_LD_LUT4c_frame_config_dffesr__07_/A
+ Inst_LD_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit9 input81/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput120 N2MID[6] vssd1 vssd1 vccd1 vccd1 input120/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix__079__A input120/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput131 N4END[3] vssd1 vssd1 vccd1 vccd1 input131/X sky130_fd_sc_hd__buf_2
Xinput142 NN4END[13] vssd1 vssd1 vccd1 vccd1 input142/X sky130_fd_sc_hd__clkbuf_1
Xinput153 NN4END[9] vssd1 vssd1 vccd1 vccd1 input153/X sky130_fd_sc_hd__clkbuf_1
Xinput164 S2END[6] vssd1 vssd1 vccd1 vccd1 input164/X sky130_fd_sc_hd__buf_2
Xinput186 S4END[6] vssd1 vssd1 vccd1 vccd1 input186/X sky130_fd_sc_hd__clkbuf_1
Xinput175 S4END[10] vssd1 vssd1 vccd1 vccd1 input175/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput197 SS4END[1] vssd1 vssd1 vccd1 vccd1 input197/X sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit11_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit20_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_outbuf_14__0_ strobe_inbuf_14__0_/X vssd1 vssd1 vccd1 vccd1 output340/A sky130_fd_sc_hd__clkbuf_1
XInst_LB_LUT4c_frame_config_dffesr_cus_mux21_O__0_ Inst_LB_LUT4c_frame_config_dffesr__13_/A0
+ hold9/A Inst_LUT4AB_ConfigMem_Inst_Frame16_bit4/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__033_/A
+ sky130_fd_sc_hd__mux2_8
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_9__0_ data_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output334/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG1_A3 input213/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit12 input53/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit23 input65/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG0 input120/X input20/X
+ input172/X Inst_LUT4AB_switch_matrix__071_/A Inst_LUT4AB_ConfigMem_Inst_Frame9_bit9/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit8/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG0 input131/X input9/X input213/X
+ Inst_LUT4AB_switch_matrix__068_/A Inst_LUT4AB_ConfigMem_Inst_Frame12_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A3 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LA_SR__0__508 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LA_SR__0__508/HI
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LA_SR__0_/A0 sky130_fd_sc_hd__conb_1
XFILLER_0_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0 input104/X
+ input112/X input4/X input12/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit13/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit16_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S3_A0 Inst_LUT4AB_switch_matrix__072_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit25_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XWW4END_inbuf_5__0_ input253/X vssd1 vssd1 vccd1 vccd1 WW4END_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_WW4BEG_outbuf_8__0__A ANTENNA_9/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4_S1
+ Inst_LE_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LC_EN__0__518 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LC_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LC_EN__0__518/LO sky130_fd_sc_hd__conb_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4 Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X Inst_LE_LUT4c_frame_config_dffesr__09_/A
+ Inst_LE_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__13_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit27 input69/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit16 input57/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput402 output402/A vssd1 vssd1 vccd1 vccd1 NN4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput424 output424/A vssd1 vssd1 vccd1 vccd1 S2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput413 output413/A vssd1 vssd1 vccd1 vccd1 S2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput435 output435/A vssd1 vssd1 vccd1 vccd1 S4BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput468 output468/A vssd1 vssd1 vccd1 vccd1 W2BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput457 output457/A vssd1 vssd1 vccd1 vccd1 SS4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput446 output446/A vssd1 vssd1 vccd1 vccd1 SS4BEG[12] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput479 output479/A vssd1 vssd1 vccd1 vccd1 W2BEGb[7] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG1_A3 Inst_LUT4AB_switch_matrix__054_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit13_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit22_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit3 input75/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit31_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit24/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_S4BEG_outbuf_2__0__A S4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__092__A input169/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit22 input64/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit11 input52/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0_A3
+ input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit18_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__050_ input18/X vssd1 vssd1 vccd1 vccd1 output271/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit27_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG3_A3 input247/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0_A1
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0 input103/X
+ input111/X input3/X input11/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput254 output254/A vssd1 vssd1 vccd1 vccd1 Co sky130_fd_sc_hd__buf_2
Xoutput276 output276/A vssd1 vssd1 vccd1 vccd1 E6BEG[10] sky130_fd_sc_hd__buf_2
Xoutput265 output265/A vssd1 vssd1 vccd1 vccd1 E2BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput287 output287/A vssd1 vssd1 vccd1 vccd1 EE4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput298 output298/A vssd1 vssd1 vccd1 vccd1 EE4BEG[5] sky130_fd_sc_hd__clkbuf_4
XANTENNA_data_inbuf_10__0__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S0_A1 Inst_LUT4AB_switch_matrix__042_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit19 input60/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG3_A3 Inst_LUT4AB_switch_matrix__101_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG2_A1 input183/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_data_inbuf_25__0__A input67/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG3_A0 input114/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_11__0_ input84/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_11__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit15 input56/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit26 input68/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix__087__A Inst_LUT4AB_switch_matrix__087_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XE6END_inbuf_5__0_ input31/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__102_ Inst_LUT4AB_switch_matrix__102_/A vssd1 vssd1 vccd1
+ vccd1 output469/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__033_ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__033_/X sky130_fd_sc_hd__buf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit2_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit3_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0_A2
+ input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit6 input78/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG2_A3 Inst_LUT4AB_switch_matrix__084_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit10 input51/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit21 input63/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit7 input79/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit19 input60/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XSS4END_inbuf_7__0_ input192/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1 input22/X
+ input162/X input214/X input226/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit13_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit18 input59/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit29 input71/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit31_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_9__0_ strobe_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output354/A sky130_fd_sc_hd__clkbuf_1
XInst_LH_LUT4c_frame_config_dffesr__07_ Inst_LH_LUT4c_frame_config_dffesr__07_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__07_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit14 input55/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit25 input67/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG1_A1 input17/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit18_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1_A0
+ input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit27_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG0_A1 input172/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XEE4END_inbuf_6__0_ input35/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_2
Xdata_inbuf_3__0_ input75/X vssd1 vssd1 vccd1 vccd1 data_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_6 ANTENNA_6/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I1_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit6_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XWW4BEG_outbuf_7__0_ ANTENNA_8/DIODE vssd1 vssd1 vccd1 vccd1 output505/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit7_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit18 input59/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit29 input71/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit1 input61/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit15_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit24_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit13/Q Inst_LD_LUT4c_frame_config_dffesr__07_/A
+ Inst_LD_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_W6BEG_outbuf_7__0__A W6END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A0
+ ANTENNA_21/DIODE Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A3
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit1/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/X sky130_fd_sc_hd__mux4_1
Xinput110 N2END[4] vssd1 vssd1 vccd1 vccd1 input110/X sky130_fd_sc_hd__clkbuf_2
Xinput154 S1END[0] vssd1 vssd1 vccd1 vccd1 input154/X sky130_fd_sc_hd__clkbuf_4
Xinput121 N2MID[7] vssd1 vssd1 vccd1 vccd1 input121/X sky130_fd_sc_hd__buf_2
Xinput143 NN4END[14] vssd1 vssd1 vccd1 vccd1 input143/X sky130_fd_sc_hd__clkbuf_1
Xinput132 N4END[4] vssd1 vssd1 vccd1 vccd1 input132/X sky130_fd_sc_hd__clkbuf_1
Xinput165 S2END[7] vssd1 vssd1 vccd1 vccd1 input165/X sky130_fd_sc_hd__buf_2
Xinput176 S4END[11] vssd1 vssd1 vccd1 vccd1 input176/X sky130_fd_sc_hd__clkbuf_1
Xinput187 S4END[7] vssd1 vssd1 vccd1 vccd1 input187/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG1_A0 input109/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput198 SS4END[2] vssd1 vssd1 vccd1 vccd1 input198/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix__095__A input172/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit29_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit13 input54/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit24 input66/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG1 input116/X input168/X
+ input220/X Inst_LUT4AB_switch_matrix__044_/A Inst_LUT4AB_ConfigMem_Inst_Frame10_bit5/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit4/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG1 input146/X input8/X input182/X
+ Inst_LUT4AB_switch_matrix__041_/A Inst_LUT4AB_ConfigMem_Inst_Frame7_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A3 sky130_fd_sc_hd__mux4_2
XFILLER_0_43_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1 input154/X
+ input156/X input164/X input208/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit13/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XN4END_inbuf_9__0_ input126/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S3_A1 Inst_LUT4AB_switch_matrix__045_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG2_A0 Inst_LUT4AB_switch_matrix__054_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_SS4BEG_outbuf_3__0__A SS4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit17 input58/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit28 input70/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XN4BEG_outbuf_1__0_ N4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output382/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput403 output403/A vssd1 vssd1 vccd1 vccd1 NN4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput425 output425/A vssd1 vssd1 vccd1 vccd1 S2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput414 output414/A vssd1 vssd1 vccd1 vccd1 S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput469 output469/A vssd1 vssd1 vccd1 vccd1 W2BEG[5] sky130_fd_sc_hd__buf_2
Xoutput458 output458/A vssd1 vssd1 vccd1 vccd1 SS4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput447 output447/A vssd1 vssd1 vccd1 vccd1 SS4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput436 output436/A vssd1 vssd1 vccd1 vccd1 S4BEG[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0 input102/X
+ input106/X input2/X input34/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit6/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XSS4BEG_outbuf_0__0_ SS4END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 output443/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LB_LUT4c_frame_config_dffesr_cus_mux21_I0mux__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/X
+ Inst_LUT4AB_switch_matrix__058_/X Inst_LUT4AB_ConfigMem_Inst_Frame15_bit9/Q vssd1
+ vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__07_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_49_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit4 input76/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit10_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit28/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit26/Q vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__08_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_68_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit12 input53/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit23 input65/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_ Inst_LUT4AB_switch_matrix__032_/X
+ Inst_LUT4AB_switch_matrix__033_/X Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X sky130_fd_sc_hd__mux2_8
XFILLER_0_75_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XW6BEG_outbuf_1__0_ W6END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output483/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0_A2
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit15_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit24_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit2 input72/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1 input155/X
+ input163/X input207/X input209/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_WW4BEG_outbuf_7__0__A ANTENNA_8/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput277 output277/A vssd1 vssd1 vccd1 vccd1 E6BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_0_10_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput255 output255/A vssd1 vssd1 vccd1 vccd1 E1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput266 output266/A vssd1 vssd1 vccd1 vccd1 E2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput299 output299/A vssd1 vssd1 vccd1 vccd1 EE4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput288 output288/A vssd1 vssd1 vccd1 vccd1 EE4BEG[10] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S0_A2 Inst_LUT4AB_switch_matrix__085_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG2_A2 input229/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_cus_mux41_buf_inst0_A3
+ ANTENNA_21/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG3_A1 input14/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit29_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit27 input69/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit16 input57/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__101_ Inst_LUT4AB_switch_matrix__101_/A vssd1 vssd1 vccd1
+ vccd1 output468/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix__032_ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__032_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit12_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit21_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit2_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xdata_outbuf_30__0_ data_inbuf_30__0_/X vssd1 vssd1 vccd1 vccd1 output326/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit30_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0_A3
+ input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit3_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit7 input79/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_S4BEG_outbuf_1__0__A S4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xdata_outbuf_21__0_ data_inbuf_21__0_/X vssd1 vssd1 vccd1 vccd1 output316/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit11 input52/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit22 input64/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit17_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit8 input80/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_12__0_ data_inbuf_12__0_/X vssd1 vssd1 vccd1 vccd1 output306/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix__098__A ANTENNA_2/DIODE vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XS4BEG_outbuf_1__0_ S4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output434/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit19 input60/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_data_inbuf_24__0__A input66/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LF_SR__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LF_SR__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit2/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__13_/S sky130_fd_sc_hd__mux2_1
XInst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit8/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit19/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit19/Q Inst_LC_LUT4c_frame_config_dffesr__07_/A
+ Inst_LC_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit26 input68/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit15 input56/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG0_A0 Inst_LUT4AB_switch_matrix__034_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG1_A2 input169/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1_A1
+ input165/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG0_A2 input224/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_7 ANTENNA_7/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit6_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit1_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit7_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XNN4END_inbuf_7__0_ input140/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit19 input60/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XW6END_inbuf_3__0_ input233/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit2_GATE input93/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XEE4BEG_outbuf_0__0_ EE4END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 output287/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LA_LUT4c_frame_config_dffesr_cus_mux21_O__0_ Inst_LA_LUT4c_frame_config_dffesr__13_/A0
+ hold1/A Inst_LUT4AB_ConfigMem_Inst_Frame15_bit7/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__032_/A
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_67_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit2 input72/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit14/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit12/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit26/Q Inst_LD_LUT4c_frame_config_dffesr__07_/A
+ Inst_LD_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit2/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit3/Q vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__08_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput100 FrameStrobe[8] vssd1 vssd1 vccd1 vccd1 input100/X sky130_fd_sc_hd__clkbuf_16
Xinput111 N2END[5] vssd1 vssd1 vccd1 vccd1 input111/X sky130_fd_sc_hd__buf_2
Xinput122 N4END[0] vssd1 vssd1 vccd1 vccd1 input122/X sky130_fd_sc_hd__clkbuf_4
Xinput144 NN4END[15] vssd1 vssd1 vccd1 vccd1 input144/X sky130_fd_sc_hd__clkbuf_1
Xinput133 N4END[5] vssd1 vssd1 vccd1 vccd1 input133/X sky130_fd_sc_hd__clkbuf_1
Xinput177 S4END[12] vssd1 vssd1 vccd1 vccd1 input177/X sky130_fd_sc_hd__clkbuf_1
Xinput166 S2MID[0] vssd1 vssd1 vccd1 vccd1 input166/X sky130_fd_sc_hd__clkbuf_4
Xinput155 S1END[1] vssd1 vssd1 vccd1 vccd1 input155/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG1_A1 input9/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput199 SS4END[3] vssd1 vssd1 vccd1 vccd1 input199/X sky130_fd_sc_hd__clkbuf_2
Xinput188 S4END[8] vssd1 vssd1 vccd1 vccd1 input188/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit21_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit30_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_output479_A output479/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1_A0
+ input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit25 input67/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit14 input55/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG2 input18/X input170/X
+ input222/X Inst_LUT4AB_switch_matrix__087_/A Inst_LUT4AB_ConfigMem_Inst_Frame9_bit7/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit6/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_49_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG0 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1 Inst_LUT4AB_switch_matrix__041_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame5_bit30/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit29/Q vssd1 vssd1 vccd1 vccd1 output407/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG2 input129/X input197/X input214/X
+ Inst_LUT4AB_switch_matrix__084_/A Inst_LUT4AB_ConfigMem_Inst_Frame8_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit17_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit13/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit0 input50/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit26_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S3_A2 Inst_LUT4AB_switch_matrix__088_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_NN4BEG_outbuf_11__0__A NN4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG2_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LC_EN__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LC_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame8_bit27/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__14_/S sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst0 input104/X
+ input4/X input208/X Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_ConfigMem_Inst_Frame6_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit22/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit29 input71/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit18 input59/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit5_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput404 output404/A vssd1 vssd1 vccd1 vccd1 NN4BEG[7] sky130_fd_sc_hd__buf_2
XFILLER_0_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput426 output426/A vssd1 vssd1 vccd1 vccd1 S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput415 output415/A vssd1 vssd1 vccd1 vccd1 S2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput459 output459/A vssd1 vssd1 vccd1 vccd1 UserCLKo sky130_fd_sc_hd__buf_1
XFILLER_0_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput448 output448/A vssd1 vssd1 vccd1 vccd1 SS4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput437 output437/A vssd1 vssd1 vccd1 vccd1 S4BEG[4] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit14_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1 input154/X
+ input158/X input206/X input208/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit6/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit6_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_W6BEG_outbuf_6__0__A W6END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit5 input77/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A3 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit29/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit27/Q vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__09_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XEE4BEG_outbuf_10__0_ EE4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 output288/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit13 input54/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit19_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit24 input66/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit28_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit3 input75/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput256 output256/A vssd1 vssd1 vccd1 vccd1 E1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput267 output267/A vssd1 vssd1 vccd1 vccd1 E2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput289 output289/A vssd1 vssd1 vccd1 vccd1 EE4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput278 output278/A vssd1 vssd1 vccd1 vccd1 E6BEG[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S0_A3 Inst_LUT4AB_switch_matrix__101_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG2_A3 Inst_LUT4AB_switch_matrix__034_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_SS4BEG_outbuf_2__0__A SS4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG3_A0 Inst_LUT4AB_switch_matrix__054_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LB_EN__0__517 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LB_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LB_EN__0__517/LO sky130_fd_sc_hd__conb_1
XFILLER_0_37_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG3_A2 input166/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit17 input58/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit28 input70/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit11/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit13/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__066_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_64_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__100_ ANTENNA_3/DIODE vssd1 vssd1 vccd1 vccd1 output467/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_23__0_ input65/X vssd1 vssd1 vccd1 vccd1 data_inbuf_23__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG2_A1 input41/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit8 input80/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit23 input65/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit12 input53/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_2__0_ input94/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_14__0_ input55/X vssd1 vssd1 vccd1 vccd1 data_inbuf_14__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0 input5/X
+ input209/X Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame19_bit21/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit9 input81/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit14_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit23_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_WW4BEG_outbuf_6__0__A WW4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XWW4BEG_outbuf_11__0_ WW4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 output494/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit14/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit13/Q Inst_LC_LUT4c_frame_config_dffesr__07_/A
+ Inst_LC_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit19_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame9_bit23/Q
+ vssd1 vssd1 vccd1 vccd1 output291/A sky130_fd_sc_hd__mux2_1
XFILLER_0_7_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit16 input57/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG0_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit27 input69/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG1_A3 input221/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit28_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1_A2
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG0_A3 Inst_LUT4AB_switch_matrix__068_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG1_A0 input117/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit20_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit11_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_8 ANTENNA_8/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_S4BEG_outbuf_0__0__A ANTENNA_6/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_outbuf_17__0_ strobe_inbuf_17__0_/X vssd1 vssd1 vccd1 vccd1 output343/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit1_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG1_A0 input116/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1_A0
+ input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit2_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit16_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit25_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit3 input75/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4 Inst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ Inst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X Inst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ Inst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X Inst_LD_LUT4c_frame_config_dffesr__09_/A
+ Inst_LD_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__13_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit2/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit0/Q vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__09_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput101 FrameStrobe[9] vssd1 vssd1 vccd1 vccd1 input101/X sky130_fd_sc_hd__clkbuf_16
Xinput145 NN4END[1] vssd1 vssd1 vccd1 vccd1 input145/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput112 N2END[6] vssd1 vssd1 vccd1 vccd1 input112/X sky130_fd_sc_hd__clkbuf_4
Xinput134 N4END[6] vssd1 vssd1 vccd1 vccd1 input134/X sky130_fd_sc_hd__clkbuf_1
Xinput123 N4END[10] vssd1 vssd1 vccd1 vccd1 input123/X sky130_fd_sc_hd__clkbuf_1
Xinput167 S2MID[1] vssd1 vssd1 vccd1 vccd1 input167/X sky130_fd_sc_hd__clkbuf_4
Xinput156 S1END[2] vssd1 vssd1 vccd1 vccd1 input156/X sky130_fd_sc_hd__clkbuf_4
Xinput178 S4END[13] vssd1 vssd1 vccd1 vccd1 input178/X sky130_fd_sc_hd__clkbuf_1
XWW4END_inbuf_8__0_ input241/X vssd1 vssd1 vccd1 vccd1 ANTENNA_9/DIODE sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG1_A2 input161/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput189 S4END[9] vssd1 vssd1 vccd1 vccd1 input189/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_data_inbuf_23__0__A input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1_A1
+ input163/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit15 input56/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit26 input68/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG3 input114/X input14/X
+ input218/X ANTENNA_4/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame9_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit1/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A0 sky130_fd_sc_hd__mux4_2
XFILLER_0_57_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG3 input43/X input174/X input245/X
+ ANTENNA_3/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame8_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A3 sky130_fd_sc_hd__mux4_1
XFILLER_0_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG1 Inst_LUT4AB_switch_matrix__054_/A
+ ANTENNA_21/DIODE Inst_LUT4AB_switch_matrix__038_/A Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit27/Q
+ vssd1 vssd1 vccd1 vccd1 output408/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit13/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit1 input61/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG1_A0 Inst_LUT4AB_switch_matrix__055_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG2_A2 Inst_LUT4AB_switch_matrix__066_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A2 Inst_LUT4AB_ConfigMem_Inst_Frame6_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit22/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit19 input60/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG0 input113/X input42/X input165/X
+ input217/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit5/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A2 sky130_fd_sc_hd__mux4_2
Xoutput405 output405/A vssd1 vssd1 vccd1 vccd1 NN4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput416 output416/A vssd1 vssd1 vccd1 vccd1 S2BEG[5] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit5_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xoutput427 output427/A vssd1 vssd1 vccd1 vccd1 S4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput438 output438/A vssd1 vssd1 vccd1 vccd1 S4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput449 output449/A vssd1 vssd1 vccd1 vccd1 SS4BEG[15] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst0 input102/X
+ input154/X input206/X Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame19_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit23/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit6/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit6_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1_A0
+ input161/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit6 input78/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit11_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit20_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A3 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit28/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit30/Q vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__10_/A
+ sky130_fd_sc_hd__mux4_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit14 input55/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit25 input67/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_14__0_ input87/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_14__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit16_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XE6END_inbuf_8__0_ input23/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame5_bit26/Q
+ vssd1 vssd1 vccd1 vccd1 output396/A sky130_fd_sc_hd__mux2_1
XANTENNA_NN4BEG_outbuf_10__0__A NN4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LH_LUT4c_frame_config_dffesr__12__A1 Inst_LH_LUT4c_frame_config_dffesr__09_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I2_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit4 input76/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput257 output257/A vssd1 vssd1 vccd1 vccd1 E1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput268 output268/A vssd1 vssd1 vccd1 vccd1 E2BEGb[1] sky130_fd_sc_hd__buf_2
XFILLER_0_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput279 output279/A vssd1 vssd1 vccd1 vccd1 E6BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_0_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG3_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG3_A3 ANTENNA_3/DIODE
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit18 input59/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit29 input71/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XE6BEG_outbuf_0__0_ E6END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 output275/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_W6BEG_outbuf_5__0__A W6END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit9_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit22_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit31_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG2_A2 input181/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit9 input81/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst0 input104/X
+ input4/X input208/X Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_ConfigMem_Inst_Frame13_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit21/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LD_SR__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit13 input54/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit24 input66/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit18_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit27_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit20/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit15/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit14/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__041_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XEE4END_inbuf_9__0_ input38/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_6__0_ input78/X vssd1 vssd1 vccd1 vccd1 data_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_SS4BEG_outbuf_1__0__A SS4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2 Inst_LUT4AB_ConfigMem_Inst_Frame18_bit14/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit12/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit12/Q Inst_LC_LUT4c_frame_config_dffesr__07_/A
+ Inst_LC_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit17 input58/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG0_A2 ANTENNA_3/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit28 input70/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1_A3
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG1_A1 input17/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0 input105/X
+ input107/X input7/X input25/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 ANTENNA_9/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG1_A1 input168/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1_A1
+ input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit4 input76/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG1_A0 Inst_LUT4AB_switch_matrix__054_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit2_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit13_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit22_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A3 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit2/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit0/Q vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__10_/A
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame2_bit27/Q
+ vssd1 vssd1 vccd1 vccd1 output498/A sky130_fd_sc_hd__mux2_1
XANTENNA_WW4BEG_outbuf_5__0__A WW4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput102 N1END[0] vssd1 vssd1 vccd1 vccd1 input102/X sky130_fd_sc_hd__buf_4
Xinput124 N4END[11] vssd1 vssd1 vccd1 vccd1 input124/X sky130_fd_sc_hd__clkbuf_1
Xinput113 N2END[7] vssd1 vssd1 vccd1 vccd1 input113/X sky130_fd_sc_hd__clkbuf_4
Xinput135 N4END[7] vssd1 vssd1 vccd1 vccd1 input135/X sky130_fd_sc_hd__clkbuf_1
Xinput168 S2MID[2] vssd1 vssd1 vccd1 vccd1 input168/X sky130_fd_sc_hd__buf_2
Xinput157 S1END[3] vssd1 vssd1 vccd1 vccd1 input157/X sky130_fd_sc_hd__clkbuf_4
Xinput146 NN4END[2] vssd1 vssd1 vccd1 vccd1 input146/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput179 S4END[14] vssd1 vssd1 vccd1 vccd1 input179/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit31_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG1_A3 input245/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1_A2
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit16 input57/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit27 input69/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XNN4BEG_outbuf_0__0_ NN4END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 output391/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XN4BEG_outbuf_4__0_ N4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output385/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit18_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG2 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 Inst_LUT4AB_switch_matrix__039_/A
+ ANTENNA_5/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame6_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit23/Q
+ vssd1 vssd1 vccd1 vccd1 output409/A sky130_fd_sc_hd__mux4_1
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit27_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit12/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit23/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__102_/A
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit2 input72/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG1_A1 ANTENNA_21/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XSS4BEG_outbuf_3__0_ SS4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output452/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG2_A3 ANTENNA_5/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit10_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1_A0
+ input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XSS4BEG_outbuf_11__0_ SS4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 output445/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG1 input109/X input9/X input161/X
+ input245/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A2 sky130_fd_sc_hd__mux4_2
Xoutput406 output406/A vssd1 vssd1 vccd1 vccd1 NN4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput417 output417/A vssd1 vssd1 vccd1 vccd1 S2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput428 output428/A vssd1 vssd1 vccd1 vccd1 S4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput439 output439/A vssd1 vssd1 vccd1 vccd1 S4BEG[6] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A2 Inst_LUT4AB_ConfigMem_Inst_Frame19_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit23/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit15_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit24_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit5_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_switch_matrix__055_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit6/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XW6BEG_outbuf_4__0_ W6END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output486/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit0_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit6_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1_A1
+ input183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit7 input79/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2_A2
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LH_LUT4c_frame_config_dffesr__10__A Inst_LH_LUT4c_frame_config_dffesr__10_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit1_GATE input94/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_22__0__A input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit26 input68/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit15 input56/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG0 input121/X input21/X
+ input173/X input225/X Inst_LUT4AB_ConfigMem_Inst_Frame11_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A1 sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit5 input77/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit24/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__085_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput258 output258/A vssd1 vssd1 vccd1 vccd1 E1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput269 output269/A vssd1 vssd1 vccd1 vccd1 E2BEGb[2] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__101__A Inst_LUT4AB_switch_matrix__101_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG3_A2 ANTENNA_14/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_outbuf_24__0_ data_inbuf_24__0_/X vssd1 vssd1 vccd1 vccd1 output319/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit19 input60/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1_A0
+ input159/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit10/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit11/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit10/Q Inst_LB_LUT4c_frame_config_dffesr__07_/A
+ Inst_LB_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_15__0_ data_inbuf_15__0_/X vssd1 vssd1 vccd1 vccd1 output309/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit9_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XS4BEG_outbuf_4__0_ S4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output437/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit10_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG2_A3 Inst_LUT4AB_switch_matrix__083_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit4_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A2 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit21/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit5_GATE input93/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__089_ input166/X vssd1 vssd1 vccd1 vccd1 output419/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit14 input55/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit21/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XS4END_inbuf_2__0_ input186/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_2__0_/X sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit24_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LA_EN__0__516 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LA_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LA_EN__0__516/LO sky130_fd_sc_hd__conb_1
XInst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit17/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit16/Q Inst_LC_LUT4c_frame_config_dffesr__07_/A
+ Inst_LC_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit0 input50/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit29_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit29 input71/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG0_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit18 input59/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XW6END_inbuf_6__0_ input236/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XEE4BEG_outbuf_3__0_ EE4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output296/A sky130_fd_sc_hd__clkbuf_1
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_W6BEG_outbuf_4__0__A W6END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG1_A2 input169/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit12_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit21_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1 input159/X
+ input181/X input211/X input229/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit30_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit8_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit17_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG1_A2 input220/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit9_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1_A2
+ input190/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit5 input77/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG0 input25/X input160/X input181/X
+ Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_ConfigMem_Inst_Frame9_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 output430/A sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG1_A1 ANTENNA_21/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG1_A0 input108/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0 input109/X
+ input131/X input3/X input9/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
Xinput136 N4END[8] vssd1 vssd1 vccd1 vccd1 input136/X sky130_fd_sc_hd__clkbuf_1
Xinput125 N4END[12] vssd1 vssd1 vccd1 vccd1 input125/X sky130_fd_sc_hd__clkbuf_1
Xinput114 N2MID[0] vssd1 vssd1 vccd1 vccd1 input114/X sky130_fd_sc_hd__clkbuf_4
Xinput103 N1END[1] vssd1 vssd1 vccd1 vccd1 input103/X sky130_fd_sc_hd__buf_4
Xinput169 S2MID[3] vssd1 vssd1 vccd1 vccd1 input169/X sky130_fd_sc_hd__clkbuf_4
Xinput158 S2END[0] vssd1 vssd1 vccd1 vccd1 input158/X sky130_fd_sc_hd__clkbuf_4
Xinput147 NN4END[3] vssd1 vssd1 vccd1 vccd1 input147/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_SS4BEG_outbuf_0__0__A SS4END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1_A0
+ input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst1_A3
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit17 input58/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit28 input70/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG3 Inst_LUT4AB_switch_matrix__056_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1 Inst_LUT4AB_switch_matrix__040_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame4_bit30/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit24/Q vssd1 vssd1 vccd1 vccd1 output410/A sky130_fd_sc_hd__mux4_1
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit3 input75/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG1_A2 Inst_LUT4AB_switch_matrix__081_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame6_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 output447/A sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1_A1
+ input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG0_A0 input131/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG2 input111/X input11/X input197/X
+ input215/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A2 sky130_fd_sc_hd__mux4_2
XANTENNA_output477_A output477/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput407 output407/A vssd1 vssd1 vccd1 vccd1 S1BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput418 output418/A vssd1 vssd1 vccd1 vccd1 S2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput429 output429/A vssd1 vssd1 vccd1 vccd1 S4BEG[11] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG0 input120/X input172/X
+ input224/X Inst_LUT4AB_switch_matrix__068_/A Inst_LUT4AB_ConfigMem_Inst_Frame9_bit0/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit5/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit7/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit5/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__072_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit12_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_WW4BEG_outbuf_4__0__A WW4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XN4END_inbuf_10__0_ input127/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_10__0_/X sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1_A2
+ input213/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit8 input80/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit0_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit21_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit30_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_strobe_inbuf_9__0__A input101/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit1_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit16 input57/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit27 input69/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xdata_outbuf_2__0_ data_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output325/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit17_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit26_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1_A0
+ input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG1 input117/X input17/X
+ input169/X input221/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit1/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I2_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput259 output259/A vssd1 vssd1 vccd1 vccd1 E2BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xdata_inbuf_26__0_ input68/X vssd1 vssd1 vccd1 vccd1 data_inbuf_26__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG3_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_5__0_ input97/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1_A1
+ input181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_inbuf_17__0_ input58/X vssd1 vssd1 vccd1 vccd1 data_inbuf_17__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit12/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit10/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit12/Q Inst_LB_LUT4c_frame_config_dffesr__07_/A
+ Inst_LB_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_49_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit14_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit23_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG2_A0 input129/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_21__0__A input63/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit4_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__112__A input225/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__088_ Inst_LUT4AB_switch_matrix__088_/A vssd1 vssd1 vccd1
+ vccd1 output418/A sky130_fd_sc_hd__buf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LA_SR__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LA_SR__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__13_/S sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit5_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit15 input56/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit19_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit28_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 Inst_LUT4AB_ConfigMem_Inst_Frame19_bit21/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit0 input50/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4 Inst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ Inst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X Inst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ Inst_LC_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X Inst_LC_LUT4c_frame_config_dffesr__09_/A
+ Inst_LC_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__13_/A0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XS4END_inbuf_10__0_ input179/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_10__0_/X sky130_fd_sc_hd__buf_2
XFILLER_0_1_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit1 input61/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix__107__A input220/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit19 input60/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG1_A3 input221/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__033_/A
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG3_A0 input138/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit8_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG1_A3 Inst_LUT4AB_switch_matrix__044_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit9_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG2_A0 input119/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1_A3
+ input238/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit6 input78/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG1 input22/X input161/X input182/X
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame10_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit24/Q
+ vssd1 vssd1 vccd1 vccd1 output431/A sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG1_A2 Inst_LUT4AB_switch_matrix__038_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG1_A0 input116/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit14_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit23_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG1_A1 input8/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I2_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XSS4END_inbuf_0__0_ input200/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_0__0_/X sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1 input25/X
+ input161/X input213/X input245/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput126 N4END[13] vssd1 vssd1 vccd1 vccd1 input126/X sky130_fd_sc_hd__clkbuf_1
Xinput115 N2MID[1] vssd1 vssd1 vccd1 vccd1 input115/X sky130_fd_sc_hd__clkbuf_4
Xinput104 N1END[2] vssd1 vssd1 vccd1 vccd1 input104/X sky130_fd_sc_hd__buf_4
Xinput159 S2END[1] vssd1 vssd1 vccd1 vccd1 input159/X sky130_fd_sc_hd__clkbuf_4
Xinput148 NN4END[4] vssd1 vssd1 vccd1 vccd1 input148/X sky130_fd_sc_hd__clkbuf_1
Xinput137 N4END[9] vssd1 vssd1 vccd1 vccd1 input137/X sky130_fd_sc_hd__clkbuf_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1_A1
+ input158/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit19_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit18 input59/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_2__0_ strobe_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output347/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_346 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit4 input76/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_W6BEG_outbuf_3__0__A W6END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG1_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit11_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit20_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0 input103/X
+ input111/X input3/X input11/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1_A2
+ input164/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG0_A1 input34/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XWW4BEG_outbuf_0__0_ ANTENNA_20/DIODE vssd1 vssd1 vccd1 vccd1 output492/A sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_17__0_ input90/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_17__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG3 input146/X input7/X input159/X
+ input211/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A2 sky130_fd_sc_hd__mux4_2
Xoutput408 output408/A vssd1 vssd1 vccd1 vccd1 S1BEG[1] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit25_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xoutput419 output419/A vssd1 vssd1 vccd1 vccd1 S2BEGb[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG1 input16/X input168/X
+ input220/X Inst_LUT4AB_switch_matrix__041_/A Inst_LUT4AB_ConfigMem_Inst_Frame14_bit11/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit10/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1_A0
+ input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit9 input81/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1_A3
+ input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit28 input70/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit17 input58/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XE6BEG_outbuf_3__0_ E6END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output280/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1_A1
+ input162/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG2 input119/X input19/X
+ input171/X input223/X Inst_LUT4AB_ConfigMem_Inst_Frame10_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit14/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A1 sky130_fd_sc_hd__mux4_1
XInst_MUX8LUT_frame_config_mux_cus_mux21_sEF__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S2/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/S Inst_LUT4AB_ConfigMem_Inst_Frame3_bit29/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/S sky130_fd_sc_hd__mux2_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit7 input79/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XN4END_inbuf_2__0_ input134/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_2__0_/X sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_cus_mux41_buf_inst0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A1
+ ANTENNA_21/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame11_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit30/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1_A2
+ input211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit8/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit7/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit17/Q Inst_LB_LUT4c_frame_config_dffesr__07_/A
+ Inst_LB_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG2_A1 input25/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0 input105/X
+ input113/X input5/X input13/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_WW4BEG_outbuf_3__0__A WW4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit11_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit20_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_9__0_ input81/X vssd1 vssd1 vccd1 vccd1 data_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_strobe_inbuf_8__0__A input100/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit4_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__087_ Inst_LUT4AB_switch_matrix__087_/A vssd1 vssd1 vccd1
+ vccd1 output417/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit16 input57/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit5_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1_A0
+ input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit27/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit19/Q vssd1 vssd1 vccd1 vccd1 output481/A sky130_fd_sc_hd__mux4_1
XFILLER_0_65_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit16_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit25_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_WW4BEG_outbuf_11__0__A WW4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit1 input61/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit2 input72/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit13_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit22_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit31_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LC_LUT4c_frame_config_dffesr_cus_mux21_I0mux__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I0/X
+ Inst_LUT4AB_switch_matrix__059_/X Inst_LUT4AB_ConfigMem_Inst_Frame13_bit13/Q vssd1
+ vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__07_/A sky130_fd_sc_hd__mux2_2
XANTENNA_Inst_LUT4AB_switch_matrix__033__A Inst_LUT4AB_switch_matrix__033_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_20__0__A input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0 input104/X
+ input112/X input4/X input12/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG3_A1 input22/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit18_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit27_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit8_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XNN4BEG_outbuf_3__0_ NN4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output400/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG2_A1 input19/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit3_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XN4BEG_outbuf_7__0_ N4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output388/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit9_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG2 input158/X input183/X input229/X
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_ConfigMem_Inst_Frame10_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit24/Q
+ vssd1 vssd1 vccd1 vccd1 output432/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit7 input79/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG1_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG1_A1 input16/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG1_A2 input160/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit4_GATE input94/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0_A1
+ input106/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LA_LUT4c_frame_config_dffesr__15_ UserCLK hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XSS4BEG_outbuf_6__0_ SS4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output455/A sky130_fd_sc_hd__clkbuf_1
Xinput127 N4END[14] vssd1 vssd1 vccd1 vccd1 input127/X sky130_fd_sc_hd__clkbuf_1
Xinput116 N2MID[2] vssd1 vssd1 vccd1 vccd1 input116/X sky130_fd_sc_hd__clkbuf_4
Xinput105 N1END[3] vssd1 vssd1 vccd1 vccd1 input105/X sky130_fd_sc_hd__buf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput138 NN4END[0] vssd1 vssd1 vccd1 vccd1 input138/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput149 NN4END[5] vssd1 vssd1 vccd1 vccd1 input149/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XS4BEG_outbuf_10__0_ S4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 output428/A sky130_fd_sc_hd__clkbuf_1
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1_A2
+ input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst0_A1
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit19 input60/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit5 input77/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux_cus_mux21_AH__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_AD__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EH__0_/X Inst_MUX8LUT_frame_config_mux_cus_mux21_AH__0_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_AH__0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_4_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XW6BEG_outbuf_7__0_ W6END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output489/A sky130_fd_sc_hd__clkbuf_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1_A0
+ input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1 input155/X
+ input157/X input163/X input207/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1_A3
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG0_A2 input183/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput409 output409/A vssd1 vssd1 vccd1 vccd1 S1BEG[2] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG2 input118/X input18/X
+ input222/X Inst_LUT4AB_switch_matrix__084_/A Inst_LUT4AB_ConfigMem_Inst_Frame4_bit0/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit0/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0
+ sky130_fd_sc_hd__mux4_2
XNN4END_inbuf_0__0_ input148/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_0__0_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit13_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit22_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit7_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1_A1
+ input164/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit31_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit7/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit5/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit6/Q Inst_LA_LUT4c_frame_config_dffesr__07_/A
+ Inst_LA_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit8_GATE input93/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit29 input71/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit18 input59/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_27__0_ data_inbuf_27__0_/X vssd1 vssd1 vccd1 vccd1 output322/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix__041__A Inst_LUT4AB_switch_matrix__041_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit27_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_W6BEG_outbuf_2__0__A W6END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit10_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG3 input115/X input15/X
+ input167/X input219/X Inst_LUT4AB_ConfigMem_Inst_Frame11_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1_A2
+ input214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit8 input80/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_18__0_ data_inbuf_18__0_/X vssd1 vssd1 vccd1 vccd1 output312/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XS4BEG_outbuf_7__0_ S4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output440/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__066_/A
+ Inst_LUT4AB_switch_matrix__039_/A Inst_LUT4AB_switch_matrix__082_/A ANTENNA_2/DIODE
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit30/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1_A0
+ input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1_A3
+ input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit24_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit15_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit6/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit9/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit8/Q Inst_LB_LUT4c_frame_config_dffesr__07_/A
+ Inst_LB_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix__036__A Inst_LUT4AB_switch_matrix__036_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XS4END_inbuf_5__0_ input189/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1 input155/X
+ input157/X input165/X input209/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG2_A2 input229/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__086_ Inst_LUT4AB_switch_matrix__086_/A vssd1 vssd1 vccd1
+ vccd1 output416/A sky130_fd_sc_hd__buf_1
XFILLER_0_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LC_EN__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit17 input58/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1_A1
+ input160/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XW6END_inbuf_9__0_ input228/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XEE4BEG_outbuf_6__0_ EE4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output299/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit0_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit2 input72/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit3 input75/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__069_ Inst_LUT4AB_switch_matrix__069_/A vssd1 vssd1 vccd1
+ vccd1 output363/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit19/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit21/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__097_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_WW4BEG_outbuf_2__0__A WW4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit10_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_strobe_inbuf_7__0__A input99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1 input156/X
+ input164/X input206/X input208/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG3_A2 input210/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG2_A2 input171/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit15_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_WW4BEG_outbuf_10__0__A WW4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG3 input159/X input174/X input226/X
+ Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_ConfigMem_Inst_Frame12_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 output433/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit8 input80/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit3_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit24_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG1_A2 input168/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG1_A3 input246/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0_A2
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I2_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LA_LUT4c_frame_config_dffesr__14_ hold1/X Inst_LA_LUT4c_frame_config_dffesr__13_/X
+ Inst_LA_LUT4c_frame_config_dffesr__14_/S vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit4_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput106 N2END[0] vssd1 vssd1 vccd1 vccd1 input106/X sky130_fd_sc_hd__buf_4
Xinput117 N2MID[3] vssd1 vssd1 vccd1 vccd1 input117/X sky130_fd_sc_hd__clkbuf_4
Xinput139 NN4END[10] vssd1 vssd1 vccd1 vccd1 input139/X sky130_fd_sc_hd__clkbuf_1
Xinput128 N4END[15] vssd1 vssd1 vccd1 vccd1 input128/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__044__A Inst_LUT4AB_switch_matrix__044_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst1_A3
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst0_A2
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit29_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XNN4BEG_outbuf_10__0_ NN4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 output392/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit6 input78/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit21_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit12_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit30_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1_A1
+ input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LG_SR__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LG_SR__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit0/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__13_/S sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__039__A Inst_LUT4AB_switch_matrix__039_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit26_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit17_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0_A1
+ input112/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG0_A3 Inst_LUT4AB_switch_matrix__069_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_outbuf_10__0_ strobe_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 output336/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_5__0_ data_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output330/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_output358_A output358/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG3 input114/X input14/X
+ input166/X ANTENNA_3/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame10_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A0 sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1_A2
+ input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit7_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst0_A1
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit4/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit2/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit15/Q Inst_LA_LUT4c_frame_config_dffesr__07_/A
+ Inst_LA_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_13_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit8_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_inbuf_29__0_ input71/X vssd1 vssd1 vccd1 vccd1 data_inbuf_29__0_/X sky130_fd_sc_hd__clkbuf_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XWW4END_inbuf_1__0_ input249/X vssd1 vssd1 vccd1 vccd1 ANTENNA_7/DIODE sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit19 input60/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1_A0
+ input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_8__0_ input100/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit0 input50/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst1_A3
+ input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit9 input81/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2_A2
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1_A1
+ input162/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4 Inst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ Inst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X Inst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ Inst_LB_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X Inst_LB_LUT4c_frame_config_dffesr__09_/A
+ Inst_LB_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__13_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__052__A input20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit12_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I2_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG2_A3 Inst_LUT4AB_switch_matrix__082_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit21_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit30_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LD_EN__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LD_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit2/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__14_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_15_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix__085_ Inst_LUT4AB_switch_matrix__085_/A vssd1 vssd1 vccd1
+ vccd1 output415/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit18 input59/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LG_EN__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1_A2
+ input212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit17_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit26_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst0 input105/X
+ input5/X input209/X Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_ConfigMem_Inst_Frame5_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit23/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_W6BEG_outbuf_1__0__A W6END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__047__A input15/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XE6END_inbuf_1__0_ input27/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_1__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit3 input75/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LB_LUT4c_frame_config_dffesr__15_ UserCLK hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1_A0
+ input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit4 input76/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__068_ Inst_LUT4AB_switch_matrix__068_/A vssd1 vssd1 vccd1
+ vccd1 output362/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit23_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit14_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_strobe_inbuf_19__0__A input92/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XSS4END_inbuf_3__0_ input203/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput390 output390/A vssd1 vssd1 vccd1 vccd1 N4BEG[9] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst0_A1
+ input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG3_A3 Inst_LUT4AB_switch_matrix__101_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit28_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG1_A0 input138/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG2_A3 input223/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_outbuf_5__0_ strobe_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output350/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit9 input81/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG1_A3 Inst_LUT4AB_switch_matrix__043_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0_A3
+ input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I2_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LA_LUT4c_frame_config_dffesr__13_ Inst_LA_LUT4c_frame_config_dffesr__13_/A0
+ Inst_LA_LUT4c_frame_config_dffesr__13_/A1 Inst_LA_LUT4c_frame_config_dffesr__13_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__13_/X sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG2_A0 input119/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit7/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit9/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__067_/A
+ sky130_fd_sc_hd__mux4_2
Xinput118 N2MID[4] vssd1 vssd1 vccd1 vccd1 input118/X sky130_fd_sc_hd__buf_2
Xinput107 N2END[1] vssd1 vssd1 vccd1 vccd1 input107/X sky130_fd_sc_hd__clkbuf_2
Xinput129 N4END[1] vssd1 vssd1 vccd1 vccd1 input129/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG1_A0 input116/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XEE4END_inbuf_2__0_ input46/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XWW4BEG_outbuf_3__0_ WW4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output501/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit7 input79/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_13_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0 input4/X
+ input208/X Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame1_bit26/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit18/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_WW4BEG_outbuf_1__0__A ANTENNA_7/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1_A2
+ input158/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_strobe_inbuf_6__0__A input98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_7_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG0_A0 input131/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0__515 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0__515/HI
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A0 sky130_fd_sc_hd__conb_1
XANTENNA_Inst_LG_LUT4c_frame_config_dffesr__09__A Inst_LG_LUT4c_frame_config_dffesr__09_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0_A2
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix__055__A Inst_LUT4AB_switch_matrix__055_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XE6BEG_outbuf_6__0_ E6END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output283/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit23_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit14_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1_A3
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst0_A2
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit7_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2 Inst_LUT4AB_ConfigMem_Inst_Frame18_bit11/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit9/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit7/Q Inst_LA_LUT4c_frame_config_dffesr__07_/A
+ Inst_LA_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XN4END_inbuf_5__0_ input137/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_5__0_/X sky130_fd_sc_hd__buf_2
XFILLER_0_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit2_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit8_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit19_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit3_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1_A1
+ input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit1 input61/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit11_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit20_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0_A1
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst2_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit16_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1_A2
+ input214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG2_A0 input106/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit25_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1_A0
+ input162/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__084_ Inst_LUT4AB_switch_matrix__084_/A vssd1 vssd1 vccd1
+ vccd1 output414/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit6_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit19 input60/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1_A3
+ input247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__056_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A2 Inst_LUT4AB_ConfigMem_Inst_Frame5_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit23/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit7_GATE input94/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0_A0
+ input146/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst0 input103/X
+ input155/X input207/X Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_ConfigMem_Inst_Frame1_bit29/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit28/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit4 input76/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LB_LUT4c_frame_config_dffesr__14_ hold9/X Inst_LB_LUT4c_frame_config_dffesr__13_/X
+ Inst_LB_LUT4c_frame_config_dffesr__14_/S vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__mux2_1
XFILLER_0_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1_A1
+ input160/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit5 input77/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix__067_ Inst_LUT4AB_switch_matrix__067_/A vssd1 vssd1 vccd1
+ vccd1 output361/A sky130_fd_sc_hd__buf_1
XNN4BEG_outbuf_6__0_ NN4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output403/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit11_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit20_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG3_A0 input43/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XSS4BEG_outbuf_9__0_ SS4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output458/A sky130_fd_sc_hd__clkbuf_1
Xoutput380 output380/A vssd1 vssd1 vccd1 vccd1 N4BEG[14] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput391 output391/A vssd1 vssd1 vccd1 vccd1 NN4BEG[0] sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst0_A2
+ input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit25_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit16_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG1_A1 input8/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_W6BEG_outbuf_0__0__A W6END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LA_LUT4c_frame_config_dffesr__12_ Inst_LA_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__057_/X
+ Inst_LA_LUT4c_frame_config_dffesr__11_/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__058_/A
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG2_A1 input19/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput108 N2END[2] vssd1 vssd1 vccd1 vccd1 input108/X sky130_fd_sc_hd__buf_2
Xinput119 N2MID[5] vssd1 vssd1 vccd1 vccd1 input119/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG1_A1 input16/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst0 input105/X
+ input5/X input209/X Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_ConfigMem_Inst_Frame5_bit28/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit21/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit13_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit8 input80/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit18/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit22_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst0_A1
+ input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XNN4END_inbuf_3__0_ input151/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit31_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_strobe_inbuf_18__0__A input91/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1_A3
+ input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit19/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__042_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_75_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_data_inbuf_9__0__A input81/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput90 FrameStrobe[17] vssd1 vssd1 vccd1 vccd1 input90/X sky130_fd_sc_hd__buf_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG0_A1 input9/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit18_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit27_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0_A3
+ input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix__071__A Inst_LUT4AB_switch_matrix__071_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG2_A1 input11/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3 Inst_LUT4AB_ConfigMem_Inst_Frame18_bit6/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit4/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit3/Q Inst_LA_LUT4c_frame_config_dffesr__07_/A
+ Inst_LA_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0 input102/X
+ input108/X input8/X input22/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit18/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XN4BEG_outbuf_10__0_ N4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 output376/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit2_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_442 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0_A1
+ input113/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit3_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1_A2
+ input164/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__066__A Inst_LUT4AB_switch_matrix__066_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame7_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 output394/A sky130_fd_sc_hd__mux2_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit2 input72/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_WW4BEG_outbuf_0__0__A ANTENNA_20/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XS4END_inbuf_8__0_ input177/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_strobe_inbuf_5__0__A input97/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LC_LUT4c_frame_config_dffesr__15_ UserCLK hold16/X vssd1 vssd1 vccd1 vccd1 hold15/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1_A3
+ input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG2_A1 input131/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XEE4BEG_outbuf_9__0_ EE4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output302/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit13_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit0 input50/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I2_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit22_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit19/Q vssd1 vssd1 vccd1 vccd1 ANTENNA_4/DIODE
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1_A1
+ input174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__083_ Inst_LUT4AB_switch_matrix__083_/A vssd1 vssd1 vccd1
+ vccd1 output413/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0 input145/X
+ input5/X input7/X input25/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit18_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit6_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_EE4BEG_outbuf_9__0__A EE4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit27_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst0_A1
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit1_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit7_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0_A1
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit10_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__066_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A2 Inst_LUT4AB_ConfigMem_Inst_Frame1_bit29/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit28/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit5 input77/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LB_LUT4c_frame_config_dffesr__13_ Inst_LB_LUT4c_frame_config_dffesr__13_/A0
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit8/Q Inst_LB_LUT4c_frame_config_dffesr__13_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__13_/X sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1_A2
+ input212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit6 input78/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__066_ Inst_LUT4AB_switch_matrix__066_/A vssd1 vssd1 vccd1
+ vccd1 output360/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit24_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit15_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LG_LUT4c_frame_config_dffesr__11__A1 Inst_LG_LUT4c_frame_config_dffesr__09_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1_A0
+ input160/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_10__0_ input51/X vssd1 vssd1 vccd1 vccd1 data_inbuf_10__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG3_A1 input174/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput370 output370/A vssd1 vssd1 vccd1 vccd1 N2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput392 output392/A vssd1 vssd1 vccd1 vccd1 NN4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput381 output381/A vssd1 vssd1 vccd1 vccd1 N4BEG[15] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit13/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__086_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit29_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__074__A input115/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG1_A2 input160/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LA_LUT4c_frame_config_dffesr__11_ Inst_LA_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__057_/X
+ Inst_LA_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__11_/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG2_A2 input171/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput109 N2END[3] vssd1 vssd1 vccd1 vccd1 input109/X sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix__049_ input17/X vssd1 vssd1 vccd1 vccd1 output270/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame2_bit28/Q
+ vssd1 vssd1 vccd1 vccd1 output496/A sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG0_A0 input25/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG1_A2 input220/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__069__A Inst_LUT4AB_switch_matrix__069_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__056_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A2 Inst_LUT4AB_ConfigMem_Inst_Frame5_bit28/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit21/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit0 input50/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_13__0_ strobe_inbuf_13__0_/X vssd1 vssd1 vccd1 vccd1 output339/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit9 input81/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_8__0_ data_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output333/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit26/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit18/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst0_A2
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I2_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit10_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput80 FrameData[8] vssd1 vssd1 vccd1 vccd1 input80/X sky130_fd_sc_hd__buf_8
Xinput91 FrameStrobe[18] vssd1 vssd1 vccd1 vccd1 input91/X sky130_fd_sc_hd__buf_8
XFILLER_0_12_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG0_A2 input213/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XWW4END_inbuf_4__0_ input252/X vssd1 vssd1 vccd1 vccd1 WW4END_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit15_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit24_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG2_A2 input163/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4 Inst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ Inst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X Inst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ Inst_LA_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X Inst_LA_LUT4c_frame_config_dffesr__09_/A
+ Inst_LA_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__13_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1 input160/X
+ input182/X input212/X input226/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit18/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG0 input131/X input34/X input183/X
+ Inst_LUT4AB_switch_matrix__069_/A Inst_LUT4AB_ConfigMem_Inst_Frame11_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit30/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A3 sky130_fd_sc_hd__mux4_1
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit29_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0_A2
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst1_A3
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit12_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit21_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit3 input75/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit30_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__082__A Inst_LUT4AB_switch_matrix__082_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_strobe_inbuf_17__0__A input90/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output356_A output356/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0_A3
+ input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_8__0__A input80/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0 input110/X
+ input122/X input4/X input10/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit5/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LG_SR__0__514 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LG_SR__0__514/HI
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LG_SR__0_/A0 sky130_fd_sc_hd__conb_1
XInst_LC_LUT4c_frame_config_dffesr__14_ hold15/X Inst_LC_LUT4c_frame_config_dffesr__13_/X
+ Inst_LC_LUT4c_frame_config_dffesr__14_/S vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__mux2_1
XFILLER_0_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit17_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit26_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG2_A2 input229/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit1 input61/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xstrobe_inbuf_10__0_ input83/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_10__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__077__A input118/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0_A1
+ input111/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XE6END_inbuf_4__0_ input30/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1_A2
+ input214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output473_A output473/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__082_ Inst_LUT4AB_switch_matrix__082_/A vssd1 vssd1 vccd1
+ vccd1 output412/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1 input159/X
+ input181/X input211/X input229/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst0_A2
+ input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0_A2
+ input42/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit1_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG3_A0 input159/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix__039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit2_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XSS4END_inbuf_6__0_ input191/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_strobe_inbuf_4__0__A input96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit6 input78/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LB_LUT4c_frame_config_dffesr__12_ Inst_LB_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__058_/X
+ Inst_LB_LUT4c_frame_config_dffesr__11_/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__059_/A
+ sky130_fd_sc_hd__a21o_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst1_A3
+ input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit7 input79/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__065_ ANTENNA_13/DIODE vssd1 vssd1 vccd1 vccd1 output359/A
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_outbuf_8__0_ strobe_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output353/A sky130_fd_sc_hd__clkbuf_1
Xinput1 Ci vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit12_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1_A1
+ input182/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit30_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG3_A2 input245/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput371 output371/A vssd1 vssd1 vccd1 vccd1 N2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput360 output360/A vssd1 vssd1 vccd1 vccd1 N2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput393 output393/A vssd1 vssd1 vccd1 vccd1 NN4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput382 output382/A vssd1 vssd1 vccd1 vccd1 N4BEG[1] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst0_A1
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit23/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit27/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XEE4END_inbuf_5__0_ input49/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_2__0_ input72/X vssd1 vssd1 vccd1 vccd1 data_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__090__A input167/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_EE4BEG_outbuf_8__0__A EE4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit17_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit26_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG1_A3 input212/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XWW4BEG_outbuf_6__0_ WW4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output504/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LA_LUT4c_frame_config_dffesr__10_ Inst_LA_LUT4c_frame_config_dffesr__10_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__10_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_24_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG2_A3 input223/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit5_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__048_ input16/X vssd1 vssd1 vccd1 vccd1 output269/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG0_A1 input160/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG1_A3 Inst_LUT4AB_switch_matrix__042_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_31__0__A input74/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit6_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG2_A0 input119/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG1_A0 input16/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LB_SR__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LB_SR__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__13_/S sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit1 input61/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix__085__A Inst_LUT4AB_switch_matrix__085_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit14_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit23_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XE6BEG_outbuf_9__0_ E6END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output286/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0 Inst_LUT4AB_ConfigMem_Inst_Frame1_bit26/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit18/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I2_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XN4END_inbuf_8__0_ input125/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_2
Xinput70 FrameData[28] vssd1 vssd1 vccd1 vccd1 input70/X sky130_fd_sc_hd__buf_8
Xinput81 FrameData[9] vssd1 vssd1 vccd1 vccd1 input81/X sky130_fd_sc_hd__buf_8
Xinput92 FrameStrobe[19] vssd1 vssd1 vccd1 vccd1 input92/X sky130_fd_sc_hd__buf_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit19_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG0_A3 Inst_LUT4AB_switch_matrix__068_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit28_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LD_LUT4c_frame_config_dffesr__15_ UserCLK hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG2_A3 input215/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XN4BEG_outbuf_0__0_ N4END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 output375/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit18/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit9_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG1 input130/X input198/X input212/X
+ Inst_LUT4AB_switch_matrix__042_/A Inst_LUT4AB_ConfigMem_Inst_Frame4_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A3 sky130_fd_sc_hd__mux4_1
XFILLER_0_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0_A3
+ input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LC_SR__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit4 input76/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LD_LUT4c_frame_config_dffesr_cus_mux21_I0mux__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/X
+ Inst_LUT4AB_switch_matrix__060_/X Inst_LUT4AB_ConfigMem_Inst_Frame15_bit21/Q vssd1
+ vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__07_/A sky130_fd_sc_hd__mux2_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst0_A1
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0_A1
+ input113/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1 input22/X
+ input162/X input214/X input226/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit5/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XW6BEG_outbuf_0__0_ W6END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 output480/A sky130_fd_sc_hd__clkbuf_1
XInst_MUX8LUT_frame_config_mux_cus_mux21_GH__0_ Inst_LUT4AB_switch_matrix__055_/X
+ Inst_LUT4AB_switch_matrix__056_/X Inst_MUX8LUT_frame_config_mux_cus_mux21_GH__0_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_GH__0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LC_LUT4c_frame_config_dffesr__13_ Inst_LC_LUT4c_frame_config_dffesr__13_/A0
+ Inst_LC_LUT4c_frame_config_dffesr__13_/A1 Inst_LC_LUT4c_frame_config_dffesr__13_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__13_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG2_A3 Inst_LUT4AB_switch_matrix__055_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit14_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit23_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame12_bit1/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit4/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0_A2
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix__093__A input170/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1_A3
+ input246/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0 input104/X
+ input112/X input4/X input12/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit14/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix__081_ Inst_LUT4AB_switch_matrix__081_/A vssd1 vssd1 vccd1
+ vccd1 output411/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit28_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit19_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__033_/A
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XNN4BEG_outbuf_9__0_ NN4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output406/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0_A3
+ input22/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG3_A1 input174/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit11_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1_A1 Inst_LUT4AB_switch_matrix__043_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_outbuf_20__0_ data_inbuf_20__0_/X vssd1 vssd1 vccd1 vccd1 output315/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit20_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit1_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_strobe_inbuf_16__0__A input89/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG0_A0 Inst_LUT4AB_switch_matrix__036_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix__082_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit2_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit7 input79/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LB_LUT4c_frame_config_dffesr__11_ Inst_LB_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__058_/X
+ Inst_LB_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__11_/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_data_inbuf_7__0__A input79/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xdata_outbuf_11__0_ data_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 output305/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix__088__A Inst_LUT4AB_switch_matrix__088_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit16_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XS4BEG_outbuf_0__0_ ANTENNA_6/DIODE vssd1 vssd1 vccd1 vccd1 output427/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit8 input80/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_43_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XInst_LUT4AB_switch_matrix__064_ Inst_LUT4AB_switch_matrix__064_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__064_/X sky130_fd_sc_hd__buf_1
XFILLER_0_60_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0_A1
+ input109/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput2 E1END[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_4
XANTENNA_Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4_S0
+ Inst_LH_LUT4c_frame_config_dffesr__09_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1_A2
+ input212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG3_A3 ANTENNA_3/DIODE
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput350 output350/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput361 output361/A vssd1 vssd1 vccd1 vccd1 N2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput394 output394/A vssd1 vssd1 vccd1 vccd1 NN4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput383 output383/A vssd1 vssd1 vccd1 vccd1 N4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput372 output372/A vssd1 vssd1 vccd1 vccd1 N2BEGb[5] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst0_A2
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame12_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit29/Q vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__08_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XNN4END_inbuf_6__0_ input139/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_11_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__047_ input15/X vssd1 vssd1 vccd1 vccd1 output268/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XW6END_inbuf_2__0_ input232/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_strobe_inbuf_3__0__A input95/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit5_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG0_A2 input181/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0 input102/X
+ input138/X input2/X input6/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit0_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG2_A1 input19/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit6_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG1_A1 input168/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit2 input72/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit31/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit30/Q vssd1 vssd1 vccd1 vccd1 output482/A sky130_fd_sc_hd__mux4_1
XFILLER_0_68_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I2_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit20_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG0_A0 input9/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput60 FrameData[19] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__buf_8
Xinput71 FrameData[29] vssd1 vssd1 vccd1 vccd1 input71/X sky130_fd_sc_hd__buf_8
Xinput82 FrameStrobe[0] vssd1 vssd1 vccd1 vccd1 input82/X sky130_fd_sc_hd__buf_8
XFILLER_0_3_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput93 FrameStrobe[1] vssd1 vssd1 vccd1 vccd1 input93/X sky130_fd_sc_hd__clkbuf_16
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_EE4BEG_outbuf_7__0__A EE4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LD_LUT4c_frame_config_dffesr__14_ hold11/X Inst_LD_LUT4c_frame_config_dffesr__13_/X
+ Inst_LD_LUT4c_frame_config_dffesr__14_/S vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit16_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit25_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame12_bit0/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit3/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG2_A0 input111/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__096__A input173/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_data_inbuf_30__0__A input73/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit18/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit9_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG2 input25/X input181/X input247/X
+ Inst_LUT4AB_switch_matrix__085_/A Inst_LUT4AB_ConfigMem_Inst_Frame6_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit28/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A3 sky130_fd_sc_hd__mux4_1
XFILLER_0_48_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0 input105/X
+ input113/X input5/X input13/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit4_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG3_A0 Inst_LUT4AB_switch_matrix__055_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit13_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit5_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LG_SR__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit31_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit5 input77/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst0_A2
+ input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0_A2
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput250 WW4END[6] vssd1 vssd1 vccd1 vccd1 input250/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit5/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LC_LUT4c_frame_config_dffesr__12_ Inst_LC_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__059_/X
+ Inst_LC_LUT4c_frame_config_dffesr__11_/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__060_/A
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit27_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit18_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit3 input75/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_cus_mux41_buf_inst0_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit1/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit1/Q vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__08_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst0_A3
+ input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_inbuf_31__0_ input74/X vssd1 vssd1 vccd1 vccd1 data_inbuf_31__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__080_ input121/X vssd1 vssd1 vccd1 vccd1 output374/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1 input154/X
+ input156/X input164/X input208/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit14/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG0 Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1 Inst_LUT4AB_switch_matrix__068_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit24/Q vssd1 vssd1 vccd1 vccd1 output255/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_inbuf_22__0_ input64/X vssd1 vssd1 vccd1 vccd1 data_inbuf_22__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst0_A1
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG0 input147/X input183/X input238/X
+ Inst_LUT4AB_switch_matrix__066_/A Inst_LUT4AB_ConfigMem_Inst_Frame1_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit20/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3 sky130_fd_sc_hd__mux4_2
XFILLER_0_14_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0_A1
+ input111/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG3_A2 input226/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1_A2 Inst_LUT4AB_switch_matrix__086_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG0_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_cus_mux41_buf_inst1_A3
+ ANTENNA_2/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_1__0_ input93/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_1__0_/X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_13__0_ input54/X vssd1 vssd1 vccd1 vccd1 data_inbuf_13__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LB_LUT4c_frame_config_dffesr__10_ Inst_LB_LUT4c_frame_config_dffesr__10_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__10_/Y sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit8 input80/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LF_SR__0__513 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LF_SR__0__513/HI
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LF_SR__0_/A0 sky130_fd_sc_hd__conb_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/A0
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AH__0_/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit29/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_55_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit9 input81/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XWW4BEG_outbuf_10__0_ WW4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 output493/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__063_ Inst_LUT4AB_switch_matrix__063_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__063_/X sky130_fd_sc_hd__buf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0_A2
+ input131/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4_S1
+ Inst_LH_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput3 E1END[1] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_4
XFILLER_0_36_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit13_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit22_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG3_A0 input122/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1_A3
+ input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0__523 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0__523/LO sky130_fd_sc_hd__conb_1
XFILLER_0_34_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0_A0
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput362 output362/A vssd1 vssd1 vccd1 vccd1 N2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput340 output340/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput351 output351/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[6] sky130_fd_sc_hd__clkbuf_4
Xoutput384 output384/A vssd1 vssd1 vccd1 vccd1 N4BEG[3] sky130_fd_sc_hd__buf_2
Xoutput373 output373/A vssd1 vssd1 vccd1 vccd1 N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput395 output395/A vssd1 vssd1 vccd1 vccd1 NN4BEG[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A3 Inst_LUT4AB_ConfigMem_Inst_Frame10_bit28/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit27/Q vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__09_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit18_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0_A0
+ input109/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit27_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix__099__A ANTENNA_14/DIODE vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_16__0_ strobe_inbuf_16__0_/X vssd1 vssd1 vccd1 vccd1 output342/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LE_LUT4c_frame_config_dffesr__15_ UserCLK hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_28_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit10_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_strobe_inbuf_15__0__A input88/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__046_ input14/X vssd1 vssd1 vccd1 vccd1 output267/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_data_inbuf_6__0__A input78/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG0_A3 Inst_LUT4AB_switch_matrix__032_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1 input154/X
+ input156/X input158/X input206/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG1_A0 Inst_LUT4AB_switch_matrix__036_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG2_A2 input171/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit0_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0_A1
+ input107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinst_clk_buf UserCLK vssd1 vssd1 vccd1 vccd1 output459/A sky130_fd_sc_hd__clkbuf_16
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG1_A2 input220/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XWW4END_inbuf_7__0_ input240/X vssd1 vssd1 vccd1 vccd1 ANTENNA_8/DIODE sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit1_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit15_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst0 input104/X
+ input4/X input156/X Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_ConfigMem_Inst_Frame13_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit3 input75/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit24_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG0_A1 input199/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput50 FrameData[0] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_8
Xinput61 FrameData[1] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__buf_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit29_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput72 FrameData[2] vssd1 vssd1 vccd1 vccd1 input72/X sky130_fd_sc_hd__buf_8
Xinput94 FrameStrobe[2] vssd1 vssd1 vccd1 vccd1 input94/X sky130_fd_sc_hd__buf_12
Xinput83 FrameStrobe[10] vssd1 vssd1 vccd1 vccd1 input83/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LD_LUT4c_frame_config_dffesr__13_ Inst_LD_LUT4c_frame_config_dffesr__13_/A0
+ Inst_LD_LUT4c_frame_config_dffesr__13_/A1 Inst_LD_LUT4c_frame_config_dffesr__13_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__13_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_74_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit1 input61/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame8_bit1/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit0/Q vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__08_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG2_A1 input11/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_strobe_inbuf_2__0__A input94/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit17/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit16/Q vssd1 vssd1 vccd1 vccd1 ANTENNA_2/DIODE
+ sky130_fd_sc_hd__mux4_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG3 input138/X input22/X input210/X
+ Inst_LUT4AB_switch_matrix__101_/A Inst_LUT4AB_ConfigMem_Inst_Frame7_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit29/Q
+ vssd1 vssd1 vccd1 vccd1 ANTENNA_5/DIODE sky130_fd_sc_hd__mux4_2
XFILLER_0_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1 input157/X
+ input165/X input207/X input209/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit4_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG3_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit5_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit6 input78/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit10_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_13__0_ input86/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_13__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0_A3
+ input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput251 WW4END[7] vssd1 vssd1 vccd1 vccd1 input251/X sky130_fd_sc_hd__clkbuf_1
Xinput240 WW4END[11] vssd1 vssd1 vccd1 vccd1 input240/X sky130_fd_sc_hd__clkbuf_1
XE6END_inbuf_7__0_ input33/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit5/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_416 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LH_LUT4c_frame_config_dffesr__11__A1 Inst_LH_LUT4c_frame_config_dffesr__09_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG0 input113/X input13/X input165/X
+ input238/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit6/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A2 sky130_fd_sc_hd__mux4_2
XInst_LC_LUT4c_frame_config_dffesr__11_ Inst_LC_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__059_/X
+ Inst_LC_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__11_/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_EE4BEG_outbuf_6__0__A EE4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit15_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0_A1
+ input113/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit4 input76/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A3 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit0/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit0/Q vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__09_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XSS4END_inbuf_9__0_ input194/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit1/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__13_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit14/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit29_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG1 Inst_LUT4AB_switch_matrix__037_/A
+ ANTENNA_21/DIODE ANTENNA_13/DIODE Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 output256/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit14/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit15/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__081_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst0_A2
+ input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput500 output500/A vssd1 vssd1 vccd1 vccd1 WW4BEG[2] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG1 input42/X input182/X input217/X
+ Inst_LUT4AB_switch_matrix__039_/A Inst_LUT4AB_ConfigMem_Inst_Frame8_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit13/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A3 sky130_fd_sc_hd__mux4_1
XFILLER_0_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0_A2
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit8_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit21_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit30_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG3_A3 Inst_LUT4AB_switch_matrix__036_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1_A3 Inst_LUT4AB_switch_matrix__102_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG0_A2 Inst_LUT4AB_switch_matrix__068_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit9_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG0 input121/X input21/X
+ input173/X input225/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit13/Q
+ vssd1 vssd1 vccd1 vccd1 ANTENNA_21/DIODE sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit9 input81/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux_cus_mux21_sCD__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_AD__0_/S
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/S Inst_LUT4AB_ConfigMem_Inst_Frame4_bit24/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_CD__0_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit26_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit17_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XEE4END_inbuf_8__0_ input37/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_inbuf_5__0_ input77/X vssd1 vssd1 vccd1 vccd1 data_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__062_ Inst_LUT4AB_switch_matrix__062_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__062_/X sky130_fd_sc_hd__buf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0_A3
+ input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XWW4BEG_outbuf_9__0_ WW4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output507/A sky130_fd_sc_hd__clkbuf_1
Xinput4 E1END[2] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__buf_4
XFILLER_0_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG3_A1 input190/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0_A1
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput341 output341/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput352 output352/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
Xoutput330 output330/A vssd1 vssd1 vccd1 vccd1 FrameData_O[5] sky130_fd_sc_hd__buf_2
Xoutput396 output396/A vssd1 vssd1 vccd1 vccd1 NN4BEG[14] sky130_fd_sc_hd__buf_2
Xoutput385 output385/A vssd1 vssd1 vccd1 vccd1 N4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput374 output374/A vssd1 vssd1 vccd1 vccd1 N2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput363 output363/A vssd1 vssd1 vccd1 vccd1 N2BEG[4] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A3 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit26/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit31/Q vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__10_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0_A1
+ input131/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LE_LUT4c_frame_config_dffesr__14_ hold5/X Inst_LE_LUT4c_frame_config_dffesr__13_/X
+ Inst_LE_LUT4c_frame_config_dffesr__14_/S vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__mux2_1
XFILLER_0_16_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix__045_ Inst_LUT4AB_switch_matrix__045_/A vssd1 vssd1 vccd1
+ vccd1 output266/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG1_A1 ANTENNA_21/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_20 ANTENNA_20/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG2_A3 input223/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LE_EN__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LE_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit4/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__14_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_6_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0_A2
+ input129/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG1_A3 Inst_LUT4AB_switch_matrix__041_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG2_A0 input119/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit1_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A2 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit4 input76/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit12_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit21_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst0 input102/X
+ input2/X input206/X Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame4_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit21/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit30_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0_A0
+ input107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XN4BEG_outbuf_3__0_ N4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output384/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0 input5/X
+ input209/X Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame5_bit29/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit29/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG0_A2 input246/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput40 EE4END[15] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__clkbuf_1
Xinput73 FrameData[30] vssd1 vssd1 vccd1 vccd1 input73/X sky130_fd_sc_hd__buf_8
Xinput62 FrameData[20] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__buf_8
Xinput51 FrameData[10] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_8
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG2_A0 input18/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput95 FrameStrobe[3] vssd1 vssd1 vccd1 vccd1 input95/X sky130_fd_sc_hd__clkbuf_16
Xinput84 FrameStrobe[11] vssd1 vssd1 vccd1 vccd1 input84/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XSS4BEG_outbuf_2__0_ SS4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output451/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit17_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LD_LUT4c_frame_config_dffesr__12_ Inst_LD_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__060_/X
+ Inst_LD_LUT4c_frame_config_dffesr__11_/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__061_/A
+ sky130_fd_sc_hd__a21o_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit26_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit2 input72/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A3 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit4/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit3/Q vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__09_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG2_A2 input197/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XSS4BEG_outbuf_10__0_ SS4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 output444/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_strobe_inbuf_14__0__A input87/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_data_inbuf_5__0__A input77/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux_cus_mux21_AD__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_CD__0_/X Inst_MUX8LUT_frame_config_mux_cus_mux21_AD__0_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_AD__0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_21_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XW6BEG_outbuf_3__0_ W6END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output485/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_71_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG2_A0 Inst_LUT4AB_switch_matrix__056_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit14_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit23_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG3_A2 Inst_LUT4AB_switch_matrix__067_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit4_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit7 input79/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit5_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput252 WW4END[8] vssd1 vssd1 vccd1 vccd1 input252/X sky130_fd_sc_hd__clkbuf_1
Xinput241 WW4END[12] vssd1 vssd1 vccd1 vccd1 input241/X sky130_fd_sc_hd__clkbuf_1
Xinput230 W6END[2] vssd1 vssd1 vccd1 vccd1 input230/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit19_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit8/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit11/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__068_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_14_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XInst_LC_LUT4c_frame_config_dffesr__10_ Inst_LC_LUT4c_frame_config_dffesr__10_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__10_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG1 input109/X input9/X input190/X
+ input213/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit14/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A2 sky130_fd_sc_hd__mux4_2
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0_A2
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG0 input20/X input172/X
+ input224/X Inst_LUT4AB_switch_matrix__069_/A Inst_LUT4AB_ConfigMem_Inst_Frame12_bit5/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit2/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit5 input77/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_23__0_ data_inbuf_23__0_/X vssd1 vssd1 vccd1 vccd1 output318/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A3 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit1/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit0/Q vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__10_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_strobe_inbuf_1__0__A input93/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit14/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xdata_outbuf_14__0_ data_inbuf_14__0_/X vssd1 vssd1 vccd1 vccd1 output308/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG2 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 Inst_LUT4AB_switch_matrix__066_/A
+ ANTENNA_5/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame3_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit24/Q
+ vssd1 vssd1 vccd1 vccd1 output257/A sky130_fd_sc_hd__mux4_1
XS4BEG_outbuf_3__0_ S4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output436/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG2 input129/X input25/X input229/X
+ Inst_LUT4AB_switch_matrix__082_/A Inst_LUT4AB_ConfigMem_Inst_Frame7_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit19/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A3 sky130_fd_sc_hd__mux4_2
Xoutput501 output501/A vssd1 vssd1 vccd1 vccd1 WW4BEG[3] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0_A3
+ input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_MUX8LUT_frame_config_mux_cus_mux21_EH_GH__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_GH__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EH__0_/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit24/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/A0 sky130_fd_sc_hd__mux2_1
XFILLER_0_5_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit8_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG0_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG1 input117/X input17/X
+ input169/X input221/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit4/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 sky130_fd_sc_hd__mux4_2
XInst_LF_LUT4c_frame_config_dffesr__15_ UserCLK hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit3_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit9_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit4_GATE input93/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XS4END_inbuf_1__0_ input185/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_1__0_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit2 input72/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0_A1
+ input111/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_EE4BEG_outbuf_5__0__A EE4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__061_ Inst_LUT4AB_switch_matrix__061_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__061_/X sky130_fd_sc_hd__buf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit23_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xinput5 E1END[3] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_4
XFILLER_0_36_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG3_A2 input226/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LE_LUT4c_frame_config_dffesr__10__A Inst_LE_LUT4c_frame_config_dffesr__10_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XNN4END_inbuf_9__0_ input142/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0_A2
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput353 output353/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[8] sky130_fd_sc_hd__clkbuf_4
Xoutput342 output342/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput320 output320/A vssd1 vssd1 vccd1 vccd1 FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput331 output331/A vssd1 vssd1 vccd1 vccd1 FrameData_O[6] sky130_fd_sc_hd__clkbuf_4
XW6END_inbuf_5__0_ input235/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_2
Xoutput386 output386/A vssd1 vssd1 vccd1 vccd1 N4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput375 output375/A vssd1 vssd1 vccd1 vccd1 N4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput364 output364/A vssd1 vssd1 vccd1 vccd1 N2BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XEE4BEG_outbuf_2__0_ EE4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output295/A sky130_fd_sc_hd__clkbuf_1
Xoutput397 output397/A vssd1 vssd1 vccd1 vccd1 NN4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit0 input50/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit28_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit19_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0_A2
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LE_LUT4c_frame_config_dffesr__13_ Inst_LE_LUT4c_frame_config_dffesr__13_/A0
+ Inst_LE_LUT4c_frame_config_dffesr__13_/A1 Inst_LE_LUT4c_frame_config_dffesr__13_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__13_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_28_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit11_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit20_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix__044_ Inst_LUT4AB_switch_matrix__044_/A vssd1 vssd1 vccd1
+ vccd1 output265/A sky130_fd_sc_hd__buf_1
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_44_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_switch_matrix__055_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_10 input62/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit7_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_21 ANTENNA_21/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LE_SR__0__512 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LE_SR__0__512/HI
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LE_SR__0_/A0 sky130_fd_sc_hd__conb_1
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0_A3
+ input41/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit16_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit8_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG2_A1 input19/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit5 input77/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LG_EN__0__522 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LG_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LG_EN__0__522/LO sky130_fd_sc_hd__conb_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A2 Inst_LUT4AB_ConfigMem_Inst_Frame4_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit21/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0_A1
+ input129/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit29/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG0_A3 Inst_LUT4AB_switch_matrix__067_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput30 E6END[6] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
Xinput63 FrameData[21] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__buf_8
Xinput52 FrameData[11] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__buf_8
XFILLER_0_12_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput41 EE4END[1] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__clkbuf_2
Xinput74 FrameData[31] vssd1 vssd1 vccd1 vccd1 input74/X sky130_fd_sc_hd__buf_8
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG2_A1 input170/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput96 FrameStrobe[4] vssd1 vssd1 vccd1 vccd1 input96/X sky130_fd_sc_hd__buf_12
Xinput85 FrameStrobe[12] vssd1 vssd1 vccd1 vccd1 input85/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG2_A0 Inst_LUT4AB_switch_matrix__055_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LD_LUT4c_frame_config_dffesr__11_ Inst_LD_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__060_/X
+ Inst_LD_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__11_/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit3 input75/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A2
+ ANTENNA_5/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame12_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__10_/A sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit20 input62/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG2_A3 input215/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0 input105/X
+ input107/X input129/X input41/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG2_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG3_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LB_EN__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit11_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit8 input80/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit20_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_outbuf_1__0_ data_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output314/A sky130_fd_sc_hd__clkbuf_1
Xinput220 W2MID[2] vssd1 vssd1 vccd1 vccd1 input220/X sky130_fd_sc_hd__clkbuf_4
Xinput253 WW4END[9] vssd1 vssd1 vccd1 vccd1 input253/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit0_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput242 WW4END[13] vssd1 vssd1 vccd1 vccd1 input242/X sky130_fd_sc_hd__clkbuf_1
Xinput231 W6END[3] vssd1 vssd1 vccd1 vccd1 input231/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG2 input145/X input11/X input163/X
+ input215/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A2 sky130_fd_sc_hd__mux4_2
XFILLER_0_26_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit16_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit25_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xdata_inbuf_25__0_ input67/X vssd1 vssd1 vccd1 vccd1 data_inbuf_25__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit30 input73/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst0 input102/X
+ input2/X input206/X Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame10_bit27/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit27/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst0_A3
+ input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG1 input116/X input16/X
+ input220/X Inst_LUT4AB_switch_matrix__042_/A Inst_LUT4AB_ConfigMem_Inst_Frame14_bit13/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit6/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_strobe_inbuf_13__0__A input86/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit6 input78/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_inbuf_4__0_ input96/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_16__0_ input57/X vssd1 vssd1 vccd1 vccd1 data_inbuf_16__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_data_inbuf_4__0__A input76/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit8/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit18/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__043_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG3 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1 Inst_LUT4AB_switch_matrix__067_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit23/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit21/Q vssd1 vssd1 vccd1 vccd1 output258/A sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit13_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit22_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG3 input122/X input22/X input174/X
+ ANTENNA_2/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame11_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit30/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A3 sky130_fd_sc_hd__mux4_1
XANTENNA_SS4BEG_outbuf_11__0__A SS4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput502 output502/A vssd1 vssd1 vccd1 vccd1 WW4BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_0_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit31_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__102__A Inst_LUT4AB_switch_matrix__102_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LF_LUT4c_frame_config_dffesr__14_ hold7/X Inst_LF_LUT4c_frame_config_dffesr__13_/X
+ Inst_LF_LUT4c_frame_config_dffesr__14_/S vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__mux2_1
XFILLER_0_9_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG2 input119/X input19/X
+ input171/X input223/X Inst_LUT4AB_ConfigMem_Inst_Frame13_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A1 sky130_fd_sc_hd__mux4_1
XFILLER_0_37_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit3_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit4_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit18_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit27_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit3 input75/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0 input103/X
+ input109/X input43/X input25/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0_A2
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__060_ Inst_LUT4AB_switch_matrix__060_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__060_/X sky130_fd_sc_hd__buf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG0 input112/X input12/X input199/X
+ input216/X Inst_LUT4AB_ConfigMem_Inst_Frame9_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A2 sky130_fd_sc_hd__mux4_2
Xinput6 E2END[0] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_0_36_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_19__0_ strobe_inbuf_19__0_/X vssd1 vssd1 vccd1 vccd1 output345/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG3_A3 ANTENNA_14/DIODE
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_strobe_inbuf_0__0__A input82/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput310 output310/A vssd1 vssd1 vccd1 vccd1 FrameData_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput343 output343/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput321 output321/A vssd1 vssd1 vccd1 vccd1 FrameData_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput332 output332/A vssd1 vssd1 vccd1 vccd1 FrameData_O[7] sky130_fd_sc_hd__clkbuf_4
Xoutput354 output354/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput376 output376/A vssd1 vssd1 vccd1 vccd1 N4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput387 output387/A vssd1 vssd1 vccd1 vccd1 N4BEG[6] sky130_fd_sc_hd__buf_2
Xoutput365 output365/A vssd1 vssd1 vccd1 vccd1 N2BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_0_77_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput398 output398/A vssd1 vssd1 vccd1 vccd1 NN4BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_N4BEG_outbuf_9__0__A N4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit1 input61/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst0_A3
+ input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LE_LUT4c_frame_config_dffesr__12_ Inst_LE_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__061_/X
+ Inst_LE_LUT4c_frame_config_dffesr__11_/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__062_/A
+ sky130_fd_sc_hd__a21o_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__112_ input225/X vssd1 vssd1 vccd1 vccd1 output479/A sky130_fd_sc_hd__buf_1
XFILLER_0_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__043_ Inst_LUT4AB_switch_matrix__043_/A vssd1 vssd1 vccd1
+ vccd1 output264/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0_A1
+ input109/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit11/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit10/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__104_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_11 input218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG1_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit7_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_EE4BEG_outbuf_4__0__A EE4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit8_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG2_A2 input171/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit6 input78/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0 input146/X
+ input2/X input42/X input22/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit13_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit22_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit31_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG0_A0 input147/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0_A2
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_1__0_ strobe_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output346/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit29/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit29/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput31 E6END[7] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
Xinput20 E2MID[6] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
Xinput64 FrameData[22] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_8
Xinput53 FrameData[12] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_8
XFILLER_0_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput42 EE4END[2] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__clkbuf_2
Xinput75 FrameData[3] vssd1 vssd1 vccd1 vccd1 input75/X sky130_fd_sc_hd__buf_8
Xinput86 FrameStrobe[13] vssd1 vssd1 vccd1 vccd1 input86/X sky130_fd_sc_hd__buf_12
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG2_A2 input222/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput97 FrameStrobe[5] vssd1 vssd1 vccd1 vccd1 input97/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit18_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__110__A input223/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG2_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LD_LUT4c_frame_config_dffesr__10_ Inst_LD_LUT4c_frame_config_dffesr__10_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__10_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit4 input76/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit10 input51/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit21 input63/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit10_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0_A1 ANTENNA_21/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_16__0_ input89/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_16__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 output292/A sky130_fd_sc_hd__mux2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit13/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit17/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__087_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_56_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1 input25/X
+ input159/X input211/X input229/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix__105__A input218/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG2_A2 Inst_LUT4AB_switch_matrix__082_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit24_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3_A3 ANTENNA_5/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LH_LUT4c_frame_config_dffesr__09__A Inst_LH_LUT4c_frame_config_dffesr__09_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit9 input81/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LF_EN__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_MUX8LUT_frame_config_mux_cus_mux21_EH__0__A0 Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput210 W2END[0] vssd1 vssd1 vccd1 vccd1 input210/X sky130_fd_sc_hd__clkbuf_2
XE6BEG_outbuf_2__0_ E6END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output279/A sky130_fd_sc_hd__clkbuf_1
Xinput221 W2MID[3] vssd1 vssd1 vccd1 vccd1 input221/X sky130_fd_sc_hd__buf_2
Xinput243 WW4END[14] vssd1 vssd1 vccd1 vccd1 input243/X sky130_fd_sc_hd__clkbuf_1
Xinput232 W6END[4] vssd1 vssd1 vccd1 vccd1 input232/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit29_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LG_LUT4c_frame_config_dffesr__15_ UserCLK hold14/X vssd1 vssd1 vccd1 vccd1 hold13/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG1_A0 input130/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG3 input107/X input43/X input159/X
+ input211/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit4/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A2 sky130_fd_sc_hd__mux4_2
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XN4END_inbuf_1__0_ input133/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_1__0_/X sky130_fd_sc_hd__buf_2
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit20 input62/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LE_LUT4c_frame_config_dffesr__13_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame18_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG0_A0 input121/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit31 input74/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A2 Inst_LUT4AB_ConfigMem_Inst_Frame10_bit27/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit27/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG2 input118/X input18/X
+ input170/X Inst_LUT4AB_switch_matrix__085_/A Inst_LUT4AB_ConfigMem_Inst_Frame2_bit4/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit4/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit7 input79/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I0_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_S4BEG_outbuf_11__0__A S4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_8__0_ input80/X vssd1 vssd1 vccd1 vccd1 data_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput503 output503/A vssd1 vssd1 vccd1 vccd1 WW4BEG[5] sky130_fd_sc_hd__buf_2
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit10_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LF_LUT4c_frame_config_dffesr__13_ Inst_LF_LUT4c_frame_config_dffesr__13_/A0
+ Inst_LF_LUT4c_frame_config_dffesr__13_/A1 Inst_LF_LUT4c_frame_config_dffesr__13_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__13_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG3 input115/X input15/X
+ input167/X input219/X Inst_LUT4AB_ConfigMem_Inst_Frame12_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A1 sky130_fd_sc_hd__mux4_1
XFILLER_0_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit3_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit4 input76/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit4_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1 input183/X
+ input199/X input213/X input229/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0_A3
+ input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit15_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit24_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG3_A0 input122/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit30 input73/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG1 input138/X input8/X input160/X
+ input212/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit2/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A2 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput7 E2END[1] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_strobe_inbuf_12__0__A input85/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput300 output300/A vssd1 vssd1 vccd1 vccd1 EE4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput344 output344/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput322 output322/A vssd1 vssd1 vccd1 vccd1 FrameData_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput311 output311/A vssd1 vssd1 vccd1 vccd1 FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput333 output333/A vssd1 vssd1 vccd1 vccd1 FrameData_O[8] sky130_fd_sc_hd__buf_2
Xoutput355 output355/A vssd1 vssd1 vccd1 vccd1 N1BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_77_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput377 output377/A vssd1 vssd1 vccd1 vccd1 N4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput366 output366/A vssd1 vssd1 vccd1 vccd1 N2BEG[7] sky130_fd_sc_hd__clkbuf_4
XANTENNA_data_inbuf_3__0__A input75/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput399 output399/A vssd1 vssd1 vccd1 vccd1 NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput388 output388/A vssd1 vssd1 vccd1 vccd1 N4BEG[7] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit29_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame6_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 output397/A sky130_fd_sc_hd__mux2_1
XFILLER_0_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit2 input72/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0 input103/X
+ input111/X input3/X input11/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit12_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_SS4BEG_outbuf_10__0__A SS4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LE_LUT4c_frame_config_dffesr__11_ Inst_LE_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__061_/X
+ Inst_LE_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__11_/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit21_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit30_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_cus_mux41_buf_inst0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A1 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit29/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit31/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix__111_ input224/X vssd1 vssd1 vccd1 vccd1 output478/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__042_ Inst_LUT4AB_switch_matrix__042_/A vssd1 vssd1 vccd1
+ vccd1 output263/A sky130_fd_sc_hd__clkbuf_1
XInst_LE_LUT4c_frame_config_dffesr_cus_mux21_I0mux__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I0/X
+ Inst_LUT4AB_switch_matrix__061_/X Inst_LUT4AB_ConfigMem_Inst_Frame16_bit25/Q vssd1
+ vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__07_/A sky130_fd_sc_hd__mux2_2
XFILLER_0_47_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0_A2
+ input43/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XNN4BEG_outbuf_2__0_ NN4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output399/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XN4BEG_outbuf_6__0_ N4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output387/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix__108__A input221/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_12 output473/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0_A0
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit17_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit7_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit26_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XSS4BEG_outbuf_5__0_ SS4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output454/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit2_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG2_A3 input223/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit7 input79/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit8_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1 input182/X
+ input198/X input212/X input226/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG0_A1 input183/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0_A3
+ input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 Inst_LUT4AB_ConfigMem_Inst_Frame5_bit29/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit29/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput21 E2MID[7] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__buf_2
Xinput10 E2END[4] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__clkbuf_2
Xinput54 FrameData[13] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__buf_8
Xinput32 E6END[8] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput43 EE4END[3] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__clkbuf_2
Xinput65 FrameData[23] vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_16
Xinput76 FrameData[4] vssd1 vssd1 vccd1 vccd1 input76/X sky130_fd_sc_hd__buf_8
Xinput98 FrameStrobe[6] vssd1 vssd1 vccd1 vccd1 input98/X sky130_fd_sc_hd__clkbuf_16
Xinput87 FrameStrobe[14] vssd1 vssd1 vccd1 vccd1 input87/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG2_A3 Inst_LUT4AB_switch_matrix__087_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_N4BEG_outbuf_8__0__A N4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG3_A0 input115/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XW6BEG_outbuf_6__0_ W6END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output488/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG2_A2 Inst_LUT4AB_switch_matrix__039_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG2_A0 input118/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit5 input77/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1_A0
+ input154/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0_A1
+ input107/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit11 input52/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit22 input64/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LD_SR__0__511 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LD_SR__0__511/HI
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LD_SR__0_/A0 sky130_fd_sc_hd__conb_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_EE4BEG_outbuf_3__0__A EE4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_E6BEG_outbuf_9__0__A E6END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__033_/A
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG2_A3 ANTENNA_5/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit12_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit21_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit6_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LF_EN__0__521 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LF_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LF_EN__0__521/LO sky130_fd_sc_hd__conb_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit30_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xdata_outbuf_26__0_ data_inbuf_26__0_/X vssd1 vssd1 vccd1 vccd1 output321/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit7_GATE input93/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput200 SS4END[4] vssd1 vssd1 vccd1 vccd1 input200/X sky130_fd_sc_hd__clkbuf_1
Xinput211 W2END[1] vssd1 vssd1 vccd1 vccd1 input211/X sky130_fd_sc_hd__buf_2
Xinput222 W2MID[4] vssd1 vssd1 vccd1 vccd1 input222/X sky130_fd_sc_hd__buf_2
Xinput244 WW4END[15] vssd1 vssd1 vccd1 vccd1 input244/X sky130_fd_sc_hd__clkbuf_1
Xinput233 W6END[5] vssd1 vssd1 vccd1 vccd1 input233/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LG_LUT4c_frame_config_dffesr__14_ hold13/X Inst_LG_LUT4c_frame_config_dffesr__13_/X
+ Inst_LG_LUT4c_frame_config_dffesr__14_/S vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__mux2_1
XFILLER_0_73_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG1_A1 input198/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_17__0_ data_inbuf_17__0_/X vssd1 vssd1 vccd1 vccd1 output311/A sky130_fd_sc_hd__clkbuf_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LC_SR__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LC_SR__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit30/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__13_/S sky130_fd_sc_hd__mux2_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit26_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XS4BEG_outbuf_6__0_ S4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output439/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit10 input51/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG0_A1 input21/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit21 input63/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG3 input114/X input166/X
+ input218/X Inst_LUT4AB_switch_matrix__101_/A Inst_LUT4AB_ConfigMem_Inst_Frame9_bit4/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit2/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_4_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit8 input80/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I0_A1 ANTENNA_21/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit0 input50/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XS4END_inbuf_4__0_ input188/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_4__0_/X sky130_fd_sc_hd__buf_2
XFILLER_0_58_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit14_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit23_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I3_A3 ANTENNA_5/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput504 output504/A vssd1 vssd1 vccd1 vccd1 WW4BEG[6] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LF_LUT4c_frame_config_dffesr__12_ Inst_LF_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__062_/X
+ Inst_LF_LUT4c_frame_config_dffesr__11_/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__063_/A
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XW6END_inbuf_8__0_ input227/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit19_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XEE4BEG_outbuf_5__0_ EE4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output298/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit5 input77/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG3_A1 input22/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit31 input74/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit20 input62/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG2 input110/X input34/X input162/X
+ input214/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit6/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A2 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 E2END[2] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_0_36_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_S4BEG_outbuf_10__0__A S4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput301 output301/A vssd1 vssd1 vccd1 vccd1 EE4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput323 output323/A vssd1 vssd1 vccd1 vccd1 FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput312 output312/A vssd1 vssd1 vccd1 vccd1 FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput334 output334/A vssd1 vssd1 vccd1 vccd1 FrameData_O[9] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput345 output345/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput378 output378/A vssd1 vssd1 vccd1 vccd1 N4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput367 output367/A vssd1 vssd1 vccd1 vccd1 N2BEGb[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput356 output356/A vssd1 vssd1 vccd1 vccd1 N1BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput389 output389/A vssd1 vssd1 vccd1 vccd1 N4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit3 input75/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_33_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1 input155/X
+ input163/X input207/X input209/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LE_LUT4c_frame_config_dffesr__10_ Inst_LE_LUT4c_frame_config_dffesr__10_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__10_/Y sky130_fd_sc_hd__inv_2
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__067_/A
+ Inst_LUT4AB_switch_matrix__040_/A Inst_LUT4AB_switch_matrix__083_/A ANTENNA_14/DIODE
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix__110_ input223/X vssd1 vssd1 vccd1 vccd1 output477/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_51_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix__041_ Inst_LUT4AB_switch_matrix__041_/A vssd1 vssd1 vccd1
+ vccd1 output262/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0_A3
+ input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_13 ANTENNA_13/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0_A1
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0 input105/X
+ input113/X input5/X input13/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit14_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit8 input80/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit30 input73/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit2_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix__034__A Inst_LUT4AB_switch_matrix__034_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit23_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_strobe_inbuf_11__0__A input84/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit3_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG0_A2 input238/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_data_inbuf_2__0__A input72/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit27/Q vssd1 vssd1 vccd1 vccd1 output276/A sky130_fd_sc_hd__mux4_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput11 E2END[5] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__buf_2
Xinput22 E6END[0] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__buf_4
Xinput55 FrameData[14] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_8
Xinput33 E6END[9] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput44 EE4END[4] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__clkbuf_1
Xinput66 FrameData[24] vssd1 vssd1 vccd1 vccd1 input66/X sky130_fd_sc_hd__clkbuf_16
Xinput77 FrameData[5] vssd1 vssd1 vccd1 vccd1 input77/X sky130_fd_sc_hd__clkbuf_16
Xinput88 FrameStrobe[15] vssd1 vssd1 vccd1 vccd1 input88/X sky130_fd_sc_hd__buf_8
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput99 FrameStrobe[7] vssd1 vssd1 vccd1 vccd1 input99/X sky130_fd_sc_hd__clkbuf_16
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit19_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit28_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG3_A1 input15/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr__15_ UserCLK hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG2_A3 ANTENNA_5/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG2_A1 input170/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG2_A2 input198/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit6 input78/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1_A1
+ input158/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0_A2
+ input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit12 input53/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit23 input65/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XSS4END_inbuf_11__0_ input196/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_11__0_/X sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit20_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit11_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xdata_outbuf_4__0_ data_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output329/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit16_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit25_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_28__0_ input70/X vssd1 vssd1 vccd1 vccd1 data_inbuf_28__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit6_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XWW4END_inbuf_0__0_ input248/X vssd1 vssd1 vccd1 vccd1 ANTENNA_20/DIODE sky130_fd_sc_hd__clkbuf_2
XFILLER_0_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput201 SS4END[5] vssd1 vssd1 vccd1 vccd1 input201/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit7_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_7__0_ input99/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_19__0_ input60/X vssd1 vssd1 vccd1 vccd1 data_inbuf_19__0_/X sky130_fd_sc_hd__clkbuf_1
Xinput223 W2MID[5] vssd1 vssd1 vccd1 vccd1 input223/X sky130_fd_sc_hd__clkbuf_2
Xinput212 W2END[2] vssd1 vssd1 vccd1 vccd1 input212/X sky130_fd_sc_hd__buf_2
Xinput245 WW4END[1] vssd1 vssd1 vccd1 vccd1 input245/X sky130_fd_sc_hd__clkbuf_2
Xinput234 W6END[6] vssd1 vssd1 vccd1 vccd1 input234/X sky130_fd_sc_hd__clkbuf_1
XInst_LG_LUT4c_frame_config_dffesr__13_ Inst_LG_LUT4c_frame_config_dffesr__13_/A0
+ Inst_LG_LUT4c_frame_config_dffesr__13_/A1 Inst_LG_LUT4c_frame_config_dffesr__13_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__13_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1_A0
+ input156/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG1_A2 input212/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_N4BEG_outbuf_7__0__A N4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit11 input52/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG0_A2 input173/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit22 input64/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit0 input50/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame0_bit9 input81/X input82/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit1 input61/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix__042__A Inst_LUT4AB_switch_matrix__042_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_E6BEG_outbuf_8__0__A E6END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_EE4BEG_outbuf_2__0__A EE4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput505 output505/A vssd1 vssd1 vccd1 vccd1 WW4BEG[7] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit11_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit26/Q
+ vssd1 vssd1 vccd1 vccd1 output448/A sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit20_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LF_LUT4c_frame_config_dffesr__11_ Inst_LF_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__062_/X
+ Inst_LF_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__11_/X
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_1_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit6 input78/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix__037__A Inst_LUT4AB_switch_matrix__037_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XE6END_inbuf_0__0_ input26/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_0__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit16_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit25_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG3_A2 input174/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit10 input51/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit21 input63/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG3 input106/X input6/X input158/X
+ input247/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit5/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A2 sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0 input102/X
+ input106/X input2/X input6/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput9 E2END[3] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_2
XFILLER_0_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput335 output335/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput324 output324/A vssd1 vssd1 vccd1 vccd1 FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput313 output313/A vssd1 vssd1 vccd1 vccd1 FrameData_O[19] sky130_fd_sc_hd__buf_2
Xoutput302 output302/A vssd1 vssd1 vccd1 vccd1 EE4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput346 output346/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
Xoutput357 output357/A vssd1 vssd1 vccd1 vccd1 N1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput368 output368/A vssd1 vssd1 vccd1 vccd1 N2BEGb[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput379 output379/A vssd1 vssd1 vccd1 vccd1 N4BEG[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit4 input76/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XSS4END_inbuf_2__0_ input202/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_2
XEE4END_inbuf_11__0_ input40/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_11__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit13_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit22_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__040_ Inst_LUT4AB_switch_matrix__040_/A vssd1 vssd1 vccd1
+ vccd1 output261/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_4__0_ strobe_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output349/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_14 ANTENNA_14/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit27_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0_A2
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1 input155/X
+ input157/X input165/X input209/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit9 input81/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit31 input74/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit20 input62/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XEE4END_inbuf_1__0_ input45/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_1__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__050__A input18/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG0_A3 Inst_LUT4AB_switch_matrix__066_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XWW4BEG_outbuf_2__0_ WW4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output500/A sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_19__0_ input92/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_19__0_/X sky130_fd_sc_hd__clkbuf_1
Xinput12 E2END[6] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__buf_2
Xinput23 E6END[10] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 EE4END[0] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__clkbuf_2
Xinput45 EE4END[5] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__clkbuf_1
Xinput67 FrameData[25] vssd1 vssd1 vccd1 vccd1 input67/X sky130_fd_sc_hd__buf_8
Xinput56 FrameData[15] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_8
Xinput78 FrameData[6] vssd1 vssd1 vccd1 vccd1 input78/X sky130_fd_sc_hd__buf_8
Xinput89 FrameStrobe[16] vssd1 vssd1 vccd1 vccd1 input89/X sky130_fd_sc_hd__buf_8
XFILLER_0_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG3_A2 input167/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr__14_ hold3/X Inst_LH_LUT4c_frame_config_dffesr__13_/X
+ Inst_LH_LUT4c_frame_config_dffesr__14_/S vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__mux2_1
XFILLER_0_74_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG2_A2 input222/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG2_A3 input214/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1_A2
+ input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit7 input79/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst0_A3
+ input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit24 input66/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit13 input54/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__045__A Inst_LUT4AB_switch_matrix__045_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4_S0
+ Inst_LG_LUT4c_frame_config_dffesr__09_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XE6BEG_outbuf_5__0_ E6END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output282/A sky130_fd_sc_hd__clkbuf_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux_cus_mux21_sEH__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_AH__0_/S
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AD__0_/S Inst_LUT4AB_ConfigMem_Inst_Frame3_bit29/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_EH__0_/S sky130_fd_sc_hd__mux2_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit10/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit9/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__038_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XN4END_inbuf_4__0_ input136/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit30 input73/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit13_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit22_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit31_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_strobe_inbuf_10__0__A input83/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit6_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput202 SS4END[6] vssd1 vssd1 vccd1 vccd1 input202/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_data_inbuf_1__0__A input61/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput224 W2MID[6] vssd1 vssd1 vccd1 vccd1 input224/X sky130_fd_sc_hd__clkbuf_4
Xinput213 W2END[3] vssd1 vssd1 vccd1 vccd1 input213/X sky130_fd_sc_hd__buf_2
Xinput235 W6END[7] vssd1 vssd1 vccd1 vccd1 input235/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit1_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xinput246 WW4END[2] vssd1 vssd1 vccd1 vccd1 input246/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit7_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LG_LUT4c_frame_config_dffesr__12_ Inst_LG_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__063_/X
+ Inst_LG_LUT4c_frame_config_dffesr__11_/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__064_/A
+ sky130_fd_sc_hd__a21o_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1_A1
+ input164/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG1_A3 Inst_LUT4AB_switch_matrix__042_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit18_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit2_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output270_A output270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit12 input53/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit23 input65/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG0_A3 input225/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit1 input61/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit10_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst0 input105/X
+ input5/X input157/X Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_ConfigMem_Inst_Frame8_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit17/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG0_A0 input121/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit2 input72/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LC_SR__0__510 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LC_SR__0__510/HI
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LC_SR__0_/A0 sky130_fd_sc_hd__conb_1
XFILLER_0_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit15_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit24_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput506 output506/A vssd1 vssd1 vccd1 vccd1 WW4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LE_EN__0__520 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LE_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LE_EN__0__520/LO sky130_fd_sc_hd__conb_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1_A0
+ input162/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LF_LUT4c_frame_config_dffesr__10_ Inst_LF_LUT4c_frame_config_dffesr__10_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__10_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit29_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_N4BEG_outbuf_6__0__A N4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit5_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit7 input79/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame9_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit12/Q vssd1 vssd1 vccd1 vccd1 ANTENNA_14/DIODE
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XInst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_ Inst_LUT4AB_switch_matrix__037_/X
+ Inst_LUT4AB_switch_matrix__054_/X Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_23_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit6_GATE input94/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I3_A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A0
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__053__A input21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG3_A3 ANTENNA_2/DIODE
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit11 input52/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit22 input64/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1 input154/X
+ input158/X input206/X input208/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG0_A0 input113/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput325 output325/A vssd1 vssd1 vccd1 vccd1 FrameData_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput314 output314/A vssd1 vssd1 vccd1 vccd1 FrameData_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput303 output303/A vssd1 vssd1 vccd1 vccd1 FrameData_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput347 output347/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput369 output369/A vssd1 vssd1 vccd1 vccd1 N2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput336 output336/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput358 output358/A vssd1 vssd1 vccd1 vccd1 N1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XNN4BEG_outbuf_5__0_ NN4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output402/A sky130_fd_sc_hd__clkbuf_1
XN4BEG_outbuf_9__0_ N4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output390/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit5 input77/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_EE4BEG_outbuf_1__0__A EE4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_E6BEG_outbuf_7__0__A E6END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit10/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XSS4BEG_outbuf_8__0_ SS4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output457/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix__048__A input16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit10_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_15 ANTENNA_4/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__099_ ANTENNA_14/DIODE vssd1 vssd1 vccd1 vccd1 output466/A
+ sky130_fd_sc_hd__clkbuf_1
XW6BEG_outbuf_9__0_ W6END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output491/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit15_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit24_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit9_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit10 input51/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG0_A0 input108/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit11/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit14/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__082_/A
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit21 input63/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LB_SR__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput13 E2END[7] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_2
Xinput24 E6END[11] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput46 EE4END[6] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__clkbuf_1
Xinput35 EE4END[10] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_1
Xinput68 FrameData[26] vssd1 vssd1 vccd1 vccd1 input68/X sky130_fd_sc_hd__buf_8
Xinput79 FrameData[7] vssd1 vssd1 vccd1 vccd1 input79/X sky130_fd_sc_hd__buf_8
Xinput57 FrameData[16] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__buf_8
XFILLER_0_3_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XNN4END_inbuf_2__0_ input150/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit29_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG3_A3 input219/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr__13_ Inst_LH_LUT4c_frame_config_dffesr__13_/A0
+ Inst_LH_LUT4c_frame_config_dffesr__13_/A1 Inst_LH_LUT4c_frame_config_dffesr__13_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__13_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_59_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG2_A3 Inst_LUT4AB_switch_matrix__086_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit12_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1_A3
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit8 input80/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG3_A0 input115/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit14 input55/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit25 input67/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit21_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit30_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG2_A0 input118/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_38_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xdata_outbuf_29__0_ data_inbuf_29__0_/X vssd1 vssd1 vccd1 vccd1 output324/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4_S1
+ Inst_LG_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_N4BEG_outbuf_11__0__A N4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit17_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit26_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit31 input74/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XS4BEG_outbuf_9__0_ S4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 output442/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit20 input62/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG1_A0 input146/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput203 SS4END[7] vssd1 vssd1 vccd1 vccd1 input203/X sky130_fd_sc_hd__clkbuf_1
Xinput225 W2MID[7] vssd1 vssd1 vccd1 vccd1 input225/X sky130_fd_sc_hd__clkbuf_2
Xinput214 W2END[4] vssd1 vssd1 vccd1 vccd1 input214/X sky130_fd_sc_hd__clkbuf_4
Xinput236 W6END[8] vssd1 vssd1 vccd1 vccd1 input236/X sky130_fd_sc_hd__clkbuf_1
Xinput247 WW4END[3] vssd1 vssd1 vccd1 vccd1 input247/X sky130_fd_sc_hd__dlymetal6s2s_1
XInst_LG_LUT4c_frame_config_dffesr__11_ Inst_LG_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__063_/X
+ Inst_LG_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__11_/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit1_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__056__A Inst_LUT4AB_switch_matrix__056_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1_A2
+ input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LF_EN__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LF_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit4/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__14_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XS4END_inbuf_7__0_ input176/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit2_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit13 input54/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit24 input66/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG3_A0 input107/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit2 input72/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG1_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__056_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A2 Inst_LUT4AB_ConfigMem_Inst_Frame8_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit17/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG0_A1 input21/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst0 input103/X
+ input3/X input207/X Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_ConfigMem_Inst_Frame4_bit27/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit23/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit3 input75/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1_A0
+ input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XEE4BEG_outbuf_8__0_ EE4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output301/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0 input4/X
+ input208/X Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame6_bit23/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit30 input73/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG0 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1 ANTENNA_3/DIODE Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 output355/A sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit12_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xoutput507 output507/A vssd1 vssd1 vccd1 vccd1 WW4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_0_34_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit21_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1_A1
+ input174/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2_A2
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst3_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_0__0__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit17_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG3_A0 input107/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit8 input80/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit5_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit26_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I3_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit0_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit12 input53/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit6_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit23 input65/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit1_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG0_A1 input13/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput326 output326/A vssd1 vssd1 vccd1 vccd1 FrameData_O[30] sky130_fd_sc_hd__buf_2
Xoutput315 output315/A vssd1 vssd1 vccd1 vccd1 FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput304 output304/A vssd1 vssd1 vccd1 vccd1 FrameData_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput359 output359/A vssd1 vssd1 vccd1 vccd1 N2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput348 output348/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
Xoutput337 output337/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit6 input78/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit13/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit12/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__069_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_60_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1_A0
+ input182/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit14_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit23_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_CD__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AD__0_/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit24/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X sky130_fd_sc_hd__mux2_4
XFILLER_0_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit19_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit28_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_16 input118/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_N4BEG_outbuf_5__0__A N4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix__098_ ANTENNA_2/DIODE vssd1 vssd1 vccd1 vccd1 output465/A
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XNN4END_inbuf_11__0_ input144/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_11__0_/X sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit9_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG0_A1 input129/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit11 input52/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LA_LUT4c_frame_config_dffesr__13_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit22 input64/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LF_SR__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_outbuf_12__0_ strobe_inbuf_12__0_/X vssd1 vssd1 vccd1 vccd1 output338/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput14 E2MID[0] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_4
Xinput36 EE4END[11] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_1
Xinput25 E6END[1] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_4
Xinput69 FrameData[27] vssd1 vssd1 vccd1 vccd1 input69/X sky130_fd_sc_hd__buf_8
Xinput58 FrameData[17] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__buf_8
Xdata_outbuf_7__0_ data_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output332/A sky130_fd_sc_hd__clkbuf_1
Xinput47 EE4END[7] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr__12_ Inst_LH_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__064_/X
+ Inst_LH_LUT4c_frame_config_dffesr__11_/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__035_/A
+ sky130_fd_sc_hd__a21o_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG2_A1 input34/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_EE4BEG_outbuf_0__0__A EE4END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_E6BEG_outbuf_6__0__A E6END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit0 input50/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit9 input81/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG3_A1 input15/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit15 input56/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG2_A1 input18/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XWW4END_inbuf_3__0_ input251/X vssd1 vssd1 vccd1 vccd1 WW4END_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit14_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit21 input63/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit10 input51/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit23_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG1_A1 input8/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput204 SS4END[8] vssd1 vssd1 vccd1 vccd1 input204/X sky130_fd_sc_hd__clkbuf_1
Xinput215 W2END[5] vssd1 vssd1 vccd1 vccd1 input215/X sky130_fd_sc_hd__clkbuf_2
Xinput226 W6END[0] vssd1 vssd1 vccd1 vccd1 input226/X sky130_fd_sc_hd__clkbuf_4
Xinput248 WW4END[4] vssd1 vssd1 vccd1 vccd1 input248/X sky130_fd_sc_hd__clkbuf_1
Xinput237 W6END[9] vssd1 vssd1 vccd1 vccd1 input237/X sky130_fd_sc_hd__clkbuf_1
XInst_LG_LUT4c_frame_config_dffesr__10_ Inst_LG_LUT4c_frame_config_dffesr__10_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__10_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst1_A3
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit19_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit28_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix__072__A Inst_LUT4AB_switch_matrix__072_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit14 input55/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit25 input67/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG3_A1 input43/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit20_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit11_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit3 input75/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG0_A2 input173/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_N4BEG_outbuf_10__0__A N4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A2 Inst_LUT4AB_ConfigMem_Inst_Frame4_bit27/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit23/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit4 input76/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1_A1
+ input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit16_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit20/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit25_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LA_LUT4c_frame_config_dffesr__09_ Inst_LA_LUT4c_frame_config_dffesr__09_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__09_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix__067__A Inst_LUT4AB_switch_matrix__067_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XE6END_inbuf_3__0_ input29/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_39_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit20 input62/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit31 input74/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG1 Inst_LUT4AB_switch_matrix__036_/A
+ ANTENNA_21/DIODE Inst_LUT4AB_switch_matrix__097_/A Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 output356/A sky130_fd_sc_hd__mux4_2
XFILLER_0_26_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1_A2
+ input214/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG3_A1 input122/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit9 input81/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_NN4BEG_outbuf_9__0__A NN4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XSS4END_inbuf_5__0_ input205/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I3_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit13 input54/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit0_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit24 input66/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_switch_matrix__055_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0 input102/X
+ input108/X input130/X input8/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1_A0
+ input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit1_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG0_A2 input165/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput316 output316/A vssd1 vssd1 vccd1 vccd1 FrameData_O[21] sky130_fd_sc_hd__buf_2
Xoutput305 output305/A vssd1 vssd1 vccd1 vccd1 FrameData_O[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput349 output349/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput338 output338/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput327 output327/A vssd1 vssd1 vccd1 vccd1 FrameData_O[31] sky130_fd_sc_hd__buf_2
XFILLER_0_10_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_7__0_ strobe_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output352/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit7 input79/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_33_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1_A1
+ input198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit30 input73/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit11_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XEE4END_inbuf_4__0_ input48/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_2
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__080__A input121/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_inbuf_1__0_ input61/X vssd1 vssd1 vccd1 vccd1 data_inbuf_1__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst0 input103/X
+ input3/X input207/X Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_ConfigMem_Inst_Frame8_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit25/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_2_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XWW4BEG_outbuf_5__0_ WW4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output503/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_17 input198/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__097_ Inst_LUT4AB_switch_matrix__097_/A vssd1 vssd1 vccd1
+ vccd1 output464/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit16_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit25_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit11/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit18/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__044_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG0_A2 input25/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit12 input53/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit23 input65/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit9_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit4_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__075__A input116/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit30 input73/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit5_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_49_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput15 E2MID[1] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_4
Xinput37 EE4END[12] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_1
Xinput26 E6END[2] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__clkbuf_1
Xinput59 FrameData[18] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_8
XFILLER_0_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput48 EE4END[8] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
XE6BEG_outbuf_8__0_ E6END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output285/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr__11_ Inst_LH_LUT4c_frame_config_dffesr__09_/A Inst_LUT4AB_switch_matrix__064_/X
+ Inst_LH_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__11_/X
+ sky130_fd_sc_hd__o21a_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG2_A2 input162/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit1 input61/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit13_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit22_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0 input104/X
+ input110/X input10/X input22/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG3_A2 input167/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XN4END_inbuf_7__0_ input124/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit16 input57/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_3_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG1_A0 input22/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG2_A2 input170/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit18_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_N4BEG_outbuf_4__0__A N4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit27_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit11 input52/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit22 input64/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG1_A2 input182/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput205 SS4END[9] vssd1 vssd1 vccd1 vccd1 input205/X sky130_fd_sc_hd__clkbuf_1
Xinput216 W2END[6] vssd1 vssd1 vccd1 vccd1 input216/X sky130_fd_sc_hd__clkbuf_2
Xinput227 W6END[10] vssd1 vssd1 vccd1 vccd1 input227/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_SR_BEG0_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame12_bit29/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 sky130_fd_sc_hd__mux2_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit8_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xinput238 WW4END[0] vssd1 vssd1 vccd1 vccd1 input238/X sky130_fd_sc_hd__clkbuf_2
Xinput249 WW4END[5] vssd1 vssd1 vccd1 vccd1 input249/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit9_GATE input94/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_E6BEG_outbuf_5__0__A E6END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit15 input56/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit26 input68/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG3_A2 input159/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit4 input76/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0 input147/X
+ input3/X input9/X input25/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG0_A3 input225/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LF_LUT4c_frame_config_dffesr_cus_mux21_I0mux__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/X
+ Inst_LUT4AB_switch_matrix__062_/X Inst_LUT4AB_ConfigMem_Inst_Frame15_bit22/Q vssd1
+ vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__07_/A sky130_fd_sc_hd__mux2_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit5 input77/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1_A2
+ input165/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG0_A0 input121/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LA_LUT4c_frame_config_dffesr__08_ Inst_LA_LUT4c_frame_config_dffesr__08_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__08_/Y sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit23/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit21 input63/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix__083__A Inst_LUT4AB_switch_matrix__083_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit10 input51/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG2 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 ANTENNA_2/DIODE ANTENNA_5/DIODE
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit13/Q
+ vssd1 vssd1 vccd1 vccd1 output357/A sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit22_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit13_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit31_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1_A0
+ input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1_A3
+ input246/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XNN4BEG_outbuf_8__0_ NN4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output405/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit18_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit27_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG3_A2 input226/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame10_bit30/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 sky130_fd_sc_hd__mux2_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit14 input55/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__067_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit25 input67/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit19/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit23/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__088_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit10_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1 input22/X
+ input160/X input212/X input247/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix__078__A input119/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_outbuf_10__0_ data_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 output304/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit0_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1_A1
+ input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit1_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG0_A3 input238/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput317 output317/A vssd1 vssd1 vccd1 vccd1 FrameData_O[22] sky130_fd_sc_hd__clkbuf_4
Xoutput306 output306/A vssd1 vssd1 vccd1 vccd1 FrameData_O[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput339 output339/A vssd1 vssd1 vccd1 vccd1 FrameStrobe_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput328 output328/A vssd1 vssd1 vccd1 vccd1 FrameData_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_10_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG2_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit15_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit8 input80/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1_A2
+ input212/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit24_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S2_A0 Inst_LUT4AB_switch_matrix__071_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0 Inst_LUT4AB_ConfigMem_Inst_Frame10_bit15/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit12/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit21/Q Inst_LH_LUT4c_frame_config_dffesr__07_/A
+ Inst_LH_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit20 input62/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit31 input74/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A2 Inst_LUT4AB_ConfigMem_Inst_Frame8_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit25/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit29_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LF_LUT4c_frame_config_dffesr__10__A Inst_LF_LUT4c_frame_config_dffesr__10_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 input224/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XNN4END_inbuf_5__0_ input153/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_5__0_/X sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix__096_ input173/X vssd1 vssd1 vccd1 vccd1 output426/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1_A0
+ input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XW6END_inbuf_1__0_ input231/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_1__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_NN4BEG_outbuf_8__0__A NN4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG0_A3 Inst_LUT4AB_switch_matrix__037_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit13 input54/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit24 input66/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit26/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit30/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit4_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit20 input62/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_68_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit31 input74/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput27 E6END[3] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix__091__A input168/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput16 E2MID[2] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__buf_2
XFILLER_0_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit5_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput49 EE4END[9] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__clkbuf_1
Xinput38 EE4END[13] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr__10_ Inst_LH_LUT4c_frame_config_dffesr__10_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__10_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG2_A3 input214/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XWW4END_inbuf_11__0_ input244/X vssd1 vssd1 vccd1 vccd1 WW4END_inbuf_11__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit2 input72/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit30 input73/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1 input162/X
+ input174/X input214/X input246/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG3_A3 input219/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit17 input58/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__079_ input120/X vssd1 vssd1 vccd1 vccd1 output373/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG1_A1 input161/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG2_A3 Inst_LUT4AB_switch_matrix__085_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG3_A0 input115/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG2_A0 input118/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit23/Q
+ vssd1 vssd1 vccd1 vccd1 output290/A sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_switch_matrix__086__A Inst_LUT4AB_switch_matrix__086_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit15_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit24_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LB_LUT4c_frame_config_dffesr__09_ Inst_LB_LUT4c_frame_config_dffesr__09_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__09_/Y sky130_fd_sc_hd__inv_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit12 input53/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit23 input65/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0 input104/X
+ input112/X input4/X input12/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit30 input73/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG1_A3 Inst_LUT4AB_switch_matrix__041_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput206 W1END[0] vssd1 vssd1 vccd1 vccd1 input206/X sky130_fd_sc_hd__buf_4
Xinput217 W2END[7] vssd1 vssd1 vccd1 vccd1 input217/X sky130_fd_sc_hd__clkbuf_2
Xinput239 WW4END[10] vssd1 vssd1 vccd1 vccd1 input239/X sky130_fd_sc_hd__clkbuf_1
Xinput228 W6END[11] vssd1 vssd1 vccd1 vccd1 input228/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit8_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit29_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit3_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit9_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit12_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit4_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit16 input57/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit27 input69/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG3_A3 input211/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit30_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG0 input108/X input129/X input25/X
+ Inst_LUT4AB_switch_matrix__037_/A Inst_LUT4AB_ConfigMem_Inst_Frame3_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit26/Q
+ vssd1 vssd1 vccd1 vccd1 output378/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit5 input77/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr_cus_mux21_O__0_ Inst_LH_LUT4c_frame_config_dffesr__13_/A0
+ hold3/A Inst_LUT4AB_ConfigMem_Inst_Frame13_bit19/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__056_/A
+ sky130_fd_sc_hd__mux2_8
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1 input161/X
+ input183/X input213/X input229/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit6 input78/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst1_A3
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit17_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG0_A1 input21/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_N4BEG_outbuf_3__0__A N4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit26_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LA_LUT4c_frame_config_dffesr__07_ Inst_LA_LUT4c_frame_config_dffesr__07_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__07_/Y sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0 Inst_LUT4AB_ConfigMem_Inst_Frame6_bit23/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_inbuf_30__0_ input73/X vssd1 vssd1 vccd1 vccd1 data_inbuf_30__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit22 input64/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit11 input52/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1 ANTENNA_14/DIODE Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 output358/A sky130_fd_sc_hd__mux4_2
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1_A1
+ input165/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xdata_inbuf_21__0_ input63/X vssd1 vssd1 vccd1 vccd1 data_inbuf_21__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG3_A3 Inst_LUT4AB_switch_matrix__056_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_E6BEG_outbuf_4__0__A E6END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_0__0_ input82/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_0__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_12__0_ input53/X vssd1 vssd1 vccd1 vccd1 data_inbuf_12__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit15 input56/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix__040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit26 input68/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A0
+ ANTENNA_21/DIODE Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A3
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I0/X sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1_A2
+ input163/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG0_A0 input113/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__094__A input171/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput307 output307/A vssd1 vssd1 vccd1 vccd1 FrameData_O[13] sky130_fd_sc_hd__buf_2
XFILLER_0_22_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput318 output318/A vssd1 vssd1 vccd1 vccd1 FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput329 output329/A vssd1 vssd1 vccd1 vccd1 FrameData_O[4] sky130_fd_sc_hd__buf_2
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit0 input50/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit9 input81/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG0 input9/X input199/X input246/X
+ Inst_LUT4AB_switch_matrix__067_/A Inst_LUT4AB_ConfigMem_Inst_Frame12_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit28/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A3 sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1_A0
+ input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame5_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 output395/A sky130_fd_sc_hd__mux2_1
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst1_A3
+ input226/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S2_A1 Inst_LUT4AB_switch_matrix__044_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1 Inst_LUT4AB_ConfigMem_Inst_Frame8_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit19/Q Inst_LH_LUT4c_frame_config_dffesr__07_/A
+ Inst_LH_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LD_SR__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LD_SR__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit0/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__13_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_67_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit10 input51/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit21 input63/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG1_A0 Inst_LUT4AB_switch_matrix__037_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_19__0__A input60/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit12_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit21_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__089__A input166/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG0 input121/X input21/X
+ input173/X input225/X Inst_LUT4AB_ConfigMem_Inst_Frame11_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A1 sky130_fd_sc_hd__mux4_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_15__0_ strobe_inbuf_15__0_/X vssd1 vssd1 vccd1 vccd1 output341/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_19 output479/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit17_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__095_ input172/X vssd1 vssd1 vccd1 vccd1 output425/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1_A1
+ input161/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit26_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit14 input55/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit25 input67/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_53_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG0_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit30/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit26/Q vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__08_/A
+ sky130_fd_sc_hd__mux4_2
XWW4END_inbuf_6__0_ input239/X vssd1 vssd1 vccd1 vccd1 WW4END_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit10 input51/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit21 input63/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LA_EN__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 E2MID[3] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__clkbuf_2
Xinput28 E6END[4] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
Xinput39 EE4END[14] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit0_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit14_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit23_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit3 input75/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit20 input62/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit31 input74/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_11_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit18 input59/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix__078_ input119/X vssd1 vssd1 vccd1 vccd1 output372/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG1_A2 input182/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG3_A1 input15/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_73_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1_A0
+ input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit19_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit28_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG2_A1 input18/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput490 output490/A vssd1 vssd1 vccd1 vccd1 W6BEG[8] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_NN4BEG_outbuf_7__0__A NN4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit1 input61/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LB_LUT4c_frame_config_dffesr__08_ Inst_LB_LUT4c_frame_config_dffesr__08_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__08_/Y sky130_fd_sc_hd__inv_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LA_EN__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LA_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame12_bit26/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__14_/S sky130_fd_sc_hd__mux2_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit13 input54/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit24 input66/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1 input156/X
+ input164/X input206/X input208/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG1_A0 input130/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit20 input62/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit31 input74/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput218 W2MID[0] vssd1 vssd1 vccd1 vccd1 input218/X sky130_fd_sc_hd__buf_2
Xinput207 W1END[1] vssd1 vssd1 vccd1 vccd1 input207/X sky130_fd_sc_hd__buf_4
Xinput229 W6END[1] vssd1 vssd1 vccd1 vccd1 input229/X sky130_fd_sc_hd__buf_4
XFILLER_0_75_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_66_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame12_bit2/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit1/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit3_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_12__0_ input85/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_12__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG3_A0 input146/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XE6END_inbuf_6__0_ input32/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit30 input73/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit17 input58/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit4_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit28 input70/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG2_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame19_bit22/Q
+ vssd1 vssd1 vccd1 vccd1 output497/A sky130_fd_sc_hd__mux2_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG1 input109/X input130/X input22/X
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_ConfigMem_Inst_Frame3_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit23/Q
+ vssd1 vssd1 vccd1 vccd1 output379/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit6 input78/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0 input102/X
+ input106/X input2/X input6/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit7 input79/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG0_A2 input173/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit19/Q vssd1 vssd1 vccd1 vccd1 output277/A sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0_A1
+ input113/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit14_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XSS4END_inbuf_8__0_ input193/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit23 input65/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit12 input53/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I0_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1_A2
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst0_A1
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit30 input73/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit19_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit28_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1_A0
+ input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit16 input57/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix__083_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit5/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit6/Q vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__08_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit7_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit27 input69/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LF_LUT4c_frame_config_dffesr__13_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit20_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst1_A3
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG0_A1 input42/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XEE4END_inbuf_7__0_ input36/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit8_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_27_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG0 input120/X input20/X
+ input224/X Inst_LUT4AB_switch_matrix__070_/A Inst_LUT4AB_ConfigMem_Inst_Frame4_bit5/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit4/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I0/A0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_54_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_4__0_ input76/X vssd1 vssd1 vccd1 vccd1 data_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput308 output308/A vssd1 vssd1 vccd1 vccd1 FrameData_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput319 output319/A vssd1 vssd1 vccd1 vccd1 FrameData_O[24] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XWW4BEG_outbuf_8__0_ ANTENNA_9/DIODE vssd1 vssd1 vccd1 vccd1 output506/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2_A2
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_N4BEG_outbuf_2__0__A N4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit1 input61/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit25_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit16_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG1 input130/X input8/X input217/X
+ Inst_LUT4AB_switch_matrix__040_/A Inst_LUT4AB_ConfigMem_Inst_Frame7_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit31/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3 sky130_fd_sc_hd__mux4_2
XFILLER_0_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1_A1
+ input163/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit17/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit21/Q Inst_LH_LUT4c_frame_config_dffesr__07_/A
+ Inst_LH_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S2_A2 Inst_LUT4AB_switch_matrix__087_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit11 input52/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit22 input64/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG1_A1 ANTENNA_21/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG1 input117/X input17/X
+ input169/X input221/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit3/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 sky130_fd_sc_hd__mux4_2
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_E6BEG_outbuf_3__0__A E6END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__094_ input171/X vssd1 vssd1 vccd1 vccd1 output424/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1_A2
+ input213/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit26 input68/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit15 input56/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LC_LUT4c_frame_config_dffesr__09_ Inst_LC_LUT4c_frame_config_dffesr__09_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__09_/Y sky130_fd_sc_hd__inv_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A3 Inst_LUT4AB_ConfigMem_Inst_Frame9_bit28/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit29/Q vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__09_/A
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit11 input52/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit22 input64/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1_A0
+ input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput18 E2MID[4] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput29 E6END[5] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LE_EN__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit4 input76/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit0_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XN4BEG_outbuf_2__0_ N4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output383/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit10 input51/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit21 input63/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_data_inbuf_18__0__A input59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame19_bit19 input60/X input92/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit11_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit20_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__077_ input118/X vssd1 vssd1 vccd1 vccd1 output371/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XSS4BEG_outbuf_1__0_ SS4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output450/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S4BEG1_A3 Inst_LUT4AB_switch_matrix__033_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG2_A0 Inst_LUT4AB_switch_matrix__037_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG3_A2 input167/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1_A1
+ input159/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst0_A1
+ input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG2_A2 input222/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput480 output480/A vssd1 vssd1 vccd1 vccd1 W6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput491 output491/A vssd1 vssd1 vccd1 vccd1 W6BEG[9] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit16_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit25_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LB_LUT4c_frame_config_dffesr__07_ Inst_LB_LUT4c_frame_config_dffesr__07_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__07_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_20_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit25 input67/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LG_LUT4c_frame_config_dffesr__13_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit14 input55/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst0 input104/X
+ input156/X input208/X Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_ConfigMem_Inst_Frame19_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit22/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XW6BEG_outbuf_2__0_ W6END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output484/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG1_A1 input8/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit10 input51/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit21 input63/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput208 W1END[2] vssd1 vssd1 vccd1 vccd1 input208/X sky130_fd_sc_hd__buf_4
Xinput219 W2MID[1] vssd1 vssd1 vccd1 vccd1 input219/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LG_LUT4c_frame_config_dffesr_cus_mux21_O__0_ Inst_LG_LUT4c_frame_config_dffesr__13_/A0
+ hold13/A Inst_LUT4AB_ConfigMem_Inst_Frame14_bit20/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__055_/A
+ sky130_fd_sc_hd__mux2_8
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit6/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit0/Q vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__08_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit13_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit22_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG3_A1 input7/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit3_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit31_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit20 input62/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit31 input74/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit18 input59/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit29 input71/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG2 input106/X input131/X input229/X
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_ConfigMem_Inst_Frame3_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 output380/A sky130_fd_sc_hd__mux4_1
XFILLER_0_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit7 input79/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit4_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1 input154/X
+ input156/X input190/X input238/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_31__0_ data_inbuf_31__0_/X vssd1 vssd1 vccd1 vccd1 output327/A sky130_fd_sc_hd__clkbuf_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_45_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit18_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit8 input80/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG0_A3 input225/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xdata_outbuf_22__0_ data_inbuf_22__0_/X vssd1 vssd1 vccd1 vccd1 output317/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0_A2
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_NN4BEG_outbuf_6__0__A NN4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG0_A0 input121/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit24 input66/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit13 input54/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_13__0_ data_inbuf_13__0_/X vssd1 vssd1 vccd1 vccd1 output307/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1_A3
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst0_A2
+ input206/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XS4BEG_outbuf_2__0_ S4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 output435/A sky130_fd_sc_hd__clkbuf_1
XInst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit18/Q Inst_LG_LUT4c_frame_config_dffesr__07_/A
+ Inst_LG_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit26/Q
+ vssd1 vssd1 vccd1 vccd1 output446/A sky130_fd_sc_hd__mux2_1
XFILLER_0_9_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit20 input62/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit31 input74/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG0_A0 input120/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1_A1
+ input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit30 input73/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit17 input58/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LC_LUT4c_frame_config_dffesr__13_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame17_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_J_EN_BEG0_cus_mux41_buf_inst1_A3
+ ANTENNA_14/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3 Inst_LUT4AB_ConfigMem_Inst_Frame6_bit0/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit5/Q vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__09_/A
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit28 input70/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit12/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit19/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__039_/A
+ sky130_fd_sc_hd__mux4_2
XS4END_inbuf_0__0_ input184/X vssd1 vssd1 vccd1 vccd1 ANTENNA_6/DIODE sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit7_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG0_A2 input165/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG1 input116/X input16/X
+ input168/X Inst_LUT4AB_switch_matrix__043_/A Inst_LUT4AB_ConfigMem_Inst_Frame12_bit6/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit7/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit2_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit8_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput309 output309/A vssd1 vssd1 vccd1 vccd1 FrameData_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_10_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0_A1
+ input111/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit3_GATE input93/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG1_cus_mux41_buf_inst2_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit2 input72/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG2 input145/X input41/X input181/X
+ Inst_LUT4AB_switch_matrix__083_/A Inst_LUT4AB_ConfigMem_Inst_Frame7_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit29/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A3 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG0_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XNN4END_inbuf_8__0_ input141/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_8__0_/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1_A2
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit19/Q Inst_LH_LUT4c_frame_config_dffesr__07_/A
+ Inst_LH_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S2_A3 ANTENNA_4/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst0_A1
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG0_A0 Inst_LUT4AB_switch_matrix__054_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XW6END_inbuf_4__0_ input234/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_2
XEE4BEG_outbuf_1__0_ EE4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output294/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit12 input53/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit23 input65/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG1_A2 ANTENNA_13/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit22_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit31_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit30 input73/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst0 input102/X
+ input2/X input154/X Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_ConfigMem_Inst_Frame10_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit22/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG2 input119/X input19/X
+ input171/X input223/X Inst_LUT4AB_ConfigMem_Inst_Frame9_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit2/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A1 sky130_fd_sc_hd__mux4_1
XFILLER_0_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1_A0
+ input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit0 input50/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit18_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit27_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__093_ input170/X vssd1 vssd1 vccd1 vccd1 output423/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1_A3
+ input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit16 input57/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit27 input69/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit10_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0_A0
+ input147/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LC_LUT4c_frame_config_dffesr__08_ Inst_LC_LUT4c_frame_config_dffesr__08_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__08_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_5_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A3 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit30/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit31/Q vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__10_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_68_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit12 input53/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit23 input65/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1_A1
+ input161/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit6_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput19 E2MID[5] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_2
XFILLER_0_64_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_N4BEG_outbuf_1__0__A N4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit15_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit7_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit5 input77/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit11 input52/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit22 input64/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit23/Q vssd1 vssd1 vccd1 vccd1 ANTENNA_3/DIODE
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__076_ input117/X vssd1 vssd1 vccd1 vccd1 output370/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG2_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDb_BEG3_A3 input219/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1_A2
+ input211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit29_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst0_A2
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABa_BEG2_A3 Inst_LUT4AB_switch_matrix__084_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput470 output470/A vssd1 vssd1 vccd1 vccd1 W2BEG[6] sky130_fd_sc_hd__buf_2
Xoutput492 output492/A vssd1 vssd1 vccd1 vccd1 WW4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput481 output481/A vssd1 vssd1 vccd1 vccd1 W6BEG[10] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG3_A0 input115/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_E6BEG_outbuf_2__0__A E6END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XEE4BEG_outbuf_11__0_ EE4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 output289/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_output277_A output277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit15 input56/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit26 input68/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__055_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A2 Inst_LUT4AB_ConfigMem_Inst_Frame19_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit22/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame19_bit8/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1_A0
+ input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_S4BEG_outbuf_9__0__A S4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG1_A2 input217/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG3_A0 input114/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit22 input64/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit11 input52/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput209 W1END[3] vssd1 vssd1 vccd1 vccd1 input209/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__059_ Inst_LUT4AB_switch_matrix__059_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__059_/X sky130_fd_sc_hd__buf_1
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A3 Inst_LUT4AB_ConfigMem_Inst_Frame9_bit2/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit4/Q vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__09_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xdata_outbuf_0__0_ data_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 output303/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG3_A2 input159/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit10 input51/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit21 input63/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LH_LUT4c_frame_config_dffesr__13_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_data_inbuf_17__0__A input58/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit10_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit19 input60/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LD_LUT4c_frame_config_dffesr__13_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame18_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst0_A1
+ input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit8 input80/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG3 input107/X input122/X input226/X
+ Inst_LUT4AB_switch_matrix__056_/A Inst_LUT4AB_ConfigMem_Inst_Frame3_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit28/Q
+ vssd1 vssd1 vccd1 vccd1 output381/A sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame9_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit15/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__083_/A
+ sky130_fd_sc_hd__mux4_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_24__0_ input66/X vssd1 vssd1 vccd1 vccd1 data_inbuf_24__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit9 input81/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG3_A0 Inst_LUT4AB_switch_matrix__032_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst0_A3
+ input13/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit15_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit24_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_inbuf_3__0_ input95/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xdata_inbuf_15__0_ input56/X vssd1 vssd1 vccd1 vccd1 data_inbuf_15__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG0_A1 input21/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit14 input55/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit25 input67/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_19_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG2_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1 Inst_LUT4AB_ConfigMem_Inst_Frame10_bit17/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit17/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit18/Q Inst_LG_LUT4c_frame_config_dffesr__07_/A
+ Inst_LG_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit10 input51/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit21 input63/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit29_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG0_A1 input20/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0_A1
+ input106/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG0_A0 Inst_LUT4AB_switch_matrix__037_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit12_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1_A2
+ input165/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit21_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit20 input62/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit31 input74/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_31_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit18 input59/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit29 input71/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A3 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit3/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit2/Q vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__10_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit30_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG0_A3 input217/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG2 input118/X input170/X
+ input222/X Inst_LUT4AB_switch_matrix__086_/A Inst_LUT4AB_ConfigMem_Inst_Frame2_bit5/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit3/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0
+ sky130_fd_sc_hd__mux4_2
XInst_LD_LUT4c_frame_config_dffesr__09_ Inst_LD_LUT4c_frame_config_dffesr__09_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__09_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit2_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0_A2
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit3_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit17_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xstrobe_outbuf_18__0_ strobe_inbuf_18__0_/X vssd1 vssd1 vccd1 vccd1 output344/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit26_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit3 input75/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LG_EN__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LG_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit1/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__14_/S sky130_fd_sc_hd__mux2_1
XFILLER_0_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG3 input122/X input190/X input226/X
+ ANTENNA_14/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame13_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit27/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A3 sky130_fd_sc_hd__mux4_1
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_NN4BEG_outbuf_5__0__A NN4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG4_cus_mux41_buf_inst1_A3
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4 Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ Inst_LH_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X Inst_LH_LUT4c_frame_config_dffesr__09_/A
+ Inst_LH_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__13_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst0_A2
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG0_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit24 input66/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit13 input54/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_E1BEG1_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit20 input62/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit31 input74/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XWW4END_inbuf_9__0_ input242/X vssd1 vssd1 vccd1 vccd1 WW4END_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__034_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A2 Inst_LUT4AB_ConfigMem_Inst_Frame10_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit22/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG2_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG3 input115/X input15/X
+ input167/X input219/X Inst_LUT4AB_ConfigMem_Inst_Frame11_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A1 sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1_A1
+ input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit1 input61/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__092_ input169/X vssd1 vssd1 vccd1 vccd1 output422/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG0 input147/X input12/X input164/X
+ input216/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit4/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I0/A2 sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst0_A1
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit17 input58/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_53_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit28 input70/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0_A1
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LC_LUT4c_frame_config_dffesr__07_ Inst_LC_LUT4c_frame_config_dffesr__07_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LC_LUT4c_frame_config_dffesr__07_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0 input107/X
+ input129/X input5/X input7/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit24 input66/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit13 input54/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1_A2
+ input213/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit6_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit7_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_74_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit6 input78/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xstrobe_outbuf_0__0_ strobe_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 output335/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit12 input53/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit23 input65/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit12_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I1_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit21_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit30_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__075_ input116/X vssd1 vssd1 vccd1 vccd1 output369/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1_A0
+ input183/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__100__A ANTENNA_3/DIODE vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG2_A2 ANTENNA_2/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit30 input73/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG0_cus_mux41_buf_inst1_A3
+ input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG3_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG6_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput471 output471/A vssd1 vssd1 vccd1 vccd1 W2BEG[7] sky130_fd_sc_hd__buf_2
Xoutput460 output460/A vssd1 vssd1 vccd1 vccd1 W1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput493 output493/A vssd1 vssd1 vccd1 vccd1 WW4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput482 output482/A vssd1 vssd1 vccd1 vccd1 W6BEG[11] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit17_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG3_A1 input15/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit20_D input62/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit4 input76/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_15__0_ input88/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_15__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit27 input69/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit16 input57/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XE6END_inbuf_9__0_ input24/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame0_bit7/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit6/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__070_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1_A1
+ input197/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_CD_BEG1_A3 Inst_LUT4AB_switch_matrix__040_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LF_LUT4c_frame_config_dffesr_cus_mux21_O__0_ Inst_LF_LUT4c_frame_config_dffesr__13_/A0
+ hold7/A Inst_LUT4AB_ConfigMem_Inst_Frame16_bit27/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__054_/A
+ sky130_fd_sc_hd__mux2_8
XFILLER_0_28_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG3_A1 input14/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit12 input53/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit23 input65/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix__058_ Inst_LUT4AB_switch_matrix__058_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__058_/X sky130_fd_sc_hd__buf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG3_A0 Inst_LUT4AB_switch_matrix__056_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_N4BEG_outbuf_0__0__A N4END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I3/A2
+ ANTENNA_5/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame13_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit12/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__10_/A sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit23_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_EF_BEG3_A3 input211/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput290 output290/A vssd1 vssd1 vccd1 vccd1 EE4BEG[12] sky130_fd_sc_hd__buf_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit11 input52/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit22 input64/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XE6BEG_outbuf_1__0_ E6END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output278/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst0_A2
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit9 input81/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_switch_matrix__055_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit15/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XN4END_inbuf_0__0_ input132/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_0__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit19_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit28_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_MUX8LUT_frame_config_mux_cus_mux21_AD__0__A0 Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG3_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_E6BEG_outbuf_1__0__A E6END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG0_A2 input173/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit15 input56/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit26 input68/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_S4BEG_outbuf_8__0__A S4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2 Inst_LUT4AB_ConfigMem_Inst_Frame12_bit15/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit15/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit14/Q Inst_LG_LUT4c_frame_config_dffesr__07_/A
+ Inst_LG_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit11 input52/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_7__0_ input79/X vssd1 vssd1 vccd1 vccd1 data_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit22 input64/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG0_A2 input172/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0_A2
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4_S1
+ Inst_LF_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG0_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG6_cus_mux41_buf_inst1_A3
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit10 input51/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit21 input63/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG0_A0 input147/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_16__0__A input57/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame17_bit19 input60/X input90/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_12_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG3 input14/X input166/X
+ input218/X Inst_LUT4AB_switch_matrix__102_/A Inst_LUT4AB_ConfigMem_Inst_Frame10_bit7/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit6/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I3/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LD_LUT4c_frame_config_dffesr__08_ Inst_LD_LUT4c_frame_config_dffesr__08_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__08_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst0_A0
+ input103/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst0_A3
+ input11/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit2_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit4 input76/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit3_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit14_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit23_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix__103__A ANTENNA_4/DIODE vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG0_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG0_A2 Inst_LUT4AB_switch_matrix__084_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit14 input55/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit25 input67/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_17_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit21 input63/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0_A1
+ input112/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit10 input51/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit19_D input60/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1_A2
+ input163/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit19_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit28_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit2 input72/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix__091_ input168/X vssd1 vssd1 vccd1 vccd1 output421/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG1 input108/X input8/X input160/X
+ input246/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit3/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A2 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit11_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xinput190 SS4END[0] vssd1 vssd1 vccd1 vccd1 input190/X sky130_fd_sc_hd__clkbuf_2
XNN4BEG_outbuf_1__0_ NN4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 output398/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst0_A2
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XN4BEG_outbuf_5__0_ N4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output386/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit18 input59/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit29 input71/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit20_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0_A2
+ input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG0_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_MUX8LUT_frame_config_mux_cus_mux21_CD__0_ Inst_LUT4AB_switch_matrix__034_/X
+ Inst_LUT4AB_switch_matrix__036_/X Inst_MUX8LUT_frame_config_mux_cus_mux21_CD__0_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_CD__0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XSS4BEG_outbuf_4__0_ SS4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output453/A sky130_fd_sc_hd__clkbuf_1
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1 input25/X
+ input197/X input211/X input229/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit25 input67/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit14 input55/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LG_LUT4c_frame_config_dffesr_cus_mux21_I0mux__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LG_I0/X
+ Inst_LUT4AB_switch_matrix__063_/X Inst_LUT4AB_ConfigMem_Inst_Frame12_bit13/Q vssd1
+ vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__07_/A sky130_fd_sc_hd__mux2_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG2_cus_mux41_buf_inst1_A3
+ input245/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit25_D input67/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit25_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit16_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit6_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_NN4BEG_outbuf_4__0__A NN4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit1_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit7 input79/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit7_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit13 input54/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit24 input66/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__074_ input115/X vssd1 vssd1 vccd1 vccd1 output368/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1_A1
+ input199/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XW6BEG_outbuf_5__0_ W6END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output487/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N1BEG2_A3 ANTENNA_5/DIODE vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0 input103/X
+ input109/X input131/X input9/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit20 input62/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit31 input74/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst0_A1
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput461 output461/A vssd1 vssd1 vccd1 vccd1 W1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput450 output450/A vssd1 vssd1 vccd1 vccd1 SS4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput472 output472/A vssd1 vssd1 vccd1 vccd1 W2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput494 output494/A vssd1 vssd1 vccd1 vccd1 WW4BEG[11] sky130_fd_sc_hd__buf_2
Xoutput483 output483/A vssd1 vssd1 vccd1 vccd1 W6BEG[1] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG3_A2 input167/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0_A1
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_64_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit13_D input54/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit5 input77/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit17 input58/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit28 input70/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG1_A0 input42/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1_A2
+ input211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG3_A2 input218/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit13 input54/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix__111__A input224/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__057_ input1/X vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__057_/X
+ sky130_fd_sc_hd__buf_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit24 input66/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG3_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG3_A0 input106/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1_A0
+ input159/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit23/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit23/Q Inst_LF_LUT4c_frame_config_dffesr__07_/A
+ Inst_LF_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xdata_outbuf_25__0_ data_inbuf_25__0_/X vssd1 vssd1 vccd1 vccd1 output320/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput280 output280/A vssd1 vssd1 vccd1 vccd1 E6BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput291 output291/A vssd1 vssd1 vccd1 vccd1 EE4BEG[13] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit23 input65/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit12 input53/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit11_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit20_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit5_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_SS4BEG_outbuf_9__0__A SS4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame7_bit10/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit13/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__045_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG4_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xdata_outbuf_16__0_ data_inbuf_16__0_/X vssd1 vssd1 vccd1 vccd1 output310/A sky130_fd_sc_hd__clkbuf_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit30 input73/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XS4BEG_outbuf_5__0_ S4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 output438/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LE_LUT4c_frame_config_dffesr__09_ Inst_LE_LUT4c_frame_config_dffesr__09_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__09_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix__106__A input219/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG3_A2 Inst_LUT4AB_switch_matrix__083_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__109_ input222/X vssd1 vssd1 vccd1 vccd1 output476/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit25_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit16 input57/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG0_A3 input225/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit27 input69/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_34_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XS4END_inbuf_3__0_ input187/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_4
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0 input103/X
+ input111/X input3/X input11/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG0 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A1 Inst_LUT4AB_switch_matrix__084_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3 Inst_LUT4AB_ConfigMem_Inst_Frame19_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit19/Q vssd1 vssd1 vccd1 vccd1 output460/A sky130_fd_sc_hd__mux4_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3 Inst_LUT4AB_ConfigMem_Inst_Frame5_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit14/Q Inst_LG_LUT4c_frame_config_dffesr__07_/A
+ Inst_LG_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG2_A0 input25/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit0 input50/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit23 input65/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit12 input53/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG0_A3 Inst_LUT4AB_switch_matrix__071_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst0_A3
+ input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG1_A0 input117/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG0_A2 Inst_LUT4AB_switch_matrix__041_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit13_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit22_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit31_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit22 input64/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit11 input52/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG0_A0 input120/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XW6END_inbuf_7__0_ input237/X vssd1 vssd1 vccd1 vccd1 W6END_inbuf_7__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XEE4BEG_outbuf_4__0_ EE4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output297/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG0_A1 input12/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit9_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LD_LUT4c_frame_config_dffesr__07_ Inst_LD_LUT4c_frame_config_dffesr__07_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr__07_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst0_A1
+ input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0_A1
+ input106/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit18_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit5 input77/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_E6BEG_outbuf_0__0__A E6END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LA_SR__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG0_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit15 input56/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit26 input68/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_S4BEG_outbuf_7__0__A S4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0_A2
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit22 input64/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit11 input52/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0 input110/X
+ input4/X input10/X input22/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1_A3
+ input207/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit3 input75/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix__090_ input167/X vssd1 vssd1 vccd1 vccd1 output420/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG2 input110/X input10/X input198/X
+ input214/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit5/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A2 sky130_fd_sc_hd__mux4_2
XFILLER_0_10_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput180 S4END[15] vssd1 vssd1 vccd1 vccd1 input180/X sky130_fd_sc_hd__clkbuf_1
Xinput191 SS4END[10] vssd1 vssd1 vccd1 vccd1 input191/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG3_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_data_inbuf_15__0__A input56/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst0_A0
+ input105/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame16_bit19 input60/X input89/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst0_A3
+ input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__033_/A
+ Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit26 input68/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit15 input56/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG0 input121/X input21/X
+ input173/X input225/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A1 sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit18_D input59/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit31_D input74/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit13_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit8 input80/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit1_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit14 input55/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit25 input67/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit22_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit31_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__073_ input114/X vssd1 vssd1 vccd1 vccd1 output367/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit2_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_3_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1_A2
+ input213/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__109__A input222/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XN4END_inbuf_11__0_ input128/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_11__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1 input25/X
+ input161/X input213/X input229/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit21 input63/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit10 input51/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1_A0
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst0_A2
+ input209/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput462 output462/A vssd1 vssd1 vccd1 vccd1 W1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput451 output451/A vssd1 vssd1 vccd1 vccd1 SS4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput440 output440/A vssd1 vssd1 vccd1 vccd1 S4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput473 output473/A vssd1 vssd1 vccd1 vccd1 W2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput495 output495/A vssd1 vssd1 vccd1 vccd1 WW4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput484 output484/A vssd1 vssd1 vccd1 vccd1 W6BEG[2] sky130_fd_sc_hd__clkbuf_4
XSS4END_inbuf_10__0_ input195/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_10__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit18_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit27_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG3_A3 input219/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LE_LUT4c_frame_config_dffesr_cus_mux21_O__0_ Inst_LE_LUT4c_frame_config_dffesr__13_/A0
+ hold5/A Inst_LUT4AB_ConfigMem_Inst_Frame17_bit24/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__037_/A
+ sky130_fd_sc_hd__mux2_8
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0_A2
+ input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit6 input78/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xdata_outbuf_3__0_ data_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output328/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit29 input71/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit18 input59/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit10_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG1_A1 input182/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1_A3
+ input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHa_BEG3_A3 ANTENNA_4/DIODE
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix__056_ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__056_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit14 input55/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit25 input67/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG7_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_27__0_ input69/X vssd1 vssd1 vccd1 vccd1 data_inbuf_27__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG3_A2 Inst_LUT4AB_switch_matrix__040_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit15_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG3_A0 input14/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit24_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG3_A1 input41/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1_A1
+ input181/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_NN4BEG_outbuf_3__0__A NN4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1 Inst_LUT4AB_ConfigMem_Inst_Frame15_bit19/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit17/Q Inst_LF_LUT4c_frame_config_dffesr__07_/A
+ Inst_LF_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
Xoutput270 output270/A vssd1 vssd1 vccd1 vccd1 E2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput281 output281/A vssd1 vssd1 vccd1 vccd1 E6BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput292 output292/A vssd1 vssd1 vccd1 vccd1 EE4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xstrobe_inbuf_6__0_ input98/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_18__0_ input59/X vssd1 vssd1 vccd1 vccd1 data_inbuf_18__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit24 input66/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit13 input54/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit5_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit6_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit20 input62/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit31 input74/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit29_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LE_LUT4c_frame_config_dffesr__08_ Inst_LE_LUT4c_frame_config_dffesr__08_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__08_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG3_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__108_ input221/X vssd1 vssd1 vccd1 vccd1 output475/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix__039_ Inst_LUT4AB_switch_matrix__039_/A vssd1 vssd1 vccd1
+ vccd1 output260/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit17 input58/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit28 input70/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit0 input50/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__032__A Inst_LUT4AB_switch_matrix__032_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1 input155/X
+ input157/X input163/X input207/X Inst_LUT4AB_ConfigMem_Inst_Frame19_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG1 Inst_LUT4AB_switch_matrix__055_/A
+ ANTENNA_21/DIODE Inst_LUT4AB_switch_matrix__081_/A Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A3
+ Inst_LUT4AB_ConfigMem_Inst_Frame0_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit16/Q
+ vssd1 vssd1 vccd1 vccd1 output461/A sky130_fd_sc_hd__mux4_1
XInst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4 Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ Inst_LG_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X Inst_LG_LUT4c_frame_config_dffesr__09_/A
+ Inst_LG_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__13_/A0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG2_A1 input181/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit13 input54/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit1 input61/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit24 input66/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XS4END_inbuf_11__0_ input180/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_11__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG2_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG1_A1 input17/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG0_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit23 input65/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit12 input53/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG0_A1 input20/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I1_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG0_A2 input164/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit10_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_SS4BEG_outbuf_8__0__A SS4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0 input105/X
+ input113/X input5/X input13/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit9_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit30 input73/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst0_A2
+ input155/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0_A2
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit6 input78/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit15_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit24_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LE_SR__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit16 input57/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit27 input69/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XSS4END_inbuf_1__0_ input201/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_1__0_/X sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XEE4END_inbuf_10__0_ input39/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_10__0_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst0_A3
+ input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit12 input53/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit23 input65/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1 input162/X
+ input174/X input214/X input246/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit4 input76/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG3 input106/X input41/X input158/X
+ input210/X Inst_LUT4AB_ConfigMem_Inst_Frame8_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit3/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I3/A2 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit12_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit21_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput181 S4END[1] vssd1 vssd1 vccd1 vccd1 input181/X sky130_fd_sc_hd__buf_2
Xinput170 S2MID[4] vssd1 vssd1 vccd1 vccd1 input170/X sky130_fd_sc_hd__buf_4
Xinput192 SS4END[11] vssd1 vssd1 vccd1 vccd1 input192/X sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_3__0_ strobe_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 output348/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst0_A1
+ input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0_A1
+ input112/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit16 input57/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit27 input69/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XEE4END_inbuf_0__0_ input44/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_0__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit26_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG1 input117/X input17/X
+ input169/X input221/X Inst_LUT4AB_ConfigMem_Inst_Frame1_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit0/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1 sky130_fd_sc_hd__mux4_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__040__A Inst_LUT4AB_switch_matrix__040_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit24_D input66/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit9 input81/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XWW4BEG_outbuf_1__0_ ANTENNA_7/DIODE vssd1 vssd1 vccd1 vccd1 output499/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit15 input56/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_18__0_ input91/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_18__0_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit26 input68/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst0_A2
+ input122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__072_ Inst_LUT4AB_switch_matrix__072_/A vssd1 vssd1 vccd1
+ vccd1 output366/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_S4BEG_outbuf_6__0__A S4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG2_cus_mux41_buf_inst1_A3
+ input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0_A0
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit22 input64/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit11 input52/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1_A1
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput441 output441/A vssd1 vssd1 vccd1 vccd1 S4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput430 output430/A vssd1 vssd1 vccd1 vccd1 S4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput452 output452/A vssd1 vssd1 vccd1 vccd1 SS4BEG[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_NN4BEG1_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput474 output474/A vssd1 vssd1 vccd1 vccd1 W2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput463 output463/A vssd1 vssd1 vccd1 vccd1 W1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput496 output496/A vssd1 vssd1 vccd1 vccd1 WW4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput485 output485/A vssd1 vssd1 vccd1 vccd1 W6BEG[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit29_D input71/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst0_A3
+ input25/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LF_LUT4c_frame_config_dffesr__09_ Inst_LF_LUT4c_frame_config_dffesr__09_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__09_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit7 input79/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit12_D input53/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit30_D input73/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_14__0__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LE_SR__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LE_SR__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_SR__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame18_bit1/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__13_/S sky130_fd_sc_hd__mux2_1
XInst_LUT4AB_ConfigMem_Inst_Frame15_bit19 input60/X input88/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame15_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XE6BEG_outbuf_4__0_ E6END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output281/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG1_A2 input217/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_data_inbuf_29__0__A input71/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix__055_ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__055_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XN4END_inbuf_3__0_ input135/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit15 input56/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit26 input68/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1BEG3_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG3_A1 input166/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0_A1
+ input108/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG3_A2 input158/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1_A2
+ input211/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit22/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit29/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit28/Q Inst_LF_LUT4c_frame_config_dffesr__07_/A
+ Inst_LF_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput260 output260/A vssd1 vssd1 vccd1 vccd1 E2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput271 output271/A vssd1 vssd1 vccd1 vccd1 E2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput282 output282/A vssd1 vssd1 vccd1 vccd1 E6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput293 output293/A vssd1 vssd1 vccd1 vccd1 EE4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit14 input55/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit25 input67/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit12_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit30_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit21_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit5_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit21 input63/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit10 input51/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit0_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit6_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LE_LUT4c_frame_config_dffesr__07_ Inst_LE_LUT4c_frame_config_dffesr__07_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr__07_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit17_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit1_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__107_ input220/X vssd1 vssd1 vccd1 vccd1 output474/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix__038_ Inst_LUT4AB_switch_matrix__038_/A vssd1 vssd1 vccd1
+ vccd1 output259/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit29 input71/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit18 input59/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_19_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit1 input61/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG5_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG2 Inst_LUT4AB_switch_matrix__056_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I1/A1 Inst_LUT4AB_switch_matrix__082_/A
+ ANTENNA_5/DIODE Inst_LUT4AB_ConfigMem_Inst_Frame0_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame0_bit23/Q
+ vssd1 vssd1 vccd1 vccd1 output462/A sky130_fd_sc_hd__mux4_1
XFILLER_0_15_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG2_A2 input247/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit2 input72/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit25 input67/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit14 input55/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_53_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_40_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit14_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LA_LUT4c_frame_config_dffesr_cus_mux21_I0mux__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LA_I0/X
+ Inst_LUT4AB_switch_matrix__057_/X Inst_LUT4AB_ConfigMem_Inst_Frame16_bit3/Q vssd1
+ vssd1 vccd1 vccd1 Inst_LA_LUT4c_frame_config_dffesr__07_/A sky130_fd_sc_hd__mux2_2
XANTENNA_NN4BEG_outbuf_2__0__A NN4END_inbuf_2__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG1_A2 input169/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit23_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit13 input54/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit24 input66/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG0_A2 input224/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LB_EN__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LB_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame13_bit27/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LB_LUT4c_frame_config_dffesr__14_/S sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LE_I1_A2 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I1/A2
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG0_A3 input216/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame11_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 output293/A sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1 input157/X
+ input165/X input207/X input209/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit20 input62/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit31 input74/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__043__A Inst_LUT4AB_switch_matrix__043_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst0_A3
+ input34/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit19_GATE input95/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit28_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit9_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit4_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit7 input79/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_1 ANTENNA_2/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit5_GATE input94/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_21_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit17 input58/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit28 input70/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XNN4BEG_outbuf_4__0_ NN4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output401/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XN4BEG_outbuf_8__0_ N4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output389/A sky130_fd_sc_hd__clkbuf_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0_A1
+ input138/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XSS4BEG_outbuf_7__0_ SS4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output456/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit24 input66/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG0_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit13 input54/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix__038__A Inst_LUT4AB_switch_matrix__038_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XS4BEG_outbuf_11__0_ S4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 output429/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit5 input77/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput171 S2MID[5] vssd1 vssd1 vccd1 vccd1 input171/X sky130_fd_sc_hd__buf_2
Xinput160 S2END[2] vssd1 vssd1 vccd1 vccd1 input160/X sky130_fd_sc_hd__buf_2
Xinput182 S4END[2] vssd1 vssd1 vccd1 vccd1 input182/X sky130_fd_sc_hd__buf_2
Xinput193 SS4END[12] vssd1 vssd1 vccd1 vccd1 input193/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst0_A2
+ input157/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0_A2
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_SS4BEG_outbuf_7__0__A SS4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_41_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XW6BEG_outbuf_8__0_ W6END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output490/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG0_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame4_bit8/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit5/Q vssd1 vssd1 vccd1 vccd1 ANTENNA_13/DIODE
+ sky130_fd_sc_hd__mux4_2
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit30 input73/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit17 input58/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit28 input70/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG2 input119/X input19/X
+ input171/X input223/X Inst_LUT4AB_ConfigMem_Inst_Frame10_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit2/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1 sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LG_LUT4c_frame_config_dffesr__10__A Inst_LG_LUT4c_frame_config_dffesr__10_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit14_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit17_D input58/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit8_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit23_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit16 input57/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit27 input69/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit9_GATE input93/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__071_ Inst_LUT4AB_switch_matrix__071_/A vssd1 vssd1 vccd1
+ vccd1 output365/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LD_LUT4c_frame_config_dffesr_cus_mux21_O__0_ Inst_LD_LUT4c_frame_config_dffesr__13_/A0
+ hold11/A Inst_LUT4AB_ConfigMem_Inst_Frame18_bit29/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__036_/A
+ sky130_fd_sc_hd__mux2_8
XNN4END_inbuf_1__0_ input149/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_1__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit21/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit21/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit20/Q Inst_LE_LUT4c_frame_config_dffesr__07_/A
+ Inst_LE_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0_A1
+ input208/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit23 input65/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit12 input53/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit17/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1_A2
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput420 output420/A vssd1 vssd1 vccd1 vccd1 S2BEGb[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit2_D input72/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xoutput431 output431/A vssd1 vssd1 vccd1 vccd1 S4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput442 output442/A vssd1 vssd1 vccd1 vccd1 S4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput453 output453/A vssd1 vssd1 vccd1 vccd1 SS4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput464 output464/A vssd1 vssd1 vccd1 vccd1 W2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput475 output475/A vssd1 vssd1 vccd1 vccd1 W2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput486 output486/A vssd1 vssd1 vccd1 vccd1 W6BEG[4] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit28_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xoutput497 output497/A vssd1 vssd1 vccd1 vccd1 WW4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0_A1
+ input122/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LF_LUT4c_frame_config_dffesr__08_ Inst_LF_LUT4c_frame_config_dffesr__08_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__08_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_64_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit11_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_28__0_ data_inbuf_28__0_/X vssd1 vssd1 vccd1 vccd1 output323/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit6_D input78/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit8 input80/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix__051__A input19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit23_D input65/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_AB_BEG1_A3 Inst_LUT4AB_switch_matrix__039_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit20_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_outbuf_19__0_ data_inbuf_19__0_/X vssd1 vssd1 vccd1 vccd1 output313/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_switch_matrix__054_ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__054_/X sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit16 input57/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit27 input69/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XS4BEG_outbuf_8__0_ S4END_inbuf_8__0_/X vssd1 vssd1 vccd1 vccd1 output441/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit16_GATE input94/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG3_A2 input218/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0_A2
+ input130/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit25_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_CD_BEG3_A3 input210/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG0_cus_mux41_buf_inst1_A3
+ input229/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3 Inst_LUT4AB_ConfigMem_Inst_Frame14_bit19/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame16_bit28/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit23/Q Inst_LF_LUT4c_frame_config_dffesr__07_/A
+ Inst_LF_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
Xoutput261 output261/A vssd1 vssd1 vccd1 vccd1 E2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput283 output283/A vssd1 vssd1 vccd1 vccd1 E6BEG[6] sky130_fd_sc_hd__buf_2
Xoutput272 output272/A vssd1 vssd1 vccd1 vccd1 E2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput294 output294/A vssd1 vssd1 vccd1 vccd1 EE4BEG[1] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit15 input56/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit26 input68/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix__046__A input14/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG7_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_S4BEG_outbuf_5__0__A S4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit11_D input52/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_52_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG0_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame0_bit21/Q
+ vssd1 vssd1 vccd1 vccd1 output495/A sky130_fd_sc_hd__mux2_1
XS4END_inbuf_6__0_ input175/X vssd1 vssd1 vccd1 vccd1 S4END_inbuf_6__0_/X sky130_fd_sc_hd__clkbuf_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0_A0
+ input108/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit11 input52/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit22 input64/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit0_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix__106_ input219/X vssd1 vssd1 vccd1 vccd1 output473/A sky130_fd_sc_hd__buf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit1_GATE input99/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__037_ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__037_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit1_D input61/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_data_inbuf_13__0__A input54/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit19 input60/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit2 input72/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit2/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_19_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_data_inbuf_28__0__A input70/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XEE4BEG_outbuf_7__0_ EE4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output300/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit5_D input77/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame19_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_W1BEG3 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A1 Inst_LUT4AB_switch_matrix__083_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A3 Inst_LUT4AB_ConfigMem_Inst_Frame8_bit25/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit26/Q vssd1 vssd1 vccd1 vccd1 output463/A sky130_fd_sc_hd__mux4_1
XFILLER_0_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_GH_BEG2_A3 Inst_LUT4AB_switch_matrix__085_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit15 input56/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit3 input75/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit26 input68/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit9_D input81/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_GHb_BEG1_A3 input221/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG0_A0 input112/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit14 input55/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit25 input67/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit11_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit20_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG1_A0 input117/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG0_A0 input20/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst0 input105/X
+ input157/X input209/X Inst_LUT4AB_switch_matrix__032_/A Inst_LUT4AB_ConfigMem_Inst_Frame1_bit31/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit30/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2 Inst_LUT4AB_switch_matrix__032_/A
+ Inst_LUT4AB_switch_matrix__033_/A Inst_LUT4AB_switch_matrix__034_/A Inst_LUT4AB_switch_matrix__036_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit21 input63/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit10 input51/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__037_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_30_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit16_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit8 input80/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S0 Inst_LUT4AB_switch_matrix__069_/A
+ Inst_LUT4AB_switch_matrix__042_/A Inst_LUT4AB_switch_matrix__085_/A Inst_LUT4AB_switch_matrix__101_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit1/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/S sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit4_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG3_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit25_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_2 ANTENNA_2/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit5_GATE input98/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit18 input59/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit29 input71/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit0_GATE input82/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0_A2
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_4_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit25 input67/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit14 input55/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__054_/A
+ Inst_LUT4AB_switch_matrix__055_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit9/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix__054__A Inst_LUT4AB_switch_matrix__054_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit6 input78/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit6/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_NN4BEG_outbuf_1__0__A NN4END_inbuf_1__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit13_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit31_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit22_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XNN4BEG_outbuf_11__0_ NN4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 output393/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xinput172 S2MID[6] vssd1 vssd1 vccd1 vccd1 input172/X sky130_fd_sc_hd__clkbuf_2
Xinput161 S2END[3] vssd1 vssd1 vccd1 vccd1 input161/X sky130_fd_sc_hd__buf_2
Xinput150 NN4END[6] vssd1 vssd1 vccd1 vccd1 input150/X sky130_fd_sc_hd__clkbuf_1
Xinput183 S4END[3] vssd1 vssd1 vccd1 vccd1 input183/X sky130_fd_sc_hd__buf_2
Xinput194 SS4END[13] vssd1 vssd1 vccd1 vccd1 input194/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG1_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LG_LUT4c_frame_config_dffesr__09_ Inst_LG_LUT4c_frame_config_dffesr__09_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__09_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst0_A3
+ input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG1_A0 input109/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XNN4END_inbuf_10__0_ input143/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_10__0_/X sky130_fd_sc_hd__clkbuf_4
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit20 input62/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit31 input74/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit18_GATE input98/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit27_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit29 input71/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit18 input59/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_ABb_BEG3 input115/X input15/X
+ input167/X input219/X Inst_LUT4AB_ConfigMem_Inst_Frame12_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I3/A1 sky130_fd_sc_hd__mux4_1
XFILLER_0_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0_A1
+ input112/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__049__A input17/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit28_D input70/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit8_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit17 input58/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit28 input70/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xstrobe_outbuf_11__0_ strobe_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 output337/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__070_ Inst_LUT4AB_switch_matrix__070_/A vssd1 vssd1 vccd1
+ vccd1 output364/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xdata_outbuf_6__0_ data_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output331/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit9_GATE input97/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit20/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame15_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit26/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit25/Q Inst_LE_LUT4c_frame_config_dffesr__07_/A
+ Inst_LE_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0_A2
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit24 input66/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG2_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame6_bit12/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit8/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__040_/A
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit13 input54/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_W6BEG0_cus_mux41_buf_inst1_A3
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput410 output410/A vssd1 vssd1 vccd1 vccd1 S1BEG[3] sky130_fd_sc_hd__buf_2
Xoutput421 output421/A vssd1 vssd1 vccd1 vccd1 S2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput443 output443/A vssd1 vssd1 vccd1 vccd1 SS4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput432 output432/A vssd1 vssd1 vccd1 vccd1 S4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput465 output465/A vssd1 vssd1 vccd1 vccd1 W2BEG[1] sky130_fd_sc_hd__buf_2
Xoutput454 output454/A vssd1 vssd1 vccd1 vccd1 SS4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput476 output476/A vssd1 vssd1 vccd1 vccd1 W2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput487 output487/A vssd1 vssd1 vccd1 vccd1 W6BEG[5] sky130_fd_sc_hd__buf_2
Xoutput498 output498/A vssd1 vssd1 vccd1 vccd1 WW4BEG[15] sky130_fd_sc_hd__buf_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst0_A2
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG1_A0 input109/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XWW4END_inbuf_2__0_ input250/X vssd1 vssd1 vccd1 vccd1 WW4END_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LF_LUT4c_frame_config_dffesr__07_ Inst_LF_LUT4c_frame_config_dffesr__07_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__07_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_49_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit0 input50/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit0/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit9 input81/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LC_I1_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_9__0_ input101/X vssd1 vssd1 vccd1 vccd1 strobe_inbuf_9__0_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit16_D input57/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_SS4BEG_outbuf_6__0__A SS4END_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit30 input73/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit30/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst0_A0
+ input104/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__053_ input21/X vssd1 vssd1 vccd1 vccd1 output274/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit28 input70/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit17 input58/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG3_A0 input106/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFa_BEG3_A3 Inst_LUT4AB_switch_matrix__102_/A
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst0_A3
+ input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG7_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst0 input103/X
+ input3/X input155/X Inst_LUT4AB_switch_matrix__036_/A Inst_LUT4AB_ConfigMem_Inst_Frame10_bit21/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit26/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__0_/A0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit13_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst4 Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst1/X Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ Inst_LF_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst3/X Inst_LF_LUT4c_frame_config_dffesr__09_/A
+ Inst_LF_LUT4c_frame_config_dffesr__10_/A vssd1 vssd1 vccd1 vccd1 Inst_LF_LUT4c_frame_config_dffesr__13_/A0
+ sky130_fd_sc_hd__mux4_1
Xoutput262 output262/A vssd1 vssd1 vccd1 vccd1 E2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput284 output284/A vssd1 vssd1 vccd1 vccd1 E6BEG[7] sky130_fd_sc_hd__buf_2
Xoutput273 output273/A vssd1 vssd1 vccd1 vccd1 E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput295 output295/A vssd1 vssd1 vccd1 vccd1 EE4BEG[2] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit16 input57/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG3_A0 input114/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit27 input69/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit22_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit31_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_25_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0_A1
+ input130/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit12 input53/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit23 input65/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit18_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit27_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix__105_ input218/X vssd1 vssd1 vccd1 vccd1 output472/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix__036_ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1
+ vccd1 Inst_LUT4AB_switch_matrix__036_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_EE4BEG_outbuf_11__0__A EE4END_inbuf_11__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit10_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit3 input75/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit3/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG2_A0 input129/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG4_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit24/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit24/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__101_/A
+ sky130_fd_sc_hd__mux4_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit16 input57/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XE6END_inbuf_2__0_ input28/X vssd1 vssd1 vccd1 vccd1 E6END_inbuf_2__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit27 input69/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit4 input76/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit15_GATE input97/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit24_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG5_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AD__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG0_A1 input12/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit15 input56/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit26 input68/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG1_A1 input17/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_S4BEG_outbuf_4__0__A S4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG0_A1 input172/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__056_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A2 Inst_LUT4AB_ConfigMem_Inst_Frame1_bit31/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit30/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_WW4BEG1_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix__054_/A Inst_LUT4AB_switch_matrix__056_/A Inst_MUX8LUT_frame_config_mux_cus_mux21_M_AH__0_/X
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit11/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit22 input64/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit22/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit11 input52/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit11/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XSS4END_inbuf_4__0_ input204/X vssd1 vssd1 vccd1 vccd1 SS4END_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LB_SR__0__509 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LB_SR__0__509/HI
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LB_SR__0_/A0 sky130_fd_sc_hd__conb_1
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame18_bit9 input81/X input91/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit9/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S1 Inst_LUT4AB_switch_matrix__070_/A
+ Inst_LUT4AB_switch_matrix__043_/A Inst_LUT4AB_switch_matrix__086_/A Inst_LUT4AB_switch_matrix__102_/A
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit3/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_AD__0_/S sky130_fd_sc_hd__mux4_2
XFILLER_0_53_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_3 ANTENNA_3/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_data_inbuf_12__0__A input53/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame13_bit19 input60/X input86/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame13_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame13_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_6__0_ strobe_inbuf_6__0_/X vssd1 vssd1 vccd1 vccd1 output351/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_data_inbuf_27__0__A input69/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst0_A3
+ input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LD_EN__0__519 vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LD_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LD_EN__0__519/LO sky130_fd_sc_hd__conb_1
XFILLER_0_8_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit0_GATE input96/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit15 input56/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit15/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit26 input68/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit26/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame2_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit17/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__084_/A
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XEE4END_inbuf_3__0_ input47/X vssd1 vssd1 vccd1 vccd1 EE4END_inbuf_3__0_/X sky130_fd_sc_hd__clkbuf_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit7 input79/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit7/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_23_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xdata_inbuf_0__0_ input50/X vssd1 vssd1 vccd1 vccd1 data_inbuf_0__0_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput162 S2END[4] vssd1 vssd1 vccd1 vccd1 input162/X sky130_fd_sc_hd__buf_2
Xinput151 NN4END[7] vssd1 vssd1 vccd1 vccd1 input151/X sky130_fd_sc_hd__clkbuf_1
Xinput140 NN4END[11] vssd1 vssd1 vccd1 vccd1 input140/X sky130_fd_sc_hd__clkbuf_1
Xinput184 S4END[4] vssd1 vssd1 vccd1 vccd1 input184/X sky130_fd_sc_hd__clkbuf_1
Xinput195 SS4END[14] vssd1 vssd1 vccd1 vccd1 input195/X sky130_fd_sc_hd__clkbuf_1
Xinput173 S2MID[7] vssd1 vssd1 vccd1 vccd1 input173/X sky130_fd_sc_hd__buf_2
XFILLER_0_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1_A3 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LD_I1/A3
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XWW4BEG_outbuf_4__0_ WW4END_inbuf_4__0_/X vssd1 vssd1 vccd1 vccd1 output502/A sky130_fd_sc_hd__clkbuf_1
XInst_LG_LUT4c_frame_config_dffesr__08_ Inst_LG_LUT4c_frame_config_dffesr__08_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__08_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit10_GATE input90/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3_A0
+ Inst_LUT4AB_switch_matrix__054_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG1_A1 input9/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit10 input51/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit10/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame2_bit21 input63/X input94/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame2_bit21/Q Inst_LUT4AB_ConfigMem_Inst_Frame2_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG1_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame9_bit19 input60/X input101/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit19/Q Inst_LUT4AB_ConfigMem_Inst_Frame9_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_MUX8LUT_frame_config_mux_cus_mux21_sGH__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_EH__0_/S
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/S Inst_LUT4AB_ConfigMem_Inst_Frame4_bit24/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_GH__0_/S sky130_fd_sc_hd__mux2_1
XInst_LC_LUT4c_frame_config_dffesr_cus_mux21_O__0_ Inst_LC_LUT4c_frame_config_dffesr__13_/A0
+ hold15/A Inst_LUT4AB_ConfigMem_Inst_Frame18_bit15/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__034_/A
+ sky130_fd_sc_hd__mux2_8
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG1_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst0_A2
+ input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit15_GATE input84/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame14_bit24_GATE input87/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__065__A ANTENNA_13/DIODE vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_SS4BEG3_my_mux2_inst__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame9_bit25/Q
+ vssd1 vssd1 vccd1 vccd1 output449/A sky130_fd_sc_hd__mux2_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit18 input59/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame12_bit29 input71/X input85/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame12_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame12_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit8_GATE input92/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XE6BEG_outbuf_7__0_ E6END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output284/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit3_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit9_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2 Inst_LUT4AB_ConfigMem_Inst_Frame18_bit28/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame18_bit26/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame18_bit25/Q Inst_LE_LUT4c_frame_config_dffesr__07_/A
+ Inst_LE_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LE_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst0_A3
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit14 input55/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit14/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit25 input67/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit25/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame3_bit4_GATE input95/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput400 output400/A vssd1 vssd1 vccd1 vccd1 NN4BEG[3] sky130_fd_sc_hd__clkbuf_4
XN4END_inbuf_6__0_ input123/X vssd1 vssd1 vccd1 vccd1 N4END_inbuf_6__0_/X sky130_fd_sc_hd__buf_2
Xoutput411 output411/A vssd1 vssd1 vccd1 vccd1 S2BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_14_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput422 output422/A vssd1 vssd1 vccd1 vccd1 S2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput433 output433/A vssd1 vssd1 vccd1 vccd1 S4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput444 output444/A vssd1 vssd1 vccd1 vccd1 SS4BEG[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput466 output466/A vssd1 vssd1 vccd1 vccd1 W2BEG[2] sky130_fd_sc_hd__buf_2
Xoutput455 output455/A vssd1 vssd1 vccd1 vccd1 SS4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput477 output477/A vssd1 vssd1 vccd1 vccd1 W2BEGb[5] sky130_fd_sc_hd__buf_2
Xoutput499 output499/A vssd1 vssd1 vccd1 vccd1 WW4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput488 output488/A vssd1 vssd1 vccd1 vccd1 W6BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_0_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_N4BEG1_A1 input130/X vssd1 vssd1
+ vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_NN4BEG_outbuf_0__0__A NN4END_inbuf_0__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1 Inst_LUT4AB_ConfigMem_Inst_Frame3_bit1/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__14_/S sky130_fd_sc_hd__mux2_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame4_bit12_GATE input96/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame14_bit1 input61/X input87/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame14_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame14_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit21_GATE input99/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame6_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit22_D input64/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_28_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit20 input62/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit20/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame1_bit31 input74/X input93/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame1_bit31/Q Inst_LUT4AB_ConfigMem_Inst_Frame1_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix__052_ input20/X vssd1 vssd1 vccd1 vccd1 output273/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame9_bit17_GATE input101/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit29 input71/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit29/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit18 input59/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit18/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG3_A1 input6/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame1_bit26_GATE input93/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_W6BEG_outbuf_9__0__A W6END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_cus_mux41_buf_inst1 Inst_LUT4AB_switch_matrix__037_/A
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LF_I2/A0 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I0/A2 Inst_LUT4AB_ConfigMem_Inst_Frame10_bit21/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit26/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux81_buf_EE4BEG3_my_mux2_inst__0_/A1
+ sky130_fd_sc_hd__mux4_1
Xoutput285 output285/A vssd1 vssd1 vccd1 vccd1 E6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput263 output263/A vssd1 vssd1 vccd1 vccd1 E2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput274 output274/A vssd1 vssd1 vccd1 vccd1 E2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput296 output296/A vssd1 vssd1 vccd1 vccd1 EE4BEG[3] sky130_fd_sc_hd__buf_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit17 input58/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG3_A1 input166/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit28 input70/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit27_D input69/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame17_bit0_D input50/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_18_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame5_bit15_D input56/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit10_D input51/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0_A2
+ input2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit13 input54/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit13/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame4_bit24 input66/X input96/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame4_bit24/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame12_bit7_GATE input85/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit4_D input76/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0 input108/X
+ input130/X input2/X input8/X Inst_LUT4AB_ConfigMem_Inst_Frame5_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame4_bit7/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG1_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame2_bit8_GATE input94/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix__104_ Inst_LUT4AB_switch_matrix__104_/A vssd1 vssd1 vccd1
+ vccd1 output471/A sky130_fd_sc_hd__clkbuf_1
XInst_LUT4AB_switch_matrix__035_ Inst_LUT4AB_switch_matrix__035_/A vssd1 vssd1 vccd1
+ vccd1 output254/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG7_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_AB__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame19_bit8_D input80/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1_A1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LB_I1/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG1_cus_mux41_buf_inst0_A0
+ input102/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame11_bit4 input76/X input84/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame11_bit4/Q Inst_LUT4AB_ConfigMem_Inst_Frame11_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_SS4BEG_outbuf_5__0__A SS4END_inbuf_5__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J_l_EF_BEG2_A1 input197/X vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG5_cus_mux41_buf_inst2_A3
+ Inst_LUT4AB_switch_matrix__036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame7_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit28 input70/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit28/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XInst_LUT4AB_ConfigMem_Inst_Frame7_bit17 input58/X input99/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame7_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame7_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame8_bit5 input77/X input100/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame8_bit5/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix__073__A input114/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_MUX8LUT_frame_config_mux_cus_mux21_EH__0_ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_GH__0_/X Inst_MUX8LUT_frame_config_mux_cus_mux21_EH__0_/S
+ vssd1 vssd1 vccd1 vccd1 Inst_MUX8LUT_frame_config_mux_cus_mux21_EH__0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr_cus_mux21_I0mux__0_ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I0/X
+ Inst_LUT4AB_switch_matrix__064_/X Inst_LUT4AB_ConfigMem_Inst_Frame12_bit18/Q vssd1
+ vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__07_/A sky130_fd_sc_hd__mux2_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_AB_BEG0_A2 input199/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit16 input57/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LUT4AB_ConfigMem_Inst_Frame10_bit27 input69/X input83/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame10_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame10_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame10_bit12_GATE input83/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame13_bit21_GATE input86/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit30_GATE input89/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XNN4BEG_outbuf_7__0_ NN4END_inbuf_7__0_/X vssd1 vssd1 vccd1 vccd1 output404/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_EFb_BEG1_A2 input169/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LH_LUT4c_frame_config_dffesr__09_ Inst_LH_LUT4c_frame_config_dffesr__09_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LH_LUT4c_frame_config_dffesr__09_/Y sky130_fd_sc_hd__inv_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2MID_CDa_BEG0_A2 input224/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG6_cus_mux41_buf_inst2_A1
+ Inst_LUT4AB_switch_matrix__033_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit26_D input68/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_47_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame11_bit21_D input63/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst4 Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst0/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst1/X Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst2/X
+ Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG6_cus_mux41_buf_inst3/X Inst_LUT4AB_ConfigMem_Inst_Frame3_bit13/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit12/Q vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix__071_/A
+ sky130_fd_sc_hd__mux4_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit12 input53/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit12/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LUT4AB_ConfigMem_Inst_Frame3_bit23 input65/X input95/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame3_bit23/Q Inst_LUT4AB_ConfigMem_Inst_Frame3_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG5_cus_mux41_buf_inst3_A2
+ Inst_LUT4AB_switch_matrix__056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit17_GATE input88/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame18_bit26_GATE input91/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_switch_matrix__068__A Inst_LUT4AB_switch_matrix__068_/A vssd1
+ vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S2 Inst_LUT4AB_switch_matrix__071_/A
+ Inst_LUT4AB_switch_matrix__044_/A Inst_LUT4AB_switch_matrix__087_/A ANTENNA_4/DIODE
+ Inst_LUT4AB_ConfigMem_Inst_Frame9_bit1/Q Inst_LUT4AB_ConfigMem_Inst_Frame8_bit0/Q
+ vssd1 vssd1 vccd1 vccd1 Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_S2/X sky130_fd_sc_hd__mux4_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit3_D input75/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_EE4BEG_outbuf_10__0__A EE4END_inbuf_10__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_4 ANTENNA_4/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_WW4BEG_outbuf_9__0__A WW4END_inbuf_9__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux21_LD_EN__0__A1 Inst_LUT4AB_switch_matrix_inst_cus_mux21_LH_EN__0_/A1
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JS2BEG3_cus_mux41_buf_inst2_A2
+ Inst_LUT4AB_switch_matrix__034_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_E6BEG1_cus_mux41_buf_inst3_A3
+ Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_LH_I2/A0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame16_bit7_D input79/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit0_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit27 input69/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit27/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JN2BEG3_cus_mux41_buf_inst3_A3
+ Inst_MUX8LUT_frame_config_mux_cus_mux21_EF__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame6_bit16 input57/X input98/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame6_bit16/Q Inst_LUT4AB_ConfigMem_Inst_Frame6_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame15_bit14_D input55/X vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame8_bit14_GATE input100/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
XInst_LUT4AB_ConfigMem_Inst_Frame5_bit8 input80/X input97/X vssd1 vssd1 vccd1 vccd1
+ Inst_LUT4AB_ConfigMem_Inst_Frame5_bit8/Q Inst_LUT4AB_ConfigMem_Inst_Frame5_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XInst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0 Inst_LUT4AB_ConfigMem_Inst_Frame16_bit18/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame16_bit17/Q Inst_LUT4AB_ConfigMem_Inst_Frame17_bit16/Q
+ Inst_LUT4AB_ConfigMem_Inst_Frame17_bit15/Q Inst_LD_LUT4c_frame_config_dffesr__07_/A
+ Inst_LD_LUT4c_frame_config_dffesr__08_/A vssd1 vssd1 vccd1 vccd1 Inst_LD_LUT4c_frame_config_dffesr_inst_cus_mux161_buf_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_ConfigMem_Inst_Frame0_bit23_GATE input82/X vssd1 vssd1 vccd1
+ vccd1 sky130_fd_sc_hd__diode_2
Xinput163 S2END[5] vssd1 vssd1 vccd1 vccd1 input163/X sky130_fd_sc_hd__clkbuf_4
Xinput141 NN4END[12] vssd1 vssd1 vccd1 vccd1 input141/X sky130_fd_sc_hd__clkbuf_1
Xinput152 NN4END[8] vssd1 vssd1 vccd1 vccd1 input152/X sky130_fd_sc_hd__clkbuf_1
Xinput130 N4END[2] vssd1 vssd1 vccd1 vccd1 input130/X sky130_fd_sc_hd__buf_2
Xinput185 S4END[5] vssd1 vssd1 vccd1 vccd1 input185/X sky130_fd_sc_hd__clkbuf_1
Xinput174 S4END[0] vssd1 vssd1 vccd1 vccd1 input174/X sky130_fd_sc_hd__buf_2
Xinput196 SS4END[15] vssd1 vssd1 vccd1 vccd1 input196/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JE2BEG4_cus_mux41_buf_inst2_A0
+ Inst_LUT4AB_switch_matrix__032_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XInst_LG_LUT4c_frame_config_dffesr__07_ Inst_LG_LUT4c_frame_config_dffesr__07_/A vssd1
+ vssd1 vccd1 vccd1 Inst_LG_LUT4c_frame_config_dffesr__07_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_73_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux161_buf_JW2BEG3_cus_mux41_buf_inst3_A1
+ Inst_LUT4AB_switch_matrix__055_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_S4BEG_outbuf_3__0__A S4END_inbuf_3__0_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_Inst_LUT4AB_switch_matrix_inst_cus_mux41_buf_J2END_GH_BEG1_A2 input190/X
+ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XNN4END_inbuf_4__0_ input152/X vssd1 vssd1 vccd1 vccd1 NN4END_inbuf_4__0_/X sky130_fd_sc_hd__clkbuf_4
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

