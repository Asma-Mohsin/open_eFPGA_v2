VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO BlockRAM_1KB
  CLASS BLOCK ;
  FOREIGN BlockRAM_1KB ;
  ORIGIN 0.000 0.000 ;
  SIZE 570.000 BY 450.000 ;
  PIN mem_dout\[9\]
    PORT
      LAYER met1 ;
        RECT 50.500 441.420 227.770 441.560 ;
    END
  END mem_dout\[9\]
  PIN _017_
    PORT
      LAYER met1 ;
        RECT 47.080 341.615 47.220 341.940 ;
    END
  END _017_
  PIN _021_
    PORT
      LAYER met1 ;
        RECT 49.380 352.000 49.520 352.325 ;
    END
  END _021_
  PIN _023_
    PORT
      LAYER met1 ;
        RECT 46.620 335.340 46.760 336.005 ;
    END
  END _023_
  PIN _024_
    PORT
      LAYER met1 ;
        RECT 30.675 336.700 39.200 336.840 ;
    END
  END _024_
  PIN _037_
    PORT
      LAYER met1 ;
        RECT 50.760 352.340 51.205 352.480 ;
    END
  END _037_
  PIN _038_
    PORT
      LAYER met1 ;
        RECT 47.540 343.160 47.680 343.825 ;
    END
  END _038_
  PIN _039_
    PORT
      LAYER met1 ;
        RECT 44.520 343.160 45.225 343.300 ;
    END
  END _039_
  PIN _040_
    PORT
      LAYER met1 ;
        RECT 51.680 352.340 54.425 352.480 ;
    END
  END _040_
  PIN _041_
    PORT
      LAYER met1 ;
        RECT 55.820 352.000 55.960 352.325 ;
    END
  END _041_
  PIN _049_
    PORT
      LAYER met1 ;
        RECT 48.460 347.070 48.600 347.720 ;
    END
  END _049_
  PIN _058_
    PORT
      LAYER met1 ;
        RECT 48.660 353.020 52.125 353.160 ;
    END
  END _058_
  PIN _060_
    PORT
      LAYER met1 ;
        RECT 39.000 359.820 45.380 359.960 ;
    END
  END _060_
  PIN _066_
    PORT
      LAYER met1 ;
        RECT 48.000 352.495 48.140 353.160 ;
    END
  END _066_
  PIN _074_
    PORT
      LAYER met1 ;
        RECT 45.855 336.020 46.100 336.160 ;
    END
  END _074_
  PIN _076_
    PORT
      LAYER met1 ;
        RECT 53.675 351.660 57.600 351.800 ;
    END
  END _076_
  PIN _096_
    PORT
      LAYER met1 ;
        RECT 54.640 357.100 56.420 357.240 ;
    END
  END _096_
  PIN _104_
    PORT
      LAYER met1 ;
        RECT 29.800 370.360 47.220 370.500 ;
    END
  END _104_
  PIN _127_
    PORT
      LAYER met1 ;
        RECT 54.900 366.095 55.040 366.760 ;
    END
  END _127_
  PIN _128_
    PORT
      LAYER met1 ;
        RECT 21.980 353.020 41.545 353.160 ;
    END
  END _128_
  PIN _129_
    PORT
      LAYER met1 ;
        RECT 33.020 354.040 40.165 354.180 ;
    END
  END _129_
  PIN _130_
    PORT
      LAYER met1 ;
        RECT 22.440 359.480 44.765 359.620 ;
    END
  END _130_
  PIN _131_
    PORT
      LAYER met1 ;
        RECT 21.520 362.200 45.685 362.340 ;
    END
  END _131_
  PIN _132_
    PORT
      LAYER met1 ;
        RECT 27.040 364.920 46.760 365.060 ;
    END
  END _132_
  PIN mem_dout\[4\]
    PORT
      LAYER met1 ;
        RECT 67.320 339.420 67.460 339.700 ;
    END
  END mem_dout\[4\]
  PIN mem_dout\[5\]
    PORT
      LAYER met1 ;
        RECT 53.215 433.600 70.680 433.740 ;
    END
  END mem_dout\[5\]
  PIN mem_dout\[7\]
    PORT
      LAYER met1 ;
        RECT 56.435 431.560 59.440 431.700 ;
    END
  END mem_dout\[7\]
  PIN _014_
    PORT
      LAYER met1 ;
        RECT 41.560 346.560 41.700 346.885 ;
    END
  END _014_
  PIN net38
    PORT
      LAYER met1 ;
        RECT 8.595 389.740 10.680 389.880 ;
    END
  END net38
  PIN net40
    PORT
      LAYER met1 ;
        RECT 8.135 400.280 11.600 400.420 ;
    END
  END net40
  PIN net42
    PORT
      LAYER met1 ;
        RECT 8.595 408.780 10.220 408.920 ;
    END
  END net42
  PIN net44
    PORT
      LAYER met1 ;
        RECT 8.595 419.660 12.060 419.800 ;
    END
  END net44
  PIN net46
    PORT
      LAYER met1 ;
        RECT 8.595 422.380 11.140 422.520 ;
    END
  END net46
  PIN net47
    PORT
      LAYER met1 ;
        RECT 8.595 427.820 9.760 427.960 ;
    END
  END net47
  PIN rd_dout_additional_register\[27\]
    PORT
      LAYER met1 ;
        RECT 42.635 354.040 43.540 354.180 ;
    END
  END rd_dout_additional_register\[27\]
  PIN rd_dout_additional_register\[29\]
    PORT
      LAYER met1 ;
        RECT 48.155 363.900 52.080 364.040 ;
    END
  END rd_dout_additional_register\[29\]
  PIN _064_
    PORT
      LAYER met1 ;
        RECT 50.300 281.280 54.380 281.420 ;
    END
  END _064_
  PIN _007_
    PORT
      LAYER met1 ;
        RECT 38.800 332.620 41.085 332.760 ;
    END
  END _007_
  PIN _070_
    PORT
      LAYER met1 ;
        RECT 52.140 238.255 52.280 238.580 ;
    END
  END _070_
  PIN _008_
    PORT
      LAYER met1 ;
        RECT 42.175 333.300 49.780 333.440 ;
    END
  END _008_
  PIN _075_
    PORT
      LAYER met1 ;
        RECT 47.145 319.770 47.155 319.780 ;
    END
  END _075_
  PIN _011_
    PORT
      LAYER met1 ;
        RECT 42.175 276.180 42.620 276.320 ;
    END
  END _011_
  PIN _078_
    PORT
      LAYER met1 ;
        RECT 30.675 240.480 31.120 240.620 ;
    END
  END _078_
  PIN _080_
    PORT
      LAYER met1 ;
        RECT 48.155 273.120 50.700 273.260 ;
    END
  END _080_
  PIN _082_
    PORT
      LAYER met1 ;
        RECT 43.600 314.940 43.845 315.080 ;
    END
  END _082_
  PIN _083_
    PORT
      LAYER met1 ;
        RECT 52.800 311.200 53.040 311.340 ;
    END
  END _083_
  PIN _084_
    PORT
      LAYER met1 ;
        RECT 52.140 311.540 53.505 311.680 ;
    END
  END _084_
  PIN _086_
    PORT
      LAYER met1 ;
        RECT 30.215 232.660 31.120 232.800 ;
    END
  END _086_
  PIN _088_
    PORT
      LAYER met1 ;
        RECT 47.540 273.460 53.460 273.600 ;
    END
  END _088_
  PIN _090_
    PORT
      LAYER met1 ;
        RECT 49.120 314.940 54.885 315.080 ;
    END
  END _090_
  PIN _092_
    PORT
      LAYER met1 ;
        RECT 52.140 309.500 53.920 309.640 ;
    END
  END _092_
  PIN _094_
    PORT
      LAYER met1 ;
        RECT 31.640 240.480 31.885 240.620 ;
    END
  END _094_
  PIN _025_
    PORT
      LAYER met1 ;
        RECT 51.680 319.855 51.820 320.320 ;
    END
  END _025_
  PIN _098_
    PORT
      LAYER met1 ;
        RECT 62.030 289.100 62.660 289.240 ;
    END
  END _098_
  PIN _100_
    PORT
      LAYER met1 ;
        RECT 51.220 289.100 58.980 289.240 ;
    END
  END _100_
  PIN _026_
    PORT
      LAYER met1 ;
        RECT 44.320 276.520 44.460 276.845 ;
    END
  END _026_
  PIN _111_
    PORT
      LAYER met1 ;
        RECT 62.030 286.720 63.580 286.860 ;
    END
  END _111_
  PIN _113_
    PORT
      LAYER met1 ;
        RECT 51.835 281.620 58.060 281.760 ;
    END
  END _113_
  PIN _115_
    PORT
      LAYER met1 ;
        RECT 54.900 294.540 55.040 295.205 ;
    END
  END _115_
  PIN _116_
    PORT
      LAYER met1 ;
        RECT 22.855 265.300 32.960 265.440 ;
    END
  END _116_
  PIN _117_
    PORT
      LAYER met1 ;
        RECT 23.315 270.740 37.560 270.880 ;
    END
  END _117_
  PIN _118_
    PORT
      LAYER met1 ;
        RECT 16.260 279.240 28.160 279.380 ;
    END
  END _118_
  PIN _119_
    PORT
      LAYER met1 ;
        RECT 19.940 278.900 27.700 279.040 ;
    END
  END _119_
  PIN _120_
    PORT
      LAYER met1 ;
        RECT 16.720 286.380 37.820 286.520 ;
    END
  END _120_
  PIN _122_
    PORT
      LAYER met1 ;
        RECT 18.255 287.060 27.240 287.200 ;
    END
  END _122_
  PIN _123_
    PORT
      LAYER met1 ;
        RECT 24.235 278.560 36.900 278.700 ;
    END
  END _123_
  PIN _124_
    PORT
      LAYER met1 ;
        RECT 23.775 284.000 38.480 284.140 ;
    END
  END _124_
  PIN _125_
    PORT
      LAYER met1 ;
        RECT 20.140 329.900 36.180 330.040 ;
    END
  END _125_
  PIN _126_
    PORT
      LAYER met1 ;
        RECT 23.775 300.320 26.780 300.460 ;
    END
  END _126_
  PIN _027_
    PORT
      LAYER met1 ;
        RECT 50.300 319.020 50.440 319.685 ;
    END
  END _027_
  PIN _029_
    PORT
      LAYER met1 ;
        RECT 43.860 229.755 44.000 230.760 ;
    END
  END _029_
  PIN _032_
    PORT
      LAYER met1 ;
        RECT 45.240 283.320 45.380 283.645 ;
    END
  END _032_
  PIN _012_
    PORT
      LAYER met1 ;
        RECT 53.520 314.415 53.660 314.740 ;
    END
  END _012_
  PIN _013_
    PORT
      LAYER met1 ;
        RECT 40.840 314.260 41.085 314.400 ;
    END
  END _013_
  PIN _005_
    PORT
      LAYER met1 ;
        RECT 30.675 238.780 42.880 238.920 ;
    END
  END _005_
  PIN _133_
    PORT
      LAYER met1 ;
        RECT 22.240 300.475 22.380 300.800 ;
    END
  END _133_
  PIN clknet_2_0__leaf_clk
    PORT
      LAYER met1 ;
        RECT 45.700 292.655 45.840 292.980 ;
    END
  END clknet_2_0__leaf_clk
  PIN clknet_2_3__leaf_clk
    PORT
      LAYER met1 ;
        RECT 41.760 262.920 55.805 263.060 ;
    END
  END clknet_2_3__leaf_clk
  PIN mem_dout\[23\]
    PORT
      LAYER met1 ;
        RECT 65.480 315.960 65.620 316.580 ;
    END
  END mem_dout\[23\]
  PIN _015_
    PORT
      LAYER met1 ;
        RECT 36.960 316.640 39.705 316.780 ;
    END
  END _015_
  PIN _016_
    PORT
      LAYER met1 ;
        RECT 44.320 324.800 45.685 324.940 ;
    END
  END _016_
  PIN _042_
    PORT
      LAYER met1 ;
        RECT 28.880 268.700 30.045 268.840 ;
    END
  END _042_
  PIN _047_
    PORT
      LAYER met1 ;
        RECT 47.540 281.960 60.820 282.100 ;
    END
  END _047_
  PIN net16
    PORT
      LAYER met1 ;
        RECT 8.440 324.120 8.580 325.125 ;
    END
  END net16
  PIN net29
    PORT
      LAYER met1 ;
        RECT 8.135 228.920 9.760 229.060 ;
    END
  END net29
  PIN _006_
    PORT
      LAYER met1 ;
        RECT 47.280 281.280 49.365 281.420 ;
    END
  END _006_
  PIN net39
    PORT
      LAYER met1 ;
        RECT 43.050 287.060 46.760 287.200 ;
    END
  END net39
  PIN _050_
    PORT
      LAYER met1 ;
        RECT 55.420 322.145 55.430 322.155 ;
    END
  END _050_
  PIN _051_
    PORT
      LAYER met1 ;
        RECT 55.975 322.420 60.360 322.560 ;
    END
  END _051_
  PIN _053_
    PORT
      LAYER met1 ;
        RECT 33.435 240.480 36.440 240.620 ;
    END
  END _053_
  PIN _018_
    PORT
      LAYER met1 ;
        RECT 51.280 319.795 51.290 319.805 ;
    END
  END _018_
  PIN _059_
    PORT
      LAYER met1 ;
        RECT 46.680 327.585 46.690 327.595 ;
    END
  END _059_
  PIN net6
    PORT
      LAYER met1 ;
        RECT 32.100 281.960 32.345 282.100 ;
    END
  END net6
  PIN net62
    PORT
      LAYER met1 ;
        RECT 21.520 264.280 21.765 264.420 ;
    END
  END net62
  PIN net63
    PORT
      LAYER met1 ;
        RECT 7.675 238.440 22.180 238.580 ;
    END
  END net63
  PIN net65
    PORT
      LAYER met1 ;
        RECT 7.675 249.320 18.960 249.460 ;
    END
  END net65
  PIN net67
    PORT
      LAYER met1 ;
        RECT 14.160 286.040 15.785 286.180 ;
    END
  END net67
  PIN net70
    PORT
      LAYER met1 ;
        RECT 7.675 267.680 13.440 267.820 ;
    END
  END net70
  PIN net73
    PORT
      LAYER met1 ;
        RECT 7.675 281.960 12.980 282.100 ;
    END
  END net73
  PIN net74
    PORT
      LAYER met1 ;
        RECT 7.675 287.400 21.260 287.540 ;
    END
  END net74
  PIN net75
    PORT
      LAYER met1 ;
        RECT 7.675 289.440 22.180 289.580 ;
    END
  END net75
  PIN net76
    PORT
      LAYER met1 ;
        RECT 7.675 294.880 23.100 295.020 ;
    END
  END net76
  PIN net78
    PORT
      LAYER met1 ;
        RECT 7.520 300.475 7.660 300.800 ;
    END
  END net78
  PIN rd_dout_additional_register\[16\]
    PORT
      LAYER met1 ;
        RECT 51.880 295.220 54.425 295.360 ;
    END
  END rd_dout_additional_register\[16\]
  PIN rd_dout_additional_register\[17\]
    PORT
      LAYER met1 ;
        RECT 43.555 303.380 50.240 303.520 ;
    END
  END rd_dout_additional_register\[17\]
  PIN rd_dout_additional_register\[18\]
    PORT
      LAYER met1 ;
        RECT 38.035 314.940 39.200 315.080 ;
    END
  END rd_dout_additional_register\[18\]
  PIN rd_dout_additional_register\[19\]
    PORT
      LAYER met1 ;
        RECT 39.000 309.500 42.005 309.640 ;
    END
  END rd_dout_additional_register\[19\]
  PIN rd_dout_additional_register\[20\]
    PORT
      LAYER met1 ;
        RECT 38.540 322.420 38.785 322.560 ;
    END
  END rd_dout_additional_register\[20\]
  PIN rd_dout_additional_register\[22\]
    PORT
      LAYER met1 ;
        RECT 45.900 295.900 51.665 296.040 ;
    END
  END rd_dout_additional_register\[22\]
  PIN rd_dout_additional_register\[24\]
    PORT
      LAYER met1 ;
        RECT 38.495 330.920 39.660 331.060 ;
    END
  END rd_dout_additional_register\[24\]
  PIN rd_dout_additional_register\[25\]
    PORT
      LAYER met1 ;
        RECT 40.840 327.860 41.545 328.000 ;
    END
  END rd_dout_additional_register\[25\]
  PIN _019_
    PORT
      LAYER met1 ;
        RECT 41.560 319.020 41.700 319.640 ;
    END
  END _019_
  PIN _062_
    PORT
      LAYER met1 ;
        RECT 37.115 240.480 39.200 240.620 ;
    END
  END _062_
  PIN rd_dout_additional_register\[31\]
    PORT
      LAYER met1 ;
        RECT 49.580 293.180 52.585 293.320 ;
    END
  END rd_dout_additional_register\[31\]
  PIN rd_dout_muxed\[11\]
    PORT
      LAYER met1 ;
        RECT 46.270 240.480 53.000 240.620 ;
    END
  END rd_dout_muxed\[11\]
  PIN rd_dout_muxed\[14\]
    PORT
      LAYER met1 ;
        RECT 49.995 286.040 53.920 286.180 ;
    END
  END rd_dout_muxed\[14\]
  PIN rd_dout_muxed\[15\]
    PORT
      LAYER met1 ;
        RECT 46.270 235.040 52.540 235.180 ;
    END
  END rd_dout_muxed\[15\]
  PIN rd_dout_muxed\[2\]
    PORT
      LAYER met1 ;
        RECT 29.250 234.700 32.300 234.840 ;
    END
  END rd_dout_muxed\[2\]
  PIN rd_dout_muxed\[3\]
    PORT
      LAYER met1 ;
        RECT 33.390 232.660 36.640 232.800 ;
    END
  END rd_dout_muxed\[3\]
  PIN rd_dout_muxed\[4\]
    PORT
      LAYER met1 ;
        RECT 44.430 233.000 47.480 233.140 ;
    END
  END rd_dout_muxed\[4\]
  PIN rd_dout_muxed\[5\]
    PORT
      LAYER met1 ;
        RECT 28.330 229.260 29.540 229.400 ;
    END
  END rd_dout_muxed\[5\]
  PIN rd_dout_muxed\[7\]
    PORT
      LAYER met1 ;
        RECT 35.690 229.600 37.360 229.740 ;
    END
  END rd_dout_muxed\[7\]
  PIN rd_dout_muxed\[8\]
    PORT
      LAYER met1 ;
        RECT 43.050 238.100 44.260 238.240 ;
    END
  END rd_dout_muxed\[8\]
  PIN rd_dout_sel\[0\]
    PORT
      LAYER met1 ;
        RECT 33.480 286.040 48.445 286.180 ;
    END
  END rd_dout_sel\[0\]
  PIN rd_dout_sel\[1\]
    PORT
      LAYER met1 ;
        RECT 32.975 317.320 34.140 317.460 ;
    END
  END rd_dout_sel\[1\]
  PIN _148_
    PORT
      LAYER met1 ;
        RECT 28.880 189.820 30.000 189.960 ;
    END
  END _148_
  PIN _150_
    PORT
      LAYER met1 ;
        RECT 51.220 194.580 52.125 194.720 ;
    END
  END _150_
  PIN _151_
    PORT
      LAYER met1 ;
        RECT 46.775 196.280 48.860 196.420 ;
    END
  END _151_
  PIN _152_
    PORT
      LAYER met1 ;
        RECT 43.140 200.360 46.975 200.500 ;
    END
  END _152_
  PIN _153_
    PORT
      LAYER met1 ;
        RECT 53.060 202.740 65.420 202.880 ;
    END
  END _153_
  PIN _155_
    PORT
      LAYER met1 ;
        RECT 49.535 209.880 59.440 210.020 ;
    END
  END _155_
  PIN _156_
    PORT
      LAYER met1 ;
        RECT 48.660 212.600 49.735 212.740 ;
    END
  END _156_
  PIN _157_
    PORT
      LAYER met1 ;
        RECT 52.295 185.740 52.540 185.880 ;
    END
  END _157_
  PIN _158_
    PORT
      LAYER met1 ;
        RECT 49.995 204.440 65.880 204.580 ;
    END
  END _158_
  PIN _161_
    PORT
      LAYER met1 ;
        RECT 50.040 184.380 66.340 184.520 ;
    END
  END _161_
  PIN _162_
    PORT
      LAYER met1 ;
        RECT 53.625 185.400 67.720 185.540 ;
    END
  END _162_
  PIN _167_
    PORT
      LAYER met1 ;
        RECT 33.940 142.560 46.605 142.700 ;
    END
  END _167_
  PIN _169_
    PORT
      LAYER met1 ;
        RECT 43.600 142.220 45.225 142.360 ;
    END
  END _169_
  PIN _089_
    PORT
      LAYER met1 ;
        RECT 23.820 203.080 24.985 203.220 ;
    END
  END _089_
  PIN _010_
    PORT
      LAYER met1 ;
        RECT 33.895 189.140 34.140 189.280 ;
    END
  END _010_
  PIN _093_
    PORT
      LAYER met1 ;
        RECT 23.160 202.740 25.445 202.880 ;
    END
  END _093_
  PIN _095_
    PORT
      LAYER met1 ;
        RECT 26.075 202.400 27.240 202.540 ;
    END
  END _095_
  PIN _061_
    PORT
      LAYER met1 ;
        RECT 32.820 199.000 32.960 199.480 ;
    END
  END _061_
  PIN muxedDataIn\[10\]
    PORT
      LAYER met1 ;
        RECT 50.960 184.040 60.820 184.180 ;
    END
  END muxedDataIn\[10\]
  PIN muxedDataIn\[11\]
    PORT
      LAYER met1 ;
        RECT 55.975 186.420 57.600 186.560 ;
    END
  END muxedDataIn\[11\]
  PIN muxedDataIn\[12\]
    PORT
      LAYER met1 ;
        RECT 51.680 193.900 53.000 194.040 ;
    END
  END muxedDataIn\[12\]
  PIN muxedDataIn\[13\]
    PORT
      LAYER met1 ;
        RECT 53.215 197.300 61.280 197.440 ;
    END
  END muxedDataIn\[13\]
  PIN muxedDataIn\[14\]
    PORT
      LAYER met1 ;
        RECT 55.820 193.900 60.360 194.040 ;
    END
  END muxedDataIn\[14\]
  PIN net1
    PORT
      LAYER met1 ;
        RECT 36.700 140.180 40.625 140.320 ;
    END
  END net1
  PIN _001_
    PORT
      LAYER met1 ;
        RECT 45.395 143.240 47.020 143.380 ;
    END
  END _001_
  PIN net24
    PORT
      LAYER met1 ;
        RECT 8.135 204.440 38.740 204.580 ;
    END
  END net24
  PIN net25
    PORT
      LAYER met1 ;
        RECT 8.135 209.880 10.680 210.020 ;
    END
  END net25
  PIN net26
    PORT
      LAYER met1 ;
        RECT 8.135 212.600 11.140 212.740 ;
    END
  END net26
  PIN net27
    PORT
      LAYER met1 ;
        RECT 8.135 218.040 11.600 218.180 ;
    END
  END net27
  PIN net28
    PORT
      LAYER met1 ;
        RECT 17.380 162.620 46.145 162.760 ;
    END
  END net28
  PIN _099_
    PORT
      LAYER met1 ;
        RECT 16.260 137.275 16.400 137.600 ;
    END
  END _099_
  PIN net30
    PORT
      LAYER met1 ;
        RECT 41.760 184.040 43.340 184.180 ;
    END
  END net30
  PIN net32
    PORT
      LAYER met1 ;
        RECT 42.220 200.700 49.365 200.840 ;
    END
  END net32
  PIN net33
    PORT
      LAYER met1 ;
        RECT 17.840 203.420 34.570 203.560 ;
    END
  END net33
  PIN _063_
    PORT
      LAYER met1 ;
        RECT 30.520 200.175 30.660 200.500 ;
    END
  END _063_
  PIN _103_
    PORT
      LAYER met1 ;
        RECT 15.495 145.620 16.660 145.760 ;
    END
  END _103_
  PIN _028_
    PORT
      LAYER met1 ;
        RECT 34.355 188.460 54.380 188.600 ;
    END
  END _028_
  PIN _106_
    PORT
      LAYER met1 ;
        RECT 19.635 148.000 20.800 148.140 ;
    END
  END _106_
  PIN _110_
    PORT
      LAYER met1 ;
        RECT 19.220 219.400 40.165 219.540 ;
    END
  END _110_
  PIN _065_
    PORT
      LAYER met1 ;
        RECT 33.740 199.680 33.880 200.005 ;
    END
  END _065_
  PIN _112_
    PORT
      LAYER met1 ;
        RECT 17.180 151.215 17.320 151.540 ;
    END
  END _112_
  PIN net5
    PORT
      LAYER met1 ;
        RECT 21.980 222.120 30.200 222.260 ;
    END
  END net5
  PIN net53
    PORT
      LAYER met1 ;
        RECT 8.135 193.560 17.580 193.700 ;
    END
  END net53
  PIN net54
    PORT
      LAYER met1 ;
        RECT 8.135 200.700 9.300 200.840 ;
    END
  END net54
  PIN _114_
    PORT
      LAYER met1 ;
        RECT 19.175 156.500 19.420 156.640 ;
    END
  END _114_
  PIN _069_
    PORT
      LAYER met1 ;
        RECT 34.355 199.340 47.940 199.480 ;
    END
  END _069_
  PIN _045_
    PORT
      LAYER met1 ;
        RECT 32.975 227.220 37.100 227.360 ;
    END
  END _045_
  PIN _071_
    PORT
      LAYER met1 ;
        RECT 34.660 200.175 34.800 200.500 ;
    END
  END _071_
  PIN _073_
    PORT
      LAYER met1 ;
        RECT 28.680 202.740 30.460 202.880 ;
    END
  END _073_
  PIN _046_
    PORT
      LAYER met1 ;
        RECT 31.440 191.180 31.580 191.505 ;
    END
  END _046_
  PIN _030_
    PORT
      LAYER met1 ;
        RECT 31.900 205.615 32.040 205.940 ;
    END
  END _030_
  PIN _048_
    PORT
      LAYER met1 ;
        RECT 30.980 197.115 31.120 197.440 ;
    END
  END _048_
  PIN _079_
    PORT
      LAYER met1 ;
        RECT 29.755 202.400 30.920 202.540 ;
    END
  END _079_
  PIN rd_dout_additional_register\[0\]
    PORT
      LAYER met1 ;
        RECT 37.115 208.860 42.880 209.000 ;
    END
  END rd_dout_additional_register\[0\]
  PIN rd_dout_additional_register\[10\]
    PORT
      LAYER met1 ;
        RECT 33.480 222.460 34.185 222.600 ;
    END
  END rd_dout_additional_register\[10\]
  PIN rd_dout_additional_register\[11\]
    PORT
      LAYER met1 ;
        RECT 47.235 218.720 49.520 218.860 ;
    END
  END rd_dout_additional_register\[11\]
  PIN rd_dout_additional_register\[12\]
    PORT
      LAYER met1 ;
        RECT 41.715 222.460 50.240 222.600 ;
    END
  END rd_dout_additional_register\[12\]
  PIN rd_dout_additional_register\[13\]
    PORT
      LAYER met1 ;
        RECT 42.635 218.380 49.980 218.520 ;
    END
  END rd_dout_additional_register\[13\]
  PIN rd_dout_additional_register\[14\]
    PORT
      LAYER met1 ;
        RECT 42.175 211.580 48.860 211.720 ;
    END
  END rd_dout_additional_register\[14\]
  PIN rd_dout_additional_register\[15\]
    PORT
      LAYER met1 ;
        RECT 47.235 213.280 51.820 213.420 ;
    END
  END rd_dout_additional_register\[15\]
  PIN _033_
    PORT
      LAYER met1 ;
        RECT 35.580 207.500 35.720 207.825 ;
    END
  END _033_
  PIN _081_
    PORT
      LAYER met1 ;
        RECT 24.080 199.680 25.905 199.820 ;
    END
  END _081_
  PIN _034_
    PORT
      LAYER met1 ;
        RECT 34.815 189.140 37.820 189.280 ;
    END
  END _034_
  PIN _052_
    PORT
      LAYER met1 ;
        RECT 31.595 197.640 40.120 197.780 ;
    END
  END _052_
  PIN rd_dout_additional_register\[1\]
    PORT
      LAYER met1 ;
        RECT 29.295 208.860 34.140 209.000 ;
    END
  END rd_dout_additional_register\[1\]
  PIN _036_
    PORT
      LAYER met1 ;
        RECT 30.520 191.675 30.660 192.000 ;
    END
  END _036_
  PIN _085_
    PORT
      LAYER met1 ;
        RECT 22.240 199.340 26.365 199.480 ;
    END
  END _085_
  PIN _054_
    PORT
      LAYER met1 ;
        RECT 32.820 216.495 32.960 217.160 ;
    END
  END _054_
  PIN _087_
    PORT
      LAYER met1 ;
        RECT 27.040 212.600 28.205 212.740 ;
    END
  END _087_
  PIN _055_
    PORT
      LAYER met1 ;
        RECT 31.640 196.960 31.885 197.100 ;
    END
  END _055_
  PIN rd_dout_additional_register\[2\]
    PORT
      LAYER met1 ;
        RECT 30.060 215.475 30.200 215.800 ;
    END
  END rd_dout_additional_register\[2\]
  PIN rd_dout_additional_register\[3\]
    PORT
      LAYER met1 ;
        RECT 31.135 219.740 38.740 219.880 ;
    END
  END rd_dout_additional_register\[3\]
  PIN rd_dout_additional_register\[4\]
    PORT
      LAYER met1 ;
        RECT 34.355 215.320 34.800 215.460 ;
    END
  END rd_dout_additional_register\[4\]
  PIN rd_dout_additional_register\[6\]
    PORT
      LAYER met1 ;
        RECT 27.455 214.300 29.540 214.440 ;
    END
  END rd_dout_additional_register\[6\]
  PIN rd_dout_additional_register\[7\]
    PORT
      LAYER met1 ;
        RECT 26.840 215.475 26.980 216.140 ;
    END
  END rd_dout_additional_register\[7\]
  PIN rd_dout_additional_register\[8\]
    PORT
      LAYER met1 ;
        RECT 34.355 211.240 49.520 211.380 ;
    END
  END rd_dout_additional_register\[8\]
  PIN rd_dout_additional_register\[9\]
    PORT
      LAYER met1 ;
        RECT 32.975 207.840 35.260 207.980 ;
    END
  END rd_dout_additional_register\[9\]
  PIN rd_dout_muxed\[0\]
    PORT
      LAYER met1 ;
        RECT 43.140 222.120 44.610 222.260 ;
    END
  END rd_dout_muxed\[0\]
  PIN _136_
    PORT
      LAYER met1 ;
        RECT 46.315 150.040 46.560 150.180 ;
    END
  END _136_
  PIN _137_
    PORT
      LAYER met1 ;
        RECT 49.840 145.620 56.680 145.760 ;
    END
  END _137_
  PIN _138_
    PORT
      LAYER met1 ;
        RECT 55.360 134.895 55.500 135.560 ;
    END
  END _138_
  PIN rd_dout_muxed\[1\]
    PORT
      LAYER met1 ;
        RECT 32.100 223.820 35.410 223.960 ;
    END
  END rd_dout_muxed\[1\]
  PIN _139_
    PORT
      LAYER met1 ;
        RECT 56.895 131.680 57.140 131.820 ;
    END
  END _139_
  PIN _140_
    PORT
      LAYER met1 ;
        RECT 48.200 137.120 53.505 137.260 ;
    END
  END _140_
  PIN _141_
    PORT
      LAYER met1 ;
        RECT 56.280 142.715 56.420 143.720 ;
    END
  END _141_
  PIN _142_
    PORT
      LAYER met1 ;
        RECT 47.540 136.780 56.265 136.920 ;
    END
  END _142_
  PIN rd_dout_muxed\[6\]
    PORT
      LAYER met1 ;
        RECT 28.330 223.820 29.080 223.960 ;
    END
  END rd_dout_muxed\[6\]
  PIN _143_
    PORT
      LAYER met1 ;
        RECT 50.500 145.960 54.885 146.100 ;
    END
  END _143_
  PIN _144_
    PORT
      LAYER met1 ;
        RECT 44.475 183.020 50.700 183.160 ;
    END
  END _144_
  PIN rd_dout_muxed\[9\]
    PORT
      LAYER met1 ;
        RECT 42.220 227.220 42.825 227.360 ;
    END
  END rd_dout_muxed\[9\]
  PIN _145_
    PORT
      LAYER met1 ;
        RECT 40.795 139.160 49.780 139.300 ;
    END
  END _145_
  PIN _146_
    PORT
      LAYER met1 ;
        RECT 50.915 131.340 54.380 131.480 ;
    END
  END _146_
  PIN _003_
    PORT
      LAYER met1 ;
        RECT 52.295 110.600 53.000 110.740 ;
    END
  END _003_
  PIN _134_
    PORT
      LAYER met1 ;
        RECT 44.935 118.420 47.680 118.560 ;
    END
  END _134_
  PIN net77
    PORT
      LAYER met1 ;
        RECT 7.675 33.760 29.540 33.900 ;
    END
  END net77
  PIN _135_
    PORT
      LAYER met1 ;
        RECT 52.800 115.360 56.725 115.500 ;
    END
  END _135_
  PIN _004_
    PORT
      LAYER met1 ;
        RECT 53.260 23.220 89.845 23.360 ;
    END
  END _004_
  PIN net80
    PORT
      LAYER met1 ;
        RECT 7.720 47.360 28.160 47.500 ;
    END
  END net80
  PIN net82
    PORT
      LAYER met1 ;
        RECT 7.675 48.040 20.340 48.180 ;
    END
  END net82
  PIN net84
    PORT
      LAYER met1 ;
        RECT 7.675 58.920 23.560 59.060 ;
    END
  END net84
  PIN net85
    PORT
      LAYER met1 ;
        RECT 7.675 60.960 17.120 61.100 ;
    END
  END net85
  PIN net55
    PORT
      LAYER met1 ;
        RECT 7.675 22.880 8.840 23.020 ;
    END
  END net55
  PIN net57
    PORT
      LAYER met1 ;
        RECT 7.675 77.280 10.680 77.420 ;
    END
  END net57
  PIN net58
    PORT
      LAYER met1 ;
        RECT 7.675 80.680 21.260 80.820 ;
    END
  END net58
  PIN net59
    PORT
      LAYER met1 ;
        RECT 7.675 86.120 10.220 86.260 ;
    END
  END net59
  PIN _002_
    PORT
      LAYER met1 ;
        RECT 65.220 22.880 91.225 23.020 ;
    END
  END _002_
  PIN net60
    PORT
      LAYER met1 ;
        RECT 7.675 91.560 11.600 91.700 ;
    END
  END net60
  PIN net61
    PORT
      LAYER met1 ;
        RECT 7.675 97.000 19.880 97.140 ;
    END
  END net61
  PIN _170_
    PORT
      LAYER met1 ;
        RECT 51.375 111.960 56.680 112.100 ;
    END
  END _170_
  PIN _000_
    PORT
      LAYER met1 ;
        RECT 50.960 60.620 54.580 60.760 ;
    END
  END _000_
  PIN _171_
    PORT
      LAYER met1 ;
        RECT 45.855 117.400 49.780 117.540 ;
    END
  END _171_
  PIN net66
    PORT
      LAYER met1 ;
        RECT 7.675 28.320 18.040 28.460 ;
    END
  END net66
  PIN _147_
    PORT
      LAYER met1 ;
        RECT 63.840 29.680 70.480 29.820 ;
    END
  END _147_
  PIN net3
    PORT
      LAYER met1 ;
        RECT 8.135 109.240 9.300 109.380 ;
    END
  END net3
  PIN mem_wr_mask\[0\]
    PORT
      LAYER met1 ;
        RECT 58.275 60.280 60.820 60.420 ;
    END
  END mem_wr_mask\[0\]
  PIN net2
    PORT
      LAYER met1 ;
        RECT 41.760 118.080 43.800 118.220 ;
    END
  END net2
  PIN _154_
    PORT
      LAYER met1 ;
        RECT 64.300 58.580 67.260 58.720 ;
    END
  END _154_
  PIN net9
    PORT
      LAYER met1 ;
        RECT 39.000 13.020 559.000 13.160 ;
    END
  END net9
  PIN muxedDataIn\[26\]
    PORT
      LAYER met1 ;
        RECT 165.915 23.900 166.160 24.040 ;
    END
  END muxedDataIn\[26\]
  PIN muxedDataIn\[31\]
    PORT
      LAYER met1 ;
        RECT 183.395 23.900 183.640 24.040 ;
    END
  END muxedDataIn\[31\]
  PIN _166_
    PORT
      LAYER met1 ;
        RECT 182.520 22.540 182.765 22.680 ;
    END
  END _166_
  PIN _159_
    PORT
      LAYER met1 ;
        RECT 166.680 19.820 166.820 20.145 ;
    END
  END _159_
  PIN _165_
    PORT
      LAYER met1 ;
        RECT 182.060 22.880 184.605 23.020 ;
    END
  END _165_
  PIN muxedDataIn\[24\]
    PORT
      LAYER met1 ;
        RECT 200.260 19.820 200.400 20.300 ;
    END
  END muxedDataIn\[24\]
  PIN _020_
    PORT
      LAYER met2 ;
        RECT 36.040 336.220 36.180 337.660 ;
    END
  END _020_
  PIN _022_
    PORT
      LAYER met2 ;
        RECT 42.940 336.900 43.080 338.340 ;
    END
  END _022_
  PIN _031_
    PORT
      LAYER met2 ;
        RECT 33.280 200.220 33.420 205.060 ;
    END
  END _031_
  PIN _035_
    PORT
      LAYER met2 ;
        RECT 63.180 274.000 63.320 328.140 ;
    END
  END _035_
  PIN _043_
    PORT
      LAYER met2 ;
        RECT 59.500 332.110 60.100 332.250 ;
    END
  END _043_
  PIN _044_
    PORT
      LAYER met2 ;
        RECT 30.980 192.400 31.120 192.640 ;
    END
  END _044_
  PIN _057_
    PORT
      LAYER met2 ;
        RECT 29.600 198.180 29.740 199.960 ;
    END
  END _057_
  PIN _067_
    PORT
      LAYER met2 ;
        RECT 43.860 332.960 44.460 333.100 ;
    END
  END _067_
  PIN _077_
    PORT
      LAYER met2 ;
        RECT 29.140 203.280 29.280 206.240 ;
    END
  END _077_
  PIN _091_
    PORT
      LAYER met2 ;
        RECT 39.720 309.360 39.860 318.620 ;
    END
  END _091_
  PIN _097_
    PORT
      LAYER met2 ;
        RECT 57.200 371.580 57.340 376.760 ;
    END
  END _097_
  PIN _101_
    PORT
      LAYER met2 ;
        RECT 22.700 193.390 23.300 193.530 ;
    END
  END _101_
  PIN _105_
    PORT
      LAYER met2 ;
        RECT 42.020 221.640 42.160 224.130 ;
    END
  END _105_
  PIN _107_
    PORT
      LAYER met2 ;
        RECT 69.160 309.020 69.300 377.100 ;
    END
  END _107_
  PIN _108_
    PORT
      LAYER met2 ;
        RECT 21.780 192.030 22.840 192.170 ;
    END
  END _108_
  PIN _109_
    PORT
      LAYER met2 ;
        RECT 56.280 295.390 57.340 295.530 ;
    END
  END _109_
  PIN _121_
    PORT
      LAYER met2 ;
        RECT 39.720 297.800 39.860 301.280 ;
    END
  END _121_
  PIN _149_
    PORT
      LAYER met2 ;
        RECT 163.460 23.080 163.600 33.360 ;
    END
  END _149_
  PIN _160_
    PORT
      LAYER met2 ;
        RECT 174.040 15.940 174.180 20.100 ;
    END
  END _160_
  PIN _168_
    PORT
      LAYER met2 ;
        RECT 49.840 146.500 49.980 153.380 ;
    END
  END _168_
  PIN clk
    PORT
      LAYER met2 ;
        RECT 283.520 0.270 285.040 0.410 ;
    END
  END clk
  PIN clknet_0_clk
    PORT
      LAYER met2 ;
        RECT 279.380 20.700 279.520 22.140 ;
    END
  END clknet_0_clk
  PIN clknet_2_2__leaf_clk
    PORT
      LAYER met2 ;
        RECT 98.600 30.900 98.740 32.160 ;
    END
  END clknet_2_2__leaf_clk
  PIN mem_dout\[19\]
    PORT
      LAYER met2 ;
        RECT 67.780 351.520 67.920 445.440 ;
    END
  END mem_dout\[19\]
  PIN mem_dout\[21\]
    PORT
      LAYER met2 ;
        RECT 66.860 330.960 67.000 444.760 ;
    END
  END mem_dout\[21\]
  PIN mem_dout\[22\]
    PORT
      LAYER met2 ;
        RECT 65.940 317.180 66.080 437.960 ;
    END
  END mem_dout\[22\]
  PIN mem_dout\[3\]
    PORT
      LAYER met2 ;
        RECT 207.160 437.540 207.300 442.040 ;
    END
  END mem_dout\[3\]
  PIN mem_wr_mask\[1\]
    PORT
      LAYER met2 ;
        RECT 159.320 18.660 159.460 23.320 ;
    END
  END mem_wr_mask\[1\]
  PIN mem_wr_mask\[2\]
    PORT
      LAYER met2 ;
        RECT 94.920 21.380 95.060 22.140 ;
    END
  END mem_wr_mask\[2\]
  PIN mem_wr_mask\[3\]
    PORT
      LAYER met2 ;
        RECT 166.680 12.880 166.820 23.320 ;
    END
  END mem_wr_mask\[3\]
  PIN muxedDataIn\[15\]
    PORT
      LAYER met2 ;
        RECT 203.480 18.160 203.620 20.780 ;
    END
  END muxedDataIn\[15\]
  PIN muxedDataIn\[16\]
    PORT
      LAYER met2 ;
        RECT 269.260 16.960 269.400 24.680 ;
    END
  END muxedDataIn\[16\]
  PIN muxedDataIn\[18\]
    PORT
      LAYER met2 ;
        RECT 278.920 17.300 279.060 24.680 ;
    END
  END muxedDataIn\[18\]
  PIN muxedDataIn\[19\]
    PORT
      LAYER met2 ;
        RECT 283.060 17.980 283.200 24.680 ;
    END
  END muxedDataIn\[19\]
  PIN muxedDataIn\[20\]
    PORT
      LAYER met2 ;
        RECT 289.960 18.660 290.100 27.400 ;
    END
  END muxedDataIn\[20\]
  PIN muxedDataIn\[21\]
    PORT
      LAYER met2 ;
        RECT 296.860 27.680 297.000 28.260 ;
    END
  END muxedDataIn\[21\]
  PIN muxedDataIn\[22\]
    PORT
      LAYER met2 ;
        RECT 303.760 27.680 303.900 28.600 ;
    END
  END muxedDataIn\[22\]
  PIN muxedDataIn\[23\]
    PORT
      LAYER met2 ;
        RECT 310.660 27.680 310.800 27.920 ;
    END
  END muxedDataIn\[23\]
  PIN muxedDataIn\[25\]
    PORT
      LAYER met2 ;
        RECT 199.865 20.140 199.875 20.150 ;
    END
  END muxedDataIn\[25\]
  PIN muxedDataIn\[27\]
    PORT
      LAYER met2 ;
        RECT 331.360 19.680 331.500 27.400 ;
    END
  END muxedDataIn\[27\]
  PIN muxedDataIn\[28\]
    PORT
      LAYER met2 ;
        RECT 172.660 21.380 172.800 22.480 ;
    END
  END muxedDataIn\[28\]
  PIN muxedDataIn\[29\]
    PORT
      LAYER met2 ;
        RECT 345.160 23.420 345.300 27.400 ;
    END
  END muxedDataIn\[29\]
  PIN muxedDataIn\[30\]
    PORT
      LAYER met2 ;
        RECT 352.520 23.080 352.660 24.680 ;
    END
  END muxedDataIn\[30\]
  PIN muxedDataIn\[8\]
    PORT
      LAYER met2 ;
        RECT 220.960 18.320 221.100 27.400 ;
    END
  END muxedDataIn\[8\]
  PIN net15
    PORT
      LAYER met2 ;
        RECT 8.440 289.270 9.040 289.410 ;
    END
  END net15
  PIN net21
    PORT
      LAYER met2 ;
        RECT 13.500 345.920 13.640 346.160 ;
    END
  END net21
  PIN net23
    PORT
      LAYER met2 ;
        RECT 21.780 134.940 21.920 155.760 ;
    END
  END net23
  PIN net31
    PORT
      LAYER met2 ;
        RECT 24.080 279.070 26.980 279.210 ;
    END
  END net31
  PIN net34
    PORT
      LAYER met2 ;
        RECT 180.940 25.800 181.080 27.400 ;
    END
  END net34
  PIN net35
    PORT
      LAYER met2 ;
        RECT 52.140 202.230 53.200 202.370 ;
    END
  END net35
  PIN net36
    PORT
      LAYER met2 ;
        RECT 8.440 379.920 8.580 381.520 ;
    END
  END net36
  PIN net37
    PORT
      LAYER met2 ;
        RECT 8.440 382.640 8.580 384.240 ;
    END
  END net37
  PIN net4
    PORT
      LAYER met2 ;
        RECT 7.980 116.580 8.120 220.700 ;
    END
  END net4
  PIN net41
    PORT
      LAYER met2 ;
        RECT 8.440 387.870 9.500 388.010 ;
    END
  END net41
  PIN net43
    PORT
      LAYER met2 ;
        RECT 7.060 287.910 8.580 288.050 ;
    END
  END net43
  PIN net45
    PORT
      LAYER met2 ;
        RECT 186.460 26.140 186.600 27.400 ;
    END
  END net45
  PIN net48
    PORT
      LAYER met2 ;
        RECT 193.360 26.820 193.500 27.400 ;
    END
  END net48
  PIN net49
    PORT
      LAYER met2 ;
        RECT 200.260 27.160 200.400 27.400 ;
    END
  END net49
  PIN net50
    PORT
      LAYER met2 ;
        RECT 201.640 26.480 201.780 27.400 ;
    END
  END net50
  PIN net52
    PORT
      LAYER met2 ;
        RECT 214.060 12.720 214.200 22.640 ;
    END
  END net52
  PIN net56
    PORT
      LAYER met2 ;
        RECT 16.460 145.110 16.860 145.250 ;
    END
  END net56
  PIN net64
    PORT
      LAYER met2 ;
        RECT 7.520 244.080 7.660 277.820 ;
    END
  END net64
  PIN net68
    PORT
      LAYER met2 ;
        RECT 17.180 257.000 17.320 285.980 ;
    END
  END net68
  PIN net69
    PORT
      LAYER met2 ;
        RECT 23.160 262.100 23.300 277.820 ;
    END
  END net69
  PIN net71
    PORT
      LAYER met2 ;
        RECT 16.720 271.280 16.860 299.580 ;
    END
  END net71
  PIN net72
    PORT
      LAYER met2 ;
        RECT 22.700 276.720 22.840 299.580 ;
    END
  END net72
  PIN net79
    PORT
      LAYER met2 ;
        RECT 7.520 301.540 7.660 305.360 ;
    END
  END net79
  PIN net81
    PORT
      LAYER met2 ;
        RECT 31.900 189.310 32.500 189.450 ;
    END
  END net81
  PIN net83
    PORT
      LAYER met2 ;
        RECT 24.080 196.790 24.680 196.930 ;
    END
  END net83
  PIN net86
    PORT
      LAYER met2 ;
        RECT 7.520 66.600 7.660 136.380 ;
    END
  END net86
  PIN rd_dout_additional_register\[21\]
    PORT
      LAYER met2 ;
        RECT 37.880 317.180 38.020 326.780 ;
    END
  END rd_dout_additional_register\[21\]
  PIN rd_dout_additional_register\[23\]
    PORT
      LAYER met2 ;
        RECT 47.540 298.820 47.680 302.980 ;
    END
  END rd_dout_additional_register\[23\]
  PIN rd_dout_additional_register\[26\]
    PORT
      LAYER met2 ;
        RECT 43.860 353.220 44.000 354.320 ;
    END
  END rd_dout_additional_register\[26\]
  PIN rd_dout_additional_register\[28\]
    PORT
      LAYER met2 ;
        RECT 47.080 360.700 47.220 380.160 ;
    END
  END rd_dout_additional_register\[28\]
  PIN rd_dout_additional_register\[30\]
    PORT
      LAYER met2 ;
        RECT 54.440 365.800 54.580 373.020 ;
    END
  END rd_dout_additional_register\[30\]
  PIN rd_dout_additional_register\[5\]
    PORT
      LAYER met2 ;
        RECT 30.060 214.500 30.200 228.860 ;
    END
  END rd_dout_additional_register\[5\]
  PIN rd_dout_muxed\[10\]
    PORT
      LAYER met2 ;
        RECT 48.460 279.070 49.060 279.210 ;
    END
  END rd_dout_muxed\[10\]
  PIN rd_dout_muxed\[12\]
    PORT
      LAYER met2 ;
        RECT 48.920 238.270 49.060 245.520 ;
    END
  END rd_dout_muxed\[12\]
  PIN rd_dout_muxed\[13\]
    PORT
      LAYER met2 ;
        RECT 51.220 281.110 52.740 281.250 ;
    END
  END rd_dout_muxed\[13\]
  PIN net87
    PORT
      LAYER met3 ;
        RECT 535.800 417.200 551.630 417.500 ;
    END
  END net87
  PIN C5
    PORT
      LAYER met3 ;
        RECT 0.000 312.990 3.770 313.290 ;
    END
  END C5
  PIN _056_
    PORT
      LAYER met3 ;
        RECT 48.670 282.390 49.060 282.690 ;
    END
  END _056_
  PIN _068_
    PORT
      LAYER met3 ;
        RECT 49.330 353.935 49.340 353.945 ;
    END
  END _068_
  PIN _072_
    PORT
      LAYER met3 ;
        RECT 43.860 281.710 45.170 282.010 ;
    END
  END _072_
  PIN _102_
    PORT
      LAYER met3 ;
        RECT 53.270 366.710 53.660 367.010 ;
    END
  END _102_
  PIN mem_dout\[25\]
    PORT
      LAYER met3 ;
        RECT 51.220 434.030 70.010 434.330 ;
    END
  END mem_dout\[25\]
  PIN C4
    PORT
      LAYER met3 ;
        RECT 0.000 308.230 3.770 308.530 ;
    END
  END C4
  PIN rd_data[16]
    PORT
      LAYER met3 ;
        RECT 0.000 232.070 4.230 232.370 ;
    END
  END rd_data[16]
  PIN rd_data[17]
    PORT
      LAYER met3 ;
        RECT 0.000 236.830 4.230 237.130 ;
    END
  END rd_data[17]
  PIN rd_data[18]
    PORT
      LAYER met3 ;
        RECT 0.000 241.590 4.230 241.890 ;
    END
  END rd_data[18]
  PIN rd_data[19]
    PORT
      LAYER met3 ;
        RECT 0.000 246.350 7.910 246.650 ;
    END
  END rd_data[19]
  PIN rd_data[20]
    PORT
      LAYER met3 ;
        RECT 0.000 251.110 4.230 251.410 ;
    END
  END rd_data[20]
  PIN rd_data[21]
    PORT
      LAYER met3 ;
        RECT 0.000 255.870 4.230 256.170 ;
    END
  END rd_data[21]
  PIN rd_data[22]
    PORT
      LAYER met3 ;
        RECT 0.000 260.630 4.290 260.930 ;
    END
  END rd_data[22]
  PIN rd_data[23]
    PORT
      LAYER met3 ;
        RECT 0.000 265.390 4.230 265.690 ;
    END
  END rd_data[23]
  PIN rd_data[24]
    PORT
      LAYER met3 ;
        RECT 0.000 270.150 4.230 270.450 ;
    END
  END rd_data[24]
  PIN rd_data[25]
    PORT
      LAYER met3 ;
        RECT 0.000 274.910 4.230 275.210 ;
    END
  END rd_data[25]
  PIN rd_data[26]
    PORT
      LAYER met3 ;
        RECT 0.000 279.670 4.230 279.970 ;
    END
  END rd_data[26]
  PIN rd_data[27]
    PORT
      LAYER met3 ;
        RECT 0.000 284.430 4.230 284.730 ;
    END
  END rd_data[27]
  PIN rd_data[28]
    PORT
      LAYER met3 ;
        RECT 0.000 289.190 7.910 289.490 ;
    END
  END rd_data[28]
  PIN rd_data[29]
    PORT
      LAYER met3 ;
        RECT 0.000 293.950 4.230 294.250 ;
    END
  END rd_data[29]
  PIN rd_data[30]
    PORT
      LAYER met3 ;
        RECT 0.000 298.710 4.230 299.010 ;
    END
  END rd_data[30]
  PIN rd_data[31]
    PORT
      LAYER met3 ;
        RECT 0.000 303.470 4.230 303.770 ;
    END
  END rd_data[31]
  PIN wr_addr[0]
    PORT
      LAYER met3 ;
        RECT 0.000 317.750 3.770 318.050 ;
    END
  END wr_addr[0]
  PIN wr_addr[1]
    PORT
      LAYER met3 ;
        RECT 0.000 322.510 4.290 322.810 ;
    END
  END wr_addr[1]
  PIN wr_addr[2]
    PORT
      LAYER met3 ;
        RECT 0.000 327.270 3.770 327.570 ;
    END
  END wr_addr[2]
  PIN wr_addr[3]
    PORT
      LAYER met3 ;
        RECT 0.000 332.030 3.770 332.330 ;
    END
  END wr_addr[3]
  PIN wr_addr[4]
    PORT
      LAYER met3 ;
        RECT 0.000 336.790 7.740 337.090 ;
    END
  END wr_addr[4]
  PIN wr_addr[5]
    PORT
      LAYER met3 ;
        RECT 0.000 341.550 3.770 341.850 ;
    END
  END wr_addr[5]
  PIN wr_addr[6]
    PORT
      LAYER met3 ;
        RECT 0.000 346.310 3.770 346.610 ;
    END
  END wr_addr[6]
  PIN wr_addr[7]
    PORT
      LAYER met3 ;
        RECT 0.000 351.070 7.740 351.370 ;
    END
  END wr_addr[7]
  PIN wr_data[16]
    PORT
      LAYER met3 ;
        RECT 0.000 355.830 3.770 356.130 ;
    END
  END wr_data[16]
  PIN wr_data[17]
    PORT
      LAYER met3 ;
        RECT 0.000 360.590 3.770 360.890 ;
    END
  END wr_data[17]
  PIN wr_data[18]
    PORT
      LAYER met3 ;
        RECT 0.000 365.350 3.770 365.650 ;
    END
  END wr_data[18]
  PIN wr_data[19]
    PORT
      LAYER met3 ;
        RECT 0.000 370.110 3.770 370.410 ;
    END
  END wr_data[19]
  PIN wr_data[20]
    PORT
      LAYER met3 ;
        RECT 0.000 374.870 3.770 375.170 ;
    END
  END wr_data[20]
  PIN wr_data[21]
    PORT
      LAYER met3 ;
        RECT 0.000 379.630 3.770 379.930 ;
    END
  END wr_data[21]
  PIN wr_data[22]
    PORT
      LAYER met3 ;
        RECT 0.000 384.390 3.770 384.690 ;
    END
  END wr_data[22]
  PIN wr_data[23]
    PORT
      LAYER met3 ;
        RECT 0.000 389.150 3.770 389.450 ;
    END
  END wr_data[23]
  PIN wr_data[24]
    PORT
      LAYER met3 ;
        RECT 0.000 393.910 3.770 394.210 ;
    END
  END wr_data[24]
  PIN wr_data[25]
    PORT
      LAYER met3 ;
        RECT 0.000 398.670 4.060 398.970 ;
    END
  END wr_data[25]
  PIN wr_data[26]
    PORT
      LAYER met3 ;
        RECT 0.000 403.430 3.770 403.730 ;
    END
  END wr_data[26]
  PIN wr_data[27]
    PORT
      LAYER met3 ;
        RECT 0.000 408.190 3.770 408.490 ;
    END
  END wr_data[27]
  PIN wr_data[28]
    PORT
      LAYER met3 ;
        RECT 0.000 412.950 4.060 413.250 ;
    END
  END wr_data[28]
  PIN wr_data[29]
    PORT
      LAYER met3 ;
        RECT 0.000 417.710 3.770 418.010 ;
    END
  END wr_data[29]
  PIN wr_data[30]
    PORT
      LAYER met3 ;
        RECT 0.000 422.470 3.770 422.770 ;
    END
  END wr_data[30]
  PIN wr_data[31]
    PORT
      LAYER met3 ;
        RECT 0.000 427.230 7.450 427.530 ;
    END
  END wr_data[31]
  PIN net18
    PORT
      LAYER met3 ;
        RECT 59.250 178.350 70.310 178.650 ;
    END
  END net18
  PIN wr_data[2]
    PORT
      LAYER met3 ;
        RECT 0.000 165.430 7.450 165.730 ;
    END
  END wr_data[2]
  PIN net19
    PORT
      LAYER met3 ;
        RECT 58.790 185.150 70.310 185.450 ;
    END
  END net19
  PIN net20
    PORT
      LAYER met3 ;
        RECT 60.170 192.630 70.310 192.930 ;
    END
  END net20
  PIN wr_data[3]
    PORT
      LAYER met3 ;
        RECT 0.000 170.190 1.530 170.490 ;
    END
  END wr_data[3]
  PIN wr_data[4]
    PORT
      LAYER met3 ;
        RECT 0.000 174.950 3.770 175.250 ;
    END
  END wr_data[4]
  PIN wr_data[5]
    PORT
      LAYER met3 ;
        RECT 0.000 179.710 3.770 180.010 ;
    END
  END wr_data[5]
  PIN wr_data[6]
    PORT
      LAYER met3 ;
        RECT 0.000 184.470 3.770 184.770 ;
    END
  END wr_data[6]
  PIN wr_data[7]
    PORT
      LAYER met3 ;
        RECT 0.000 189.230 3.770 189.530 ;
    END
  END wr_data[7]
  PIN wr_data[8]
    PORT
      LAYER met3 ;
        RECT 0.000 193.990 3.770 194.290 ;
    END
  END wr_data[8]
  PIN wr_data[9]
    PORT
      LAYER met3 ;
        RECT 0.000 198.750 4.290 199.050 ;
    END
  END wr_data[9]
  PIN C0
    PORT
      LAYER met3 ;
        RECT 0.000 98.790 3.770 99.090 ;
    END
  END C0
  PIN C1
    PORT
      LAYER met3 ;
        RECT 0.000 103.550 3.770 103.850 ;
    END
  END C1
  PIN C2
    PORT
      LAYER met3 ;
        RECT 0.000 108.310 3.770 108.610 ;
    END
  END C2
  PIN C3
    PORT
      LAYER met3 ;
        RECT 0.000 113.070 3.770 113.370 ;
    END
  END C3
  PIN net22
    PORT
      LAYER met3 ;
        RECT 60.630 205.550 70.310 205.850 ;
    END
  END net22
  PIN rd_addr[0]
    PORT
      LAYER met3 ;
        RECT 0.000 117.830 3.770 118.130 ;
    END
  END rd_addr[0]
  PIN rd_addr[1]
    PORT
      LAYER met3 ;
        RECT 0.000 122.590 3.770 122.890 ;
    END
  END rd_addr[1]
  PIN rd_addr[2]
    PORT
      LAYER met3 ;
        RECT 0.000 127.350 3.770 127.650 ;
    END
  END rd_addr[2]
  PIN rd_addr[3]
    PORT
      LAYER met3 ;
        RECT 0.000 132.110 3.770 132.410 ;
    END
  END rd_addr[3]
  PIN rd_addr[4]
    PORT
      LAYER met3 ;
        RECT 0.000 136.870 3.770 137.170 ;
    END
  END rd_addr[4]
  PIN rd_addr[5]
    PORT
      LAYER met3 ;
        RECT 0.000 141.630 3.770 141.930 ;
    END
  END rd_addr[5]
  PIN rd_addr[6]
    PORT
      LAYER met3 ;
        RECT 0.000 146.390 3.770 146.690 ;
    END
  END rd_addr[6]
  PIN rd_addr[7]
    PORT
      LAYER met3 ;
        RECT 0.000 151.150 6.990 151.450 ;
    END
  END rd_addr[7]
  PIN rd_data[0]
    PORT
      LAYER met3 ;
        RECT 0.000 22.630 4.230 22.930 ;
    END
  END rd_data[0]
  PIN rd_data[10]
    PORT
      LAYER met3 ;
        RECT 0.000 70.230 4.230 70.530 ;
    END
  END rd_data[10]
  PIN rd_data[11]
    PORT
      LAYER met3 ;
        RECT 0.000 74.990 4.290 75.290 ;
    END
  END rd_data[11]
  PIN rd_data[12]
    PORT
      LAYER met3 ;
        RECT 0.000 79.750 4.230 80.050 ;
    END
  END rd_data[12]
  PIN rd_data[13]
    PORT
      LAYER met3 ;
        RECT 0.000 84.510 4.230 84.810 ;
    END
  END rd_data[13]
  PIN rd_data[14]
    PORT
      LAYER met3 ;
        RECT 0.000 89.270 7.910 89.570 ;
    END
  END rd_data[14]
  PIN rd_data[15]
    PORT
      LAYER met3 ;
        RECT 0.000 94.030 4.230 94.330 ;
    END
  END rd_data[15]
  PIN rd_data[2]
    PORT
      LAYER met3 ;
        RECT 0.000 32.150 4.230 32.450 ;
    END
  END rd_data[2]
  PIN rd_data[1]
    PORT
      LAYER met3 ;
        RECT 0.000 27.390 7.910 27.690 ;
    END
  END rd_data[1]
  PIN rd_data[3]
    PORT
      LAYER met3 ;
        RECT 0.000 36.910 4.230 37.210 ;
    END
  END rd_data[3]
  PIN rd_data[4]
    PORT
      LAYER met3 ;
        RECT 0.000 41.670 4.230 41.970 ;
    END
  END rd_data[4]
  PIN rd_data[5]
    PORT
      LAYER met3 ;
        RECT 0.000 46.430 4.230 46.730 ;
    END
  END rd_data[5]
  PIN rd_data[6]
    PORT
      LAYER met3 ;
        RECT 0.000 51.190 4.230 51.490 ;
    END
  END rd_data[6]
  PIN rd_data[7]
    PORT
      LAYER met3 ;
        RECT 0.000 55.950 4.230 56.250 ;
    END
  END rd_data[7]
  PIN rd_data[8]
    PORT
      LAYER met3 ;
        RECT 0.000 60.710 4.230 61.010 ;
    END
  END rd_data[8]
  PIN rd_data[9]
    PORT
      LAYER met3 ;
        RECT 0.000 65.470 4.230 65.770 ;
    END
  END rd_data[9]
  PIN wr_data[0]
    PORT
      LAYER met3 ;
        RECT 0.000 155.910 3.770 156.210 ;
    END
  END wr_data[0]
  PIN wr_data[10]
    PORT
      LAYER met3 ;
        RECT 0.000 203.510 3.770 203.810 ;
    END
  END wr_data[10]
  PIN wr_data[11]
    PORT
      LAYER met3 ;
        RECT 0.000 208.270 3.770 208.570 ;
    END
  END wr_data[11]
  PIN wr_data[12]
    PORT
      LAYER met3 ;
        RECT 0.000 213.030 3.770 213.330 ;
    END
  END wr_data[12]
  PIN wr_data[13]
    PORT
      LAYER met3 ;
        RECT 0.000 217.790 3.770 218.090 ;
    END
  END wr_data[13]
  PIN wr_data[14]
    PORT
      LAYER met3 ;
        RECT 0.000 222.550 3.770 222.850 ;
    END
  END wr_data[14]
  PIN wr_data[15]
    PORT
      LAYER met3 ;
        RECT 0.000 227.310 6.990 227.610 ;
    END
  END wr_data[15]
  PIN wr_data[1]
    PORT
      LAYER met3 ;
        RECT 0.000 160.670 3.770 160.970 ;
    END
  END wr_data[1]
  PIN _163_
    PORT
      LAYER met3 ;
        RECT 49.590 194.670 65.620 194.970 ;
    END
  END _163_
  PIN _164_
    PORT
      LAYER met3 ;
        RECT 96.910 32.150 97.210 33.130 ;
    END
  END _164_
  PIN memWriteEnable
    PORT
      LAYER met3 ;
        RECT 70.010 62.880 70.310 73.250 ;
    END
  END memWriteEnable
  PIN muxedDataIn\[17\]
    PORT
      LAYER met3 ;
        RECT 186.065 23.540 186.075 23.550 ;
    END
  END muxedDataIn\[17\]
  PIN net17
    PORT
      LAYER met3 ;
        RECT 55.425 172.290 55.435 172.300 ;
    END
  END net17
  PIN net8
    PORT
      LAYER met3 ;
        RECT 484.910 118.000 552.610 118.300 ;
    END
  END net8
  PIN net10
    PORT
      LAYER met3 ;
        RECT 484.120 103.040 552.610 103.340 ;
    END
  END net10
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 563.100 21.520 563.900 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.720 -5.460 546.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 524.720 -5.460 526.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.720 -5.460 506.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.720 -5.460 486.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 464.720 -5.460 466.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 444.720 -5.460 446.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 424.720 -5.460 426.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.720 -5.460 406.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 384.720 -5.460 386.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.720 -5.460 366.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 344.720 -5.460 346.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 324.720 -5.460 326.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 304.720 -5.460 306.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 284.720 -5.460 286.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 264.720 -5.460 266.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 244.720 -5.460 246.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.720 -5.460 226.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 204.720 -5.460 206.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 184.720 -5.460 186.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 164.720 -5.460 166.320 24.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 144.720 -5.460 146.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 124.720 -5.460 126.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 104.720 -5.460 106.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.720 -5.460 86.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.720 -5.460 66.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 44.720 -5.460 46.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.720 -5.460 26.320 454.260 ;
    END
  END VGND
  PIN VPWR
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 561.260 21.520 562.060 443.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 554.720 -5.460 556.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 534.720 -5.460 536.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 514.720 -5.460 516.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 494.720 -5.460 496.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 474.720 -5.460 476.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 454.720 -5.460 456.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 434.720 -5.460 436.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 414.720 -5.460 416.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 394.720 -5.460 396.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 374.720 -5.460 376.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 354.720 -5.460 356.320 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 334.720 -5.460 336.320 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.720 -5.460 316.320 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.720 -5.460 296.320 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 274.720 -5.460 276.320 24.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 254.720 -5.460 256.320 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.720 -5.460 236.320 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 214.720 -5.460 216.320 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 194.720 -5.460 196.320 24.485 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.720 -5.460 176.320 24.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.720 -5.460 156.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 134.720 -5.460 136.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 114.720 -5.460 116.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 94.720 -5.460 96.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.720 -5.460 76.320 25.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 54.720 -5.460 56.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 34.720 -5.460 36.320 454.260 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.720 -5.460 16.320 454.260 ;
    END
  END VPWR
  PIN _009_
    PORT
      LAYER met4 ;
        RECT 48.180 298.855 48.190 298.865 ;
    END
  END _009_
  PIN clknet_2_1__leaf_clk
    PORT
      LAYER met4 ;
        RECT 520.200 417.510 520.500 433.650 ;
    END
  END clknet_2_1__leaf_clk
  PIN mem_dout\[0\]
    PORT
      LAYER met4 ;
        RECT 210.800 405.950 211.100 433.650 ;
    END
  END mem_dout\[0\]
  PIN mem_dout\[10\]
    PORT
      LAYER met4 ;
        RECT 273.360 405.950 273.660 433.650 ;
    END
  END mem_dout\[10\]
  PIN mem_dout\[11\]
    PORT
      LAYER met4 ;
        RECT 279.480 405.950 279.780 433.650 ;
    END
  END mem_dout\[11\]
  PIN mem_dout\[12\]
    PORT
      LAYER met4 ;
        RECT 286.280 405.950 286.580 433.650 ;
    END
  END mem_dout\[12\]
  PIN mem_dout\[13\]
    PORT
      LAYER met4 ;
        RECT 291.720 405.950 292.020 433.650 ;
    END
  END mem_dout\[13\]
  PIN mem_dout\[14\]
    PORT
      LAYER met4 ;
        RECT 297.840 405.950 298.140 433.650 ;
    END
  END mem_dout\[14\]
  PIN mem_dout\[15\]
    PORT
      LAYER met4 ;
        RECT 304.640 405.950 304.940 433.340 ;
    END
  END mem_dout\[15\]
  PIN mem_dout\[16\]
    PORT
      LAYER met4 ;
        RECT 310.760 405.950 311.060 433.650 ;
    END
  END mem_dout\[16\]
  PIN mem_dout\[17\]
    PORT
      LAYER met4 ;
        RECT 317.560 405.950 317.860 433.650 ;
    END
  END mem_dout\[17\]
  PIN mem_dout\[18\]
    PORT
      LAYER met4 ;
        RECT 323.000 405.950 323.300 434.020 ;
    END
  END mem_dout\[18\]
  PIN mem_dout\[1\]
    PORT
      LAYER met4 ;
        RECT 217.600 405.950 217.900 433.650 ;
    END
  END mem_dout\[1\]
  PIN mem_dout\[20\]
    PORT
      LAYER met4 ;
        RECT 335.240 405.950 335.540 434.330 ;
    END
  END mem_dout\[20\]
  PIN mem_dout\[24\]
    PORT
      LAYER met4 ;
        RECT 361.080 405.950 361.380 434.330 ;
    END
  END mem_dout\[24\]
  PIN mem_dout\[26\]
    PORT
      LAYER met4 ;
        RECT 373.320 405.950 373.620 433.650 ;
    END
  END mem_dout\[26\]
  PIN mem_dout\[27\]
    PORT
      LAYER met4 ;
        RECT 379.440 405.950 379.740 433.650 ;
    END
  END mem_dout\[27\]
  PIN mem_dout\[28\]
    PORT
      LAYER met4 ;
        RECT 386.240 405.950 386.540 433.650 ;
    END
  END mem_dout\[28\]
  PIN mem_dout\[29\]
    PORT
      LAYER met4 ;
        RECT 391.680 405.950 391.980 433.650 ;
    END
  END mem_dout\[29\]
  PIN mem_dout\[2\]
    PORT
      LAYER met4 ;
        RECT 223.040 405.950 223.340 433.650 ;
    END
  END mem_dout\[2\]
  PIN mem_dout\[30\]
    PORT
      LAYER met4 ;
        RECT 397.800 405.950 398.100 433.650 ;
    END
  END mem_dout\[30\]
  PIN mem_dout\[31\]
    PORT
      LAYER met4 ;
        RECT 404.600 405.950 404.900 433.650 ;
    END
  END mem_dout\[31\]
  PIN mem_dout\[6\]
    PORT
      LAYER met4 ;
        RECT 248.880 405.950 249.180 433.650 ;
    END
  END mem_dout\[6\]
  PIN mem_dout\[8\]
    PORT
      LAYER met4 ;
        RECT 261.120 405.950 261.420 433.650 ;
    END
  END mem_dout\[8\]
  PIN muxedDataIn\[9\]
    PORT
      LAYER met4 ;
        RECT 226.630 27.700 226.930 32.450 ;
    END
  END muxedDataIn\[9\]
  PIN net11
    PORT
      LAYER met4 ;
        RECT 486.070 27.020 486.370 34.650 ;
    END
  END net11
  PIN net12
    PORT
      LAYER met4 ;
        RECT 483.310 26.340 483.610 34.650 ;
    END
  END net12
  PIN net13
    PORT
      LAYER met4 ;
        RECT 486.990 20.900 487.290 34.180 ;
    END
  END net13
  PIN net14
    PORT
      LAYER met4 ;
        RECT 484.230 25.660 484.530 32.450 ;
    END
  END net14
  PIN net51
    PORT
      LAYER met4 ;
        RECT 210.990 20.220 211.290 34.650 ;
    END
  END net51
  PIN net7
    PORT
      LAYER met4 ;
        RECT 467.160 414.790 467.460 433.650 ;
    END
  END net7
  OBS
      LAYER li1 ;
        RECT 5.520 5.355 564.420 443.445 ;
      LAYER met1 ;
        RECT 3.750 441.840 564.420 449.100 ;
        RECT 3.750 441.140 50.220 441.840 ;
        RECT 228.050 441.140 564.420 441.840 ;
        RECT 3.750 434.020 564.420 441.140 ;
        RECT 3.750 433.320 52.935 434.020 ;
        RECT 70.960 433.320 564.420 434.020 ;
        RECT 3.750 431.980 564.420 433.320 ;
        RECT 3.750 431.280 56.155 431.980 ;
        RECT 59.720 431.280 564.420 431.980 ;
        RECT 3.750 428.240 564.420 431.280 ;
        RECT 3.750 427.540 8.315 428.240 ;
        RECT 10.040 427.540 564.420 428.240 ;
        RECT 3.750 422.800 564.420 427.540 ;
        RECT 3.750 422.100 8.315 422.800 ;
        RECT 11.420 422.100 564.420 422.800 ;
        RECT 3.750 420.080 564.420 422.100 ;
        RECT 3.750 419.380 8.315 420.080 ;
        RECT 12.340 419.380 564.420 420.080 ;
        RECT 3.750 409.200 564.420 419.380 ;
        RECT 3.750 408.500 8.315 409.200 ;
        RECT 10.500 408.500 564.420 409.200 ;
        RECT 3.750 400.700 564.420 408.500 ;
        RECT 3.750 400.000 7.855 400.700 ;
        RECT 11.880 400.000 564.420 400.700 ;
        RECT 3.750 390.160 564.420 400.000 ;
        RECT 3.750 389.460 8.315 390.160 ;
        RECT 10.960 389.460 564.420 390.160 ;
        RECT 3.750 370.780 564.420 389.460 ;
        RECT 3.750 370.080 29.520 370.780 ;
        RECT 47.500 370.080 564.420 370.780 ;
        RECT 3.750 367.040 564.420 370.080 ;
        RECT 3.750 365.815 54.620 367.040 ;
        RECT 55.320 365.815 564.420 367.040 ;
        RECT 3.750 365.340 564.420 365.815 ;
        RECT 3.750 364.640 26.760 365.340 ;
        RECT 47.040 364.640 564.420 365.340 ;
        RECT 3.750 364.320 564.420 364.640 ;
        RECT 3.750 363.620 47.875 364.320 ;
        RECT 52.360 363.620 564.420 364.320 ;
        RECT 3.750 362.620 564.420 363.620 ;
        RECT 3.750 361.920 21.240 362.620 ;
        RECT 45.965 361.920 564.420 362.620 ;
        RECT 3.750 360.240 564.420 361.920 ;
        RECT 3.750 359.900 38.720 360.240 ;
        RECT 3.750 359.200 22.160 359.900 ;
        RECT 45.660 359.540 564.420 360.240 ;
        RECT 45.045 359.200 564.420 359.540 ;
        RECT 3.750 357.520 564.420 359.200 ;
        RECT 3.750 356.820 54.360 357.520 ;
        RECT 56.700 356.820 564.420 357.520 ;
        RECT 3.750 354.460 564.420 356.820 ;
        RECT 3.750 353.760 32.740 354.460 ;
        RECT 40.445 353.760 42.355 354.460 ;
        RECT 43.820 353.760 564.420 354.460 ;
        RECT 3.750 353.440 564.420 353.760 ;
        RECT 3.750 352.740 21.700 353.440 ;
        RECT 41.825 352.740 47.720 353.440 ;
        RECT 52.405 352.760 564.420 353.440 ;
        RECT 3.750 352.215 47.720 352.740 ;
        RECT 48.420 352.605 50.480 352.740 ;
        RECT 48.420 352.215 49.100 352.605 ;
        RECT 3.750 351.720 49.100 352.215 ;
        RECT 49.800 352.060 50.480 352.605 ;
        RECT 54.705 352.605 564.420 352.760 ;
        RECT 54.705 352.080 55.540 352.605 ;
        RECT 56.240 352.080 564.420 352.605 ;
        RECT 49.800 351.720 53.395 352.060 ;
        RECT 3.750 351.380 53.395 351.720 ;
        RECT 57.880 351.380 564.420 352.080 ;
        RECT 3.750 348.000 564.420 351.380 ;
        RECT 3.750 347.165 48.180 348.000 ;
        RECT 3.750 346.280 41.280 347.165 ;
        RECT 41.980 346.790 48.180 347.165 ;
        RECT 48.880 346.790 564.420 348.000 ;
        RECT 41.980 346.280 564.420 346.790 ;
        RECT 3.750 344.105 564.420 346.280 ;
        RECT 3.750 343.580 47.260 344.105 ;
        RECT 3.750 342.880 44.240 343.580 ;
        RECT 45.505 342.880 47.260 343.580 ;
        RECT 47.960 342.880 564.420 344.105 ;
        RECT 3.750 342.220 564.420 342.880 ;
        RECT 3.750 341.335 46.800 342.220 ;
        RECT 47.500 341.335 564.420 342.220 ;
        RECT 3.750 339.980 564.420 341.335 ;
        RECT 3.750 339.140 67.040 339.980 ;
        RECT 67.740 339.140 564.420 339.980 ;
        RECT 3.750 337.120 564.420 339.140 ;
        RECT 3.750 336.420 30.395 337.120 ;
        RECT 39.480 336.440 564.420 337.120 ;
        RECT 39.480 336.420 45.575 336.440 ;
        RECT 3.750 335.740 45.575 336.420 ;
        RECT 46.380 336.285 564.420 336.440 ;
        RECT 3.750 335.060 46.340 335.740 ;
        RECT 47.040 335.060 564.420 336.285 ;
        RECT 3.750 333.720 564.420 335.060 ;
        RECT 3.750 333.040 41.895 333.720 ;
        RECT 3.750 332.340 38.520 333.040 ;
        RECT 41.365 333.020 41.895 333.040 ;
        RECT 50.060 333.020 564.420 333.720 ;
        RECT 41.365 332.340 564.420 333.020 ;
        RECT 3.750 331.340 564.420 332.340 ;
        RECT 3.750 330.640 38.215 331.340 ;
        RECT 39.940 330.640 564.420 331.340 ;
        RECT 3.750 330.320 564.420 330.640 ;
        RECT 3.750 329.620 19.860 330.320 ;
        RECT 36.460 329.620 564.420 330.320 ;
        RECT 3.750 328.280 564.420 329.620 ;
        RECT 3.750 327.580 40.560 328.280 ;
        RECT 41.825 327.875 564.420 328.280 ;
        RECT 41.825 327.580 46.400 327.875 ;
        RECT 3.750 327.305 46.400 327.580 ;
        RECT 46.970 327.305 564.420 327.875 ;
        RECT 3.750 325.405 564.420 327.305 ;
        RECT 3.750 323.840 8.160 325.405 ;
        RECT 8.860 325.220 564.420 325.405 ;
        RECT 8.860 324.520 44.040 325.220 ;
        RECT 45.965 324.520 564.420 325.220 ;
        RECT 8.860 323.840 564.420 324.520 ;
        RECT 3.750 322.840 564.420 323.840 ;
        RECT 3.750 322.140 38.260 322.840 ;
        RECT 39.065 322.435 55.695 322.840 ;
        RECT 39.065 322.140 55.140 322.435 ;
        RECT 60.640 322.140 564.420 322.840 ;
        RECT 3.750 321.865 55.140 322.140 ;
        RECT 55.710 321.865 564.420 322.140 ;
        RECT 3.750 320.600 564.420 321.865 ;
        RECT 3.750 320.085 51.400 320.600 ;
        RECT 3.750 320.060 51.000 320.085 ;
        RECT 3.750 319.920 46.865 320.060 ;
        RECT 3.750 318.740 41.280 319.920 ;
        RECT 41.980 319.490 46.865 319.920 ;
        RECT 47.435 319.965 51.000 320.060 ;
        RECT 47.435 319.490 50.020 319.965 ;
        RECT 41.980 318.740 50.020 319.490 ;
        RECT 50.720 319.515 51.000 319.965 ;
        RECT 52.100 319.575 564.420 320.600 ;
        RECT 51.570 319.515 564.420 319.575 ;
        RECT 50.720 318.740 564.420 319.515 ;
        RECT 3.750 317.740 564.420 318.740 ;
        RECT 3.750 317.040 32.695 317.740 ;
        RECT 34.420 317.060 564.420 317.740 ;
        RECT 34.420 317.040 36.680 317.060 ;
        RECT 3.750 316.360 36.680 317.040 ;
        RECT 39.985 316.860 564.420 317.060 ;
        RECT 39.985 316.360 65.200 316.860 ;
        RECT 3.750 315.680 65.200 316.360 ;
        RECT 65.900 315.680 564.420 316.860 ;
        RECT 3.750 315.360 564.420 315.680 ;
        RECT 3.750 314.660 37.755 315.360 ;
        RECT 39.480 314.680 43.320 315.360 ;
        RECT 39.480 314.660 40.560 314.680 ;
        RECT 3.750 313.980 40.560 314.660 ;
        RECT 41.365 314.660 43.320 314.680 ;
        RECT 44.125 314.660 48.840 315.360 ;
        RECT 55.165 314.660 564.420 315.360 ;
        RECT 41.365 314.135 53.240 314.660 ;
        RECT 53.940 314.135 564.420 314.660 ;
        RECT 41.365 313.980 564.420 314.135 ;
        RECT 3.750 311.960 564.420 313.980 ;
        RECT 3.750 311.260 51.860 311.960 ;
        RECT 53.785 311.260 564.420 311.960 ;
        RECT 3.750 310.920 52.520 311.260 ;
        RECT 53.320 310.920 564.420 311.260 ;
        RECT 3.750 309.920 564.420 310.920 ;
        RECT 3.750 309.220 38.720 309.920 ;
        RECT 42.285 309.220 51.860 309.920 ;
        RECT 54.200 309.220 564.420 309.920 ;
        RECT 3.750 303.800 564.420 309.220 ;
        RECT 3.750 303.100 43.275 303.800 ;
        RECT 50.520 303.100 564.420 303.800 ;
        RECT 3.750 301.080 564.420 303.100 ;
        RECT 3.750 300.195 7.240 301.080 ;
        RECT 7.940 300.195 21.960 301.080 ;
        RECT 22.660 300.740 564.420 301.080 ;
        RECT 22.660 300.195 23.495 300.740 ;
        RECT 3.750 300.040 23.495 300.195 ;
        RECT 27.060 300.040 564.420 300.740 ;
        RECT 3.750 296.320 564.420 300.040 ;
        RECT 3.750 295.620 45.620 296.320 ;
        RECT 51.945 295.640 564.420 296.320 ;
        RECT 3.750 295.300 51.600 295.620 ;
        RECT 54.705 295.485 564.420 295.640 ;
        RECT 3.750 294.600 7.395 295.300 ;
        RECT 23.380 294.940 51.600 295.300 ;
        RECT 23.380 294.600 54.620 294.940 ;
        RECT 3.750 294.260 54.620 294.600 ;
        RECT 55.320 294.260 564.420 295.485 ;
        RECT 3.750 293.600 564.420 294.260 ;
        RECT 3.750 293.260 49.300 293.600 ;
        RECT 3.750 292.375 45.420 293.260 ;
        RECT 46.120 292.900 49.300 293.260 ;
        RECT 52.865 292.900 564.420 293.600 ;
        RECT 46.120 292.375 564.420 292.900 ;
        RECT 3.750 289.860 564.420 292.375 ;
        RECT 3.750 289.160 7.395 289.860 ;
        RECT 22.460 289.520 564.420 289.860 ;
        RECT 22.460 289.160 50.940 289.520 ;
        RECT 3.750 288.820 50.940 289.160 ;
        RECT 59.260 288.820 61.750 289.520 ;
        RECT 62.940 288.820 564.420 289.520 ;
        RECT 3.750 287.820 564.420 288.820 ;
        RECT 3.750 287.120 7.395 287.820 ;
        RECT 21.540 287.480 564.420 287.820 ;
        RECT 3.750 286.800 17.975 287.120 ;
        RECT 27.520 286.800 42.770 287.480 ;
        RECT 3.750 286.460 16.440 286.800 ;
        RECT 38.100 286.780 42.770 286.800 ;
        RECT 47.040 287.140 564.420 287.480 ;
        RECT 47.040 286.780 61.750 287.140 ;
        RECT 38.100 286.460 61.750 286.780 ;
        RECT 3.750 285.760 13.880 286.460 ;
        RECT 16.065 286.100 16.440 286.460 ;
        RECT 16.065 285.760 33.200 286.100 ;
        RECT 48.725 285.760 49.715 286.460 ;
        RECT 54.200 286.440 61.750 286.460 ;
        RECT 63.860 286.440 564.420 287.140 ;
        RECT 54.200 285.760 564.420 286.440 ;
        RECT 3.750 284.420 564.420 285.760 ;
        RECT 3.750 283.720 23.495 284.420 ;
        RECT 38.760 283.925 564.420 284.420 ;
        RECT 38.760 283.720 44.960 283.925 ;
        RECT 3.750 283.040 44.960 283.720 ;
        RECT 45.660 283.040 564.420 283.925 ;
        RECT 3.750 282.380 564.420 283.040 ;
        RECT 3.750 281.680 7.395 282.380 ;
        RECT 13.260 281.680 31.820 282.380 ;
        RECT 32.625 281.700 47.260 282.380 ;
        RECT 32.625 281.680 47.000 281.700 ;
        RECT 61.100 281.680 564.420 282.380 ;
        RECT 3.750 281.000 47.000 281.680 ;
        RECT 49.645 281.000 50.020 281.680 ;
        RECT 58.340 281.340 564.420 281.680 ;
        RECT 54.660 281.000 564.420 281.340 ;
        RECT 3.750 279.660 564.420 281.000 ;
        RECT 3.750 278.960 15.980 279.660 ;
        RECT 28.440 278.980 564.420 279.660 ;
        RECT 3.750 278.620 19.660 278.960 ;
        RECT 3.750 278.280 23.955 278.620 ;
        RECT 37.180 278.280 564.420 278.980 ;
        RECT 3.750 277.125 564.420 278.280 ;
        RECT 3.750 276.600 44.040 277.125 ;
        RECT 3.750 275.900 41.895 276.600 ;
        RECT 42.900 276.240 44.040 276.600 ;
        RECT 44.740 276.240 564.420 277.125 ;
        RECT 42.900 275.900 564.420 276.240 ;
        RECT 3.750 273.880 564.420 275.900 ;
        RECT 3.750 273.180 47.260 273.880 ;
        RECT 53.740 273.180 564.420 273.880 ;
        RECT 3.750 272.840 47.875 273.180 ;
        RECT 50.980 272.840 564.420 273.180 ;
        RECT 3.750 271.160 564.420 272.840 ;
        RECT 3.750 270.460 23.035 271.160 ;
        RECT 37.840 270.460 564.420 271.160 ;
        RECT 3.750 269.120 564.420 270.460 ;
        RECT 3.750 268.420 28.600 269.120 ;
        RECT 30.325 268.420 564.420 269.120 ;
        RECT 3.750 268.100 564.420 268.420 ;
        RECT 3.750 267.400 7.395 268.100 ;
        RECT 13.720 267.400 564.420 268.100 ;
        RECT 3.750 265.720 564.420 267.400 ;
        RECT 3.750 265.020 22.575 265.720 ;
        RECT 33.240 265.020 564.420 265.720 ;
        RECT 3.750 264.700 564.420 265.020 ;
        RECT 3.750 264.000 21.240 264.700 ;
        RECT 22.045 264.000 564.420 264.700 ;
        RECT 3.750 263.340 564.420 264.000 ;
        RECT 3.750 262.640 41.480 263.340 ;
        RECT 56.085 262.640 564.420 263.340 ;
        RECT 3.750 249.740 564.420 262.640 ;
        RECT 3.750 249.040 7.395 249.740 ;
        RECT 19.240 249.040 564.420 249.740 ;
        RECT 3.750 240.900 564.420 249.040 ;
        RECT 3.750 240.200 30.395 240.900 ;
        RECT 32.165 240.200 33.155 240.900 ;
        RECT 36.720 240.200 36.835 240.900 ;
        RECT 39.480 240.200 45.990 240.900 ;
        RECT 53.280 240.200 564.420 240.900 ;
        RECT 3.750 239.200 564.420 240.200 ;
        RECT 3.750 238.860 30.395 239.200 ;
        RECT 3.750 238.160 7.395 238.860 ;
        RECT 22.460 238.500 30.395 238.860 ;
        RECT 43.160 238.860 564.420 239.200 ;
        RECT 43.160 238.520 51.860 238.860 ;
        RECT 22.460 238.160 42.770 238.500 ;
        RECT 3.750 237.820 42.770 238.160 ;
        RECT 44.540 237.975 51.860 238.520 ;
        RECT 52.560 237.975 564.420 238.860 ;
        RECT 44.540 237.820 564.420 237.975 ;
        RECT 3.750 235.460 564.420 237.820 ;
        RECT 3.750 235.120 45.990 235.460 ;
        RECT 3.750 234.420 28.970 235.120 ;
        RECT 32.580 234.760 45.990 235.120 ;
        RECT 52.820 234.760 564.420 235.460 ;
        RECT 32.580 234.420 564.420 234.760 ;
        RECT 3.750 233.420 564.420 234.420 ;
        RECT 3.750 233.080 44.150 233.420 ;
        RECT 3.750 232.380 29.935 233.080 ;
        RECT 31.400 232.380 33.110 233.080 ;
        RECT 36.920 232.720 44.150 233.080 ;
        RECT 47.760 232.720 564.420 233.420 ;
        RECT 36.920 232.380 564.420 232.720 ;
        RECT 3.750 231.040 564.420 232.380 ;
        RECT 3.750 230.020 43.580 231.040 ;
        RECT 3.750 229.680 35.410 230.020 ;
        RECT 3.750 229.340 28.050 229.680 ;
        RECT 3.750 228.640 7.855 229.340 ;
        RECT 10.040 228.980 28.050 229.340 ;
        RECT 29.820 229.320 35.410 229.680 ;
        RECT 37.640 229.475 43.580 230.020 ;
        RECT 44.280 229.475 564.420 231.040 ;
        RECT 37.640 229.320 564.420 229.475 ;
        RECT 29.820 228.980 564.420 229.320 ;
        RECT 10.040 228.640 564.420 228.980 ;
        RECT 3.750 227.640 564.420 228.640 ;
        RECT 3.750 226.940 32.695 227.640 ;
        RECT 37.380 226.940 41.940 227.640 ;
        RECT 43.105 226.940 564.420 227.640 ;
        RECT 3.750 224.240 564.420 226.940 ;
        RECT 3.750 223.540 28.050 224.240 ;
        RECT 29.360 223.540 31.820 224.240 ;
        RECT 35.690 223.540 564.420 224.240 ;
        RECT 3.750 222.880 564.420 223.540 ;
        RECT 3.750 222.540 33.200 222.880 ;
        RECT 3.750 221.840 21.700 222.540 ;
        RECT 30.480 222.180 33.200 222.540 ;
        RECT 34.465 222.180 41.435 222.880 ;
        RECT 50.520 222.180 564.420 222.880 ;
        RECT 30.480 221.840 42.860 222.180 ;
        RECT 44.890 221.840 564.420 222.180 ;
        RECT 3.750 220.160 564.420 221.840 ;
        RECT 3.750 219.820 30.855 220.160 ;
        RECT 39.020 219.820 564.420 220.160 ;
        RECT 3.750 219.120 18.940 219.820 ;
        RECT 40.445 219.140 564.420 219.820 ;
        RECT 40.445 219.120 46.955 219.140 ;
        RECT 3.750 218.800 46.955 219.120 ;
        RECT 49.800 218.800 564.420 219.140 ;
        RECT 3.750 218.460 42.355 218.800 ;
        RECT 3.750 217.760 7.855 218.460 ;
        RECT 11.880 218.100 42.355 218.460 ;
        RECT 50.260 218.100 564.420 218.800 ;
        RECT 11.880 217.760 564.420 218.100 ;
        RECT 3.750 217.440 564.420 217.760 ;
        RECT 3.750 216.420 32.540 217.440 ;
        RECT 3.750 215.195 26.560 216.420 ;
        RECT 27.260 216.215 32.540 216.420 ;
        RECT 33.240 216.215 564.420 217.440 ;
        RECT 27.260 216.080 564.420 216.215 ;
        RECT 27.260 215.195 29.780 216.080 ;
        RECT 30.480 215.740 564.420 216.080 ;
        RECT 30.480 215.195 34.075 215.740 ;
        RECT 3.750 215.040 34.075 215.195 ;
        RECT 35.080 215.040 564.420 215.740 ;
        RECT 3.750 214.720 564.420 215.040 ;
        RECT 3.750 214.020 27.175 214.720 ;
        RECT 29.820 214.020 564.420 214.720 ;
        RECT 3.750 213.700 564.420 214.020 ;
        RECT 3.750 213.020 46.955 213.700 ;
        RECT 3.750 212.320 7.855 213.020 ;
        RECT 11.420 212.320 26.760 213.020 ;
        RECT 28.485 213.000 46.955 213.020 ;
        RECT 52.100 213.000 564.420 213.700 ;
        RECT 28.485 212.320 48.380 213.000 ;
        RECT 50.015 212.320 564.420 213.000 ;
        RECT 3.750 212.000 564.420 212.320 ;
        RECT 3.750 211.660 41.895 212.000 ;
        RECT 49.140 211.660 564.420 212.000 ;
        RECT 3.750 210.960 34.075 211.660 ;
        RECT 49.800 210.960 564.420 211.660 ;
        RECT 3.750 210.300 564.420 210.960 ;
        RECT 3.750 209.600 7.855 210.300 ;
        RECT 10.960 209.600 49.255 210.300 ;
        RECT 59.720 209.600 564.420 210.300 ;
        RECT 3.750 209.280 564.420 209.600 ;
        RECT 3.750 208.580 29.015 209.280 ;
        RECT 34.420 208.580 36.835 209.280 ;
        RECT 43.160 208.580 564.420 209.280 ;
        RECT 3.750 208.260 564.420 208.580 ;
        RECT 3.750 207.560 32.695 208.260 ;
        RECT 35.540 208.105 564.420 208.260 ;
        RECT 3.750 207.220 35.300 207.560 ;
        RECT 36.000 207.220 564.420 208.105 ;
        RECT 3.750 206.220 564.420 207.220 ;
        RECT 3.750 205.335 31.620 206.220 ;
        RECT 32.320 205.335 564.420 206.220 ;
        RECT 3.750 204.860 564.420 205.335 ;
        RECT 3.750 204.160 7.855 204.860 ;
        RECT 39.020 204.160 49.715 204.860 ;
        RECT 66.160 204.160 564.420 204.860 ;
        RECT 3.750 203.840 564.420 204.160 ;
        RECT 3.750 203.140 17.560 203.840 ;
        RECT 34.850 203.160 564.420 203.840 ;
        RECT 34.850 203.140 52.780 203.160 ;
        RECT 3.750 202.460 22.880 203.140 ;
        RECT 25.725 202.820 28.400 203.140 ;
        RECT 30.740 202.820 52.780 203.140 ;
        RECT 25.725 202.460 25.795 202.820 ;
        RECT 3.750 202.120 25.795 202.460 ;
        RECT 27.520 202.460 28.400 202.820 ;
        RECT 31.200 202.460 52.780 202.820 ;
        RECT 65.700 202.460 564.420 203.160 ;
        RECT 27.520 202.120 29.475 202.460 ;
        RECT 31.200 202.120 564.420 202.460 ;
        RECT 3.750 201.120 564.420 202.120 ;
        RECT 3.750 200.420 7.855 201.120 ;
        RECT 9.580 200.780 41.940 201.120 ;
        RECT 9.580 200.420 30.240 200.780 ;
        RECT 3.750 200.100 30.240 200.420 ;
        RECT 3.750 199.760 23.800 200.100 ;
        RECT 26.185 199.895 30.240 200.100 ;
        RECT 30.940 200.285 34.380 200.780 ;
        RECT 30.940 199.895 33.460 200.285 ;
        RECT 26.185 199.760 33.460 199.895 ;
        RECT 34.160 199.895 34.380 200.285 ;
        RECT 35.080 200.420 41.940 200.780 ;
        RECT 49.645 200.420 564.420 201.120 ;
        RECT 35.080 200.080 42.860 200.420 ;
        RECT 47.255 200.080 564.420 200.420 ;
        RECT 35.080 199.895 564.420 200.080 ;
        RECT 34.160 199.760 564.420 199.895 ;
        RECT 3.750 199.060 21.960 199.760 ;
        RECT 26.645 199.060 32.540 199.760 ;
        RECT 3.750 198.720 32.540 199.060 ;
        RECT 33.240 199.400 33.460 199.760 ;
        RECT 33.240 199.060 34.075 199.400 ;
        RECT 48.220 199.060 564.420 199.760 ;
        RECT 33.240 198.720 564.420 199.060 ;
        RECT 3.750 198.060 564.420 198.720 ;
        RECT 3.750 197.720 31.315 198.060 ;
        RECT 40.400 197.720 564.420 198.060 ;
        RECT 3.750 196.835 30.700 197.720 ;
        RECT 40.400 197.360 52.935 197.720 ;
        RECT 32.165 197.020 52.935 197.360 ;
        RECT 61.560 197.020 564.420 197.720 ;
        RECT 3.750 196.680 31.360 196.835 ;
        RECT 32.165 196.700 564.420 197.020 ;
        RECT 32.165 196.680 46.495 196.700 ;
        RECT 3.750 196.000 46.495 196.680 ;
        RECT 49.140 196.000 564.420 196.700 ;
        RECT 3.750 195.000 564.420 196.000 ;
        RECT 3.750 194.300 50.940 195.000 ;
        RECT 52.405 194.320 564.420 195.000 ;
        RECT 3.750 193.980 51.400 194.300 ;
        RECT 3.750 193.280 7.855 193.980 ;
        RECT 17.860 193.620 51.400 193.980 ;
        RECT 53.280 193.620 55.540 194.320 ;
        RECT 60.640 193.620 564.420 194.320 ;
        RECT 17.860 193.280 564.420 193.620 ;
        RECT 3.750 192.280 564.420 193.280 ;
        RECT 3.750 191.395 30.240 192.280 ;
        RECT 30.940 191.785 564.420 192.280 ;
        RECT 30.940 191.395 31.160 191.785 ;
        RECT 3.750 190.900 31.160 191.395 ;
        RECT 31.860 190.900 564.420 191.785 ;
        RECT 3.750 190.240 564.420 190.900 ;
        RECT 3.750 189.540 28.600 190.240 ;
        RECT 30.280 189.560 564.420 190.240 ;
        RECT 30.280 189.540 33.615 189.560 ;
        RECT 3.750 188.860 33.615 189.540 ;
        RECT 34.420 188.880 34.535 189.560 ;
        RECT 38.100 188.880 564.420 189.560 ;
        RECT 3.750 188.180 34.075 188.860 ;
        RECT 54.660 188.180 564.420 188.880 ;
        RECT 3.750 186.840 564.420 188.180 ;
        RECT 3.750 186.160 55.695 186.840 ;
        RECT 3.750 185.460 52.015 186.160 ;
        RECT 52.820 186.140 55.695 186.160 ;
        RECT 57.880 186.140 564.420 186.840 ;
        RECT 52.820 185.820 564.420 186.140 ;
        RECT 52.820 185.460 53.345 185.820 ;
        RECT 3.750 185.120 53.345 185.460 ;
        RECT 68.000 185.120 564.420 185.820 ;
        RECT 3.750 184.800 564.420 185.120 ;
        RECT 3.750 184.460 49.760 184.800 ;
        RECT 3.750 183.760 41.480 184.460 ;
        RECT 43.620 184.100 49.760 184.460 ;
        RECT 66.620 184.100 564.420 184.800 ;
        RECT 43.620 183.760 50.680 184.100 ;
        RECT 61.100 183.760 564.420 184.100 ;
        RECT 3.750 183.440 564.420 183.760 ;
        RECT 3.750 182.740 44.195 183.440 ;
        RECT 50.980 182.740 564.420 183.440 ;
        RECT 3.750 163.040 564.420 182.740 ;
        RECT 3.750 162.340 17.100 163.040 ;
        RECT 46.425 162.340 564.420 163.040 ;
        RECT 3.750 156.920 564.420 162.340 ;
        RECT 3.750 156.220 18.895 156.920 ;
        RECT 19.700 156.220 564.420 156.920 ;
        RECT 3.750 151.820 564.420 156.220 ;
        RECT 3.750 150.935 16.900 151.820 ;
        RECT 17.600 150.935 564.420 151.820 ;
        RECT 3.750 150.460 564.420 150.935 ;
        RECT 3.750 149.760 46.035 150.460 ;
        RECT 46.840 149.760 564.420 150.460 ;
        RECT 3.750 148.420 564.420 149.760 ;
        RECT 3.750 147.720 19.355 148.420 ;
        RECT 21.080 147.720 564.420 148.420 ;
        RECT 3.750 146.380 564.420 147.720 ;
        RECT 3.750 146.040 50.220 146.380 ;
        RECT 55.165 146.040 564.420 146.380 ;
        RECT 3.750 145.340 15.215 146.040 ;
        RECT 16.940 145.340 49.560 146.040 ;
        RECT 56.960 145.340 564.420 146.040 ;
        RECT 3.750 144.000 564.420 145.340 ;
        RECT 3.750 143.660 56.000 144.000 ;
        RECT 3.750 142.980 45.115 143.660 ;
        RECT 3.750 142.280 33.660 142.980 ;
        RECT 47.300 142.960 56.000 143.660 ;
        RECT 46.885 142.435 56.000 142.960 ;
        RECT 56.700 142.435 564.420 144.000 ;
        RECT 46.885 142.280 564.420 142.435 ;
        RECT 3.750 141.940 43.320 142.280 ;
        RECT 45.505 141.940 564.420 142.280 ;
        RECT 3.750 140.600 564.420 141.940 ;
        RECT 3.750 139.900 36.420 140.600 ;
        RECT 40.905 139.900 564.420 140.600 ;
        RECT 3.750 139.580 564.420 139.900 ;
        RECT 3.750 138.880 40.515 139.580 ;
        RECT 50.060 138.880 564.420 139.580 ;
        RECT 3.750 137.880 564.420 138.880 ;
        RECT 3.750 136.995 15.980 137.880 ;
        RECT 16.680 137.540 564.420 137.880 ;
        RECT 16.680 137.200 47.920 137.540 ;
        RECT 53.785 137.200 564.420 137.540 ;
        RECT 16.680 136.995 47.260 137.200 ;
        RECT 3.750 136.500 47.260 136.995 ;
        RECT 56.545 136.500 564.420 137.200 ;
        RECT 3.750 135.840 564.420 136.500 ;
        RECT 3.750 134.615 55.080 135.840 ;
        RECT 55.780 134.615 564.420 135.840 ;
        RECT 3.750 132.100 564.420 134.615 ;
        RECT 3.750 131.760 56.615 132.100 ;
        RECT 3.750 131.060 50.635 131.760 ;
        RECT 54.660 131.400 56.615 131.760 ;
        RECT 57.420 131.400 564.420 132.100 ;
        RECT 54.660 131.060 564.420 131.400 ;
        RECT 3.750 118.840 564.420 131.060 ;
        RECT 3.750 118.500 44.655 118.840 ;
        RECT 3.750 117.800 41.480 118.500 ;
        RECT 44.080 118.140 44.655 118.500 ;
        RECT 47.960 118.140 564.420 118.840 ;
        RECT 44.080 117.820 564.420 118.140 ;
        RECT 44.080 117.800 45.575 117.820 ;
        RECT 3.750 117.120 45.575 117.800 ;
        RECT 50.060 117.120 564.420 117.820 ;
        RECT 3.750 115.780 564.420 117.120 ;
        RECT 3.750 115.080 52.520 115.780 ;
        RECT 57.005 115.080 564.420 115.780 ;
        RECT 3.750 112.380 564.420 115.080 ;
        RECT 3.750 111.680 51.095 112.380 ;
        RECT 56.960 111.680 564.420 112.380 ;
        RECT 3.750 111.020 564.420 111.680 ;
        RECT 3.750 110.320 52.015 111.020 ;
        RECT 53.280 110.320 564.420 111.020 ;
        RECT 3.750 109.660 564.420 110.320 ;
        RECT 3.750 108.960 7.855 109.660 ;
        RECT 9.580 108.960 564.420 109.660 ;
        RECT 3.750 97.420 564.420 108.960 ;
        RECT 3.750 96.720 7.395 97.420 ;
        RECT 20.160 96.720 564.420 97.420 ;
        RECT 3.750 91.980 564.420 96.720 ;
        RECT 3.750 91.280 7.395 91.980 ;
        RECT 11.880 91.280 564.420 91.980 ;
        RECT 3.750 86.540 564.420 91.280 ;
        RECT 3.750 85.840 7.395 86.540 ;
        RECT 10.500 85.840 564.420 86.540 ;
        RECT 3.750 81.100 564.420 85.840 ;
        RECT 3.750 80.400 7.395 81.100 ;
        RECT 21.540 80.400 564.420 81.100 ;
        RECT 3.750 77.700 564.420 80.400 ;
        RECT 3.750 77.000 7.395 77.700 ;
        RECT 10.960 77.000 564.420 77.700 ;
        RECT 3.750 61.380 564.420 77.000 ;
        RECT 3.750 60.680 7.395 61.380 ;
        RECT 17.400 61.040 564.420 61.380 ;
        RECT 17.400 60.680 50.680 61.040 ;
        RECT 3.750 60.340 50.680 60.680 ;
        RECT 54.860 60.700 564.420 61.040 ;
        RECT 54.860 60.340 57.995 60.700 ;
        RECT 3.750 60.000 57.995 60.340 ;
        RECT 61.100 60.000 564.420 60.700 ;
        RECT 3.750 59.340 564.420 60.000 ;
        RECT 3.750 58.640 7.395 59.340 ;
        RECT 23.840 59.000 564.420 59.340 ;
        RECT 23.840 58.640 64.020 59.000 ;
        RECT 3.750 58.300 64.020 58.640 ;
        RECT 67.540 58.300 564.420 59.000 ;
        RECT 3.750 48.460 564.420 58.300 ;
        RECT 3.750 47.760 7.395 48.460 ;
        RECT 20.620 47.780 564.420 48.460 ;
        RECT 3.750 47.080 7.440 47.760 ;
        RECT 28.440 47.080 564.420 47.780 ;
        RECT 3.750 34.180 564.420 47.080 ;
        RECT 3.750 33.480 7.395 34.180 ;
        RECT 29.820 33.480 564.420 34.180 ;
        RECT 3.750 30.100 564.420 33.480 ;
        RECT 3.750 29.400 63.560 30.100 ;
        RECT 70.760 29.400 564.420 30.100 ;
        RECT 3.750 28.740 564.420 29.400 ;
        RECT 3.750 28.040 7.395 28.740 ;
        RECT 18.320 28.040 564.420 28.740 ;
        RECT 3.750 24.320 564.420 28.040 ;
        RECT 3.750 23.640 165.635 24.320 ;
        RECT 3.750 23.300 52.980 23.640 ;
        RECT 90.125 23.620 165.635 23.640 ;
        RECT 166.440 23.620 183.115 24.320 ;
        RECT 183.920 23.620 564.420 24.320 ;
        RECT 90.125 23.300 564.420 23.620 ;
        RECT 3.750 22.600 7.395 23.300 ;
        RECT 9.120 22.940 52.980 23.300 ;
        RECT 9.120 22.600 64.940 22.940 ;
        RECT 91.505 22.600 181.780 23.300 ;
        RECT 184.885 22.600 564.420 23.300 ;
        RECT 3.750 22.260 182.240 22.600 ;
        RECT 183.045 22.260 564.420 22.600 ;
        RECT 3.750 20.580 564.420 22.260 ;
        RECT 3.750 20.425 199.980 20.580 ;
        RECT 3.750 19.540 166.400 20.425 ;
        RECT 167.100 19.540 199.980 20.425 ;
        RECT 200.680 19.540 564.420 20.580 ;
        RECT 3.750 13.440 564.420 19.540 ;
        RECT 3.750 12.740 38.720 13.440 ;
        RECT 559.280 12.740 564.420 13.440 ;
        RECT 3.750 5.200 564.420 12.740 ;
      LAYER met2 ;
        RECT 3.770 445.720 563.840 449.130 ;
        RECT 3.770 445.040 67.500 445.720 ;
        RECT 3.770 438.240 66.580 445.040 ;
        RECT 3.770 388.290 65.660 438.240 ;
        RECT 3.770 387.590 8.160 388.290 ;
        RECT 9.780 387.590 65.660 388.290 ;
        RECT 3.770 384.520 65.660 387.590 ;
        RECT 3.770 382.360 8.160 384.520 ;
        RECT 8.860 382.360 65.660 384.520 ;
        RECT 3.770 381.800 65.660 382.360 ;
        RECT 3.770 379.640 8.160 381.800 ;
        RECT 8.860 380.440 65.660 381.800 ;
        RECT 8.860 379.640 46.800 380.440 ;
        RECT 3.770 360.420 46.800 379.640 ;
        RECT 47.500 377.040 65.660 380.440 ;
        RECT 47.500 373.300 56.920 377.040 ;
        RECT 47.500 365.520 54.160 373.300 ;
        RECT 54.860 371.300 56.920 373.300 ;
        RECT 57.620 371.300 65.660 377.040 ;
        RECT 54.860 365.520 65.660 371.300 ;
        RECT 47.500 360.420 65.660 365.520 ;
        RECT 3.770 354.600 65.660 360.420 ;
        RECT 3.770 352.940 43.580 354.600 ;
        RECT 44.280 352.940 65.660 354.600 ;
        RECT 3.770 346.440 65.660 352.940 ;
        RECT 3.770 345.640 13.220 346.440 ;
        RECT 13.920 345.640 65.660 346.440 ;
        RECT 3.770 338.620 65.660 345.640 ;
        RECT 3.770 337.940 42.660 338.620 ;
        RECT 3.770 335.940 35.760 337.940 ;
        RECT 36.460 336.620 42.660 337.940 ;
        RECT 43.360 336.620 65.660 338.620 ;
        RECT 36.460 335.940 65.660 336.620 ;
        RECT 3.770 333.380 65.660 335.940 ;
        RECT 3.770 332.680 43.580 333.380 ;
        RECT 44.740 332.680 65.660 333.380 ;
        RECT 3.770 332.530 65.660 332.680 ;
        RECT 3.770 331.830 59.220 332.530 ;
        RECT 60.380 331.830 65.660 332.530 ;
        RECT 3.770 328.420 65.660 331.830 ;
        RECT 3.770 327.060 62.900 328.420 ;
        RECT 3.770 316.900 37.600 327.060 ;
        RECT 38.300 318.900 62.900 327.060 ;
        RECT 38.300 316.900 39.440 318.900 ;
        RECT 3.770 309.080 39.440 316.900 ;
        RECT 40.140 309.080 62.900 318.900 ;
        RECT 3.770 305.640 62.900 309.080 ;
        RECT 3.770 301.260 7.240 305.640 ;
        RECT 7.940 303.260 62.900 305.640 ;
        RECT 7.940 301.560 47.260 303.260 ;
        RECT 7.940 301.260 39.440 301.560 ;
        RECT 3.770 299.860 39.440 301.260 ;
        RECT 3.770 289.690 16.440 299.860 ;
        RECT 3.770 288.990 8.160 289.690 ;
        RECT 9.320 288.990 16.440 289.690 ;
        RECT 3.770 288.330 16.440 288.990 ;
        RECT 3.770 287.630 6.780 288.330 ;
        RECT 8.860 287.630 16.440 288.330 ;
        RECT 3.770 278.100 16.440 287.630 ;
        RECT 17.140 286.260 22.420 299.860 ;
        RECT 3.770 243.800 7.240 278.100 ;
        RECT 7.940 271.000 16.440 278.100 ;
        RECT 17.600 276.440 22.420 286.260 ;
        RECT 23.120 297.520 39.440 299.860 ;
        RECT 40.140 298.540 47.260 301.560 ;
        RECT 47.960 298.540 62.900 303.260 ;
        RECT 40.140 297.520 62.900 298.540 ;
        RECT 23.120 295.810 62.900 297.520 ;
        RECT 23.120 295.110 56.000 295.810 ;
        RECT 57.620 295.110 62.900 295.810 ;
        RECT 23.120 281.530 62.900 295.110 ;
        RECT 23.120 280.830 50.940 281.530 ;
        RECT 53.020 280.830 62.900 281.530 ;
        RECT 23.120 279.490 62.900 280.830 ;
        RECT 23.120 278.790 23.800 279.490 ;
        RECT 27.260 278.790 48.180 279.490 ;
        RECT 49.340 278.790 62.900 279.490 ;
        RECT 23.120 278.100 62.900 278.790 ;
        RECT 7.940 256.720 16.900 271.000 ;
        RECT 17.600 261.820 22.880 276.440 ;
        RECT 23.580 273.720 62.900 278.100 ;
        RECT 63.600 316.900 65.660 328.420 ;
        RECT 66.360 330.680 66.580 438.240 ;
        RECT 67.280 351.240 67.500 445.040 ;
        RECT 68.200 442.320 563.840 445.720 ;
        RECT 68.200 437.260 206.880 442.320 ;
        RECT 207.580 437.260 563.840 442.320 ;
        RECT 68.200 377.380 563.840 437.260 ;
        RECT 68.200 351.240 68.880 377.380 ;
        RECT 67.280 330.680 68.880 351.240 ;
        RECT 66.360 316.900 68.880 330.680 ;
        RECT 63.600 308.740 68.880 316.900 ;
        RECT 69.580 308.740 563.840 377.380 ;
        RECT 63.600 273.720 563.840 308.740 ;
        RECT 23.580 261.820 563.840 273.720 ;
        RECT 17.600 256.720 563.840 261.820 ;
        RECT 7.940 245.800 563.840 256.720 ;
        RECT 7.940 243.800 48.640 245.800 ;
        RECT 3.770 237.990 48.640 243.800 ;
        RECT 49.340 237.990 563.840 245.800 ;
        RECT 3.770 229.140 563.840 237.990 ;
        RECT 3.770 220.980 29.780 229.140 ;
        RECT 3.770 136.660 7.700 220.980 ;
        RECT 8.400 214.220 29.780 220.980 ;
        RECT 30.480 224.410 563.840 229.140 ;
        RECT 30.480 221.360 41.740 224.410 ;
        RECT 42.440 221.360 563.840 224.410 ;
        RECT 30.480 214.220 563.840 221.360 ;
        RECT 8.400 206.520 563.840 214.220 ;
        RECT 8.400 203.000 28.860 206.520 ;
        RECT 29.560 205.340 563.840 206.520 ;
        RECT 29.560 203.000 33.000 205.340 ;
        RECT 8.400 200.240 33.000 203.000 ;
        RECT 8.400 197.900 29.320 200.240 ;
        RECT 30.020 199.940 33.000 200.240 ;
        RECT 33.700 202.650 563.840 205.340 ;
        RECT 33.700 201.950 51.860 202.650 ;
        RECT 53.480 201.950 563.840 202.650 ;
        RECT 33.700 199.940 563.840 201.950 ;
        RECT 30.020 197.900 563.840 199.940 ;
        RECT 8.400 197.210 563.840 197.900 ;
        RECT 8.400 196.510 23.800 197.210 ;
        RECT 24.960 196.510 563.840 197.210 ;
        RECT 8.400 193.810 563.840 196.510 ;
        RECT 8.400 193.110 22.420 193.810 ;
        RECT 23.580 193.110 563.840 193.810 ;
        RECT 8.400 192.920 563.840 193.110 ;
        RECT 8.400 192.450 30.700 192.920 ;
        RECT 8.400 191.750 21.500 192.450 ;
        RECT 23.120 192.120 30.700 192.450 ;
        RECT 31.400 192.120 563.840 192.920 ;
        RECT 23.120 191.750 563.840 192.120 ;
        RECT 8.400 189.730 563.840 191.750 ;
        RECT 8.400 189.030 31.620 189.730 ;
        RECT 32.780 189.030 563.840 189.730 ;
        RECT 8.400 156.040 563.840 189.030 ;
        RECT 8.400 145.530 21.500 156.040 ;
        RECT 8.400 144.830 16.180 145.530 ;
        RECT 17.140 144.830 21.500 145.530 ;
        RECT 3.770 66.320 7.240 136.660 ;
        RECT 8.400 134.660 21.500 144.830 ;
        RECT 22.200 153.660 563.840 156.040 ;
        RECT 22.200 146.220 49.560 153.660 ;
        RECT 50.260 146.220 563.840 153.660 ;
        RECT 22.200 134.660 563.840 146.220 ;
        RECT 8.400 116.300 563.840 134.660 ;
        RECT 7.940 66.320 563.840 116.300 ;
        RECT 3.770 33.640 563.840 66.320 ;
        RECT 3.770 32.440 163.180 33.640 ;
        RECT 3.770 30.620 98.320 32.440 ;
        RECT 99.020 30.620 163.180 32.440 ;
        RECT 3.770 23.600 163.180 30.620 ;
        RECT 3.770 22.420 159.040 23.600 ;
        RECT 3.770 21.100 94.640 22.420 ;
        RECT 95.340 21.100 159.040 22.420 ;
        RECT 3.770 18.380 159.040 21.100 ;
        RECT 159.740 22.800 163.180 23.600 ;
        RECT 163.880 28.880 563.840 33.640 ;
        RECT 163.880 28.540 303.480 28.880 ;
        RECT 163.880 27.680 296.580 28.540 ;
        RECT 163.880 25.520 180.660 27.680 ;
        RECT 181.360 25.860 186.180 27.680 ;
        RECT 186.880 26.540 193.080 27.680 ;
        RECT 193.780 26.880 199.980 27.680 ;
        RECT 200.680 26.880 201.360 27.680 ;
        RECT 193.780 26.540 201.360 26.880 ;
        RECT 186.880 26.200 201.360 26.540 ;
        RECT 202.060 26.200 220.680 27.680 ;
        RECT 186.880 25.860 220.680 26.200 ;
        RECT 181.360 25.520 220.680 25.860 ;
        RECT 163.880 23.600 220.680 25.520 ;
        RECT 163.880 22.800 166.400 23.600 ;
        RECT 159.740 18.380 166.400 22.800 ;
        RECT 3.770 12.600 166.400 18.380 ;
        RECT 167.100 22.920 220.680 23.600 ;
        RECT 167.100 22.760 213.780 22.920 ;
        RECT 167.100 21.100 172.380 22.760 ;
        RECT 173.080 21.100 213.780 22.760 ;
        RECT 167.100 21.060 213.780 21.100 ;
        RECT 167.100 20.430 203.200 21.060 ;
        RECT 167.100 20.380 199.585 20.430 ;
        RECT 167.100 15.660 173.760 20.380 ;
        RECT 174.460 19.860 199.585 20.380 ;
        RECT 200.155 19.860 203.200 20.430 ;
        RECT 174.460 17.880 203.200 19.860 ;
        RECT 203.900 17.880 213.780 21.060 ;
        RECT 174.460 15.660 213.780 17.880 ;
        RECT 167.100 12.600 213.780 15.660 ;
        RECT 3.770 12.440 213.780 12.600 ;
        RECT 214.480 18.040 220.680 22.920 ;
        RECT 221.380 24.960 289.680 27.680 ;
        RECT 221.380 18.040 268.980 24.960 ;
        RECT 214.480 16.680 268.980 18.040 ;
        RECT 269.680 17.020 278.640 24.960 ;
        RECT 279.340 22.420 282.780 24.960 ;
        RECT 279.800 20.420 282.780 22.420 ;
        RECT 279.340 17.700 282.780 20.420 ;
        RECT 283.480 18.380 289.680 24.960 ;
        RECT 290.380 27.400 296.580 27.680 ;
        RECT 297.280 27.400 303.480 28.540 ;
        RECT 304.180 28.200 563.840 28.880 ;
        RECT 304.180 27.400 310.380 28.200 ;
        RECT 311.080 27.680 563.840 28.200 ;
        RECT 311.080 27.400 331.080 27.680 ;
        RECT 290.380 19.400 331.080 27.400 ;
        RECT 331.780 23.140 344.880 27.680 ;
        RECT 345.580 24.960 563.840 27.680 ;
        RECT 345.580 23.140 352.240 24.960 ;
        RECT 331.780 22.800 352.240 23.140 ;
        RECT 352.940 22.800 563.840 24.960 ;
        RECT 331.780 19.400 563.840 22.800 ;
        RECT 290.380 18.380 563.840 19.400 ;
        RECT 283.480 17.700 563.840 18.380 ;
        RECT 279.340 17.020 563.840 17.700 ;
        RECT 269.680 16.680 563.840 17.020 ;
        RECT 214.480 12.440 563.840 16.680 ;
        RECT 3.770 0.690 563.840 12.440 ;
        RECT 3.770 0.000 283.240 0.690 ;
        RECT 285.320 0.000 563.840 0.690 ;
      LAYER met3 ;
        RECT 0.310 434.730 563.900 443.865 ;
        RECT 0.310 433.630 50.820 434.730 ;
        RECT 70.410 433.630 563.900 434.730 ;
        RECT 0.310 427.930 563.900 433.630 ;
        RECT 7.850 426.830 563.900 427.930 ;
        RECT 0.310 423.170 563.900 426.830 ;
        RECT 4.170 422.070 563.900 423.170 ;
        RECT 0.310 418.410 563.900 422.070 ;
        RECT 4.170 417.900 563.900 418.410 ;
        RECT 4.170 417.310 535.400 417.900 ;
        RECT 0.310 416.800 535.400 417.310 ;
        RECT 552.030 416.800 563.900 417.900 ;
        RECT 0.310 413.650 563.900 416.800 ;
        RECT 4.460 412.550 563.900 413.650 ;
        RECT 0.310 408.890 563.900 412.550 ;
        RECT 4.170 407.790 563.900 408.890 ;
        RECT 0.310 404.130 563.900 407.790 ;
        RECT 4.170 403.030 563.900 404.130 ;
        RECT 0.310 399.370 563.900 403.030 ;
        RECT 4.460 398.270 563.900 399.370 ;
        RECT 0.310 394.610 563.900 398.270 ;
        RECT 4.170 393.510 563.900 394.610 ;
        RECT 0.310 389.850 563.900 393.510 ;
        RECT 4.170 388.750 563.900 389.850 ;
        RECT 0.310 385.090 563.900 388.750 ;
        RECT 4.170 383.990 563.900 385.090 ;
        RECT 0.310 380.330 563.900 383.990 ;
        RECT 4.170 379.230 563.900 380.330 ;
        RECT 0.310 375.570 563.900 379.230 ;
        RECT 4.170 374.470 563.900 375.570 ;
        RECT 0.310 370.810 563.900 374.470 ;
        RECT 4.170 369.710 563.900 370.810 ;
        RECT 0.310 367.410 563.900 369.710 ;
        RECT 0.310 366.310 52.870 367.410 ;
        RECT 54.060 366.310 563.900 367.410 ;
        RECT 0.310 366.050 563.900 366.310 ;
        RECT 4.170 364.950 563.900 366.050 ;
        RECT 0.310 361.290 563.900 364.950 ;
        RECT 4.170 360.190 563.900 361.290 ;
        RECT 0.310 356.530 563.900 360.190 ;
        RECT 4.170 355.430 563.900 356.530 ;
        RECT 0.310 354.345 563.900 355.430 ;
        RECT 0.310 353.535 48.930 354.345 ;
        RECT 49.740 353.535 563.900 354.345 ;
        RECT 0.310 351.770 563.900 353.535 ;
        RECT 8.140 350.670 563.900 351.770 ;
        RECT 0.310 347.010 563.900 350.670 ;
        RECT 4.170 345.910 563.900 347.010 ;
        RECT 0.310 342.250 563.900 345.910 ;
        RECT 4.170 341.150 563.900 342.250 ;
        RECT 0.310 337.490 563.900 341.150 ;
        RECT 8.140 336.390 563.900 337.490 ;
        RECT 0.310 332.730 563.900 336.390 ;
        RECT 4.170 331.630 563.900 332.730 ;
        RECT 0.310 327.970 563.900 331.630 ;
        RECT 4.170 326.870 563.900 327.970 ;
        RECT 0.310 323.210 563.900 326.870 ;
        RECT 4.690 322.110 563.900 323.210 ;
        RECT 0.310 318.450 563.900 322.110 ;
        RECT 4.170 317.350 563.900 318.450 ;
        RECT 0.310 313.690 563.900 317.350 ;
        RECT 4.170 312.590 563.900 313.690 ;
        RECT 0.310 308.930 563.900 312.590 ;
        RECT 4.170 307.830 563.900 308.930 ;
        RECT 0.310 304.170 563.900 307.830 ;
        RECT 4.630 303.070 563.900 304.170 ;
        RECT 0.310 299.410 563.900 303.070 ;
        RECT 4.630 298.310 563.900 299.410 ;
        RECT 0.310 294.650 563.900 298.310 ;
        RECT 4.630 293.550 563.900 294.650 ;
        RECT 0.310 289.890 563.900 293.550 ;
        RECT 8.310 288.790 563.900 289.890 ;
        RECT 0.310 285.130 563.900 288.790 ;
        RECT 4.630 284.030 563.900 285.130 ;
        RECT 0.310 283.090 563.900 284.030 ;
        RECT 0.310 282.410 48.270 283.090 ;
        RECT 0.310 281.310 43.460 282.410 ;
        RECT 45.570 281.990 48.270 282.410 ;
        RECT 49.460 281.990 563.900 283.090 ;
        RECT 45.570 281.310 563.900 281.990 ;
        RECT 0.310 280.370 563.900 281.310 ;
        RECT 4.630 279.270 563.900 280.370 ;
        RECT 0.310 275.610 563.900 279.270 ;
        RECT 4.630 274.510 563.900 275.610 ;
        RECT 0.310 270.850 563.900 274.510 ;
        RECT 4.630 269.750 563.900 270.850 ;
        RECT 0.310 266.090 563.900 269.750 ;
        RECT 4.630 264.990 563.900 266.090 ;
        RECT 0.310 261.330 563.900 264.990 ;
        RECT 4.690 260.230 563.900 261.330 ;
        RECT 0.310 256.570 563.900 260.230 ;
        RECT 4.630 255.470 563.900 256.570 ;
        RECT 0.310 251.810 563.900 255.470 ;
        RECT 4.630 250.710 563.900 251.810 ;
        RECT 0.310 247.050 563.900 250.710 ;
        RECT 8.310 245.950 563.900 247.050 ;
        RECT 0.310 242.290 563.900 245.950 ;
        RECT 4.630 241.190 563.900 242.290 ;
        RECT 0.310 237.530 563.900 241.190 ;
        RECT 4.630 236.430 563.900 237.530 ;
        RECT 0.310 232.770 563.900 236.430 ;
        RECT 4.630 231.670 563.900 232.770 ;
        RECT 0.310 228.010 563.900 231.670 ;
        RECT 7.390 226.910 563.900 228.010 ;
        RECT 0.310 223.250 563.900 226.910 ;
        RECT 4.170 222.150 563.900 223.250 ;
        RECT 0.310 218.490 563.900 222.150 ;
        RECT 4.170 217.390 563.900 218.490 ;
        RECT 0.310 213.730 563.900 217.390 ;
        RECT 4.170 212.630 563.900 213.730 ;
        RECT 0.310 208.970 563.900 212.630 ;
        RECT 4.170 207.870 563.900 208.970 ;
        RECT 0.310 206.250 563.900 207.870 ;
        RECT 0.310 205.150 60.230 206.250 ;
        RECT 70.710 205.150 563.900 206.250 ;
        RECT 0.310 204.210 563.900 205.150 ;
        RECT 4.170 203.110 563.900 204.210 ;
        RECT 0.310 199.450 563.900 203.110 ;
        RECT 4.690 198.350 563.900 199.450 ;
        RECT 0.310 195.370 563.900 198.350 ;
        RECT 0.310 194.690 49.190 195.370 ;
        RECT 4.170 194.270 49.190 194.690 ;
        RECT 66.020 194.270 563.900 195.370 ;
        RECT 4.170 193.590 563.900 194.270 ;
        RECT 0.310 193.330 563.900 193.590 ;
        RECT 0.310 192.230 59.770 193.330 ;
        RECT 70.710 192.230 563.900 193.330 ;
        RECT 0.310 189.930 563.900 192.230 ;
        RECT 4.170 188.830 563.900 189.930 ;
        RECT 0.310 185.850 563.900 188.830 ;
        RECT 0.310 185.170 58.390 185.850 ;
        RECT 4.170 184.750 58.390 185.170 ;
        RECT 70.710 184.750 563.900 185.850 ;
        RECT 4.170 184.070 563.900 184.750 ;
        RECT 0.310 180.410 563.900 184.070 ;
        RECT 4.170 179.310 563.900 180.410 ;
        RECT 0.310 179.050 563.900 179.310 ;
        RECT 0.310 177.950 58.850 179.050 ;
        RECT 70.710 177.950 563.900 179.050 ;
        RECT 0.310 175.650 563.900 177.950 ;
        RECT 4.170 174.550 563.900 175.650 ;
        RECT 0.310 172.700 563.900 174.550 ;
        RECT 0.310 171.890 55.025 172.700 ;
        RECT 55.835 171.890 563.900 172.700 ;
        RECT 0.310 170.890 563.900 171.890 ;
        RECT 1.930 169.790 563.900 170.890 ;
        RECT 0.310 166.130 563.900 169.790 ;
        RECT 7.850 165.030 563.900 166.130 ;
        RECT 0.310 161.370 563.900 165.030 ;
        RECT 4.170 160.270 563.900 161.370 ;
        RECT 0.310 156.610 563.900 160.270 ;
        RECT 4.170 155.510 563.900 156.610 ;
        RECT 0.310 151.850 563.900 155.510 ;
        RECT 7.390 150.750 563.900 151.850 ;
        RECT 0.310 147.090 563.900 150.750 ;
        RECT 4.170 145.990 563.900 147.090 ;
        RECT 0.310 142.330 563.900 145.990 ;
        RECT 4.170 141.230 563.900 142.330 ;
        RECT 0.310 137.570 563.900 141.230 ;
        RECT 4.170 136.470 563.900 137.570 ;
        RECT 0.310 132.810 563.900 136.470 ;
        RECT 4.170 131.710 563.900 132.810 ;
        RECT 0.310 128.050 563.900 131.710 ;
        RECT 4.170 126.950 563.900 128.050 ;
        RECT 0.310 123.290 563.900 126.950 ;
        RECT 4.170 122.190 563.900 123.290 ;
        RECT 0.310 118.700 563.900 122.190 ;
        RECT 0.310 118.530 484.510 118.700 ;
        RECT 4.170 117.600 484.510 118.530 ;
        RECT 553.010 117.600 563.900 118.700 ;
        RECT 4.170 117.430 563.900 117.600 ;
        RECT 0.310 113.770 563.900 117.430 ;
        RECT 4.170 112.670 563.900 113.770 ;
        RECT 0.310 109.010 563.900 112.670 ;
        RECT 4.170 107.910 563.900 109.010 ;
        RECT 0.310 104.250 563.900 107.910 ;
        RECT 4.170 103.740 563.900 104.250 ;
        RECT 4.170 103.150 483.720 103.740 ;
        RECT 0.310 102.640 483.720 103.150 ;
        RECT 553.010 102.640 563.900 103.740 ;
        RECT 0.310 99.490 563.900 102.640 ;
        RECT 4.170 98.390 563.900 99.490 ;
        RECT 0.310 94.730 563.900 98.390 ;
        RECT 4.630 93.630 563.900 94.730 ;
        RECT 0.310 89.970 563.900 93.630 ;
        RECT 8.310 88.870 563.900 89.970 ;
        RECT 0.310 85.210 563.900 88.870 ;
        RECT 4.630 84.110 563.900 85.210 ;
        RECT 0.310 80.450 563.900 84.110 ;
        RECT 4.630 79.350 563.900 80.450 ;
        RECT 0.310 75.690 563.900 79.350 ;
        RECT 4.690 74.590 563.900 75.690 ;
        RECT 0.310 73.650 563.900 74.590 ;
        RECT 0.310 70.930 69.610 73.650 ;
        RECT 4.630 69.830 69.610 70.930 ;
        RECT 0.310 66.170 69.610 69.830 ;
        RECT 4.630 65.070 69.610 66.170 ;
        RECT 0.310 62.480 69.610 65.070 ;
        RECT 70.710 62.480 563.900 73.650 ;
        RECT 0.310 61.410 563.900 62.480 ;
        RECT 4.630 60.310 563.900 61.410 ;
        RECT 0.310 56.650 563.900 60.310 ;
        RECT 4.630 55.550 563.900 56.650 ;
        RECT 0.310 51.890 563.900 55.550 ;
        RECT 4.630 50.790 563.900 51.890 ;
        RECT 0.310 47.130 563.900 50.790 ;
        RECT 4.630 46.030 563.900 47.130 ;
        RECT 0.310 42.370 563.900 46.030 ;
        RECT 4.630 41.270 563.900 42.370 ;
        RECT 0.310 37.610 563.900 41.270 ;
        RECT 4.630 36.510 563.900 37.610 ;
        RECT 0.310 33.530 563.900 36.510 ;
        RECT 0.310 32.850 96.510 33.530 ;
        RECT 4.630 31.750 96.510 32.850 ;
        RECT 97.610 31.750 563.900 33.530 ;
        RECT 0.310 28.090 563.900 31.750 ;
        RECT 8.310 26.990 563.900 28.090 ;
        RECT 0.310 23.950 563.900 26.990 ;
        RECT 0.310 23.330 185.665 23.950 ;
        RECT 4.630 23.140 185.665 23.330 ;
        RECT 186.475 23.140 563.900 23.950 ;
        RECT 4.630 22.230 563.900 23.140 ;
        RECT 0.310 5.275 563.900 22.230 ;
      LAYER met4 ;
        RECT 11.335 12.415 14.320 443.865 ;
        RECT 16.720 12.415 24.320 443.865 ;
        RECT 26.720 12.415 34.320 443.865 ;
        RECT 36.720 12.415 44.320 443.865 ;
        RECT 46.720 299.265 54.320 443.865 ;
        RECT 46.720 298.455 47.780 299.265 ;
        RECT 48.590 298.455 54.320 299.265 ;
        RECT 46.720 12.415 54.320 298.455 ;
        RECT 56.720 434.730 548.420 443.865 ;
        RECT 56.720 434.420 334.840 434.730 ;
        RECT 56.720 434.050 322.600 434.420 ;
        RECT 56.720 405.550 210.400 434.050 ;
        RECT 211.500 405.550 217.200 434.050 ;
        RECT 218.300 405.550 222.640 434.050 ;
        RECT 223.740 405.550 248.480 434.050 ;
        RECT 249.580 405.550 260.720 434.050 ;
        RECT 261.820 405.550 272.960 434.050 ;
        RECT 274.060 405.550 279.080 434.050 ;
        RECT 280.180 405.550 285.880 434.050 ;
        RECT 286.980 405.550 291.320 434.050 ;
        RECT 292.420 405.550 297.440 434.050 ;
        RECT 298.540 433.740 310.360 434.050 ;
        RECT 298.540 405.550 304.240 433.740 ;
        RECT 305.340 405.550 310.360 433.740 ;
        RECT 311.460 405.550 317.160 434.050 ;
        RECT 318.260 405.550 322.600 434.050 ;
        RECT 323.700 405.550 334.840 434.420 ;
        RECT 335.940 405.550 360.680 434.730 ;
        RECT 361.780 434.050 548.420 434.730 ;
        RECT 361.780 405.550 372.920 434.050 ;
        RECT 374.020 405.550 379.040 434.050 ;
        RECT 380.140 405.550 385.840 434.050 ;
        RECT 386.940 405.550 391.280 434.050 ;
        RECT 392.380 405.550 397.400 434.050 ;
        RECT 398.500 405.550 404.200 434.050 ;
        RECT 405.300 414.390 466.760 434.050 ;
        RECT 467.860 417.110 519.800 434.050 ;
        RECT 520.900 417.110 548.420 434.050 ;
        RECT 467.860 414.390 548.420 417.110 ;
        RECT 405.300 405.550 548.420 414.390 ;
        RECT 56.720 35.050 548.420 405.550 ;
        RECT 56.720 25.420 210.590 35.050 ;
        RECT 56.720 12.415 64.320 25.420 ;
        RECT 66.720 12.415 74.320 25.420 ;
        RECT 76.720 12.415 84.320 25.420 ;
        RECT 86.720 12.415 94.320 25.420 ;
        RECT 96.720 12.415 104.320 25.420 ;
        RECT 106.720 12.415 114.320 25.420 ;
        RECT 116.720 12.415 124.320 25.420 ;
        RECT 126.720 12.415 134.320 25.420 ;
        RECT 136.720 12.415 144.320 25.420 ;
        RECT 146.720 12.415 154.320 25.420 ;
        RECT 156.720 25.120 184.320 25.420 ;
        RECT 156.720 24.800 174.320 25.120 ;
        RECT 156.720 12.415 164.320 24.800 ;
        RECT 166.720 12.415 174.320 24.800 ;
        RECT 176.720 12.415 184.320 25.120 ;
        RECT 186.720 24.885 210.590 25.420 ;
        RECT 186.720 12.415 194.320 24.885 ;
        RECT 196.720 24.800 210.590 24.885 ;
        RECT 196.720 12.415 204.320 24.800 ;
        RECT 206.720 19.820 210.590 24.800 ;
        RECT 211.690 32.850 482.910 35.050 ;
        RECT 484.010 32.850 485.670 35.050 ;
        RECT 486.770 34.580 548.420 35.050 ;
        RECT 211.690 27.300 226.230 32.850 ;
        RECT 227.330 27.300 482.910 32.850 ;
        RECT 211.690 25.940 482.910 27.300 ;
        RECT 484.930 26.620 485.670 32.850 ;
        RECT 211.690 25.420 483.830 25.940 ;
        RECT 211.690 24.885 224.320 25.420 ;
        RECT 211.690 19.820 214.320 24.885 ;
        RECT 206.720 12.415 214.320 19.820 ;
        RECT 216.720 12.415 224.320 24.885 ;
        RECT 226.720 24.885 244.320 25.420 ;
        RECT 226.720 12.415 234.320 24.885 ;
        RECT 236.720 12.415 244.320 24.885 ;
        RECT 246.720 25.120 324.320 25.420 ;
        RECT 246.720 24.885 274.320 25.120 ;
        RECT 246.720 12.415 254.320 24.885 ;
        RECT 256.720 24.800 274.320 24.885 ;
        RECT 256.720 12.415 264.320 24.800 ;
        RECT 266.720 12.415 274.320 24.800 ;
        RECT 276.720 24.885 324.320 25.120 ;
        RECT 276.720 24.800 294.320 24.885 ;
        RECT 276.720 12.415 284.320 24.800 ;
        RECT 286.720 12.415 294.320 24.800 ;
        RECT 296.720 24.800 314.320 24.885 ;
        RECT 296.720 12.415 304.320 24.800 ;
        RECT 306.720 12.415 314.320 24.800 ;
        RECT 316.720 12.415 324.320 24.885 ;
        RECT 326.720 24.885 374.320 25.420 ;
        RECT 326.720 12.415 334.320 24.885 ;
        RECT 336.720 24.800 354.320 24.885 ;
        RECT 336.720 12.415 344.320 24.800 ;
        RECT 346.720 12.415 354.320 24.800 ;
        RECT 356.720 24.800 374.320 24.885 ;
        RECT 356.720 12.415 364.320 24.800 ;
        RECT 366.720 12.415 374.320 24.800 ;
        RECT 376.720 24.800 394.320 25.420 ;
        RECT 376.720 12.415 384.320 24.800 ;
        RECT 386.720 12.415 394.320 24.800 ;
        RECT 396.720 24.800 414.320 25.420 ;
        RECT 396.720 12.415 404.320 24.800 ;
        RECT 406.720 12.415 414.320 24.800 ;
        RECT 416.720 12.415 424.320 25.420 ;
        RECT 426.720 12.415 434.320 25.420 ;
        RECT 436.720 12.415 444.320 25.420 ;
        RECT 446.720 12.415 454.320 25.420 ;
        RECT 456.720 12.415 464.320 25.420 ;
        RECT 466.720 12.415 474.320 25.420 ;
        RECT 476.720 25.260 483.830 25.420 ;
        RECT 484.930 25.260 486.590 26.620 ;
        RECT 476.720 24.800 486.590 25.260 ;
        RECT 487.690 25.420 548.420 34.580 ;
        RECT 476.720 12.415 484.320 24.800 ;
        RECT 487.690 20.500 494.320 25.420 ;
        RECT 486.720 12.415 494.320 20.500 ;
        RECT 496.720 12.415 504.320 25.420 ;
        RECT 506.720 12.415 514.320 25.420 ;
        RECT 516.720 12.415 524.320 25.420 ;
        RECT 526.720 12.415 534.320 25.420 ;
        RECT 536.720 12.415 544.320 25.420 ;
        RECT 546.720 12.415 548.420 25.420 ;
  END
END BlockRAM_1KB
END LIBRARY

