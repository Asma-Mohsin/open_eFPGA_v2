magic
tech sky130A
magscale 1 2
timestamp 1733761843
<< obsli1 >>
rect 1104 1071 43516 88689
<< obsm1 >>
rect 14 484 44698 89820
<< metal2 >>
rect 5170 89840 5226 90040
rect 5446 89840 5502 90040
rect 5722 89840 5778 90040
rect 5998 89840 6054 90040
rect 6274 89840 6330 90040
rect 6550 89840 6606 90040
rect 6826 89840 6882 90040
rect 7102 89840 7158 90040
rect 7378 89840 7434 90040
rect 7654 89840 7710 90040
rect 7930 89840 7986 90040
rect 8206 89840 8262 90040
rect 8482 89840 8538 90040
rect 8758 89840 8814 90040
rect 9034 89840 9090 90040
rect 9310 89840 9366 90040
rect 9586 89840 9642 90040
rect 9862 89840 9918 90040
rect 10138 89840 10194 90040
rect 10414 89840 10470 90040
rect 10690 89840 10746 90040
rect 10966 89840 11022 90040
rect 11242 89840 11298 90040
rect 11518 89840 11574 90040
rect 11794 89840 11850 90040
rect 12070 89840 12126 90040
rect 12346 89840 12402 90040
rect 12622 89840 12678 90040
rect 12898 89840 12954 90040
rect 13174 89840 13230 90040
rect 13450 89840 13506 90040
rect 13726 89840 13782 90040
rect 14002 89840 14058 90040
rect 14278 89840 14334 90040
rect 14554 89840 14610 90040
rect 14830 89840 14886 90040
rect 15106 89840 15162 90040
rect 15382 89840 15438 90040
rect 15658 89840 15714 90040
rect 15934 89840 15990 90040
rect 16210 89840 16266 90040
rect 16486 89840 16542 90040
rect 16762 89840 16818 90040
rect 17038 89840 17094 90040
rect 17314 89840 17370 90040
rect 17590 89840 17646 90040
rect 17866 89840 17922 90040
rect 18142 89840 18198 90040
rect 18418 89840 18474 90040
rect 18694 89840 18750 90040
rect 18970 89840 19026 90040
rect 19246 89840 19302 90040
rect 19522 89840 19578 90040
rect 19798 89840 19854 90040
rect 20074 89840 20130 90040
rect 20350 89840 20406 90040
rect 20626 89840 20682 90040
rect 20902 89840 20958 90040
rect 21178 89840 21234 90040
rect 21454 89840 21510 90040
rect 21730 89840 21786 90040
rect 22006 89840 22062 90040
rect 22282 89840 22338 90040
rect 22558 89840 22614 90040
rect 22834 89840 22890 90040
rect 23110 89840 23166 90040
rect 23386 89840 23442 90040
rect 23662 89840 23718 90040
rect 23938 89840 23994 90040
rect 24214 89840 24270 90040
rect 24490 89840 24546 90040
rect 24766 89840 24822 90040
rect 25042 89840 25098 90040
rect 25318 89840 25374 90040
rect 25594 89840 25650 90040
rect 25870 89840 25926 90040
rect 26146 89840 26202 90040
rect 26422 89840 26478 90040
rect 26698 89840 26754 90040
rect 26974 89840 27030 90040
rect 27250 89840 27306 90040
rect 27526 89840 27582 90040
rect 27802 89840 27858 90040
rect 28078 89840 28134 90040
rect 28354 89840 28410 90040
rect 28630 89840 28686 90040
rect 28906 89840 28962 90040
rect 29182 89840 29238 90040
rect 29458 89840 29514 90040
rect 29734 89840 29790 90040
rect 30010 89840 30066 90040
rect 30286 89840 30342 90040
rect 30562 89840 30618 90040
rect 30838 89840 30894 90040
rect 31114 89840 31170 90040
rect 31390 89840 31446 90040
rect 31666 89840 31722 90040
rect 31942 89840 31998 90040
rect 32218 89840 32274 90040
rect 32494 89840 32550 90040
rect 32770 89840 32826 90040
rect 33046 89840 33102 90040
rect 33322 89840 33378 90040
rect 33598 89840 33654 90040
rect 33874 89840 33930 90040
rect 34150 89840 34206 90040
rect 34426 89840 34482 90040
rect 34702 89840 34758 90040
rect 34978 89840 35034 90040
rect 35254 89840 35310 90040
rect 35530 89840 35586 90040
rect 35806 89840 35862 90040
rect 36082 89840 36138 90040
rect 36358 89840 36414 90040
rect 36634 89840 36690 90040
rect 36910 89840 36966 90040
rect 37186 89840 37242 90040
rect 37462 89840 37518 90040
rect 37738 89840 37794 90040
rect 38014 89840 38070 90040
rect 38290 89840 38346 90040
rect 38566 89840 38622 90040
rect 38842 89840 38898 90040
rect 39118 89840 39174 90040
rect 39394 89840 39450 90040
rect 5170 -40 5226 160
rect 5446 -40 5502 160
rect 5722 -40 5778 160
rect 5998 -40 6054 160
rect 6274 -40 6330 160
rect 6550 -40 6606 160
rect 6826 -40 6882 160
rect 7102 -40 7158 160
rect 7378 -40 7434 160
rect 7654 -40 7710 160
rect 7930 -40 7986 160
rect 8206 -40 8262 160
rect 8482 -40 8538 160
rect 8758 -40 8814 160
rect 9034 -40 9090 160
rect 9310 -40 9366 160
rect 9586 -40 9642 160
rect 9862 -40 9918 160
rect 10138 -40 10194 160
rect 10414 -40 10470 160
rect 10690 -40 10746 160
rect 10966 -40 11022 160
rect 11242 -40 11298 160
rect 11518 -40 11574 160
rect 11794 -40 11850 160
rect 12070 -40 12126 160
rect 12346 -40 12402 160
rect 12622 -40 12678 160
rect 12898 -40 12954 160
rect 13174 -40 13230 160
rect 13450 -40 13506 160
rect 13726 -40 13782 160
rect 14002 -40 14058 160
rect 14278 -40 14334 160
rect 14554 -40 14610 160
rect 14830 -40 14886 160
rect 15106 -40 15162 160
rect 15382 -40 15438 160
rect 15658 -40 15714 160
rect 15934 -40 15990 160
rect 16210 -40 16266 160
rect 16486 -40 16542 160
rect 16762 -40 16818 160
rect 17038 -40 17094 160
rect 17314 -40 17370 160
rect 17590 -40 17646 160
rect 17866 -40 17922 160
rect 18142 -40 18198 160
rect 18418 -40 18474 160
rect 18694 -40 18750 160
rect 18970 -40 19026 160
rect 19246 -40 19302 160
rect 19522 -40 19578 160
rect 19798 -40 19854 160
rect 20074 -40 20130 160
rect 20350 -40 20406 160
rect 20626 -40 20682 160
rect 20902 -40 20958 160
rect 21178 -40 21234 160
rect 21454 -40 21510 160
rect 21730 -40 21786 160
rect 22006 -40 22062 160
rect 22282 -40 22338 160
rect 22558 -40 22614 160
rect 22834 -40 22890 160
rect 23110 -40 23166 160
rect 23386 -40 23442 160
rect 23662 -40 23718 160
rect 23938 -40 23994 160
rect 24214 -40 24270 160
rect 24490 -40 24546 160
rect 24766 -40 24822 160
rect 25042 -40 25098 160
rect 25318 -40 25374 160
rect 25594 -40 25650 160
rect 25870 -40 25926 160
rect 26146 -40 26202 160
rect 26422 -40 26478 160
rect 26698 -40 26754 160
rect 26974 -40 27030 160
rect 27250 -40 27306 160
rect 27526 -40 27582 160
rect 27802 -40 27858 160
rect 28078 -40 28134 160
rect 28354 -40 28410 160
rect 28630 -40 28686 160
rect 28906 -40 28962 160
rect 29182 -40 29238 160
rect 29458 -40 29514 160
rect 29734 -40 29790 160
rect 30010 -40 30066 160
rect 30286 -40 30342 160
rect 30562 -40 30618 160
rect 30838 -40 30894 160
rect 31114 -40 31170 160
rect 31390 -40 31446 160
rect 31666 -40 31722 160
rect 31942 -40 31998 160
rect 32218 -40 32274 160
rect 32494 -40 32550 160
rect 32770 -40 32826 160
rect 33046 -40 33102 160
rect 33322 -40 33378 160
rect 33598 -40 33654 160
rect 33874 -40 33930 160
rect 34150 -40 34206 160
rect 34426 -40 34482 160
rect 34702 -40 34758 160
rect 34978 -40 35034 160
rect 35254 -40 35310 160
rect 35530 -40 35586 160
rect 35806 -40 35862 160
rect 36082 -40 36138 160
rect 36358 -40 36414 160
rect 36634 -40 36690 160
rect 36910 -40 36966 160
rect 37186 -40 37242 160
rect 37462 -40 37518 160
rect 37738 -40 37794 160
rect 38014 -40 38070 160
rect 38290 -40 38346 160
rect 38566 -40 38622 160
rect 38842 -40 38898 160
rect 39118 -40 39174 160
rect 39394 -40 39450 160
<< obsm2 >>
rect 20 89784 5114 89978
rect 5282 89784 5390 89978
rect 5558 89784 5666 89978
rect 5834 89784 5942 89978
rect 6110 89784 6218 89978
rect 6386 89784 6494 89978
rect 6662 89784 6770 89978
rect 6938 89784 7046 89978
rect 7214 89784 7322 89978
rect 7490 89784 7598 89978
rect 7766 89784 7874 89978
rect 8042 89784 8150 89978
rect 8318 89784 8426 89978
rect 8594 89784 8702 89978
rect 8870 89784 8978 89978
rect 9146 89784 9254 89978
rect 9422 89784 9530 89978
rect 9698 89784 9806 89978
rect 9974 89784 10082 89978
rect 10250 89784 10358 89978
rect 10526 89784 10634 89978
rect 10802 89784 10910 89978
rect 11078 89784 11186 89978
rect 11354 89784 11462 89978
rect 11630 89784 11738 89978
rect 11906 89784 12014 89978
rect 12182 89784 12290 89978
rect 12458 89784 12566 89978
rect 12734 89784 12842 89978
rect 13010 89784 13118 89978
rect 13286 89784 13394 89978
rect 13562 89784 13670 89978
rect 13838 89784 13946 89978
rect 14114 89784 14222 89978
rect 14390 89784 14498 89978
rect 14666 89784 14774 89978
rect 14942 89784 15050 89978
rect 15218 89784 15326 89978
rect 15494 89784 15602 89978
rect 15770 89784 15878 89978
rect 16046 89784 16154 89978
rect 16322 89784 16430 89978
rect 16598 89784 16706 89978
rect 16874 89784 16982 89978
rect 17150 89784 17258 89978
rect 17426 89784 17534 89978
rect 17702 89784 17810 89978
rect 17978 89784 18086 89978
rect 18254 89784 18362 89978
rect 18530 89784 18638 89978
rect 18806 89784 18914 89978
rect 19082 89784 19190 89978
rect 19358 89784 19466 89978
rect 19634 89784 19742 89978
rect 19910 89784 20018 89978
rect 20186 89784 20294 89978
rect 20462 89784 20570 89978
rect 20738 89784 20846 89978
rect 21014 89784 21122 89978
rect 21290 89784 21398 89978
rect 21566 89784 21674 89978
rect 21842 89784 21950 89978
rect 22118 89784 22226 89978
rect 22394 89784 22502 89978
rect 22670 89784 22778 89978
rect 22946 89784 23054 89978
rect 23222 89784 23330 89978
rect 23498 89784 23606 89978
rect 23774 89784 23882 89978
rect 24050 89784 24158 89978
rect 24326 89784 24434 89978
rect 24602 89784 24710 89978
rect 24878 89784 24986 89978
rect 25154 89784 25262 89978
rect 25430 89784 25538 89978
rect 25706 89784 25814 89978
rect 25982 89784 26090 89978
rect 26258 89784 26366 89978
rect 26534 89784 26642 89978
rect 26810 89784 26918 89978
rect 27086 89784 27194 89978
rect 27362 89784 27470 89978
rect 27638 89784 27746 89978
rect 27914 89784 28022 89978
rect 28190 89784 28298 89978
rect 28466 89784 28574 89978
rect 28742 89784 28850 89978
rect 29018 89784 29126 89978
rect 29294 89784 29402 89978
rect 29570 89784 29678 89978
rect 29846 89784 29954 89978
rect 30122 89784 30230 89978
rect 30398 89784 30506 89978
rect 30674 89784 30782 89978
rect 30950 89784 31058 89978
rect 31226 89784 31334 89978
rect 31502 89784 31610 89978
rect 31778 89784 31886 89978
rect 32054 89784 32162 89978
rect 32330 89784 32438 89978
rect 32606 89784 32714 89978
rect 32882 89784 32990 89978
rect 33158 89784 33266 89978
rect 33434 89784 33542 89978
rect 33710 89784 33818 89978
rect 33986 89784 34094 89978
rect 34262 89784 34370 89978
rect 34538 89784 34646 89978
rect 34814 89784 34922 89978
rect 35090 89784 35198 89978
rect 35366 89784 35474 89978
rect 35642 89784 35750 89978
rect 35918 89784 36026 89978
rect 36194 89784 36302 89978
rect 36470 89784 36578 89978
rect 36746 89784 36854 89978
rect 37022 89784 37130 89978
rect 37298 89784 37406 89978
rect 37574 89784 37682 89978
rect 37850 89784 37958 89978
rect 38126 89784 38234 89978
rect 38402 89784 38510 89978
rect 38678 89784 38786 89978
rect 38954 89784 39062 89978
rect 39230 89784 39338 89978
rect 39506 89784 44692 89978
rect 20 216 44692 89784
rect 20 54 5114 216
rect 5282 54 5390 216
rect 5558 54 5666 216
rect 5834 54 5942 216
rect 6110 54 6218 216
rect 6386 54 6494 216
rect 6662 54 6770 216
rect 6938 54 7046 216
rect 7214 54 7322 216
rect 7490 54 7598 216
rect 7766 54 7874 216
rect 8042 54 8150 216
rect 8318 54 8426 216
rect 8594 54 8702 216
rect 8870 54 8978 216
rect 9146 54 9254 216
rect 9422 54 9530 216
rect 9698 54 9806 216
rect 9974 54 10082 216
rect 10250 54 10358 216
rect 10526 54 10634 216
rect 10802 54 10910 216
rect 11078 54 11186 216
rect 11354 54 11462 216
rect 11630 54 11738 216
rect 11906 54 12014 216
rect 12182 54 12290 216
rect 12458 54 12566 216
rect 12734 54 12842 216
rect 13010 54 13118 216
rect 13286 54 13394 216
rect 13562 54 13670 216
rect 13838 54 13946 216
rect 14114 54 14222 216
rect 14390 54 14498 216
rect 14666 54 14774 216
rect 14942 54 15050 216
rect 15218 54 15326 216
rect 15494 54 15602 216
rect 15770 54 15878 216
rect 16046 54 16154 216
rect 16322 54 16430 216
rect 16598 54 16706 216
rect 16874 54 16982 216
rect 17150 54 17258 216
rect 17426 54 17534 216
rect 17702 54 17810 216
rect 17978 54 18086 216
rect 18254 54 18362 216
rect 18530 54 18638 216
rect 18806 54 18914 216
rect 19082 54 19190 216
rect 19358 54 19466 216
rect 19634 54 19742 216
rect 19910 54 20018 216
rect 20186 54 20294 216
rect 20462 54 20570 216
rect 20738 54 20846 216
rect 21014 54 21122 216
rect 21290 54 21398 216
rect 21566 54 21674 216
rect 21842 54 21950 216
rect 22118 54 22226 216
rect 22394 54 22502 216
rect 22670 54 22778 216
rect 22946 54 23054 216
rect 23222 54 23330 216
rect 23498 54 23606 216
rect 23774 54 23882 216
rect 24050 54 24158 216
rect 24326 54 24434 216
rect 24602 54 24710 216
rect 24878 54 24986 216
rect 25154 54 25262 216
rect 25430 54 25538 216
rect 25706 54 25814 216
rect 25982 54 26090 216
rect 26258 54 26366 216
rect 26534 54 26642 216
rect 26810 54 26918 216
rect 27086 54 27194 216
rect 27362 54 27470 216
rect 27638 54 27746 216
rect 27914 54 28022 216
rect 28190 54 28298 216
rect 28466 54 28574 216
rect 28742 54 28850 216
rect 29018 54 29126 216
rect 29294 54 29402 216
rect 29570 54 29678 216
rect 29846 54 29954 216
rect 30122 54 30230 216
rect 30398 54 30506 216
rect 30674 54 30782 216
rect 30950 54 31058 216
rect 31226 54 31334 216
rect 31502 54 31610 216
rect 31778 54 31886 216
rect 32054 54 32162 216
rect 32330 54 32438 216
rect 32606 54 32714 216
rect 32882 54 32990 216
rect 33158 54 33266 216
rect 33434 54 33542 216
rect 33710 54 33818 216
rect 33986 54 34094 216
rect 34262 54 34370 216
rect 34538 54 34646 216
rect 34814 54 34922 216
rect 35090 54 35198 216
rect 35366 54 35474 216
rect 35642 54 35750 216
rect 35918 54 36026 216
rect 36194 54 36302 216
rect 36470 54 36578 216
rect 36746 54 36854 216
rect 37022 54 37130 216
rect 37298 54 37406 216
rect 37574 54 37682 216
rect 37850 54 37958 216
rect 38126 54 38234 216
rect 38402 54 38510 216
rect 38678 54 38786 216
rect 38954 54 39062 216
rect 39230 54 39338 216
rect 39506 54 44692 216
<< metal3 >>
rect -40 85416 160 85536
rect -40 85144 160 85264
rect -40 84872 160 84992
rect -40 84600 160 84720
rect -40 84328 160 84448
rect -40 84056 160 84176
rect -40 83784 160 83904
rect -40 83512 160 83632
rect -40 83240 160 83360
rect -40 82968 160 83088
rect -40 82696 160 82816
rect -40 82424 160 82544
rect -40 82152 160 82272
rect -40 81880 160 82000
rect -40 81608 160 81728
rect -40 81336 160 81456
rect -40 81064 160 81184
rect -40 80792 160 80912
rect -40 80520 160 80640
rect -40 80248 160 80368
rect -40 79976 160 80096
rect -40 79704 160 79824
rect -40 79432 160 79552
rect -40 79160 160 79280
rect -40 78888 160 79008
rect -40 78616 160 78736
rect -40 78344 160 78464
rect -40 78072 160 78192
rect -40 77800 160 77920
rect -40 77528 160 77648
rect -40 77256 160 77376
rect -40 76984 160 77104
rect -40 76712 160 76832
rect -40 76440 160 76560
rect -40 76168 160 76288
rect -40 75896 160 76016
rect -40 75624 160 75744
rect -40 75352 160 75472
rect -40 75080 160 75200
rect -40 74808 160 74928
rect -40 74536 160 74656
rect -40 74264 160 74384
rect -40 73992 160 74112
rect -40 73720 160 73840
rect -40 73448 160 73568
rect -40 73176 160 73296
rect -40 72904 160 73024
rect -40 72632 160 72752
rect -40 72360 160 72480
rect -40 72088 160 72208
rect -40 71816 160 71936
rect -40 71544 160 71664
rect -40 71272 160 71392
rect -40 71000 160 71120
rect -40 70728 160 70848
rect -40 70456 160 70576
rect -40 70184 160 70304
rect -40 69912 160 70032
rect -40 69640 160 69760
rect -40 69368 160 69488
rect -40 69096 160 69216
rect -40 68824 160 68944
rect -40 68552 160 68672
rect -40 68280 160 68400
rect -40 68008 160 68128
rect -40 67736 160 67856
rect -40 67464 160 67584
rect -40 67192 160 67312
rect -40 66920 160 67040
rect -40 66648 160 66768
rect -40 66376 160 66496
rect -40 66104 160 66224
rect -40 65832 160 65952
rect -40 65560 160 65680
rect -40 65288 160 65408
rect -40 65016 160 65136
rect -40 64744 160 64864
rect -40 64472 160 64592
rect -40 64200 160 64320
rect -40 63928 160 64048
rect -40 63656 160 63776
rect -40 63384 160 63504
rect -40 63112 160 63232
rect -40 62840 160 62960
rect -40 62568 160 62688
rect -40 62296 160 62416
rect -40 62024 160 62144
rect -40 61752 160 61872
rect -40 61480 160 61600
rect -40 61208 160 61328
rect -40 60936 160 61056
rect -40 60664 160 60784
rect -40 60392 160 60512
rect -40 60120 160 60240
rect -40 59848 160 59968
rect -40 59576 160 59696
rect -40 59304 160 59424
rect -40 59032 160 59152
rect -40 58760 160 58880
rect -40 58488 160 58608
rect -40 58216 160 58336
rect -40 57944 160 58064
rect -40 57672 160 57792
rect -40 57400 160 57520
rect -40 57128 160 57248
rect -40 56856 160 56976
rect -40 56584 160 56704
rect -40 56312 160 56432
rect -40 56040 160 56160
rect -40 55768 160 55888
rect -40 55496 160 55616
rect -40 55224 160 55344
rect -40 54952 160 55072
rect -40 54680 160 54800
rect -40 54408 160 54528
rect -40 54136 160 54256
rect -40 53864 160 53984
rect -40 53592 160 53712
rect -40 53320 160 53440
rect -40 53048 160 53168
rect -40 52776 160 52896
rect -40 52504 160 52624
rect -40 52232 160 52352
rect -40 51960 160 52080
rect -40 51688 160 51808
rect -40 51416 160 51536
rect -40 51144 160 51264
rect -40 50872 160 50992
rect 44540 85416 44740 85536
rect 44540 85144 44740 85264
rect 44540 84872 44740 84992
rect 44540 84600 44740 84720
rect 44540 84328 44740 84448
rect 44540 84056 44740 84176
rect 44540 83784 44740 83904
rect 44540 83512 44740 83632
rect 44540 83240 44740 83360
rect 44540 82968 44740 83088
rect 44540 82696 44740 82816
rect 44540 82424 44740 82544
rect 44540 82152 44740 82272
rect 44540 81880 44740 82000
rect 44540 81608 44740 81728
rect 44540 81336 44740 81456
rect 44540 81064 44740 81184
rect 44540 80792 44740 80912
rect 44540 80520 44740 80640
rect 44540 80248 44740 80368
rect 44540 79976 44740 80096
rect 44540 79704 44740 79824
rect 44540 79432 44740 79552
rect 44540 79160 44740 79280
rect 44540 78888 44740 79008
rect 44540 78616 44740 78736
rect 44540 78344 44740 78464
rect 44540 78072 44740 78192
rect 44540 77800 44740 77920
rect 44540 77528 44740 77648
rect 44540 77256 44740 77376
rect 44540 76984 44740 77104
rect 44540 76712 44740 76832
rect 44540 76440 44740 76560
rect 44540 76168 44740 76288
rect 44540 75896 44740 76016
rect 44540 75624 44740 75744
rect 44540 75352 44740 75472
rect 44540 75080 44740 75200
rect 44540 74808 44740 74928
rect 44540 74536 44740 74656
rect 44540 74264 44740 74384
rect 44540 73992 44740 74112
rect 44540 73720 44740 73840
rect 44540 73448 44740 73568
rect 44540 73176 44740 73296
rect 44540 72904 44740 73024
rect 44540 72632 44740 72752
rect 44540 72360 44740 72480
rect 44540 72088 44740 72208
rect 44540 71816 44740 71936
rect 44540 71544 44740 71664
rect 44540 71272 44740 71392
rect 44540 71000 44740 71120
rect 44540 70728 44740 70848
rect 44540 70456 44740 70576
rect 44540 70184 44740 70304
rect 44540 69912 44740 70032
rect 44540 69640 44740 69760
rect 44540 69368 44740 69488
rect 44540 69096 44740 69216
rect 44540 68824 44740 68944
rect 44540 68552 44740 68672
rect 44540 68280 44740 68400
rect 44540 68008 44740 68128
rect 44540 67736 44740 67856
rect 44540 67464 44740 67584
rect 44540 67192 44740 67312
rect 44540 66920 44740 67040
rect 44540 66648 44740 66768
rect 44540 66376 44740 66496
rect 44540 66104 44740 66224
rect 44540 65832 44740 65952
rect 44540 65560 44740 65680
rect 44540 65288 44740 65408
rect 44540 65016 44740 65136
rect 44540 64744 44740 64864
rect 44540 64472 44740 64592
rect 44540 64200 44740 64320
rect 44540 63928 44740 64048
rect 44540 63656 44740 63776
rect 44540 63384 44740 63504
rect 44540 63112 44740 63232
rect 44540 62840 44740 62960
rect 44540 62568 44740 62688
rect 44540 62296 44740 62416
rect 44540 62024 44740 62144
rect 44540 61752 44740 61872
rect 44540 61480 44740 61600
rect 44540 61208 44740 61328
rect 44540 60936 44740 61056
rect 44540 60664 44740 60784
rect 44540 60392 44740 60512
rect 44540 60120 44740 60240
rect 44540 59848 44740 59968
rect 44540 59576 44740 59696
rect 44540 59304 44740 59424
rect 44540 59032 44740 59152
rect 44540 58760 44740 58880
rect 44540 58488 44740 58608
rect 44540 58216 44740 58336
rect 44540 57944 44740 58064
rect 44540 57672 44740 57792
rect 44540 57400 44740 57520
rect 44540 57128 44740 57248
rect 44540 56856 44740 56976
rect 44540 56584 44740 56704
rect 44540 56312 44740 56432
rect 44540 56040 44740 56160
rect 44540 55768 44740 55888
rect 44540 55496 44740 55616
rect 44540 55224 44740 55344
rect 44540 54952 44740 55072
rect 44540 54680 44740 54800
rect 44540 54408 44740 54528
rect 44540 54136 44740 54256
rect 44540 53864 44740 53984
rect 44540 53592 44740 53712
rect 44540 53320 44740 53440
rect 44540 53048 44740 53168
rect 44540 52776 44740 52896
rect 44540 52504 44740 52624
rect 44540 52232 44740 52352
rect 44540 51960 44740 52080
rect 44540 51688 44740 51808
rect 44540 51416 44740 51536
rect 44540 51144 44740 51264
rect 44540 50872 44740 50992
rect -40 39448 160 39568
rect -40 39176 160 39296
rect -40 38904 160 39024
rect -40 38632 160 38752
rect -40 38360 160 38480
rect -40 38088 160 38208
rect -40 37816 160 37936
rect -40 37544 160 37664
rect -40 37272 160 37392
rect -40 37000 160 37120
rect -40 36728 160 36848
rect -40 36456 160 36576
rect -40 36184 160 36304
rect -40 35912 160 36032
rect -40 35640 160 35760
rect -40 35368 160 35488
rect -40 35096 160 35216
rect -40 34824 160 34944
rect -40 34552 160 34672
rect -40 34280 160 34400
rect -40 34008 160 34128
rect -40 33736 160 33856
rect -40 33464 160 33584
rect -40 33192 160 33312
rect -40 32920 160 33040
rect -40 32648 160 32768
rect -40 32376 160 32496
rect -40 32104 160 32224
rect -40 31832 160 31952
rect -40 31560 160 31680
rect -40 31288 160 31408
rect -40 31016 160 31136
rect -40 30744 160 30864
rect -40 30472 160 30592
rect -40 30200 160 30320
rect -40 29928 160 30048
rect -40 29656 160 29776
rect -40 29384 160 29504
rect -40 29112 160 29232
rect -40 28840 160 28960
rect -40 28568 160 28688
rect -40 28296 160 28416
rect -40 28024 160 28144
rect -40 27752 160 27872
rect -40 27480 160 27600
rect -40 27208 160 27328
rect -40 26936 160 27056
rect -40 26664 160 26784
rect -40 26392 160 26512
rect -40 26120 160 26240
rect -40 25848 160 25968
rect -40 25576 160 25696
rect -40 25304 160 25424
rect -40 25032 160 25152
rect -40 24760 160 24880
rect -40 24488 160 24608
rect -40 24216 160 24336
rect -40 23944 160 24064
rect -40 23672 160 23792
rect -40 23400 160 23520
rect -40 23128 160 23248
rect -40 22856 160 22976
rect -40 22584 160 22704
rect -40 22312 160 22432
rect -40 22040 160 22160
rect -40 21768 160 21888
rect -40 21496 160 21616
rect -40 21224 160 21344
rect -40 20952 160 21072
rect -40 20680 160 20800
rect -40 20408 160 20528
rect -40 20136 160 20256
rect -40 19864 160 19984
rect -40 19592 160 19712
rect -40 19320 160 19440
rect -40 19048 160 19168
rect -40 18776 160 18896
rect -40 18504 160 18624
rect -40 18232 160 18352
rect -40 17960 160 18080
rect -40 17688 160 17808
rect -40 17416 160 17536
rect -40 17144 160 17264
rect -40 16872 160 16992
rect -40 16600 160 16720
rect -40 16328 160 16448
rect -40 16056 160 16176
rect -40 15784 160 15904
rect -40 15512 160 15632
rect -40 15240 160 15360
rect -40 14968 160 15088
rect -40 14696 160 14816
rect -40 14424 160 14544
rect -40 14152 160 14272
rect -40 13880 160 14000
rect -40 13608 160 13728
rect -40 13336 160 13456
rect -40 13064 160 13184
rect -40 12792 160 12912
rect -40 12520 160 12640
rect -40 12248 160 12368
rect -40 11976 160 12096
rect -40 11704 160 11824
rect -40 11432 160 11552
rect -40 11160 160 11280
rect -40 10888 160 11008
rect -40 10616 160 10736
rect -40 10344 160 10464
rect -40 10072 160 10192
rect -40 9800 160 9920
rect -40 9528 160 9648
rect -40 9256 160 9376
rect -40 8984 160 9104
rect -40 8712 160 8832
rect -40 8440 160 8560
rect -40 8168 160 8288
rect -40 7896 160 8016
rect -40 7624 160 7744
rect -40 7352 160 7472
rect -40 7080 160 7200
rect -40 6808 160 6928
rect -40 6536 160 6656
rect -40 6264 160 6384
rect -40 5992 160 6112
rect -40 5720 160 5840
rect -40 5448 160 5568
rect -40 5176 160 5296
rect -40 4904 160 5024
rect 44540 39448 44740 39568
rect 44540 39176 44740 39296
rect 44540 38904 44740 39024
rect 44540 38632 44740 38752
rect 44540 38360 44740 38480
rect 44540 38088 44740 38208
rect 44540 37816 44740 37936
rect 44540 37544 44740 37664
rect 44540 37272 44740 37392
rect 44540 37000 44740 37120
rect 44540 36728 44740 36848
rect 44540 36456 44740 36576
rect 44540 36184 44740 36304
rect 44540 35912 44740 36032
rect 44540 35640 44740 35760
rect 44540 35368 44740 35488
rect 44540 35096 44740 35216
rect 44540 34824 44740 34944
rect 44540 34552 44740 34672
rect 44540 34280 44740 34400
rect 44540 34008 44740 34128
rect 44540 33736 44740 33856
rect 44540 33464 44740 33584
rect 44540 33192 44740 33312
rect 44540 32920 44740 33040
rect 44540 32648 44740 32768
rect 44540 32376 44740 32496
rect 44540 32104 44740 32224
rect 44540 31832 44740 31952
rect 44540 31560 44740 31680
rect 44540 31288 44740 31408
rect 44540 31016 44740 31136
rect 44540 30744 44740 30864
rect 44540 30472 44740 30592
rect 44540 30200 44740 30320
rect 44540 29928 44740 30048
rect 44540 29656 44740 29776
rect 44540 29384 44740 29504
rect 44540 29112 44740 29232
rect 44540 28840 44740 28960
rect 44540 28568 44740 28688
rect 44540 28296 44740 28416
rect 44540 28024 44740 28144
rect 44540 27752 44740 27872
rect 44540 27480 44740 27600
rect 44540 27208 44740 27328
rect 44540 26936 44740 27056
rect 44540 26664 44740 26784
rect 44540 26392 44740 26512
rect 44540 26120 44740 26240
rect 44540 25848 44740 25968
rect 44540 25576 44740 25696
rect 44540 25304 44740 25424
rect 44540 25032 44740 25152
rect 44540 24760 44740 24880
rect 44540 24488 44740 24608
rect 44540 24216 44740 24336
rect 44540 23944 44740 24064
rect 44540 23672 44740 23792
rect 44540 23400 44740 23520
rect 44540 23128 44740 23248
rect 44540 22856 44740 22976
rect 44540 22584 44740 22704
rect 44540 22312 44740 22432
rect 44540 22040 44740 22160
rect 44540 21768 44740 21888
rect 44540 21496 44740 21616
rect 44540 21224 44740 21344
rect 44540 20952 44740 21072
rect 44540 20680 44740 20800
rect 44540 20408 44740 20528
rect 44540 20136 44740 20256
rect 44540 19864 44740 19984
rect 44540 19592 44740 19712
rect 44540 19320 44740 19440
rect 44540 19048 44740 19168
rect 44540 18776 44740 18896
rect 44540 18504 44740 18624
rect 44540 18232 44740 18352
rect 44540 17960 44740 18080
rect 44540 17688 44740 17808
rect 44540 17416 44740 17536
rect 44540 17144 44740 17264
rect 44540 16872 44740 16992
rect 44540 16600 44740 16720
rect 44540 16328 44740 16448
rect 44540 16056 44740 16176
rect 44540 15784 44740 15904
rect 44540 15512 44740 15632
rect 44540 15240 44740 15360
rect 44540 14968 44740 15088
rect 44540 14696 44740 14816
rect 44540 14424 44740 14544
rect 44540 14152 44740 14272
rect 44540 13880 44740 14000
rect 44540 13608 44740 13728
rect 44540 13336 44740 13456
rect 44540 13064 44740 13184
rect 44540 12792 44740 12912
rect 44540 12520 44740 12640
rect 44540 12248 44740 12368
rect 44540 11976 44740 12096
rect 44540 11704 44740 11824
rect 44540 11432 44740 11552
rect 44540 11160 44740 11280
rect 44540 10888 44740 11008
rect 44540 10616 44740 10736
rect 44540 10344 44740 10464
rect 44540 10072 44740 10192
rect 44540 9800 44740 9920
rect 44540 9528 44740 9648
rect 44540 9256 44740 9376
rect 44540 8984 44740 9104
rect 44540 8712 44740 8832
rect 44540 8440 44740 8560
rect 44540 8168 44740 8288
rect 44540 7896 44740 8016
rect 44540 7624 44740 7744
rect 44540 7352 44740 7472
rect 44540 7080 44740 7200
rect 44540 6808 44740 6928
rect 44540 6536 44740 6656
rect 44540 6264 44740 6384
rect 44540 5992 44740 6112
rect 44540 5720 44740 5840
rect 44540 5448 44740 5568
rect 44540 5176 44740 5296
rect 44540 4904 44740 5024
<< obsm3 >>
rect 105 85616 44540 88909
rect 240 50792 44460 85616
rect 105 39648 44540 50792
rect 240 4824 44460 39648
rect 105 851 44540 4824
<< metal4 >>
rect 4208 1040 4528 88720
rect 19568 1040 19888 88720
rect 34928 1040 35248 88720
<< obsm4 >>
rect 611 88800 44285 88909
rect 611 960 4128 88800
rect 4608 960 19488 88800
rect 19968 960 34848 88800
rect 35328 960 44285 88800
rect 611 851 44285 960
<< labels >>
rlabel metal3 s 44540 63928 44740 64048 6 Tile_X0Y0_E1BEG[0]
port 1 nsew signal output
rlabel metal3 s 44540 64200 44740 64320 6 Tile_X0Y0_E1BEG[1]
port 2 nsew signal output
rlabel metal3 s 44540 64472 44740 64592 6 Tile_X0Y0_E1BEG[2]
port 3 nsew signal output
rlabel metal3 s 44540 64744 44740 64864 6 Tile_X0Y0_E1BEG[3]
port 4 nsew signal output
rlabel metal3 s -40 63928 160 64048 6 Tile_X0Y0_E1END[0]
port 5 nsew signal input
rlabel metal3 s -40 64200 160 64320 6 Tile_X0Y0_E1END[1]
port 6 nsew signal input
rlabel metal3 s -40 64472 160 64592 6 Tile_X0Y0_E1END[2]
port 7 nsew signal input
rlabel metal3 s -40 64744 160 64864 6 Tile_X0Y0_E1END[3]
port 8 nsew signal input
rlabel metal3 s 44540 65016 44740 65136 6 Tile_X0Y0_E2BEG[0]
port 9 nsew signal output
rlabel metal3 s 44540 65288 44740 65408 6 Tile_X0Y0_E2BEG[1]
port 10 nsew signal output
rlabel metal3 s 44540 65560 44740 65680 6 Tile_X0Y0_E2BEG[2]
port 11 nsew signal output
rlabel metal3 s 44540 65832 44740 65952 6 Tile_X0Y0_E2BEG[3]
port 12 nsew signal output
rlabel metal3 s 44540 66104 44740 66224 6 Tile_X0Y0_E2BEG[4]
port 13 nsew signal output
rlabel metal3 s 44540 66376 44740 66496 6 Tile_X0Y0_E2BEG[5]
port 14 nsew signal output
rlabel metal3 s 44540 66648 44740 66768 6 Tile_X0Y0_E2BEG[6]
port 15 nsew signal output
rlabel metal3 s 44540 66920 44740 67040 6 Tile_X0Y0_E2BEG[7]
port 16 nsew signal output
rlabel metal3 s 44540 67192 44740 67312 6 Tile_X0Y0_E2BEGb[0]
port 17 nsew signal output
rlabel metal3 s 44540 67464 44740 67584 6 Tile_X0Y0_E2BEGb[1]
port 18 nsew signal output
rlabel metal3 s 44540 67736 44740 67856 6 Tile_X0Y0_E2BEGb[2]
port 19 nsew signal output
rlabel metal3 s 44540 68008 44740 68128 6 Tile_X0Y0_E2BEGb[3]
port 20 nsew signal output
rlabel metal3 s 44540 68280 44740 68400 6 Tile_X0Y0_E2BEGb[4]
port 21 nsew signal output
rlabel metal3 s 44540 68552 44740 68672 6 Tile_X0Y0_E2BEGb[5]
port 22 nsew signal output
rlabel metal3 s 44540 68824 44740 68944 6 Tile_X0Y0_E2BEGb[6]
port 23 nsew signal output
rlabel metal3 s 44540 69096 44740 69216 6 Tile_X0Y0_E2BEGb[7]
port 24 nsew signal output
rlabel metal3 s -40 67192 160 67312 6 Tile_X0Y0_E2END[0]
port 25 nsew signal input
rlabel metal3 s -40 67464 160 67584 6 Tile_X0Y0_E2END[1]
port 26 nsew signal input
rlabel metal3 s -40 67736 160 67856 6 Tile_X0Y0_E2END[2]
port 27 nsew signal input
rlabel metal3 s -40 68008 160 68128 6 Tile_X0Y0_E2END[3]
port 28 nsew signal input
rlabel metal3 s -40 68280 160 68400 6 Tile_X0Y0_E2END[4]
port 29 nsew signal input
rlabel metal3 s -40 68552 160 68672 6 Tile_X0Y0_E2END[5]
port 30 nsew signal input
rlabel metal3 s -40 68824 160 68944 6 Tile_X0Y0_E2END[6]
port 31 nsew signal input
rlabel metal3 s -40 69096 160 69216 6 Tile_X0Y0_E2END[7]
port 32 nsew signal input
rlabel metal3 s -40 65016 160 65136 6 Tile_X0Y0_E2MID[0]
port 33 nsew signal input
rlabel metal3 s -40 65288 160 65408 6 Tile_X0Y0_E2MID[1]
port 34 nsew signal input
rlabel metal3 s -40 65560 160 65680 6 Tile_X0Y0_E2MID[2]
port 35 nsew signal input
rlabel metal3 s -40 65832 160 65952 6 Tile_X0Y0_E2MID[3]
port 36 nsew signal input
rlabel metal3 s -40 66104 160 66224 6 Tile_X0Y0_E2MID[4]
port 37 nsew signal input
rlabel metal3 s -40 66376 160 66496 6 Tile_X0Y0_E2MID[5]
port 38 nsew signal input
rlabel metal3 s -40 66648 160 66768 6 Tile_X0Y0_E2MID[6]
port 39 nsew signal input
rlabel metal3 s -40 66920 160 67040 6 Tile_X0Y0_E2MID[7]
port 40 nsew signal input
rlabel metal3 s 44540 73720 44740 73840 6 Tile_X0Y0_E6BEG[0]
port 41 nsew signal output
rlabel metal3 s 44540 76440 44740 76560 6 Tile_X0Y0_E6BEG[10]
port 42 nsew signal output
rlabel metal3 s 44540 76712 44740 76832 6 Tile_X0Y0_E6BEG[11]
port 43 nsew signal output
rlabel metal3 s 44540 73992 44740 74112 6 Tile_X0Y0_E6BEG[1]
port 44 nsew signal output
rlabel metal3 s 44540 74264 44740 74384 6 Tile_X0Y0_E6BEG[2]
port 45 nsew signal output
rlabel metal3 s 44540 74536 44740 74656 6 Tile_X0Y0_E6BEG[3]
port 46 nsew signal output
rlabel metal3 s 44540 74808 44740 74928 6 Tile_X0Y0_E6BEG[4]
port 47 nsew signal output
rlabel metal3 s 44540 75080 44740 75200 6 Tile_X0Y0_E6BEG[5]
port 48 nsew signal output
rlabel metal3 s 44540 75352 44740 75472 6 Tile_X0Y0_E6BEG[6]
port 49 nsew signal output
rlabel metal3 s 44540 75624 44740 75744 6 Tile_X0Y0_E6BEG[7]
port 50 nsew signal output
rlabel metal3 s 44540 75896 44740 76016 6 Tile_X0Y0_E6BEG[8]
port 51 nsew signal output
rlabel metal3 s 44540 76168 44740 76288 6 Tile_X0Y0_E6BEG[9]
port 52 nsew signal output
rlabel metal3 s -40 73720 160 73840 6 Tile_X0Y0_E6END[0]
port 53 nsew signal input
rlabel metal3 s -40 76440 160 76560 6 Tile_X0Y0_E6END[10]
port 54 nsew signal input
rlabel metal3 s -40 76712 160 76832 6 Tile_X0Y0_E6END[11]
port 55 nsew signal input
rlabel metal3 s -40 73992 160 74112 6 Tile_X0Y0_E6END[1]
port 56 nsew signal input
rlabel metal3 s -40 74264 160 74384 6 Tile_X0Y0_E6END[2]
port 57 nsew signal input
rlabel metal3 s -40 74536 160 74656 6 Tile_X0Y0_E6END[3]
port 58 nsew signal input
rlabel metal3 s -40 74808 160 74928 6 Tile_X0Y0_E6END[4]
port 59 nsew signal input
rlabel metal3 s -40 75080 160 75200 6 Tile_X0Y0_E6END[5]
port 60 nsew signal input
rlabel metal3 s -40 75352 160 75472 6 Tile_X0Y0_E6END[6]
port 61 nsew signal input
rlabel metal3 s -40 75624 160 75744 6 Tile_X0Y0_E6END[7]
port 62 nsew signal input
rlabel metal3 s -40 75896 160 76016 6 Tile_X0Y0_E6END[8]
port 63 nsew signal input
rlabel metal3 s -40 76168 160 76288 6 Tile_X0Y0_E6END[9]
port 64 nsew signal input
rlabel metal3 s 44540 69368 44740 69488 6 Tile_X0Y0_EE4BEG[0]
port 65 nsew signal output
rlabel metal3 s 44540 72088 44740 72208 6 Tile_X0Y0_EE4BEG[10]
port 66 nsew signal output
rlabel metal3 s 44540 72360 44740 72480 6 Tile_X0Y0_EE4BEG[11]
port 67 nsew signal output
rlabel metal3 s 44540 72632 44740 72752 6 Tile_X0Y0_EE4BEG[12]
port 68 nsew signal output
rlabel metal3 s 44540 72904 44740 73024 6 Tile_X0Y0_EE4BEG[13]
port 69 nsew signal output
rlabel metal3 s 44540 73176 44740 73296 6 Tile_X0Y0_EE4BEG[14]
port 70 nsew signal output
rlabel metal3 s 44540 73448 44740 73568 6 Tile_X0Y0_EE4BEG[15]
port 71 nsew signal output
rlabel metal3 s 44540 69640 44740 69760 6 Tile_X0Y0_EE4BEG[1]
port 72 nsew signal output
rlabel metal3 s 44540 69912 44740 70032 6 Tile_X0Y0_EE4BEG[2]
port 73 nsew signal output
rlabel metal3 s 44540 70184 44740 70304 6 Tile_X0Y0_EE4BEG[3]
port 74 nsew signal output
rlabel metal3 s 44540 70456 44740 70576 6 Tile_X0Y0_EE4BEG[4]
port 75 nsew signal output
rlabel metal3 s 44540 70728 44740 70848 6 Tile_X0Y0_EE4BEG[5]
port 76 nsew signal output
rlabel metal3 s 44540 71000 44740 71120 6 Tile_X0Y0_EE4BEG[6]
port 77 nsew signal output
rlabel metal3 s 44540 71272 44740 71392 6 Tile_X0Y0_EE4BEG[7]
port 78 nsew signal output
rlabel metal3 s 44540 71544 44740 71664 6 Tile_X0Y0_EE4BEG[8]
port 79 nsew signal output
rlabel metal3 s 44540 71816 44740 71936 6 Tile_X0Y0_EE4BEG[9]
port 80 nsew signal output
rlabel metal3 s -40 69368 160 69488 6 Tile_X0Y0_EE4END[0]
port 81 nsew signal input
rlabel metal3 s -40 72088 160 72208 6 Tile_X0Y0_EE4END[10]
port 82 nsew signal input
rlabel metal3 s -40 72360 160 72480 6 Tile_X0Y0_EE4END[11]
port 83 nsew signal input
rlabel metal3 s -40 72632 160 72752 6 Tile_X0Y0_EE4END[12]
port 84 nsew signal input
rlabel metal3 s -40 72904 160 73024 6 Tile_X0Y0_EE4END[13]
port 85 nsew signal input
rlabel metal3 s -40 73176 160 73296 6 Tile_X0Y0_EE4END[14]
port 86 nsew signal input
rlabel metal3 s -40 73448 160 73568 6 Tile_X0Y0_EE4END[15]
port 87 nsew signal input
rlabel metal3 s -40 69640 160 69760 6 Tile_X0Y0_EE4END[1]
port 88 nsew signal input
rlabel metal3 s -40 69912 160 70032 6 Tile_X0Y0_EE4END[2]
port 89 nsew signal input
rlabel metal3 s -40 70184 160 70304 6 Tile_X0Y0_EE4END[3]
port 90 nsew signal input
rlabel metal3 s -40 70456 160 70576 6 Tile_X0Y0_EE4END[4]
port 91 nsew signal input
rlabel metal3 s -40 70728 160 70848 6 Tile_X0Y0_EE4END[5]
port 92 nsew signal input
rlabel metal3 s -40 71000 160 71120 6 Tile_X0Y0_EE4END[6]
port 93 nsew signal input
rlabel metal3 s -40 71272 160 71392 6 Tile_X0Y0_EE4END[7]
port 94 nsew signal input
rlabel metal3 s -40 71544 160 71664 6 Tile_X0Y0_EE4END[8]
port 95 nsew signal input
rlabel metal3 s -40 71816 160 71936 6 Tile_X0Y0_EE4END[9]
port 96 nsew signal input
rlabel metal3 s -40 76984 160 77104 6 Tile_X0Y0_FrameData[0]
port 97 nsew signal input
rlabel metal3 s -40 79704 160 79824 6 Tile_X0Y0_FrameData[10]
port 98 nsew signal input
rlabel metal3 s -40 79976 160 80096 6 Tile_X0Y0_FrameData[11]
port 99 nsew signal input
rlabel metal3 s -40 80248 160 80368 6 Tile_X0Y0_FrameData[12]
port 100 nsew signal input
rlabel metal3 s -40 80520 160 80640 6 Tile_X0Y0_FrameData[13]
port 101 nsew signal input
rlabel metal3 s -40 80792 160 80912 6 Tile_X0Y0_FrameData[14]
port 102 nsew signal input
rlabel metal3 s -40 81064 160 81184 6 Tile_X0Y0_FrameData[15]
port 103 nsew signal input
rlabel metal3 s -40 81336 160 81456 6 Tile_X0Y0_FrameData[16]
port 104 nsew signal input
rlabel metal3 s -40 81608 160 81728 6 Tile_X0Y0_FrameData[17]
port 105 nsew signal input
rlabel metal3 s -40 81880 160 82000 6 Tile_X0Y0_FrameData[18]
port 106 nsew signal input
rlabel metal3 s -40 82152 160 82272 6 Tile_X0Y0_FrameData[19]
port 107 nsew signal input
rlabel metal3 s -40 77256 160 77376 6 Tile_X0Y0_FrameData[1]
port 108 nsew signal input
rlabel metal3 s -40 82424 160 82544 6 Tile_X0Y0_FrameData[20]
port 109 nsew signal input
rlabel metal3 s -40 82696 160 82816 6 Tile_X0Y0_FrameData[21]
port 110 nsew signal input
rlabel metal3 s -40 82968 160 83088 6 Tile_X0Y0_FrameData[22]
port 111 nsew signal input
rlabel metal3 s -40 83240 160 83360 6 Tile_X0Y0_FrameData[23]
port 112 nsew signal input
rlabel metal3 s -40 83512 160 83632 6 Tile_X0Y0_FrameData[24]
port 113 nsew signal input
rlabel metal3 s -40 83784 160 83904 6 Tile_X0Y0_FrameData[25]
port 114 nsew signal input
rlabel metal3 s -40 84056 160 84176 6 Tile_X0Y0_FrameData[26]
port 115 nsew signal input
rlabel metal3 s -40 84328 160 84448 6 Tile_X0Y0_FrameData[27]
port 116 nsew signal input
rlabel metal3 s -40 84600 160 84720 6 Tile_X0Y0_FrameData[28]
port 117 nsew signal input
rlabel metal3 s -40 84872 160 84992 6 Tile_X0Y0_FrameData[29]
port 118 nsew signal input
rlabel metal3 s -40 77528 160 77648 6 Tile_X0Y0_FrameData[2]
port 119 nsew signal input
rlabel metal3 s -40 85144 160 85264 6 Tile_X0Y0_FrameData[30]
port 120 nsew signal input
rlabel metal3 s -40 85416 160 85536 6 Tile_X0Y0_FrameData[31]
port 121 nsew signal input
rlabel metal3 s -40 77800 160 77920 6 Tile_X0Y0_FrameData[3]
port 122 nsew signal input
rlabel metal3 s -40 78072 160 78192 6 Tile_X0Y0_FrameData[4]
port 123 nsew signal input
rlabel metal3 s -40 78344 160 78464 6 Tile_X0Y0_FrameData[5]
port 124 nsew signal input
rlabel metal3 s -40 78616 160 78736 6 Tile_X0Y0_FrameData[6]
port 125 nsew signal input
rlabel metal3 s -40 78888 160 79008 6 Tile_X0Y0_FrameData[7]
port 126 nsew signal input
rlabel metal3 s -40 79160 160 79280 6 Tile_X0Y0_FrameData[8]
port 127 nsew signal input
rlabel metal3 s -40 79432 160 79552 6 Tile_X0Y0_FrameData[9]
port 128 nsew signal input
rlabel metal3 s 44540 76984 44740 77104 6 Tile_X0Y0_FrameData_O[0]
port 129 nsew signal output
rlabel metal3 s 44540 79704 44740 79824 6 Tile_X0Y0_FrameData_O[10]
port 130 nsew signal output
rlabel metal3 s 44540 79976 44740 80096 6 Tile_X0Y0_FrameData_O[11]
port 131 nsew signal output
rlabel metal3 s 44540 80248 44740 80368 6 Tile_X0Y0_FrameData_O[12]
port 132 nsew signal output
rlabel metal3 s 44540 80520 44740 80640 6 Tile_X0Y0_FrameData_O[13]
port 133 nsew signal output
rlabel metal3 s 44540 80792 44740 80912 6 Tile_X0Y0_FrameData_O[14]
port 134 nsew signal output
rlabel metal3 s 44540 81064 44740 81184 6 Tile_X0Y0_FrameData_O[15]
port 135 nsew signal output
rlabel metal3 s 44540 81336 44740 81456 6 Tile_X0Y0_FrameData_O[16]
port 136 nsew signal output
rlabel metal3 s 44540 81608 44740 81728 6 Tile_X0Y0_FrameData_O[17]
port 137 nsew signal output
rlabel metal3 s 44540 81880 44740 82000 6 Tile_X0Y0_FrameData_O[18]
port 138 nsew signal output
rlabel metal3 s 44540 82152 44740 82272 6 Tile_X0Y0_FrameData_O[19]
port 139 nsew signal output
rlabel metal3 s 44540 77256 44740 77376 6 Tile_X0Y0_FrameData_O[1]
port 140 nsew signal output
rlabel metal3 s 44540 82424 44740 82544 6 Tile_X0Y0_FrameData_O[20]
port 141 nsew signal output
rlabel metal3 s 44540 82696 44740 82816 6 Tile_X0Y0_FrameData_O[21]
port 142 nsew signal output
rlabel metal3 s 44540 82968 44740 83088 6 Tile_X0Y0_FrameData_O[22]
port 143 nsew signal output
rlabel metal3 s 44540 83240 44740 83360 6 Tile_X0Y0_FrameData_O[23]
port 144 nsew signal output
rlabel metal3 s 44540 83512 44740 83632 6 Tile_X0Y0_FrameData_O[24]
port 145 nsew signal output
rlabel metal3 s 44540 83784 44740 83904 6 Tile_X0Y0_FrameData_O[25]
port 146 nsew signal output
rlabel metal3 s 44540 84056 44740 84176 6 Tile_X0Y0_FrameData_O[26]
port 147 nsew signal output
rlabel metal3 s 44540 84328 44740 84448 6 Tile_X0Y0_FrameData_O[27]
port 148 nsew signal output
rlabel metal3 s 44540 84600 44740 84720 6 Tile_X0Y0_FrameData_O[28]
port 149 nsew signal output
rlabel metal3 s 44540 84872 44740 84992 6 Tile_X0Y0_FrameData_O[29]
port 150 nsew signal output
rlabel metal3 s 44540 77528 44740 77648 6 Tile_X0Y0_FrameData_O[2]
port 151 nsew signal output
rlabel metal3 s 44540 85144 44740 85264 6 Tile_X0Y0_FrameData_O[30]
port 152 nsew signal output
rlabel metal3 s 44540 85416 44740 85536 6 Tile_X0Y0_FrameData_O[31]
port 153 nsew signal output
rlabel metal3 s 44540 77800 44740 77920 6 Tile_X0Y0_FrameData_O[3]
port 154 nsew signal output
rlabel metal3 s 44540 78072 44740 78192 6 Tile_X0Y0_FrameData_O[4]
port 155 nsew signal output
rlabel metal3 s 44540 78344 44740 78464 6 Tile_X0Y0_FrameData_O[5]
port 156 nsew signal output
rlabel metal3 s 44540 78616 44740 78736 6 Tile_X0Y0_FrameData_O[6]
port 157 nsew signal output
rlabel metal3 s 44540 78888 44740 79008 6 Tile_X0Y0_FrameData_O[7]
port 158 nsew signal output
rlabel metal3 s 44540 79160 44740 79280 6 Tile_X0Y0_FrameData_O[8]
port 159 nsew signal output
rlabel metal3 s 44540 79432 44740 79552 6 Tile_X0Y0_FrameData_O[9]
port 160 nsew signal output
rlabel metal2 s 34150 89840 34206 90040 6 Tile_X0Y0_FrameStrobe_O[0]
port 161 nsew signal output
rlabel metal2 s 36910 89840 36966 90040 6 Tile_X0Y0_FrameStrobe_O[10]
port 162 nsew signal output
rlabel metal2 s 37186 89840 37242 90040 6 Tile_X0Y0_FrameStrobe_O[11]
port 163 nsew signal output
rlabel metal2 s 37462 89840 37518 90040 6 Tile_X0Y0_FrameStrobe_O[12]
port 164 nsew signal output
rlabel metal2 s 37738 89840 37794 90040 6 Tile_X0Y0_FrameStrobe_O[13]
port 165 nsew signal output
rlabel metal2 s 38014 89840 38070 90040 6 Tile_X0Y0_FrameStrobe_O[14]
port 166 nsew signal output
rlabel metal2 s 38290 89840 38346 90040 6 Tile_X0Y0_FrameStrobe_O[15]
port 167 nsew signal output
rlabel metal2 s 38566 89840 38622 90040 6 Tile_X0Y0_FrameStrobe_O[16]
port 168 nsew signal output
rlabel metal2 s 38842 89840 38898 90040 6 Tile_X0Y0_FrameStrobe_O[17]
port 169 nsew signal output
rlabel metal2 s 39118 89840 39174 90040 6 Tile_X0Y0_FrameStrobe_O[18]
port 170 nsew signal output
rlabel metal2 s 39394 89840 39450 90040 6 Tile_X0Y0_FrameStrobe_O[19]
port 171 nsew signal output
rlabel metal2 s 34426 89840 34482 90040 6 Tile_X0Y0_FrameStrobe_O[1]
port 172 nsew signal output
rlabel metal2 s 34702 89840 34758 90040 6 Tile_X0Y0_FrameStrobe_O[2]
port 173 nsew signal output
rlabel metal2 s 34978 89840 35034 90040 6 Tile_X0Y0_FrameStrobe_O[3]
port 174 nsew signal output
rlabel metal2 s 35254 89840 35310 90040 6 Tile_X0Y0_FrameStrobe_O[4]
port 175 nsew signal output
rlabel metal2 s 35530 89840 35586 90040 6 Tile_X0Y0_FrameStrobe_O[5]
port 176 nsew signal output
rlabel metal2 s 35806 89840 35862 90040 6 Tile_X0Y0_FrameStrobe_O[6]
port 177 nsew signal output
rlabel metal2 s 36082 89840 36138 90040 6 Tile_X0Y0_FrameStrobe_O[7]
port 178 nsew signal output
rlabel metal2 s 36358 89840 36414 90040 6 Tile_X0Y0_FrameStrobe_O[8]
port 179 nsew signal output
rlabel metal2 s 36634 89840 36690 90040 6 Tile_X0Y0_FrameStrobe_O[9]
port 180 nsew signal output
rlabel metal2 s 5170 89840 5226 90040 6 Tile_X0Y0_N1BEG[0]
port 181 nsew signal output
rlabel metal2 s 5446 89840 5502 90040 6 Tile_X0Y0_N1BEG[1]
port 182 nsew signal output
rlabel metal2 s 5722 89840 5778 90040 6 Tile_X0Y0_N1BEG[2]
port 183 nsew signal output
rlabel metal2 s 5998 89840 6054 90040 6 Tile_X0Y0_N1BEG[3]
port 184 nsew signal output
rlabel metal2 s 6274 89840 6330 90040 6 Tile_X0Y0_N2BEG[0]
port 185 nsew signal output
rlabel metal2 s 6550 89840 6606 90040 6 Tile_X0Y0_N2BEG[1]
port 186 nsew signal output
rlabel metal2 s 6826 89840 6882 90040 6 Tile_X0Y0_N2BEG[2]
port 187 nsew signal output
rlabel metal2 s 7102 89840 7158 90040 6 Tile_X0Y0_N2BEG[3]
port 188 nsew signal output
rlabel metal2 s 7378 89840 7434 90040 6 Tile_X0Y0_N2BEG[4]
port 189 nsew signal output
rlabel metal2 s 7654 89840 7710 90040 6 Tile_X0Y0_N2BEG[5]
port 190 nsew signal output
rlabel metal2 s 7930 89840 7986 90040 6 Tile_X0Y0_N2BEG[6]
port 191 nsew signal output
rlabel metal2 s 8206 89840 8262 90040 6 Tile_X0Y0_N2BEG[7]
port 192 nsew signal output
rlabel metal2 s 8482 89840 8538 90040 6 Tile_X0Y0_N2BEGb[0]
port 193 nsew signal output
rlabel metal2 s 8758 89840 8814 90040 6 Tile_X0Y0_N2BEGb[1]
port 194 nsew signal output
rlabel metal2 s 9034 89840 9090 90040 6 Tile_X0Y0_N2BEGb[2]
port 195 nsew signal output
rlabel metal2 s 9310 89840 9366 90040 6 Tile_X0Y0_N2BEGb[3]
port 196 nsew signal output
rlabel metal2 s 9586 89840 9642 90040 6 Tile_X0Y0_N2BEGb[4]
port 197 nsew signal output
rlabel metal2 s 9862 89840 9918 90040 6 Tile_X0Y0_N2BEGb[5]
port 198 nsew signal output
rlabel metal2 s 10138 89840 10194 90040 6 Tile_X0Y0_N2BEGb[6]
port 199 nsew signal output
rlabel metal2 s 10414 89840 10470 90040 6 Tile_X0Y0_N2BEGb[7]
port 200 nsew signal output
rlabel metal2 s 10690 89840 10746 90040 6 Tile_X0Y0_N4BEG[0]
port 201 nsew signal output
rlabel metal2 s 13450 89840 13506 90040 6 Tile_X0Y0_N4BEG[10]
port 202 nsew signal output
rlabel metal2 s 13726 89840 13782 90040 6 Tile_X0Y0_N4BEG[11]
port 203 nsew signal output
rlabel metal2 s 14002 89840 14058 90040 6 Tile_X0Y0_N4BEG[12]
port 204 nsew signal output
rlabel metal2 s 14278 89840 14334 90040 6 Tile_X0Y0_N4BEG[13]
port 205 nsew signal output
rlabel metal2 s 14554 89840 14610 90040 6 Tile_X0Y0_N4BEG[14]
port 206 nsew signal output
rlabel metal2 s 14830 89840 14886 90040 6 Tile_X0Y0_N4BEG[15]
port 207 nsew signal output
rlabel metal2 s 10966 89840 11022 90040 6 Tile_X0Y0_N4BEG[1]
port 208 nsew signal output
rlabel metal2 s 11242 89840 11298 90040 6 Tile_X0Y0_N4BEG[2]
port 209 nsew signal output
rlabel metal2 s 11518 89840 11574 90040 6 Tile_X0Y0_N4BEG[3]
port 210 nsew signal output
rlabel metal2 s 11794 89840 11850 90040 6 Tile_X0Y0_N4BEG[4]
port 211 nsew signal output
rlabel metal2 s 12070 89840 12126 90040 6 Tile_X0Y0_N4BEG[5]
port 212 nsew signal output
rlabel metal2 s 12346 89840 12402 90040 6 Tile_X0Y0_N4BEG[6]
port 213 nsew signal output
rlabel metal2 s 12622 89840 12678 90040 6 Tile_X0Y0_N4BEG[7]
port 214 nsew signal output
rlabel metal2 s 12898 89840 12954 90040 6 Tile_X0Y0_N4BEG[8]
port 215 nsew signal output
rlabel metal2 s 13174 89840 13230 90040 6 Tile_X0Y0_N4BEG[9]
port 216 nsew signal output
rlabel metal2 s 15106 89840 15162 90040 6 Tile_X0Y0_NN4BEG[0]
port 217 nsew signal output
rlabel metal2 s 17866 89840 17922 90040 6 Tile_X0Y0_NN4BEG[10]
port 218 nsew signal output
rlabel metal2 s 18142 89840 18198 90040 6 Tile_X0Y0_NN4BEG[11]
port 219 nsew signal output
rlabel metal2 s 18418 89840 18474 90040 6 Tile_X0Y0_NN4BEG[12]
port 220 nsew signal output
rlabel metal2 s 18694 89840 18750 90040 6 Tile_X0Y0_NN4BEG[13]
port 221 nsew signal output
rlabel metal2 s 18970 89840 19026 90040 6 Tile_X0Y0_NN4BEG[14]
port 222 nsew signal output
rlabel metal2 s 19246 89840 19302 90040 6 Tile_X0Y0_NN4BEG[15]
port 223 nsew signal output
rlabel metal2 s 15382 89840 15438 90040 6 Tile_X0Y0_NN4BEG[1]
port 224 nsew signal output
rlabel metal2 s 15658 89840 15714 90040 6 Tile_X0Y0_NN4BEG[2]
port 225 nsew signal output
rlabel metal2 s 15934 89840 15990 90040 6 Tile_X0Y0_NN4BEG[3]
port 226 nsew signal output
rlabel metal2 s 16210 89840 16266 90040 6 Tile_X0Y0_NN4BEG[4]
port 227 nsew signal output
rlabel metal2 s 16486 89840 16542 90040 6 Tile_X0Y0_NN4BEG[5]
port 228 nsew signal output
rlabel metal2 s 16762 89840 16818 90040 6 Tile_X0Y0_NN4BEG[6]
port 229 nsew signal output
rlabel metal2 s 17038 89840 17094 90040 6 Tile_X0Y0_NN4BEG[7]
port 230 nsew signal output
rlabel metal2 s 17314 89840 17370 90040 6 Tile_X0Y0_NN4BEG[8]
port 231 nsew signal output
rlabel metal2 s 17590 89840 17646 90040 6 Tile_X0Y0_NN4BEG[9]
port 232 nsew signal output
rlabel metal2 s 19522 89840 19578 90040 6 Tile_X0Y0_S1END[0]
port 233 nsew signal input
rlabel metal2 s 19798 89840 19854 90040 6 Tile_X0Y0_S1END[1]
port 234 nsew signal input
rlabel metal2 s 20074 89840 20130 90040 6 Tile_X0Y0_S1END[2]
port 235 nsew signal input
rlabel metal2 s 20350 89840 20406 90040 6 Tile_X0Y0_S1END[3]
port 236 nsew signal input
rlabel metal2 s 20626 89840 20682 90040 6 Tile_X0Y0_S2END[0]
port 237 nsew signal input
rlabel metal2 s 20902 89840 20958 90040 6 Tile_X0Y0_S2END[1]
port 238 nsew signal input
rlabel metal2 s 21178 89840 21234 90040 6 Tile_X0Y0_S2END[2]
port 239 nsew signal input
rlabel metal2 s 21454 89840 21510 90040 6 Tile_X0Y0_S2END[3]
port 240 nsew signal input
rlabel metal2 s 21730 89840 21786 90040 6 Tile_X0Y0_S2END[4]
port 241 nsew signal input
rlabel metal2 s 22006 89840 22062 90040 6 Tile_X0Y0_S2END[5]
port 242 nsew signal input
rlabel metal2 s 22282 89840 22338 90040 6 Tile_X0Y0_S2END[6]
port 243 nsew signal input
rlabel metal2 s 22558 89840 22614 90040 6 Tile_X0Y0_S2END[7]
port 244 nsew signal input
rlabel metal2 s 22834 89840 22890 90040 6 Tile_X0Y0_S2MID[0]
port 245 nsew signal input
rlabel metal2 s 23110 89840 23166 90040 6 Tile_X0Y0_S2MID[1]
port 246 nsew signal input
rlabel metal2 s 23386 89840 23442 90040 6 Tile_X0Y0_S2MID[2]
port 247 nsew signal input
rlabel metal2 s 23662 89840 23718 90040 6 Tile_X0Y0_S2MID[3]
port 248 nsew signal input
rlabel metal2 s 23938 89840 23994 90040 6 Tile_X0Y0_S2MID[4]
port 249 nsew signal input
rlabel metal2 s 24214 89840 24270 90040 6 Tile_X0Y0_S2MID[5]
port 250 nsew signal input
rlabel metal2 s 24490 89840 24546 90040 6 Tile_X0Y0_S2MID[6]
port 251 nsew signal input
rlabel metal2 s 24766 89840 24822 90040 6 Tile_X0Y0_S2MID[7]
port 252 nsew signal input
rlabel metal2 s 25042 89840 25098 90040 6 Tile_X0Y0_S4END[0]
port 253 nsew signal input
rlabel metal2 s 27802 89840 27858 90040 6 Tile_X0Y0_S4END[10]
port 254 nsew signal input
rlabel metal2 s 28078 89840 28134 90040 6 Tile_X0Y0_S4END[11]
port 255 nsew signal input
rlabel metal2 s 28354 89840 28410 90040 6 Tile_X0Y0_S4END[12]
port 256 nsew signal input
rlabel metal2 s 28630 89840 28686 90040 6 Tile_X0Y0_S4END[13]
port 257 nsew signal input
rlabel metal2 s 28906 89840 28962 90040 6 Tile_X0Y0_S4END[14]
port 258 nsew signal input
rlabel metal2 s 29182 89840 29238 90040 6 Tile_X0Y0_S4END[15]
port 259 nsew signal input
rlabel metal2 s 25318 89840 25374 90040 6 Tile_X0Y0_S4END[1]
port 260 nsew signal input
rlabel metal2 s 25594 89840 25650 90040 6 Tile_X0Y0_S4END[2]
port 261 nsew signal input
rlabel metal2 s 25870 89840 25926 90040 6 Tile_X0Y0_S4END[3]
port 262 nsew signal input
rlabel metal2 s 26146 89840 26202 90040 6 Tile_X0Y0_S4END[4]
port 263 nsew signal input
rlabel metal2 s 26422 89840 26478 90040 6 Tile_X0Y0_S4END[5]
port 264 nsew signal input
rlabel metal2 s 26698 89840 26754 90040 6 Tile_X0Y0_S4END[6]
port 265 nsew signal input
rlabel metal2 s 26974 89840 27030 90040 6 Tile_X0Y0_S4END[7]
port 266 nsew signal input
rlabel metal2 s 27250 89840 27306 90040 6 Tile_X0Y0_S4END[8]
port 267 nsew signal input
rlabel metal2 s 27526 89840 27582 90040 6 Tile_X0Y0_S4END[9]
port 268 nsew signal input
rlabel metal2 s 29458 89840 29514 90040 6 Tile_X0Y0_SS4END[0]
port 269 nsew signal input
rlabel metal2 s 32218 89840 32274 90040 6 Tile_X0Y0_SS4END[10]
port 270 nsew signal input
rlabel metal2 s 32494 89840 32550 90040 6 Tile_X0Y0_SS4END[11]
port 271 nsew signal input
rlabel metal2 s 32770 89840 32826 90040 6 Tile_X0Y0_SS4END[12]
port 272 nsew signal input
rlabel metal2 s 33046 89840 33102 90040 6 Tile_X0Y0_SS4END[13]
port 273 nsew signal input
rlabel metal2 s 33322 89840 33378 90040 6 Tile_X0Y0_SS4END[14]
port 274 nsew signal input
rlabel metal2 s 33598 89840 33654 90040 6 Tile_X0Y0_SS4END[15]
port 275 nsew signal input
rlabel metal2 s 29734 89840 29790 90040 6 Tile_X0Y0_SS4END[1]
port 276 nsew signal input
rlabel metal2 s 30010 89840 30066 90040 6 Tile_X0Y0_SS4END[2]
port 277 nsew signal input
rlabel metal2 s 30286 89840 30342 90040 6 Tile_X0Y0_SS4END[3]
port 278 nsew signal input
rlabel metal2 s 30562 89840 30618 90040 6 Tile_X0Y0_SS4END[4]
port 279 nsew signal input
rlabel metal2 s 30838 89840 30894 90040 6 Tile_X0Y0_SS4END[5]
port 280 nsew signal input
rlabel metal2 s 31114 89840 31170 90040 6 Tile_X0Y0_SS4END[6]
port 281 nsew signal input
rlabel metal2 s 31390 89840 31446 90040 6 Tile_X0Y0_SS4END[7]
port 282 nsew signal input
rlabel metal2 s 31666 89840 31722 90040 6 Tile_X0Y0_SS4END[8]
port 283 nsew signal input
rlabel metal2 s 31942 89840 31998 90040 6 Tile_X0Y0_SS4END[9]
port 284 nsew signal input
rlabel metal2 s 33874 89840 33930 90040 6 Tile_X0Y0_UserCLKo
port 285 nsew signal output
rlabel metal3 s -40 50872 160 50992 6 Tile_X0Y0_W1BEG[0]
port 286 nsew signal output
rlabel metal3 s -40 51144 160 51264 6 Tile_X0Y0_W1BEG[1]
port 287 nsew signal output
rlabel metal3 s -40 51416 160 51536 6 Tile_X0Y0_W1BEG[2]
port 288 nsew signal output
rlabel metal3 s -40 51688 160 51808 6 Tile_X0Y0_W1BEG[3]
port 289 nsew signal output
rlabel metal3 s 44540 50872 44740 50992 6 Tile_X0Y0_W1END[0]
port 290 nsew signal input
rlabel metal3 s 44540 51144 44740 51264 6 Tile_X0Y0_W1END[1]
port 291 nsew signal input
rlabel metal3 s 44540 51416 44740 51536 6 Tile_X0Y0_W1END[2]
port 292 nsew signal input
rlabel metal3 s 44540 51688 44740 51808 6 Tile_X0Y0_W1END[3]
port 293 nsew signal input
rlabel metal3 s -40 51960 160 52080 6 Tile_X0Y0_W2BEG[0]
port 294 nsew signal output
rlabel metal3 s -40 52232 160 52352 6 Tile_X0Y0_W2BEG[1]
port 295 nsew signal output
rlabel metal3 s -40 52504 160 52624 6 Tile_X0Y0_W2BEG[2]
port 296 nsew signal output
rlabel metal3 s -40 52776 160 52896 6 Tile_X0Y0_W2BEG[3]
port 297 nsew signal output
rlabel metal3 s -40 53048 160 53168 6 Tile_X0Y0_W2BEG[4]
port 298 nsew signal output
rlabel metal3 s -40 53320 160 53440 6 Tile_X0Y0_W2BEG[5]
port 299 nsew signal output
rlabel metal3 s -40 53592 160 53712 6 Tile_X0Y0_W2BEG[6]
port 300 nsew signal output
rlabel metal3 s -40 53864 160 53984 6 Tile_X0Y0_W2BEG[7]
port 301 nsew signal output
rlabel metal3 s -40 54136 160 54256 6 Tile_X0Y0_W2BEGb[0]
port 302 nsew signal output
rlabel metal3 s -40 54408 160 54528 6 Tile_X0Y0_W2BEGb[1]
port 303 nsew signal output
rlabel metal3 s -40 54680 160 54800 6 Tile_X0Y0_W2BEGb[2]
port 304 nsew signal output
rlabel metal3 s -40 54952 160 55072 6 Tile_X0Y0_W2BEGb[3]
port 305 nsew signal output
rlabel metal3 s -40 55224 160 55344 6 Tile_X0Y0_W2BEGb[4]
port 306 nsew signal output
rlabel metal3 s -40 55496 160 55616 6 Tile_X0Y0_W2BEGb[5]
port 307 nsew signal output
rlabel metal3 s -40 55768 160 55888 6 Tile_X0Y0_W2BEGb[6]
port 308 nsew signal output
rlabel metal3 s -40 56040 160 56160 6 Tile_X0Y0_W2BEGb[7]
port 309 nsew signal output
rlabel metal3 s 44540 54136 44740 54256 6 Tile_X0Y0_W2END[0]
port 310 nsew signal input
rlabel metal3 s 44540 54408 44740 54528 6 Tile_X0Y0_W2END[1]
port 311 nsew signal input
rlabel metal3 s 44540 54680 44740 54800 6 Tile_X0Y0_W2END[2]
port 312 nsew signal input
rlabel metal3 s 44540 54952 44740 55072 6 Tile_X0Y0_W2END[3]
port 313 nsew signal input
rlabel metal3 s 44540 55224 44740 55344 6 Tile_X0Y0_W2END[4]
port 314 nsew signal input
rlabel metal3 s 44540 55496 44740 55616 6 Tile_X0Y0_W2END[5]
port 315 nsew signal input
rlabel metal3 s 44540 55768 44740 55888 6 Tile_X0Y0_W2END[6]
port 316 nsew signal input
rlabel metal3 s 44540 56040 44740 56160 6 Tile_X0Y0_W2END[7]
port 317 nsew signal input
rlabel metal3 s 44540 51960 44740 52080 6 Tile_X0Y0_W2MID[0]
port 318 nsew signal input
rlabel metal3 s 44540 52232 44740 52352 6 Tile_X0Y0_W2MID[1]
port 319 nsew signal input
rlabel metal3 s 44540 52504 44740 52624 6 Tile_X0Y0_W2MID[2]
port 320 nsew signal input
rlabel metal3 s 44540 52776 44740 52896 6 Tile_X0Y0_W2MID[3]
port 321 nsew signal input
rlabel metal3 s 44540 53048 44740 53168 6 Tile_X0Y0_W2MID[4]
port 322 nsew signal input
rlabel metal3 s 44540 53320 44740 53440 6 Tile_X0Y0_W2MID[5]
port 323 nsew signal input
rlabel metal3 s 44540 53592 44740 53712 6 Tile_X0Y0_W2MID[6]
port 324 nsew signal input
rlabel metal3 s 44540 53864 44740 53984 6 Tile_X0Y0_W2MID[7]
port 325 nsew signal input
rlabel metal3 s -40 60664 160 60784 6 Tile_X0Y0_W6BEG[0]
port 326 nsew signal output
rlabel metal3 s -40 63384 160 63504 6 Tile_X0Y0_W6BEG[10]
port 327 nsew signal output
rlabel metal3 s -40 63656 160 63776 6 Tile_X0Y0_W6BEG[11]
port 328 nsew signal output
rlabel metal3 s -40 60936 160 61056 6 Tile_X0Y0_W6BEG[1]
port 329 nsew signal output
rlabel metal3 s -40 61208 160 61328 6 Tile_X0Y0_W6BEG[2]
port 330 nsew signal output
rlabel metal3 s -40 61480 160 61600 6 Tile_X0Y0_W6BEG[3]
port 331 nsew signal output
rlabel metal3 s -40 61752 160 61872 6 Tile_X0Y0_W6BEG[4]
port 332 nsew signal output
rlabel metal3 s -40 62024 160 62144 6 Tile_X0Y0_W6BEG[5]
port 333 nsew signal output
rlabel metal3 s -40 62296 160 62416 6 Tile_X0Y0_W6BEG[6]
port 334 nsew signal output
rlabel metal3 s -40 62568 160 62688 6 Tile_X0Y0_W6BEG[7]
port 335 nsew signal output
rlabel metal3 s -40 62840 160 62960 6 Tile_X0Y0_W6BEG[8]
port 336 nsew signal output
rlabel metal3 s -40 63112 160 63232 6 Tile_X0Y0_W6BEG[9]
port 337 nsew signal output
rlabel metal3 s 44540 60664 44740 60784 6 Tile_X0Y0_W6END[0]
port 338 nsew signal input
rlabel metal3 s 44540 63384 44740 63504 6 Tile_X0Y0_W6END[10]
port 339 nsew signal input
rlabel metal3 s 44540 63656 44740 63776 6 Tile_X0Y0_W6END[11]
port 340 nsew signal input
rlabel metal3 s 44540 60936 44740 61056 6 Tile_X0Y0_W6END[1]
port 341 nsew signal input
rlabel metal3 s 44540 61208 44740 61328 6 Tile_X0Y0_W6END[2]
port 342 nsew signal input
rlabel metal3 s 44540 61480 44740 61600 6 Tile_X0Y0_W6END[3]
port 343 nsew signal input
rlabel metal3 s 44540 61752 44740 61872 6 Tile_X0Y0_W6END[4]
port 344 nsew signal input
rlabel metal3 s 44540 62024 44740 62144 6 Tile_X0Y0_W6END[5]
port 345 nsew signal input
rlabel metal3 s 44540 62296 44740 62416 6 Tile_X0Y0_W6END[6]
port 346 nsew signal input
rlabel metal3 s 44540 62568 44740 62688 6 Tile_X0Y0_W6END[7]
port 347 nsew signal input
rlabel metal3 s 44540 62840 44740 62960 6 Tile_X0Y0_W6END[8]
port 348 nsew signal input
rlabel metal3 s 44540 63112 44740 63232 6 Tile_X0Y0_W6END[9]
port 349 nsew signal input
rlabel metal3 s -40 56312 160 56432 6 Tile_X0Y0_WW4BEG[0]
port 350 nsew signal output
rlabel metal3 s -40 59032 160 59152 6 Tile_X0Y0_WW4BEG[10]
port 351 nsew signal output
rlabel metal3 s -40 59304 160 59424 6 Tile_X0Y0_WW4BEG[11]
port 352 nsew signal output
rlabel metal3 s -40 59576 160 59696 6 Tile_X0Y0_WW4BEG[12]
port 353 nsew signal output
rlabel metal3 s -40 59848 160 59968 6 Tile_X0Y0_WW4BEG[13]
port 354 nsew signal output
rlabel metal3 s -40 60120 160 60240 6 Tile_X0Y0_WW4BEG[14]
port 355 nsew signal output
rlabel metal3 s -40 60392 160 60512 6 Tile_X0Y0_WW4BEG[15]
port 356 nsew signal output
rlabel metal3 s -40 56584 160 56704 6 Tile_X0Y0_WW4BEG[1]
port 357 nsew signal output
rlabel metal3 s -40 56856 160 56976 6 Tile_X0Y0_WW4BEG[2]
port 358 nsew signal output
rlabel metal3 s -40 57128 160 57248 6 Tile_X0Y0_WW4BEG[3]
port 359 nsew signal output
rlabel metal3 s -40 57400 160 57520 6 Tile_X0Y0_WW4BEG[4]
port 360 nsew signal output
rlabel metal3 s -40 57672 160 57792 6 Tile_X0Y0_WW4BEG[5]
port 361 nsew signal output
rlabel metal3 s -40 57944 160 58064 6 Tile_X0Y0_WW4BEG[6]
port 362 nsew signal output
rlabel metal3 s -40 58216 160 58336 6 Tile_X0Y0_WW4BEG[7]
port 363 nsew signal output
rlabel metal3 s -40 58488 160 58608 6 Tile_X0Y0_WW4BEG[8]
port 364 nsew signal output
rlabel metal3 s -40 58760 160 58880 6 Tile_X0Y0_WW4BEG[9]
port 365 nsew signal output
rlabel metal3 s 44540 56312 44740 56432 6 Tile_X0Y0_WW4END[0]
port 366 nsew signal input
rlabel metal3 s 44540 59032 44740 59152 6 Tile_X0Y0_WW4END[10]
port 367 nsew signal input
rlabel metal3 s 44540 59304 44740 59424 6 Tile_X0Y0_WW4END[11]
port 368 nsew signal input
rlabel metal3 s 44540 59576 44740 59696 6 Tile_X0Y0_WW4END[12]
port 369 nsew signal input
rlabel metal3 s 44540 59848 44740 59968 6 Tile_X0Y0_WW4END[13]
port 370 nsew signal input
rlabel metal3 s 44540 60120 44740 60240 6 Tile_X0Y0_WW4END[14]
port 371 nsew signal input
rlabel metal3 s 44540 60392 44740 60512 6 Tile_X0Y0_WW4END[15]
port 372 nsew signal input
rlabel metal3 s 44540 56584 44740 56704 6 Tile_X0Y0_WW4END[1]
port 373 nsew signal input
rlabel metal3 s 44540 56856 44740 56976 6 Tile_X0Y0_WW4END[2]
port 374 nsew signal input
rlabel metal3 s 44540 57128 44740 57248 6 Tile_X0Y0_WW4END[3]
port 375 nsew signal input
rlabel metal3 s 44540 57400 44740 57520 6 Tile_X0Y0_WW4END[4]
port 376 nsew signal input
rlabel metal3 s 44540 57672 44740 57792 6 Tile_X0Y0_WW4END[5]
port 377 nsew signal input
rlabel metal3 s 44540 57944 44740 58064 6 Tile_X0Y0_WW4END[6]
port 378 nsew signal input
rlabel metal3 s 44540 58216 44740 58336 6 Tile_X0Y0_WW4END[7]
port 379 nsew signal input
rlabel metal3 s 44540 58488 44740 58608 6 Tile_X0Y0_WW4END[8]
port 380 nsew signal input
rlabel metal3 s 44540 58760 44740 58880 6 Tile_X0Y0_WW4END[9]
port 381 nsew signal input
rlabel metal3 s 44540 17960 44740 18080 6 Tile_X0Y1_E1BEG[0]
port 382 nsew signal output
rlabel metal3 s 44540 18232 44740 18352 6 Tile_X0Y1_E1BEG[1]
port 383 nsew signal output
rlabel metal3 s 44540 18504 44740 18624 6 Tile_X0Y1_E1BEG[2]
port 384 nsew signal output
rlabel metal3 s 44540 18776 44740 18896 6 Tile_X0Y1_E1BEG[3]
port 385 nsew signal output
rlabel metal3 s -40 17960 160 18080 6 Tile_X0Y1_E1END[0]
port 386 nsew signal input
rlabel metal3 s -40 18232 160 18352 6 Tile_X0Y1_E1END[1]
port 387 nsew signal input
rlabel metal3 s -40 18504 160 18624 6 Tile_X0Y1_E1END[2]
port 388 nsew signal input
rlabel metal3 s -40 18776 160 18896 6 Tile_X0Y1_E1END[3]
port 389 nsew signal input
rlabel metal3 s 44540 19048 44740 19168 6 Tile_X0Y1_E2BEG[0]
port 390 nsew signal output
rlabel metal3 s 44540 19320 44740 19440 6 Tile_X0Y1_E2BEG[1]
port 391 nsew signal output
rlabel metal3 s 44540 19592 44740 19712 6 Tile_X0Y1_E2BEG[2]
port 392 nsew signal output
rlabel metal3 s 44540 19864 44740 19984 6 Tile_X0Y1_E2BEG[3]
port 393 nsew signal output
rlabel metal3 s 44540 20136 44740 20256 6 Tile_X0Y1_E2BEG[4]
port 394 nsew signal output
rlabel metal3 s 44540 20408 44740 20528 6 Tile_X0Y1_E2BEG[5]
port 395 nsew signal output
rlabel metal3 s 44540 20680 44740 20800 6 Tile_X0Y1_E2BEG[6]
port 396 nsew signal output
rlabel metal3 s 44540 20952 44740 21072 6 Tile_X0Y1_E2BEG[7]
port 397 nsew signal output
rlabel metal3 s 44540 21224 44740 21344 6 Tile_X0Y1_E2BEGb[0]
port 398 nsew signal output
rlabel metal3 s 44540 21496 44740 21616 6 Tile_X0Y1_E2BEGb[1]
port 399 nsew signal output
rlabel metal3 s 44540 21768 44740 21888 6 Tile_X0Y1_E2BEGb[2]
port 400 nsew signal output
rlabel metal3 s 44540 22040 44740 22160 6 Tile_X0Y1_E2BEGb[3]
port 401 nsew signal output
rlabel metal3 s 44540 22312 44740 22432 6 Tile_X0Y1_E2BEGb[4]
port 402 nsew signal output
rlabel metal3 s 44540 22584 44740 22704 6 Tile_X0Y1_E2BEGb[5]
port 403 nsew signal output
rlabel metal3 s 44540 22856 44740 22976 6 Tile_X0Y1_E2BEGb[6]
port 404 nsew signal output
rlabel metal3 s 44540 23128 44740 23248 6 Tile_X0Y1_E2BEGb[7]
port 405 nsew signal output
rlabel metal3 s -40 21224 160 21344 6 Tile_X0Y1_E2END[0]
port 406 nsew signal input
rlabel metal3 s -40 21496 160 21616 6 Tile_X0Y1_E2END[1]
port 407 nsew signal input
rlabel metal3 s -40 21768 160 21888 6 Tile_X0Y1_E2END[2]
port 408 nsew signal input
rlabel metal3 s -40 22040 160 22160 6 Tile_X0Y1_E2END[3]
port 409 nsew signal input
rlabel metal3 s -40 22312 160 22432 6 Tile_X0Y1_E2END[4]
port 410 nsew signal input
rlabel metal3 s -40 22584 160 22704 6 Tile_X0Y1_E2END[5]
port 411 nsew signal input
rlabel metal3 s -40 22856 160 22976 6 Tile_X0Y1_E2END[6]
port 412 nsew signal input
rlabel metal3 s -40 23128 160 23248 6 Tile_X0Y1_E2END[7]
port 413 nsew signal input
rlabel metal3 s -40 19048 160 19168 6 Tile_X0Y1_E2MID[0]
port 414 nsew signal input
rlabel metal3 s -40 19320 160 19440 6 Tile_X0Y1_E2MID[1]
port 415 nsew signal input
rlabel metal3 s -40 19592 160 19712 6 Tile_X0Y1_E2MID[2]
port 416 nsew signal input
rlabel metal3 s -40 19864 160 19984 6 Tile_X0Y1_E2MID[3]
port 417 nsew signal input
rlabel metal3 s -40 20136 160 20256 6 Tile_X0Y1_E2MID[4]
port 418 nsew signal input
rlabel metal3 s -40 20408 160 20528 6 Tile_X0Y1_E2MID[5]
port 419 nsew signal input
rlabel metal3 s -40 20680 160 20800 6 Tile_X0Y1_E2MID[6]
port 420 nsew signal input
rlabel metal3 s -40 20952 160 21072 6 Tile_X0Y1_E2MID[7]
port 421 nsew signal input
rlabel metal3 s 44540 27752 44740 27872 6 Tile_X0Y1_E6BEG[0]
port 422 nsew signal output
rlabel metal3 s 44540 30472 44740 30592 6 Tile_X0Y1_E6BEG[10]
port 423 nsew signal output
rlabel metal3 s 44540 30744 44740 30864 6 Tile_X0Y1_E6BEG[11]
port 424 nsew signal output
rlabel metal3 s 44540 28024 44740 28144 6 Tile_X0Y1_E6BEG[1]
port 425 nsew signal output
rlabel metal3 s 44540 28296 44740 28416 6 Tile_X0Y1_E6BEG[2]
port 426 nsew signal output
rlabel metal3 s 44540 28568 44740 28688 6 Tile_X0Y1_E6BEG[3]
port 427 nsew signal output
rlabel metal3 s 44540 28840 44740 28960 6 Tile_X0Y1_E6BEG[4]
port 428 nsew signal output
rlabel metal3 s 44540 29112 44740 29232 6 Tile_X0Y1_E6BEG[5]
port 429 nsew signal output
rlabel metal3 s 44540 29384 44740 29504 6 Tile_X0Y1_E6BEG[6]
port 430 nsew signal output
rlabel metal3 s 44540 29656 44740 29776 6 Tile_X0Y1_E6BEG[7]
port 431 nsew signal output
rlabel metal3 s 44540 29928 44740 30048 6 Tile_X0Y1_E6BEG[8]
port 432 nsew signal output
rlabel metal3 s 44540 30200 44740 30320 6 Tile_X0Y1_E6BEG[9]
port 433 nsew signal output
rlabel metal3 s -40 27752 160 27872 6 Tile_X0Y1_E6END[0]
port 434 nsew signal input
rlabel metal3 s -40 30472 160 30592 6 Tile_X0Y1_E6END[10]
port 435 nsew signal input
rlabel metal3 s -40 30744 160 30864 6 Tile_X0Y1_E6END[11]
port 436 nsew signal input
rlabel metal3 s -40 28024 160 28144 6 Tile_X0Y1_E6END[1]
port 437 nsew signal input
rlabel metal3 s -40 28296 160 28416 6 Tile_X0Y1_E6END[2]
port 438 nsew signal input
rlabel metal3 s -40 28568 160 28688 6 Tile_X0Y1_E6END[3]
port 439 nsew signal input
rlabel metal3 s -40 28840 160 28960 6 Tile_X0Y1_E6END[4]
port 440 nsew signal input
rlabel metal3 s -40 29112 160 29232 6 Tile_X0Y1_E6END[5]
port 441 nsew signal input
rlabel metal3 s -40 29384 160 29504 6 Tile_X0Y1_E6END[6]
port 442 nsew signal input
rlabel metal3 s -40 29656 160 29776 6 Tile_X0Y1_E6END[7]
port 443 nsew signal input
rlabel metal3 s -40 29928 160 30048 6 Tile_X0Y1_E6END[8]
port 444 nsew signal input
rlabel metal3 s -40 30200 160 30320 6 Tile_X0Y1_E6END[9]
port 445 nsew signal input
rlabel metal3 s 44540 23400 44740 23520 6 Tile_X0Y1_EE4BEG[0]
port 446 nsew signal output
rlabel metal3 s 44540 26120 44740 26240 6 Tile_X0Y1_EE4BEG[10]
port 447 nsew signal output
rlabel metal3 s 44540 26392 44740 26512 6 Tile_X0Y1_EE4BEG[11]
port 448 nsew signal output
rlabel metal3 s 44540 26664 44740 26784 6 Tile_X0Y1_EE4BEG[12]
port 449 nsew signal output
rlabel metal3 s 44540 26936 44740 27056 6 Tile_X0Y1_EE4BEG[13]
port 450 nsew signal output
rlabel metal3 s 44540 27208 44740 27328 6 Tile_X0Y1_EE4BEG[14]
port 451 nsew signal output
rlabel metal3 s 44540 27480 44740 27600 6 Tile_X0Y1_EE4BEG[15]
port 452 nsew signal output
rlabel metal3 s 44540 23672 44740 23792 6 Tile_X0Y1_EE4BEG[1]
port 453 nsew signal output
rlabel metal3 s 44540 23944 44740 24064 6 Tile_X0Y1_EE4BEG[2]
port 454 nsew signal output
rlabel metal3 s 44540 24216 44740 24336 6 Tile_X0Y1_EE4BEG[3]
port 455 nsew signal output
rlabel metal3 s 44540 24488 44740 24608 6 Tile_X0Y1_EE4BEG[4]
port 456 nsew signal output
rlabel metal3 s 44540 24760 44740 24880 6 Tile_X0Y1_EE4BEG[5]
port 457 nsew signal output
rlabel metal3 s 44540 25032 44740 25152 6 Tile_X0Y1_EE4BEG[6]
port 458 nsew signal output
rlabel metal3 s 44540 25304 44740 25424 6 Tile_X0Y1_EE4BEG[7]
port 459 nsew signal output
rlabel metal3 s 44540 25576 44740 25696 6 Tile_X0Y1_EE4BEG[8]
port 460 nsew signal output
rlabel metal3 s 44540 25848 44740 25968 6 Tile_X0Y1_EE4BEG[9]
port 461 nsew signal output
rlabel metal3 s -40 23400 160 23520 6 Tile_X0Y1_EE4END[0]
port 462 nsew signal input
rlabel metal3 s -40 26120 160 26240 6 Tile_X0Y1_EE4END[10]
port 463 nsew signal input
rlabel metal3 s -40 26392 160 26512 6 Tile_X0Y1_EE4END[11]
port 464 nsew signal input
rlabel metal3 s -40 26664 160 26784 6 Tile_X0Y1_EE4END[12]
port 465 nsew signal input
rlabel metal3 s -40 26936 160 27056 6 Tile_X0Y1_EE4END[13]
port 466 nsew signal input
rlabel metal3 s -40 27208 160 27328 6 Tile_X0Y1_EE4END[14]
port 467 nsew signal input
rlabel metal3 s -40 27480 160 27600 6 Tile_X0Y1_EE4END[15]
port 468 nsew signal input
rlabel metal3 s -40 23672 160 23792 6 Tile_X0Y1_EE4END[1]
port 469 nsew signal input
rlabel metal3 s -40 23944 160 24064 6 Tile_X0Y1_EE4END[2]
port 470 nsew signal input
rlabel metal3 s -40 24216 160 24336 6 Tile_X0Y1_EE4END[3]
port 471 nsew signal input
rlabel metal3 s -40 24488 160 24608 6 Tile_X0Y1_EE4END[4]
port 472 nsew signal input
rlabel metal3 s -40 24760 160 24880 6 Tile_X0Y1_EE4END[5]
port 473 nsew signal input
rlabel metal3 s -40 25032 160 25152 6 Tile_X0Y1_EE4END[6]
port 474 nsew signal input
rlabel metal3 s -40 25304 160 25424 6 Tile_X0Y1_EE4END[7]
port 475 nsew signal input
rlabel metal3 s -40 25576 160 25696 6 Tile_X0Y1_EE4END[8]
port 476 nsew signal input
rlabel metal3 s -40 25848 160 25968 6 Tile_X0Y1_EE4END[9]
port 477 nsew signal input
rlabel metal3 s -40 31016 160 31136 6 Tile_X0Y1_FrameData[0]
port 478 nsew signal input
rlabel metal3 s -40 33736 160 33856 6 Tile_X0Y1_FrameData[10]
port 479 nsew signal input
rlabel metal3 s -40 34008 160 34128 6 Tile_X0Y1_FrameData[11]
port 480 nsew signal input
rlabel metal3 s -40 34280 160 34400 6 Tile_X0Y1_FrameData[12]
port 481 nsew signal input
rlabel metal3 s -40 34552 160 34672 6 Tile_X0Y1_FrameData[13]
port 482 nsew signal input
rlabel metal3 s -40 34824 160 34944 6 Tile_X0Y1_FrameData[14]
port 483 nsew signal input
rlabel metal3 s -40 35096 160 35216 6 Tile_X0Y1_FrameData[15]
port 484 nsew signal input
rlabel metal3 s -40 35368 160 35488 6 Tile_X0Y1_FrameData[16]
port 485 nsew signal input
rlabel metal3 s -40 35640 160 35760 6 Tile_X0Y1_FrameData[17]
port 486 nsew signal input
rlabel metal3 s -40 35912 160 36032 6 Tile_X0Y1_FrameData[18]
port 487 nsew signal input
rlabel metal3 s -40 36184 160 36304 6 Tile_X0Y1_FrameData[19]
port 488 nsew signal input
rlabel metal3 s -40 31288 160 31408 6 Tile_X0Y1_FrameData[1]
port 489 nsew signal input
rlabel metal3 s -40 36456 160 36576 6 Tile_X0Y1_FrameData[20]
port 490 nsew signal input
rlabel metal3 s -40 36728 160 36848 6 Tile_X0Y1_FrameData[21]
port 491 nsew signal input
rlabel metal3 s -40 37000 160 37120 6 Tile_X0Y1_FrameData[22]
port 492 nsew signal input
rlabel metal3 s -40 37272 160 37392 6 Tile_X0Y1_FrameData[23]
port 493 nsew signal input
rlabel metal3 s -40 37544 160 37664 6 Tile_X0Y1_FrameData[24]
port 494 nsew signal input
rlabel metal3 s -40 37816 160 37936 6 Tile_X0Y1_FrameData[25]
port 495 nsew signal input
rlabel metal3 s -40 38088 160 38208 6 Tile_X0Y1_FrameData[26]
port 496 nsew signal input
rlabel metal3 s -40 38360 160 38480 6 Tile_X0Y1_FrameData[27]
port 497 nsew signal input
rlabel metal3 s -40 38632 160 38752 6 Tile_X0Y1_FrameData[28]
port 498 nsew signal input
rlabel metal3 s -40 38904 160 39024 6 Tile_X0Y1_FrameData[29]
port 499 nsew signal input
rlabel metal3 s -40 31560 160 31680 6 Tile_X0Y1_FrameData[2]
port 500 nsew signal input
rlabel metal3 s -40 39176 160 39296 6 Tile_X0Y1_FrameData[30]
port 501 nsew signal input
rlabel metal3 s -40 39448 160 39568 6 Tile_X0Y1_FrameData[31]
port 502 nsew signal input
rlabel metal3 s -40 31832 160 31952 6 Tile_X0Y1_FrameData[3]
port 503 nsew signal input
rlabel metal3 s -40 32104 160 32224 6 Tile_X0Y1_FrameData[4]
port 504 nsew signal input
rlabel metal3 s -40 32376 160 32496 6 Tile_X0Y1_FrameData[5]
port 505 nsew signal input
rlabel metal3 s -40 32648 160 32768 6 Tile_X0Y1_FrameData[6]
port 506 nsew signal input
rlabel metal3 s -40 32920 160 33040 6 Tile_X0Y1_FrameData[7]
port 507 nsew signal input
rlabel metal3 s -40 33192 160 33312 6 Tile_X0Y1_FrameData[8]
port 508 nsew signal input
rlabel metal3 s -40 33464 160 33584 6 Tile_X0Y1_FrameData[9]
port 509 nsew signal input
rlabel metal3 s 44540 31016 44740 31136 6 Tile_X0Y1_FrameData_O[0]
port 510 nsew signal output
rlabel metal3 s 44540 33736 44740 33856 6 Tile_X0Y1_FrameData_O[10]
port 511 nsew signal output
rlabel metal3 s 44540 34008 44740 34128 6 Tile_X0Y1_FrameData_O[11]
port 512 nsew signal output
rlabel metal3 s 44540 34280 44740 34400 6 Tile_X0Y1_FrameData_O[12]
port 513 nsew signal output
rlabel metal3 s 44540 34552 44740 34672 6 Tile_X0Y1_FrameData_O[13]
port 514 nsew signal output
rlabel metal3 s 44540 34824 44740 34944 6 Tile_X0Y1_FrameData_O[14]
port 515 nsew signal output
rlabel metal3 s 44540 35096 44740 35216 6 Tile_X0Y1_FrameData_O[15]
port 516 nsew signal output
rlabel metal3 s 44540 35368 44740 35488 6 Tile_X0Y1_FrameData_O[16]
port 517 nsew signal output
rlabel metal3 s 44540 35640 44740 35760 6 Tile_X0Y1_FrameData_O[17]
port 518 nsew signal output
rlabel metal3 s 44540 35912 44740 36032 6 Tile_X0Y1_FrameData_O[18]
port 519 nsew signal output
rlabel metal3 s 44540 36184 44740 36304 6 Tile_X0Y1_FrameData_O[19]
port 520 nsew signal output
rlabel metal3 s 44540 31288 44740 31408 6 Tile_X0Y1_FrameData_O[1]
port 521 nsew signal output
rlabel metal3 s 44540 36456 44740 36576 6 Tile_X0Y1_FrameData_O[20]
port 522 nsew signal output
rlabel metal3 s 44540 36728 44740 36848 6 Tile_X0Y1_FrameData_O[21]
port 523 nsew signal output
rlabel metal3 s 44540 37000 44740 37120 6 Tile_X0Y1_FrameData_O[22]
port 524 nsew signal output
rlabel metal3 s 44540 37272 44740 37392 6 Tile_X0Y1_FrameData_O[23]
port 525 nsew signal output
rlabel metal3 s 44540 37544 44740 37664 6 Tile_X0Y1_FrameData_O[24]
port 526 nsew signal output
rlabel metal3 s 44540 37816 44740 37936 6 Tile_X0Y1_FrameData_O[25]
port 527 nsew signal output
rlabel metal3 s 44540 38088 44740 38208 6 Tile_X0Y1_FrameData_O[26]
port 528 nsew signal output
rlabel metal3 s 44540 38360 44740 38480 6 Tile_X0Y1_FrameData_O[27]
port 529 nsew signal output
rlabel metal3 s 44540 38632 44740 38752 6 Tile_X0Y1_FrameData_O[28]
port 530 nsew signal output
rlabel metal3 s 44540 38904 44740 39024 6 Tile_X0Y1_FrameData_O[29]
port 531 nsew signal output
rlabel metal3 s 44540 31560 44740 31680 6 Tile_X0Y1_FrameData_O[2]
port 532 nsew signal output
rlabel metal3 s 44540 39176 44740 39296 6 Tile_X0Y1_FrameData_O[30]
port 533 nsew signal output
rlabel metal3 s 44540 39448 44740 39568 6 Tile_X0Y1_FrameData_O[31]
port 534 nsew signal output
rlabel metal3 s 44540 31832 44740 31952 6 Tile_X0Y1_FrameData_O[3]
port 535 nsew signal output
rlabel metal3 s 44540 32104 44740 32224 6 Tile_X0Y1_FrameData_O[4]
port 536 nsew signal output
rlabel metal3 s 44540 32376 44740 32496 6 Tile_X0Y1_FrameData_O[5]
port 537 nsew signal output
rlabel metal3 s 44540 32648 44740 32768 6 Tile_X0Y1_FrameData_O[6]
port 538 nsew signal output
rlabel metal3 s 44540 32920 44740 33040 6 Tile_X0Y1_FrameData_O[7]
port 539 nsew signal output
rlabel metal3 s 44540 33192 44740 33312 6 Tile_X0Y1_FrameData_O[8]
port 540 nsew signal output
rlabel metal3 s 44540 33464 44740 33584 6 Tile_X0Y1_FrameData_O[9]
port 541 nsew signal output
rlabel metal2 s 34150 -40 34206 160 6 Tile_X0Y1_FrameStrobe[0]
port 542 nsew signal input
rlabel metal2 s 36910 -40 36966 160 6 Tile_X0Y1_FrameStrobe[10]
port 543 nsew signal input
rlabel metal2 s 37186 -40 37242 160 6 Tile_X0Y1_FrameStrobe[11]
port 544 nsew signal input
rlabel metal2 s 37462 -40 37518 160 6 Tile_X0Y1_FrameStrobe[12]
port 545 nsew signal input
rlabel metal2 s 37738 -40 37794 160 6 Tile_X0Y1_FrameStrobe[13]
port 546 nsew signal input
rlabel metal2 s 38014 -40 38070 160 6 Tile_X0Y1_FrameStrobe[14]
port 547 nsew signal input
rlabel metal2 s 38290 -40 38346 160 6 Tile_X0Y1_FrameStrobe[15]
port 548 nsew signal input
rlabel metal2 s 38566 -40 38622 160 6 Tile_X0Y1_FrameStrobe[16]
port 549 nsew signal input
rlabel metal2 s 38842 -40 38898 160 6 Tile_X0Y1_FrameStrobe[17]
port 550 nsew signal input
rlabel metal2 s 39118 -40 39174 160 6 Tile_X0Y1_FrameStrobe[18]
port 551 nsew signal input
rlabel metal2 s 39394 -40 39450 160 6 Tile_X0Y1_FrameStrobe[19]
port 552 nsew signal input
rlabel metal2 s 34426 -40 34482 160 6 Tile_X0Y1_FrameStrobe[1]
port 553 nsew signal input
rlabel metal2 s 34702 -40 34758 160 6 Tile_X0Y1_FrameStrobe[2]
port 554 nsew signal input
rlabel metal2 s 34978 -40 35034 160 6 Tile_X0Y1_FrameStrobe[3]
port 555 nsew signal input
rlabel metal2 s 35254 -40 35310 160 6 Tile_X0Y1_FrameStrobe[4]
port 556 nsew signal input
rlabel metal2 s 35530 -40 35586 160 6 Tile_X0Y1_FrameStrobe[5]
port 557 nsew signal input
rlabel metal2 s 35806 -40 35862 160 6 Tile_X0Y1_FrameStrobe[6]
port 558 nsew signal input
rlabel metal2 s 36082 -40 36138 160 6 Tile_X0Y1_FrameStrobe[7]
port 559 nsew signal input
rlabel metal2 s 36358 -40 36414 160 6 Tile_X0Y1_FrameStrobe[8]
port 560 nsew signal input
rlabel metal2 s 36634 -40 36690 160 6 Tile_X0Y1_FrameStrobe[9]
port 561 nsew signal input
rlabel metal2 s 5170 -40 5226 160 6 Tile_X0Y1_N1END[0]
port 562 nsew signal input
rlabel metal2 s 5446 -40 5502 160 6 Tile_X0Y1_N1END[1]
port 563 nsew signal input
rlabel metal2 s 5722 -40 5778 160 6 Tile_X0Y1_N1END[2]
port 564 nsew signal input
rlabel metal2 s 5998 -40 6054 160 6 Tile_X0Y1_N1END[3]
port 565 nsew signal input
rlabel metal2 s 8482 -40 8538 160 6 Tile_X0Y1_N2END[0]
port 566 nsew signal input
rlabel metal2 s 8758 -40 8814 160 6 Tile_X0Y1_N2END[1]
port 567 nsew signal input
rlabel metal2 s 9034 -40 9090 160 6 Tile_X0Y1_N2END[2]
port 568 nsew signal input
rlabel metal2 s 9310 -40 9366 160 6 Tile_X0Y1_N2END[3]
port 569 nsew signal input
rlabel metal2 s 9586 -40 9642 160 6 Tile_X0Y1_N2END[4]
port 570 nsew signal input
rlabel metal2 s 9862 -40 9918 160 6 Tile_X0Y1_N2END[5]
port 571 nsew signal input
rlabel metal2 s 10138 -40 10194 160 6 Tile_X0Y1_N2END[6]
port 572 nsew signal input
rlabel metal2 s 10414 -40 10470 160 6 Tile_X0Y1_N2END[7]
port 573 nsew signal input
rlabel metal2 s 6274 -40 6330 160 6 Tile_X0Y1_N2MID[0]
port 574 nsew signal input
rlabel metal2 s 6550 -40 6606 160 6 Tile_X0Y1_N2MID[1]
port 575 nsew signal input
rlabel metal2 s 6826 -40 6882 160 6 Tile_X0Y1_N2MID[2]
port 576 nsew signal input
rlabel metal2 s 7102 -40 7158 160 6 Tile_X0Y1_N2MID[3]
port 577 nsew signal input
rlabel metal2 s 7378 -40 7434 160 6 Tile_X0Y1_N2MID[4]
port 578 nsew signal input
rlabel metal2 s 7654 -40 7710 160 6 Tile_X0Y1_N2MID[5]
port 579 nsew signal input
rlabel metal2 s 7930 -40 7986 160 6 Tile_X0Y1_N2MID[6]
port 580 nsew signal input
rlabel metal2 s 8206 -40 8262 160 6 Tile_X0Y1_N2MID[7]
port 581 nsew signal input
rlabel metal2 s 10690 -40 10746 160 6 Tile_X0Y1_N4END[0]
port 582 nsew signal input
rlabel metal2 s 13450 -40 13506 160 6 Tile_X0Y1_N4END[10]
port 583 nsew signal input
rlabel metal2 s 13726 -40 13782 160 6 Tile_X0Y1_N4END[11]
port 584 nsew signal input
rlabel metal2 s 14002 -40 14058 160 6 Tile_X0Y1_N4END[12]
port 585 nsew signal input
rlabel metal2 s 14278 -40 14334 160 6 Tile_X0Y1_N4END[13]
port 586 nsew signal input
rlabel metal2 s 14554 -40 14610 160 6 Tile_X0Y1_N4END[14]
port 587 nsew signal input
rlabel metal2 s 14830 -40 14886 160 6 Tile_X0Y1_N4END[15]
port 588 nsew signal input
rlabel metal2 s 10966 -40 11022 160 6 Tile_X0Y1_N4END[1]
port 589 nsew signal input
rlabel metal2 s 11242 -40 11298 160 6 Tile_X0Y1_N4END[2]
port 590 nsew signal input
rlabel metal2 s 11518 -40 11574 160 6 Tile_X0Y1_N4END[3]
port 591 nsew signal input
rlabel metal2 s 11794 -40 11850 160 6 Tile_X0Y1_N4END[4]
port 592 nsew signal input
rlabel metal2 s 12070 -40 12126 160 6 Tile_X0Y1_N4END[5]
port 593 nsew signal input
rlabel metal2 s 12346 -40 12402 160 6 Tile_X0Y1_N4END[6]
port 594 nsew signal input
rlabel metal2 s 12622 -40 12678 160 6 Tile_X0Y1_N4END[7]
port 595 nsew signal input
rlabel metal2 s 12898 -40 12954 160 6 Tile_X0Y1_N4END[8]
port 596 nsew signal input
rlabel metal2 s 13174 -40 13230 160 6 Tile_X0Y1_N4END[9]
port 597 nsew signal input
rlabel metal2 s 15106 -40 15162 160 6 Tile_X0Y1_NN4END[0]
port 598 nsew signal input
rlabel metal2 s 17866 -40 17922 160 6 Tile_X0Y1_NN4END[10]
port 599 nsew signal input
rlabel metal2 s 18142 -40 18198 160 6 Tile_X0Y1_NN4END[11]
port 600 nsew signal input
rlabel metal2 s 18418 -40 18474 160 6 Tile_X0Y1_NN4END[12]
port 601 nsew signal input
rlabel metal2 s 18694 -40 18750 160 6 Tile_X0Y1_NN4END[13]
port 602 nsew signal input
rlabel metal2 s 18970 -40 19026 160 6 Tile_X0Y1_NN4END[14]
port 603 nsew signal input
rlabel metal2 s 19246 -40 19302 160 6 Tile_X0Y1_NN4END[15]
port 604 nsew signal input
rlabel metal2 s 15382 -40 15438 160 6 Tile_X0Y1_NN4END[1]
port 605 nsew signal input
rlabel metal2 s 15658 -40 15714 160 6 Tile_X0Y1_NN4END[2]
port 606 nsew signal input
rlabel metal2 s 15934 -40 15990 160 6 Tile_X0Y1_NN4END[3]
port 607 nsew signal input
rlabel metal2 s 16210 -40 16266 160 6 Tile_X0Y1_NN4END[4]
port 608 nsew signal input
rlabel metal2 s 16486 -40 16542 160 6 Tile_X0Y1_NN4END[5]
port 609 nsew signal input
rlabel metal2 s 16762 -40 16818 160 6 Tile_X0Y1_NN4END[6]
port 610 nsew signal input
rlabel metal2 s 17038 -40 17094 160 6 Tile_X0Y1_NN4END[7]
port 611 nsew signal input
rlabel metal2 s 17314 -40 17370 160 6 Tile_X0Y1_NN4END[8]
port 612 nsew signal input
rlabel metal2 s 17590 -40 17646 160 6 Tile_X0Y1_NN4END[9]
port 613 nsew signal input
rlabel metal2 s 19522 -40 19578 160 6 Tile_X0Y1_S1BEG[0]
port 614 nsew signal output
rlabel metal2 s 19798 -40 19854 160 6 Tile_X0Y1_S1BEG[1]
port 615 nsew signal output
rlabel metal2 s 20074 -40 20130 160 6 Tile_X0Y1_S1BEG[2]
port 616 nsew signal output
rlabel metal2 s 20350 -40 20406 160 6 Tile_X0Y1_S1BEG[3]
port 617 nsew signal output
rlabel metal2 s 22834 -40 22890 160 6 Tile_X0Y1_S2BEG[0]
port 618 nsew signal output
rlabel metal2 s 23110 -40 23166 160 6 Tile_X0Y1_S2BEG[1]
port 619 nsew signal output
rlabel metal2 s 23386 -40 23442 160 6 Tile_X0Y1_S2BEG[2]
port 620 nsew signal output
rlabel metal2 s 23662 -40 23718 160 6 Tile_X0Y1_S2BEG[3]
port 621 nsew signal output
rlabel metal2 s 23938 -40 23994 160 6 Tile_X0Y1_S2BEG[4]
port 622 nsew signal output
rlabel metal2 s 24214 -40 24270 160 6 Tile_X0Y1_S2BEG[5]
port 623 nsew signal output
rlabel metal2 s 24490 -40 24546 160 6 Tile_X0Y1_S2BEG[6]
port 624 nsew signal output
rlabel metal2 s 24766 -40 24822 160 6 Tile_X0Y1_S2BEG[7]
port 625 nsew signal output
rlabel metal2 s 20626 -40 20682 160 6 Tile_X0Y1_S2BEGb[0]
port 626 nsew signal output
rlabel metal2 s 20902 -40 20958 160 6 Tile_X0Y1_S2BEGb[1]
port 627 nsew signal output
rlabel metal2 s 21178 -40 21234 160 6 Tile_X0Y1_S2BEGb[2]
port 628 nsew signal output
rlabel metal2 s 21454 -40 21510 160 6 Tile_X0Y1_S2BEGb[3]
port 629 nsew signal output
rlabel metal2 s 21730 -40 21786 160 6 Tile_X0Y1_S2BEGb[4]
port 630 nsew signal output
rlabel metal2 s 22006 -40 22062 160 6 Tile_X0Y1_S2BEGb[5]
port 631 nsew signal output
rlabel metal2 s 22282 -40 22338 160 6 Tile_X0Y1_S2BEGb[6]
port 632 nsew signal output
rlabel metal2 s 22558 -40 22614 160 6 Tile_X0Y1_S2BEGb[7]
port 633 nsew signal output
rlabel metal2 s 25042 -40 25098 160 6 Tile_X0Y1_S4BEG[0]
port 634 nsew signal output
rlabel metal2 s 27802 -40 27858 160 6 Tile_X0Y1_S4BEG[10]
port 635 nsew signal output
rlabel metal2 s 28078 -40 28134 160 6 Tile_X0Y1_S4BEG[11]
port 636 nsew signal output
rlabel metal2 s 28354 -40 28410 160 6 Tile_X0Y1_S4BEG[12]
port 637 nsew signal output
rlabel metal2 s 28630 -40 28686 160 6 Tile_X0Y1_S4BEG[13]
port 638 nsew signal output
rlabel metal2 s 28906 -40 28962 160 6 Tile_X0Y1_S4BEG[14]
port 639 nsew signal output
rlabel metal2 s 29182 -40 29238 160 6 Tile_X0Y1_S4BEG[15]
port 640 nsew signal output
rlabel metal2 s 25318 -40 25374 160 6 Tile_X0Y1_S4BEG[1]
port 641 nsew signal output
rlabel metal2 s 25594 -40 25650 160 6 Tile_X0Y1_S4BEG[2]
port 642 nsew signal output
rlabel metal2 s 25870 -40 25926 160 6 Tile_X0Y1_S4BEG[3]
port 643 nsew signal output
rlabel metal2 s 26146 -40 26202 160 6 Tile_X0Y1_S4BEG[4]
port 644 nsew signal output
rlabel metal2 s 26422 -40 26478 160 6 Tile_X0Y1_S4BEG[5]
port 645 nsew signal output
rlabel metal2 s 26698 -40 26754 160 6 Tile_X0Y1_S4BEG[6]
port 646 nsew signal output
rlabel metal2 s 26974 -40 27030 160 6 Tile_X0Y1_S4BEG[7]
port 647 nsew signal output
rlabel metal2 s 27250 -40 27306 160 6 Tile_X0Y1_S4BEG[8]
port 648 nsew signal output
rlabel metal2 s 27526 -40 27582 160 6 Tile_X0Y1_S4BEG[9]
port 649 nsew signal output
rlabel metal2 s 29458 -40 29514 160 6 Tile_X0Y1_SS4BEG[0]
port 650 nsew signal output
rlabel metal2 s 32218 -40 32274 160 6 Tile_X0Y1_SS4BEG[10]
port 651 nsew signal output
rlabel metal2 s 32494 -40 32550 160 6 Tile_X0Y1_SS4BEG[11]
port 652 nsew signal output
rlabel metal2 s 32770 -40 32826 160 6 Tile_X0Y1_SS4BEG[12]
port 653 nsew signal output
rlabel metal2 s 33046 -40 33102 160 6 Tile_X0Y1_SS4BEG[13]
port 654 nsew signal output
rlabel metal2 s 33322 -40 33378 160 6 Tile_X0Y1_SS4BEG[14]
port 655 nsew signal output
rlabel metal2 s 33598 -40 33654 160 6 Tile_X0Y1_SS4BEG[15]
port 656 nsew signal output
rlabel metal2 s 29734 -40 29790 160 6 Tile_X0Y1_SS4BEG[1]
port 657 nsew signal output
rlabel metal2 s 30010 -40 30066 160 6 Tile_X0Y1_SS4BEG[2]
port 658 nsew signal output
rlabel metal2 s 30286 -40 30342 160 6 Tile_X0Y1_SS4BEG[3]
port 659 nsew signal output
rlabel metal2 s 30562 -40 30618 160 6 Tile_X0Y1_SS4BEG[4]
port 660 nsew signal output
rlabel metal2 s 30838 -40 30894 160 6 Tile_X0Y1_SS4BEG[5]
port 661 nsew signal output
rlabel metal2 s 31114 -40 31170 160 6 Tile_X0Y1_SS4BEG[6]
port 662 nsew signal output
rlabel metal2 s 31390 -40 31446 160 6 Tile_X0Y1_SS4BEG[7]
port 663 nsew signal output
rlabel metal2 s 31666 -40 31722 160 6 Tile_X0Y1_SS4BEG[8]
port 664 nsew signal output
rlabel metal2 s 31942 -40 31998 160 6 Tile_X0Y1_SS4BEG[9]
port 665 nsew signal output
rlabel metal2 s 33874 -40 33930 160 6 Tile_X0Y1_UserCLK
port 666 nsew signal input
rlabel metal3 s -40 4904 160 5024 6 Tile_X0Y1_W1BEG[0]
port 667 nsew signal output
rlabel metal3 s -40 5176 160 5296 6 Tile_X0Y1_W1BEG[1]
port 668 nsew signal output
rlabel metal3 s -40 5448 160 5568 6 Tile_X0Y1_W1BEG[2]
port 669 nsew signal output
rlabel metal3 s -40 5720 160 5840 6 Tile_X0Y1_W1BEG[3]
port 670 nsew signal output
rlabel metal3 s 44540 4904 44740 5024 6 Tile_X0Y1_W1END[0]
port 671 nsew signal input
rlabel metal3 s 44540 5176 44740 5296 6 Tile_X0Y1_W1END[1]
port 672 nsew signal input
rlabel metal3 s 44540 5448 44740 5568 6 Tile_X0Y1_W1END[2]
port 673 nsew signal input
rlabel metal3 s 44540 5720 44740 5840 6 Tile_X0Y1_W1END[3]
port 674 nsew signal input
rlabel metal3 s -40 5992 160 6112 6 Tile_X0Y1_W2BEG[0]
port 675 nsew signal output
rlabel metal3 s -40 6264 160 6384 6 Tile_X0Y1_W2BEG[1]
port 676 nsew signal output
rlabel metal3 s -40 6536 160 6656 6 Tile_X0Y1_W2BEG[2]
port 677 nsew signal output
rlabel metal3 s -40 6808 160 6928 6 Tile_X0Y1_W2BEG[3]
port 678 nsew signal output
rlabel metal3 s -40 7080 160 7200 6 Tile_X0Y1_W2BEG[4]
port 679 nsew signal output
rlabel metal3 s -40 7352 160 7472 6 Tile_X0Y1_W2BEG[5]
port 680 nsew signal output
rlabel metal3 s -40 7624 160 7744 6 Tile_X0Y1_W2BEG[6]
port 681 nsew signal output
rlabel metal3 s -40 7896 160 8016 6 Tile_X0Y1_W2BEG[7]
port 682 nsew signal output
rlabel metal3 s -40 8168 160 8288 6 Tile_X0Y1_W2BEGb[0]
port 683 nsew signal output
rlabel metal3 s -40 8440 160 8560 6 Tile_X0Y1_W2BEGb[1]
port 684 nsew signal output
rlabel metal3 s -40 8712 160 8832 6 Tile_X0Y1_W2BEGb[2]
port 685 nsew signal output
rlabel metal3 s -40 8984 160 9104 6 Tile_X0Y1_W2BEGb[3]
port 686 nsew signal output
rlabel metal3 s -40 9256 160 9376 6 Tile_X0Y1_W2BEGb[4]
port 687 nsew signal output
rlabel metal3 s -40 9528 160 9648 6 Tile_X0Y1_W2BEGb[5]
port 688 nsew signal output
rlabel metal3 s -40 9800 160 9920 6 Tile_X0Y1_W2BEGb[6]
port 689 nsew signal output
rlabel metal3 s -40 10072 160 10192 6 Tile_X0Y1_W2BEGb[7]
port 690 nsew signal output
rlabel metal3 s 44540 8168 44740 8288 6 Tile_X0Y1_W2END[0]
port 691 nsew signal input
rlabel metal3 s 44540 8440 44740 8560 6 Tile_X0Y1_W2END[1]
port 692 nsew signal input
rlabel metal3 s 44540 8712 44740 8832 6 Tile_X0Y1_W2END[2]
port 693 nsew signal input
rlabel metal3 s 44540 8984 44740 9104 6 Tile_X0Y1_W2END[3]
port 694 nsew signal input
rlabel metal3 s 44540 9256 44740 9376 6 Tile_X0Y1_W2END[4]
port 695 nsew signal input
rlabel metal3 s 44540 9528 44740 9648 6 Tile_X0Y1_W2END[5]
port 696 nsew signal input
rlabel metal3 s 44540 9800 44740 9920 6 Tile_X0Y1_W2END[6]
port 697 nsew signal input
rlabel metal3 s 44540 10072 44740 10192 6 Tile_X0Y1_W2END[7]
port 698 nsew signal input
rlabel metal3 s 44540 5992 44740 6112 6 Tile_X0Y1_W2MID[0]
port 699 nsew signal input
rlabel metal3 s 44540 6264 44740 6384 6 Tile_X0Y1_W2MID[1]
port 700 nsew signal input
rlabel metal3 s 44540 6536 44740 6656 6 Tile_X0Y1_W2MID[2]
port 701 nsew signal input
rlabel metal3 s 44540 6808 44740 6928 6 Tile_X0Y1_W2MID[3]
port 702 nsew signal input
rlabel metal3 s 44540 7080 44740 7200 6 Tile_X0Y1_W2MID[4]
port 703 nsew signal input
rlabel metal3 s 44540 7352 44740 7472 6 Tile_X0Y1_W2MID[5]
port 704 nsew signal input
rlabel metal3 s 44540 7624 44740 7744 6 Tile_X0Y1_W2MID[6]
port 705 nsew signal input
rlabel metal3 s 44540 7896 44740 8016 6 Tile_X0Y1_W2MID[7]
port 706 nsew signal input
rlabel metal3 s -40 14696 160 14816 6 Tile_X0Y1_W6BEG[0]
port 707 nsew signal output
rlabel metal3 s -40 17416 160 17536 6 Tile_X0Y1_W6BEG[10]
port 708 nsew signal output
rlabel metal3 s -40 17688 160 17808 6 Tile_X0Y1_W6BEG[11]
port 709 nsew signal output
rlabel metal3 s -40 14968 160 15088 6 Tile_X0Y1_W6BEG[1]
port 710 nsew signal output
rlabel metal3 s -40 15240 160 15360 6 Tile_X0Y1_W6BEG[2]
port 711 nsew signal output
rlabel metal3 s -40 15512 160 15632 6 Tile_X0Y1_W6BEG[3]
port 712 nsew signal output
rlabel metal3 s -40 15784 160 15904 6 Tile_X0Y1_W6BEG[4]
port 713 nsew signal output
rlabel metal3 s -40 16056 160 16176 6 Tile_X0Y1_W6BEG[5]
port 714 nsew signal output
rlabel metal3 s -40 16328 160 16448 6 Tile_X0Y1_W6BEG[6]
port 715 nsew signal output
rlabel metal3 s -40 16600 160 16720 6 Tile_X0Y1_W6BEG[7]
port 716 nsew signal output
rlabel metal3 s -40 16872 160 16992 6 Tile_X0Y1_W6BEG[8]
port 717 nsew signal output
rlabel metal3 s -40 17144 160 17264 6 Tile_X0Y1_W6BEG[9]
port 718 nsew signal output
rlabel metal3 s 44540 14696 44740 14816 6 Tile_X0Y1_W6END[0]
port 719 nsew signal input
rlabel metal3 s 44540 17416 44740 17536 6 Tile_X0Y1_W6END[10]
port 720 nsew signal input
rlabel metal3 s 44540 17688 44740 17808 6 Tile_X0Y1_W6END[11]
port 721 nsew signal input
rlabel metal3 s 44540 14968 44740 15088 6 Tile_X0Y1_W6END[1]
port 722 nsew signal input
rlabel metal3 s 44540 15240 44740 15360 6 Tile_X0Y1_W6END[2]
port 723 nsew signal input
rlabel metal3 s 44540 15512 44740 15632 6 Tile_X0Y1_W6END[3]
port 724 nsew signal input
rlabel metal3 s 44540 15784 44740 15904 6 Tile_X0Y1_W6END[4]
port 725 nsew signal input
rlabel metal3 s 44540 16056 44740 16176 6 Tile_X0Y1_W6END[5]
port 726 nsew signal input
rlabel metal3 s 44540 16328 44740 16448 6 Tile_X0Y1_W6END[6]
port 727 nsew signal input
rlabel metal3 s 44540 16600 44740 16720 6 Tile_X0Y1_W6END[7]
port 728 nsew signal input
rlabel metal3 s 44540 16872 44740 16992 6 Tile_X0Y1_W6END[8]
port 729 nsew signal input
rlabel metal3 s 44540 17144 44740 17264 6 Tile_X0Y1_W6END[9]
port 730 nsew signal input
rlabel metal3 s -40 10344 160 10464 6 Tile_X0Y1_WW4BEG[0]
port 731 nsew signal output
rlabel metal3 s -40 13064 160 13184 6 Tile_X0Y1_WW4BEG[10]
port 732 nsew signal output
rlabel metal3 s -40 13336 160 13456 6 Tile_X0Y1_WW4BEG[11]
port 733 nsew signal output
rlabel metal3 s -40 13608 160 13728 6 Tile_X0Y1_WW4BEG[12]
port 734 nsew signal output
rlabel metal3 s -40 13880 160 14000 6 Tile_X0Y1_WW4BEG[13]
port 735 nsew signal output
rlabel metal3 s -40 14152 160 14272 6 Tile_X0Y1_WW4BEG[14]
port 736 nsew signal output
rlabel metal3 s -40 14424 160 14544 6 Tile_X0Y1_WW4BEG[15]
port 737 nsew signal output
rlabel metal3 s -40 10616 160 10736 6 Tile_X0Y1_WW4BEG[1]
port 738 nsew signal output
rlabel metal3 s -40 10888 160 11008 6 Tile_X0Y1_WW4BEG[2]
port 739 nsew signal output
rlabel metal3 s -40 11160 160 11280 6 Tile_X0Y1_WW4BEG[3]
port 740 nsew signal output
rlabel metal3 s -40 11432 160 11552 6 Tile_X0Y1_WW4BEG[4]
port 741 nsew signal output
rlabel metal3 s -40 11704 160 11824 6 Tile_X0Y1_WW4BEG[5]
port 742 nsew signal output
rlabel metal3 s -40 11976 160 12096 6 Tile_X0Y1_WW4BEG[6]
port 743 nsew signal output
rlabel metal3 s -40 12248 160 12368 6 Tile_X0Y1_WW4BEG[7]
port 744 nsew signal output
rlabel metal3 s -40 12520 160 12640 6 Tile_X0Y1_WW4BEG[8]
port 745 nsew signal output
rlabel metal3 s -40 12792 160 12912 6 Tile_X0Y1_WW4BEG[9]
port 746 nsew signal output
rlabel metal3 s 44540 10344 44740 10464 6 Tile_X0Y1_WW4END[0]
port 747 nsew signal input
rlabel metal3 s 44540 13064 44740 13184 6 Tile_X0Y1_WW4END[10]
port 748 nsew signal input
rlabel metal3 s 44540 13336 44740 13456 6 Tile_X0Y1_WW4END[11]
port 749 nsew signal input
rlabel metal3 s 44540 13608 44740 13728 6 Tile_X0Y1_WW4END[12]
port 750 nsew signal input
rlabel metal3 s 44540 13880 44740 14000 6 Tile_X0Y1_WW4END[13]
port 751 nsew signal input
rlabel metal3 s 44540 14152 44740 14272 6 Tile_X0Y1_WW4END[14]
port 752 nsew signal input
rlabel metal3 s 44540 14424 44740 14544 6 Tile_X0Y1_WW4END[15]
port 753 nsew signal input
rlabel metal3 s 44540 10616 44740 10736 6 Tile_X0Y1_WW4END[1]
port 754 nsew signal input
rlabel metal3 s 44540 10888 44740 11008 6 Tile_X0Y1_WW4END[2]
port 755 nsew signal input
rlabel metal3 s 44540 11160 44740 11280 6 Tile_X0Y1_WW4END[3]
port 756 nsew signal input
rlabel metal3 s 44540 11432 44740 11552 6 Tile_X0Y1_WW4END[4]
port 757 nsew signal input
rlabel metal3 s 44540 11704 44740 11824 6 Tile_X0Y1_WW4END[5]
port 758 nsew signal input
rlabel metal3 s 44540 11976 44740 12096 6 Tile_X0Y1_WW4END[6]
port 759 nsew signal input
rlabel metal3 s 44540 12248 44740 12368 6 Tile_X0Y1_WW4END[7]
port 760 nsew signal input
rlabel metal3 s 44540 12520 44740 12640 6 Tile_X0Y1_WW4END[8]
port 761 nsew signal input
rlabel metal3 s 44540 12792 44740 12912 6 Tile_X0Y1_WW4END[9]
port 762 nsew signal input
rlabel metal4 s 19568 1040 19888 88720 6 VGND
port 763 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 88720 6 VPWR
port 764 nsew power bidirectional
rlabel metal4 s 34928 1040 35248 88720 6 VPWR
port 764 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 44700 90000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 14339710
string GDS_FILE /home/asma/Desktop/open_eFPGA_v2/openlane/DSP/runs/24_12_09_16_26/results/signoff/DSP.magic.gds
string GDS_START 1095822
<< end >>

