magic
tech sky130A
magscale 1 2
timestamp 1733616470
<< obsli1 >>
rect 1104 1071 14536 43537
<< obsm1 >>
rect 474 1040 15700 43568
<< metal2 >>
rect 478 44540 534 45000
rect 1214 44540 1270 45000
rect 1950 44540 2006 45000
rect 2686 44540 2742 45000
rect 3422 44540 3478 45000
rect 4158 44540 4214 45000
rect 4894 44540 4950 45000
rect 5630 44540 5686 45000
rect 6366 44540 6422 45000
rect 7102 44540 7158 45000
rect 7838 44540 7894 45000
rect 8574 44540 8630 45000
rect 9310 44540 9366 45000
rect 10046 44540 10102 45000
rect 10782 44540 10838 45000
rect 11518 44540 11574 45000
rect 12254 44540 12310 45000
rect 12990 44540 13046 45000
rect 13726 44540 13782 45000
rect 14462 44540 14518 45000
rect 15198 44540 15254 45000
rect 478 -300 534 160
rect 1214 -300 1270 160
rect 1950 -300 2006 160
rect 2686 -300 2742 160
rect 3422 -300 3478 160
rect 4158 -300 4214 160
rect 4894 -300 4950 160
rect 5630 -300 5686 160
rect 6366 -300 6422 160
rect 7102 -300 7158 160
rect 7838 -300 7894 160
rect 8574 -300 8630 160
rect 9310 -300 9366 160
rect 10046 -300 10102 160
rect 10782 -300 10838 160
rect 11518 -300 11574 160
rect 12254 -300 12310 160
rect 12990 -300 13046 160
rect 13726 -300 13782 160
rect 14462 -300 14518 160
rect 15198 -300 15254 160
<< obsm2 >>
rect 590 44484 1158 44540
rect 1326 44484 1894 44540
rect 2062 44484 2630 44540
rect 2798 44484 3366 44540
rect 3534 44484 4102 44540
rect 4270 44484 4838 44540
rect 5006 44484 5574 44540
rect 5742 44484 6310 44540
rect 6478 44484 7046 44540
rect 7214 44484 7782 44540
rect 7950 44484 8518 44540
rect 8686 44484 9254 44540
rect 9422 44484 9990 44540
rect 10158 44484 10726 44540
rect 10894 44484 11462 44540
rect 11630 44484 12198 44540
rect 12366 44484 12934 44540
rect 13102 44484 13670 44540
rect 13838 44484 14406 44540
rect 14574 44484 15142 44540
rect 15310 44484 15700 44540
rect 480 216 15700 44484
rect 590 54 1158 216
rect 1326 54 1894 216
rect 2062 54 2630 216
rect 2798 54 3366 216
rect 3534 54 4102 216
rect 4270 54 4838 216
rect 5006 54 5574 216
rect 5742 54 6310 216
rect 6478 54 7046 216
rect 7214 54 7782 216
rect 7950 54 8518 216
rect 8686 54 9254 216
rect 9422 54 9990 216
rect 10158 54 10726 216
rect 10894 54 11462 216
rect 11630 54 12198 216
rect 12366 54 12934 216
rect 13102 54 13670 216
rect 13838 54 14406 216
rect 14574 54 15142 216
rect 15310 54 15700 216
<< metal3 >>
rect -300 40536 160 40656
rect -300 39720 160 39840
rect 15540 39448 16000 39568
rect 15540 39176 16000 39296
rect -300 38904 160 39024
rect 15540 38904 16000 39024
rect 15540 38632 16000 38752
rect 15540 38360 16000 38480
rect -300 38088 160 38208
rect 15540 38088 16000 38208
rect 15540 37816 16000 37936
rect 15540 37544 16000 37664
rect -300 37272 160 37392
rect 15540 37272 16000 37392
rect 15540 37000 16000 37120
rect 15540 36728 16000 36848
rect -300 36456 160 36576
rect 15540 36456 16000 36576
rect 15540 36184 16000 36304
rect 15540 35912 16000 36032
rect -300 35640 160 35760
rect 15540 35640 16000 35760
rect 15540 35368 16000 35488
rect 15540 35096 16000 35216
rect -300 34824 160 34944
rect 15540 34824 16000 34944
rect 15540 34552 16000 34672
rect 15540 34280 16000 34400
rect -300 34008 160 34128
rect 15540 34008 16000 34128
rect 15540 33736 16000 33856
rect 15540 33464 16000 33584
rect -300 33192 160 33312
rect 15540 33192 16000 33312
rect 15540 32920 16000 33040
rect 15540 32648 16000 32768
rect -300 32376 160 32496
rect 15540 32376 16000 32496
rect 15540 32104 16000 32224
rect 15540 31832 16000 31952
rect -300 31560 160 31680
rect 15540 31560 16000 31680
rect 15540 31288 16000 31408
rect 15540 31016 16000 31136
rect -300 30744 160 30864
rect 15540 30744 16000 30864
rect 15540 30472 16000 30592
rect 15540 30200 16000 30320
rect -300 29928 160 30048
rect 15540 29928 16000 30048
rect 15540 29656 16000 29776
rect 15540 29384 16000 29504
rect -300 29112 160 29232
rect 15540 29112 16000 29232
rect 15540 28840 16000 28960
rect 15540 28568 16000 28688
rect -300 28296 160 28416
rect 15540 28296 16000 28416
rect 15540 28024 16000 28144
rect 15540 27752 16000 27872
rect -300 27480 160 27600
rect 15540 27480 16000 27600
rect 15540 27208 16000 27328
rect 15540 26936 16000 27056
rect -300 26664 160 26784
rect 15540 26664 16000 26784
rect 15540 26392 16000 26512
rect 15540 26120 16000 26240
rect -300 25848 160 25968
rect 15540 25848 16000 25968
rect 15540 25576 16000 25696
rect 15540 25304 16000 25424
rect -300 25032 160 25152
rect 15540 25032 16000 25152
rect 15540 24760 16000 24880
rect 15540 24488 16000 24608
rect -300 24216 160 24336
rect 15540 24216 16000 24336
rect 15540 23944 16000 24064
rect 15540 23672 16000 23792
rect -300 23400 160 23520
rect 15540 23400 16000 23520
rect 15540 23128 16000 23248
rect 15540 22856 16000 22976
rect -300 22584 160 22704
rect 15540 22584 16000 22704
rect 15540 22312 16000 22432
rect 15540 22040 16000 22160
rect -300 21768 160 21888
rect 15540 21768 16000 21888
rect 15540 21496 16000 21616
rect 15540 21224 16000 21344
rect -300 20952 160 21072
rect 15540 20952 16000 21072
rect 15540 20680 16000 20800
rect 15540 20408 16000 20528
rect -300 20136 160 20256
rect 15540 20136 16000 20256
rect 15540 19864 16000 19984
rect 15540 19592 16000 19712
rect -300 19320 160 19440
rect 15540 19320 16000 19440
rect 15540 19048 16000 19168
rect 15540 18776 16000 18896
rect -300 18504 160 18624
rect 15540 18504 16000 18624
rect 15540 18232 16000 18352
rect 15540 17960 16000 18080
rect -300 17688 160 17808
rect 15540 17688 16000 17808
rect 15540 17416 16000 17536
rect 15540 17144 16000 17264
rect -300 16872 160 16992
rect 15540 16872 16000 16992
rect 15540 16600 16000 16720
rect 15540 16328 16000 16448
rect -300 16056 160 16176
rect 15540 16056 16000 16176
rect 15540 15784 16000 15904
rect 15540 15512 16000 15632
rect -300 15240 160 15360
rect 15540 15240 16000 15360
rect 15540 14968 16000 15088
rect 15540 14696 16000 14816
rect -300 14424 160 14544
rect 15540 14424 16000 14544
rect 15540 14152 16000 14272
rect 15540 13880 16000 14000
rect -300 13608 160 13728
rect 15540 13608 16000 13728
rect 15540 13336 16000 13456
rect 15540 13064 16000 13184
rect -300 12792 160 12912
rect 15540 12792 16000 12912
rect 15540 12520 16000 12640
rect 15540 12248 16000 12368
rect -300 11976 160 12096
rect 15540 11976 16000 12096
rect 15540 11704 16000 11824
rect 15540 11432 16000 11552
rect -300 11160 160 11280
rect 15540 11160 16000 11280
rect 15540 10888 16000 11008
rect 15540 10616 16000 10736
rect -300 10344 160 10464
rect 15540 10344 16000 10464
rect 15540 10072 16000 10192
rect 15540 9800 16000 9920
rect -300 9528 160 9648
rect 15540 9528 16000 9648
rect 15540 9256 16000 9376
rect 15540 8984 16000 9104
rect -300 8712 160 8832
rect 15540 8712 16000 8832
rect 15540 8440 16000 8560
rect 15540 8168 16000 8288
rect -300 7896 160 8016
rect 15540 7896 16000 8016
rect 15540 7624 16000 7744
rect 15540 7352 16000 7472
rect -300 7080 160 7200
rect 15540 7080 16000 7200
rect 15540 6808 16000 6928
rect 15540 6536 16000 6656
rect -300 6264 160 6384
rect 15540 6264 16000 6384
rect 15540 5992 16000 6112
rect 15540 5720 16000 5840
rect -300 5448 160 5568
rect 15540 5448 16000 5568
rect 15540 5176 16000 5296
rect 15540 4904 16000 5024
rect -300 4632 160 4752
rect -300 3816 160 3936
<< obsm3 >>
rect 160 40736 15540 43553
rect 240 40456 15540 40736
rect 160 39920 15540 40456
rect 240 39648 15540 39920
rect 240 39640 15460 39648
rect 160 39104 15460 39640
rect 240 38824 15460 39104
rect 160 38288 15460 38824
rect 240 38008 15460 38288
rect 160 37472 15460 38008
rect 240 37192 15460 37472
rect 160 36656 15460 37192
rect 240 36376 15460 36656
rect 160 35840 15460 36376
rect 240 35560 15460 35840
rect 160 35024 15460 35560
rect 240 34744 15460 35024
rect 160 34208 15460 34744
rect 240 33928 15460 34208
rect 160 33392 15460 33928
rect 240 33112 15460 33392
rect 160 32576 15460 33112
rect 240 32296 15460 32576
rect 160 31760 15460 32296
rect 240 31480 15460 31760
rect 160 30944 15460 31480
rect 240 30664 15460 30944
rect 160 30128 15460 30664
rect 240 29848 15460 30128
rect 160 29312 15460 29848
rect 240 29032 15460 29312
rect 160 28496 15460 29032
rect 240 28216 15460 28496
rect 160 27680 15460 28216
rect 240 27400 15460 27680
rect 160 26864 15460 27400
rect 240 26584 15460 26864
rect 160 26048 15460 26584
rect 240 25768 15460 26048
rect 160 25232 15460 25768
rect 240 24952 15460 25232
rect 160 24416 15460 24952
rect 240 24136 15460 24416
rect 160 23600 15460 24136
rect 240 23320 15460 23600
rect 160 22784 15460 23320
rect 240 22504 15460 22784
rect 160 21968 15460 22504
rect 240 21688 15460 21968
rect 160 21152 15460 21688
rect 240 20872 15460 21152
rect 160 20336 15460 20872
rect 240 20056 15460 20336
rect 160 19520 15460 20056
rect 240 19240 15460 19520
rect 160 18704 15460 19240
rect 240 18424 15460 18704
rect 160 17888 15460 18424
rect 240 17608 15460 17888
rect 160 17072 15460 17608
rect 240 16792 15460 17072
rect 160 16256 15460 16792
rect 240 15976 15460 16256
rect 160 15440 15460 15976
rect 240 15160 15460 15440
rect 160 14624 15460 15160
rect 240 14344 15460 14624
rect 160 13808 15460 14344
rect 240 13528 15460 13808
rect 160 12992 15460 13528
rect 240 12712 15460 12992
rect 160 12176 15460 12712
rect 240 11896 15460 12176
rect 160 11360 15460 11896
rect 240 11080 15460 11360
rect 160 10544 15460 11080
rect 240 10264 15460 10544
rect 160 9728 15460 10264
rect 240 9448 15460 9728
rect 160 8912 15460 9448
rect 240 8632 15460 8912
rect 160 8096 15460 8632
rect 240 7816 15460 8096
rect 160 7280 15460 7816
rect 240 7000 15460 7280
rect 160 6464 15460 7000
rect 240 6184 15460 6464
rect 160 5648 15460 6184
rect 240 5368 15460 5648
rect 160 4832 15460 5368
rect 240 4824 15460 4832
rect 240 4552 15540 4824
rect 160 4016 15540 4552
rect 240 3736 15540 4016
rect 160 1055 15540 3736
<< metal4 >>
rect 2623 1040 2943 43568
rect 4302 1040 4622 43568
rect 5981 1040 6301 43568
rect 7660 1040 7980 43568
rect 9339 1040 9659 43568
rect 11018 1040 11338 43568
rect 12697 1040 13017 43568
rect 14376 1040 14696 43568
<< obsm4 >>
rect 1531 1259 2543 42805
rect 3023 1259 4222 42805
rect 4702 1259 5901 42805
rect 6381 1259 7580 42805
rect 8060 1259 9259 42805
rect 9739 1259 10938 42805
rect 11418 1259 12617 42805
rect 13097 1259 14296 42805
rect 14776 1259 15397 42805
<< labels >>
rlabel metal3 s -300 11160 160 11280 4 A_I_top
port 1 nsew signal output
rlabel metal3 s -300 9528 160 9648 4 A_O_top
port 2 nsew signal input
rlabel metal3 s -300 10344 160 10464 4 A_T_top
port 3 nsew signal output
rlabel metal3 s -300 11976 160 12096 4 A_config_C_bit0
port 4 nsew signal output
rlabel metal3 s -300 12792 160 12912 4 A_config_C_bit1
port 5 nsew signal output
rlabel metal3 s -300 13608 160 13728 4 A_config_C_bit2
port 6 nsew signal output
rlabel metal3 s -300 14424 160 14544 4 A_config_C_bit3
port 7 nsew signal output
rlabel metal3 s -300 5448 160 5568 4 B_I_top
port 8 nsew signal output
rlabel metal3 s -300 3816 160 3936 4 B_O_top
port 9 nsew signal input
rlabel metal3 s -300 4632 160 4752 4 B_T_top
port 10 nsew signal output
rlabel metal3 s -300 6264 160 6384 4 B_config_C_bit0
port 11 nsew signal output
rlabel metal3 s -300 7080 160 7200 4 B_config_C_bit1
port 12 nsew signal output
rlabel metal3 s -300 7896 160 8016 4 B_config_C_bit2
port 13 nsew signal output
rlabel metal3 s -300 8712 160 8832 4 B_config_C_bit3
port 14 nsew signal output
rlabel metal3 s 15540 17960 16000 18080 6 E1BEG[0]
port 15 nsew signal output
rlabel metal3 s 15540 18232 16000 18352 6 E1BEG[1]
port 16 nsew signal output
rlabel metal3 s 15540 18504 16000 18624 6 E1BEG[2]
port 17 nsew signal output
rlabel metal3 s 15540 18776 16000 18896 6 E1BEG[3]
port 18 nsew signal output
rlabel metal3 s 15540 19048 16000 19168 6 E2BEG[0]
port 19 nsew signal output
rlabel metal3 s 15540 19320 16000 19440 6 E2BEG[1]
port 20 nsew signal output
rlabel metal3 s 15540 19592 16000 19712 6 E2BEG[2]
port 21 nsew signal output
rlabel metal3 s 15540 19864 16000 19984 6 E2BEG[3]
port 22 nsew signal output
rlabel metal3 s 15540 20136 16000 20256 6 E2BEG[4]
port 23 nsew signal output
rlabel metal3 s 15540 20408 16000 20528 6 E2BEG[5]
port 24 nsew signal output
rlabel metal3 s 15540 20680 16000 20800 6 E2BEG[6]
port 25 nsew signal output
rlabel metal3 s 15540 20952 16000 21072 6 E2BEG[7]
port 26 nsew signal output
rlabel metal3 s 15540 21224 16000 21344 6 E2BEGb[0]
port 27 nsew signal output
rlabel metal3 s 15540 21496 16000 21616 6 E2BEGb[1]
port 28 nsew signal output
rlabel metal3 s 15540 21768 16000 21888 6 E2BEGb[2]
port 29 nsew signal output
rlabel metal3 s 15540 22040 16000 22160 6 E2BEGb[3]
port 30 nsew signal output
rlabel metal3 s 15540 22312 16000 22432 6 E2BEGb[4]
port 31 nsew signal output
rlabel metal3 s 15540 22584 16000 22704 6 E2BEGb[5]
port 32 nsew signal output
rlabel metal3 s 15540 22856 16000 22976 6 E2BEGb[6]
port 33 nsew signal output
rlabel metal3 s 15540 23128 16000 23248 6 E2BEGb[7]
port 34 nsew signal output
rlabel metal3 s 15540 27752 16000 27872 6 E6BEG[0]
port 35 nsew signal output
rlabel metal3 s 15540 30472 16000 30592 6 E6BEG[10]
port 36 nsew signal output
rlabel metal3 s 15540 30744 16000 30864 6 E6BEG[11]
port 37 nsew signal output
rlabel metal3 s 15540 28024 16000 28144 6 E6BEG[1]
port 38 nsew signal output
rlabel metal3 s 15540 28296 16000 28416 6 E6BEG[2]
port 39 nsew signal output
rlabel metal3 s 15540 28568 16000 28688 6 E6BEG[3]
port 40 nsew signal output
rlabel metal3 s 15540 28840 16000 28960 6 E6BEG[4]
port 41 nsew signal output
rlabel metal3 s 15540 29112 16000 29232 6 E6BEG[5]
port 42 nsew signal output
rlabel metal3 s 15540 29384 16000 29504 6 E6BEG[6]
port 43 nsew signal output
rlabel metal3 s 15540 29656 16000 29776 6 E6BEG[7]
port 44 nsew signal output
rlabel metal3 s 15540 29928 16000 30048 6 E6BEG[8]
port 45 nsew signal output
rlabel metal3 s 15540 30200 16000 30320 6 E6BEG[9]
port 46 nsew signal output
rlabel metal3 s 15540 23400 16000 23520 6 EE4BEG[0]
port 47 nsew signal output
rlabel metal3 s 15540 26120 16000 26240 6 EE4BEG[10]
port 48 nsew signal output
rlabel metal3 s 15540 26392 16000 26512 6 EE4BEG[11]
port 49 nsew signal output
rlabel metal3 s 15540 26664 16000 26784 6 EE4BEG[12]
port 50 nsew signal output
rlabel metal3 s 15540 26936 16000 27056 6 EE4BEG[13]
port 51 nsew signal output
rlabel metal3 s 15540 27208 16000 27328 6 EE4BEG[14]
port 52 nsew signal output
rlabel metal3 s 15540 27480 16000 27600 6 EE4BEG[15]
port 53 nsew signal output
rlabel metal3 s 15540 23672 16000 23792 6 EE4BEG[1]
port 54 nsew signal output
rlabel metal3 s 15540 23944 16000 24064 6 EE4BEG[2]
port 55 nsew signal output
rlabel metal3 s 15540 24216 16000 24336 6 EE4BEG[3]
port 56 nsew signal output
rlabel metal3 s 15540 24488 16000 24608 6 EE4BEG[4]
port 57 nsew signal output
rlabel metal3 s 15540 24760 16000 24880 6 EE4BEG[5]
port 58 nsew signal output
rlabel metal3 s 15540 25032 16000 25152 6 EE4BEG[6]
port 59 nsew signal output
rlabel metal3 s 15540 25304 16000 25424 6 EE4BEG[7]
port 60 nsew signal output
rlabel metal3 s 15540 25576 16000 25696 6 EE4BEG[8]
port 61 nsew signal output
rlabel metal3 s 15540 25848 16000 25968 6 EE4BEG[9]
port 62 nsew signal output
rlabel metal3 s -300 15240 160 15360 4 FrameData[0]
port 63 nsew signal input
rlabel metal3 s -300 23400 160 23520 4 FrameData[10]
port 64 nsew signal input
rlabel metal3 s -300 24216 160 24336 4 FrameData[11]
port 65 nsew signal input
rlabel metal3 s -300 25032 160 25152 4 FrameData[12]
port 66 nsew signal input
rlabel metal3 s -300 25848 160 25968 4 FrameData[13]
port 67 nsew signal input
rlabel metal3 s -300 26664 160 26784 4 FrameData[14]
port 68 nsew signal input
rlabel metal3 s -300 27480 160 27600 4 FrameData[15]
port 69 nsew signal input
rlabel metal3 s -300 28296 160 28416 4 FrameData[16]
port 70 nsew signal input
rlabel metal3 s -300 29112 160 29232 4 FrameData[17]
port 71 nsew signal input
rlabel metal3 s -300 29928 160 30048 4 FrameData[18]
port 72 nsew signal input
rlabel metal3 s -300 30744 160 30864 4 FrameData[19]
port 73 nsew signal input
rlabel metal3 s -300 16056 160 16176 4 FrameData[1]
port 74 nsew signal input
rlabel metal3 s -300 31560 160 31680 4 FrameData[20]
port 75 nsew signal input
rlabel metal3 s -300 32376 160 32496 4 FrameData[21]
port 76 nsew signal input
rlabel metal3 s -300 33192 160 33312 4 FrameData[22]
port 77 nsew signal input
rlabel metal3 s -300 34008 160 34128 4 FrameData[23]
port 78 nsew signal input
rlabel metal3 s -300 34824 160 34944 4 FrameData[24]
port 79 nsew signal input
rlabel metal3 s -300 35640 160 35760 4 FrameData[25]
port 80 nsew signal input
rlabel metal3 s -300 36456 160 36576 4 FrameData[26]
port 81 nsew signal input
rlabel metal3 s -300 37272 160 37392 4 FrameData[27]
port 82 nsew signal input
rlabel metal3 s -300 38088 160 38208 4 FrameData[28]
port 83 nsew signal input
rlabel metal3 s -300 38904 160 39024 4 FrameData[29]
port 84 nsew signal input
rlabel metal3 s -300 16872 160 16992 4 FrameData[2]
port 85 nsew signal input
rlabel metal3 s -300 39720 160 39840 4 FrameData[30]
port 86 nsew signal input
rlabel metal3 s -300 40536 160 40656 4 FrameData[31]
port 87 nsew signal input
rlabel metal3 s -300 17688 160 17808 4 FrameData[3]
port 88 nsew signal input
rlabel metal3 s -300 18504 160 18624 4 FrameData[4]
port 89 nsew signal input
rlabel metal3 s -300 19320 160 19440 4 FrameData[5]
port 90 nsew signal input
rlabel metal3 s -300 20136 160 20256 4 FrameData[6]
port 91 nsew signal input
rlabel metal3 s -300 20952 160 21072 4 FrameData[7]
port 92 nsew signal input
rlabel metal3 s -300 21768 160 21888 4 FrameData[8]
port 93 nsew signal input
rlabel metal3 s -300 22584 160 22704 4 FrameData[9]
port 94 nsew signal input
rlabel metal3 s 15540 31016 16000 31136 6 FrameData_O[0]
port 95 nsew signal output
rlabel metal3 s 15540 33736 16000 33856 6 FrameData_O[10]
port 96 nsew signal output
rlabel metal3 s 15540 34008 16000 34128 6 FrameData_O[11]
port 97 nsew signal output
rlabel metal3 s 15540 34280 16000 34400 6 FrameData_O[12]
port 98 nsew signal output
rlabel metal3 s 15540 34552 16000 34672 6 FrameData_O[13]
port 99 nsew signal output
rlabel metal3 s 15540 34824 16000 34944 6 FrameData_O[14]
port 100 nsew signal output
rlabel metal3 s 15540 35096 16000 35216 6 FrameData_O[15]
port 101 nsew signal output
rlabel metal3 s 15540 35368 16000 35488 6 FrameData_O[16]
port 102 nsew signal output
rlabel metal3 s 15540 35640 16000 35760 6 FrameData_O[17]
port 103 nsew signal output
rlabel metal3 s 15540 35912 16000 36032 6 FrameData_O[18]
port 104 nsew signal output
rlabel metal3 s 15540 36184 16000 36304 6 FrameData_O[19]
port 105 nsew signal output
rlabel metal3 s 15540 31288 16000 31408 6 FrameData_O[1]
port 106 nsew signal output
rlabel metal3 s 15540 36456 16000 36576 6 FrameData_O[20]
port 107 nsew signal output
rlabel metal3 s 15540 36728 16000 36848 6 FrameData_O[21]
port 108 nsew signal output
rlabel metal3 s 15540 37000 16000 37120 6 FrameData_O[22]
port 109 nsew signal output
rlabel metal3 s 15540 37272 16000 37392 6 FrameData_O[23]
port 110 nsew signal output
rlabel metal3 s 15540 37544 16000 37664 6 FrameData_O[24]
port 111 nsew signal output
rlabel metal3 s 15540 37816 16000 37936 6 FrameData_O[25]
port 112 nsew signal output
rlabel metal3 s 15540 38088 16000 38208 6 FrameData_O[26]
port 113 nsew signal output
rlabel metal3 s 15540 38360 16000 38480 6 FrameData_O[27]
port 114 nsew signal output
rlabel metal3 s 15540 38632 16000 38752 6 FrameData_O[28]
port 115 nsew signal output
rlabel metal3 s 15540 38904 16000 39024 6 FrameData_O[29]
port 116 nsew signal output
rlabel metal3 s 15540 31560 16000 31680 6 FrameData_O[2]
port 117 nsew signal output
rlabel metal3 s 15540 39176 16000 39296 6 FrameData_O[30]
port 118 nsew signal output
rlabel metal3 s 15540 39448 16000 39568 6 FrameData_O[31]
port 119 nsew signal output
rlabel metal3 s 15540 31832 16000 31952 6 FrameData_O[3]
port 120 nsew signal output
rlabel metal3 s 15540 32104 16000 32224 6 FrameData_O[4]
port 121 nsew signal output
rlabel metal3 s 15540 32376 16000 32496 6 FrameData_O[5]
port 122 nsew signal output
rlabel metal3 s 15540 32648 16000 32768 6 FrameData_O[6]
port 123 nsew signal output
rlabel metal3 s 15540 32920 16000 33040 6 FrameData_O[7]
port 124 nsew signal output
rlabel metal3 s 15540 33192 16000 33312 6 FrameData_O[8]
port 125 nsew signal output
rlabel metal3 s 15540 33464 16000 33584 6 FrameData_O[9]
port 126 nsew signal output
rlabel metal2 s 1214 -300 1270 160 8 FrameStrobe[0]
port 127 nsew signal input
rlabel metal2 s 8574 -300 8630 160 8 FrameStrobe[10]
port 128 nsew signal input
rlabel metal2 s 9310 -300 9366 160 8 FrameStrobe[11]
port 129 nsew signal input
rlabel metal2 s 10046 -300 10102 160 8 FrameStrobe[12]
port 130 nsew signal input
rlabel metal2 s 10782 -300 10838 160 8 FrameStrobe[13]
port 131 nsew signal input
rlabel metal2 s 11518 -300 11574 160 8 FrameStrobe[14]
port 132 nsew signal input
rlabel metal2 s 12254 -300 12310 160 8 FrameStrobe[15]
port 133 nsew signal input
rlabel metal2 s 12990 -300 13046 160 8 FrameStrobe[16]
port 134 nsew signal input
rlabel metal2 s 13726 -300 13782 160 8 FrameStrobe[17]
port 135 nsew signal input
rlabel metal2 s 14462 -300 14518 160 8 FrameStrobe[18]
port 136 nsew signal input
rlabel metal2 s 15198 -300 15254 160 8 FrameStrobe[19]
port 137 nsew signal input
rlabel metal2 s 1950 -300 2006 160 8 FrameStrobe[1]
port 138 nsew signal input
rlabel metal2 s 2686 -300 2742 160 8 FrameStrobe[2]
port 139 nsew signal input
rlabel metal2 s 3422 -300 3478 160 8 FrameStrobe[3]
port 140 nsew signal input
rlabel metal2 s 4158 -300 4214 160 8 FrameStrobe[4]
port 141 nsew signal input
rlabel metal2 s 4894 -300 4950 160 8 FrameStrobe[5]
port 142 nsew signal input
rlabel metal2 s 5630 -300 5686 160 8 FrameStrobe[6]
port 143 nsew signal input
rlabel metal2 s 6366 -300 6422 160 8 FrameStrobe[7]
port 144 nsew signal input
rlabel metal2 s 7102 -300 7158 160 8 FrameStrobe[8]
port 145 nsew signal input
rlabel metal2 s 7838 -300 7894 160 8 FrameStrobe[9]
port 146 nsew signal input
rlabel metal2 s 1214 44540 1270 45000 6 FrameStrobe_O[0]
port 147 nsew signal output
rlabel metal2 s 8574 44540 8630 45000 6 FrameStrobe_O[10]
port 148 nsew signal output
rlabel metal2 s 9310 44540 9366 45000 6 FrameStrobe_O[11]
port 149 nsew signal output
rlabel metal2 s 10046 44540 10102 45000 6 FrameStrobe_O[12]
port 150 nsew signal output
rlabel metal2 s 10782 44540 10838 45000 6 FrameStrobe_O[13]
port 151 nsew signal output
rlabel metal2 s 11518 44540 11574 45000 6 FrameStrobe_O[14]
port 152 nsew signal output
rlabel metal2 s 12254 44540 12310 45000 6 FrameStrobe_O[15]
port 153 nsew signal output
rlabel metal2 s 12990 44540 13046 45000 6 FrameStrobe_O[16]
port 154 nsew signal output
rlabel metal2 s 13726 44540 13782 45000 6 FrameStrobe_O[17]
port 155 nsew signal output
rlabel metal2 s 14462 44540 14518 45000 6 FrameStrobe_O[18]
port 156 nsew signal output
rlabel metal2 s 15198 44540 15254 45000 6 FrameStrobe_O[19]
port 157 nsew signal output
rlabel metal2 s 1950 44540 2006 45000 6 FrameStrobe_O[1]
port 158 nsew signal output
rlabel metal2 s 2686 44540 2742 45000 6 FrameStrobe_O[2]
port 159 nsew signal output
rlabel metal2 s 3422 44540 3478 45000 6 FrameStrobe_O[3]
port 160 nsew signal output
rlabel metal2 s 4158 44540 4214 45000 6 FrameStrobe_O[4]
port 161 nsew signal output
rlabel metal2 s 4894 44540 4950 45000 6 FrameStrobe_O[5]
port 162 nsew signal output
rlabel metal2 s 5630 44540 5686 45000 6 FrameStrobe_O[6]
port 163 nsew signal output
rlabel metal2 s 6366 44540 6422 45000 6 FrameStrobe_O[7]
port 164 nsew signal output
rlabel metal2 s 7102 44540 7158 45000 6 FrameStrobe_O[8]
port 165 nsew signal output
rlabel metal2 s 7838 44540 7894 45000 6 FrameStrobe_O[9]
port 166 nsew signal output
rlabel metal2 s 478 -300 534 160 8 UserCLK
port 167 nsew signal input
rlabel metal2 s 478 44540 534 45000 6 UserCLKo
port 168 nsew signal output
rlabel metal4 s 4302 1040 4622 43568 6 VGND
port 169 nsew ground bidirectional
rlabel metal4 s 7660 1040 7980 43568 6 VGND
port 169 nsew ground bidirectional
rlabel metal4 s 11018 1040 11338 43568 6 VGND
port 169 nsew ground bidirectional
rlabel metal4 s 14376 1040 14696 43568 6 VGND
port 169 nsew ground bidirectional
rlabel metal4 s 2623 1040 2943 43568 6 VPWR
port 170 nsew power bidirectional
rlabel metal4 s 5981 1040 6301 43568 6 VPWR
port 170 nsew power bidirectional
rlabel metal4 s 9339 1040 9659 43568 6 VPWR
port 170 nsew power bidirectional
rlabel metal4 s 12697 1040 13017 43568 6 VPWR
port 170 nsew power bidirectional
rlabel metal3 s 15540 4904 16000 5024 6 W1END[0]
port 171 nsew signal input
rlabel metal3 s 15540 5176 16000 5296 6 W1END[1]
port 172 nsew signal input
rlabel metal3 s 15540 5448 16000 5568 6 W1END[2]
port 173 nsew signal input
rlabel metal3 s 15540 5720 16000 5840 6 W1END[3]
port 174 nsew signal input
rlabel metal3 s 15540 8168 16000 8288 6 W2END[0]
port 175 nsew signal input
rlabel metal3 s 15540 8440 16000 8560 6 W2END[1]
port 176 nsew signal input
rlabel metal3 s 15540 8712 16000 8832 6 W2END[2]
port 177 nsew signal input
rlabel metal3 s 15540 8984 16000 9104 6 W2END[3]
port 178 nsew signal input
rlabel metal3 s 15540 9256 16000 9376 6 W2END[4]
port 179 nsew signal input
rlabel metal3 s 15540 9528 16000 9648 6 W2END[5]
port 180 nsew signal input
rlabel metal3 s 15540 9800 16000 9920 6 W2END[6]
port 181 nsew signal input
rlabel metal3 s 15540 10072 16000 10192 6 W2END[7]
port 182 nsew signal input
rlabel metal3 s 15540 5992 16000 6112 6 W2MID[0]
port 183 nsew signal input
rlabel metal3 s 15540 6264 16000 6384 6 W2MID[1]
port 184 nsew signal input
rlabel metal3 s 15540 6536 16000 6656 6 W2MID[2]
port 185 nsew signal input
rlabel metal3 s 15540 6808 16000 6928 6 W2MID[3]
port 186 nsew signal input
rlabel metal3 s 15540 7080 16000 7200 6 W2MID[4]
port 187 nsew signal input
rlabel metal3 s 15540 7352 16000 7472 6 W2MID[5]
port 188 nsew signal input
rlabel metal3 s 15540 7624 16000 7744 6 W2MID[6]
port 189 nsew signal input
rlabel metal3 s 15540 7896 16000 8016 6 W2MID[7]
port 190 nsew signal input
rlabel metal3 s 15540 14696 16000 14816 6 W6END[0]
port 191 nsew signal input
rlabel metal3 s 15540 17416 16000 17536 6 W6END[10]
port 192 nsew signal input
rlabel metal3 s 15540 17688 16000 17808 6 W6END[11]
port 193 nsew signal input
rlabel metal3 s 15540 14968 16000 15088 6 W6END[1]
port 194 nsew signal input
rlabel metal3 s 15540 15240 16000 15360 6 W6END[2]
port 195 nsew signal input
rlabel metal3 s 15540 15512 16000 15632 6 W6END[3]
port 196 nsew signal input
rlabel metal3 s 15540 15784 16000 15904 6 W6END[4]
port 197 nsew signal input
rlabel metal3 s 15540 16056 16000 16176 6 W6END[5]
port 198 nsew signal input
rlabel metal3 s 15540 16328 16000 16448 6 W6END[6]
port 199 nsew signal input
rlabel metal3 s 15540 16600 16000 16720 6 W6END[7]
port 200 nsew signal input
rlabel metal3 s 15540 16872 16000 16992 6 W6END[8]
port 201 nsew signal input
rlabel metal3 s 15540 17144 16000 17264 6 W6END[9]
port 202 nsew signal input
rlabel metal3 s 15540 10344 16000 10464 6 WW4END[0]
port 203 nsew signal input
rlabel metal3 s 15540 13064 16000 13184 6 WW4END[10]
port 204 nsew signal input
rlabel metal3 s 15540 13336 16000 13456 6 WW4END[11]
port 205 nsew signal input
rlabel metal3 s 15540 13608 16000 13728 6 WW4END[12]
port 206 nsew signal input
rlabel metal3 s 15540 13880 16000 14000 6 WW4END[13]
port 207 nsew signal input
rlabel metal3 s 15540 14152 16000 14272 6 WW4END[14]
port 208 nsew signal input
rlabel metal3 s 15540 14424 16000 14544 6 WW4END[15]
port 209 nsew signal input
rlabel metal3 s 15540 10616 16000 10736 6 WW4END[1]
port 210 nsew signal input
rlabel metal3 s 15540 10888 16000 11008 6 WW4END[2]
port 211 nsew signal input
rlabel metal3 s 15540 11160 16000 11280 6 WW4END[3]
port 212 nsew signal input
rlabel metal3 s 15540 11432 16000 11552 6 WW4END[4]
port 213 nsew signal input
rlabel metal3 s 15540 11704 16000 11824 6 WW4END[5]
port 214 nsew signal input
rlabel metal3 s 15540 11976 16000 12096 6 WW4END[6]
port 215 nsew signal input
rlabel metal3 s 15540 12248 16000 12368 6 WW4END[7]
port 216 nsew signal input
rlabel metal3 s 15540 12520 16000 12640 6 WW4END[8]
port 217 nsew signal input
rlabel metal3 s 15540 12792 16000 12912 6 WW4END[9]
port 218 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 15700 44700
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1897612
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/W_IO/runs/24_12_08_00_06/results/signoff/W_IO.magic.gds
string GDS_START 151184
<< end >>

