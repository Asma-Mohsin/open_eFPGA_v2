magic
tech sky130A
magscale 1 2
timestamp 1733608735
<< obsli1 >>
rect 460 1071 44160 43537
<< obsm1 >>
rect 14 212 44698 44600
<< metal2 >>
rect 5078 44540 5134 45000
rect 5354 44540 5410 45000
rect 5630 44540 5686 45000
rect 5906 44540 5962 45000
rect 6182 44540 6238 45000
rect 6458 44540 6514 45000
rect 6734 44540 6790 45000
rect 7010 44540 7066 45000
rect 7286 44540 7342 45000
rect 7562 44540 7618 45000
rect 7838 44540 7894 45000
rect 8114 44540 8170 45000
rect 8390 44540 8446 45000
rect 8666 44540 8722 45000
rect 8942 44540 8998 45000
rect 9218 44540 9274 45000
rect 9494 44540 9550 45000
rect 9770 44540 9826 45000
rect 10046 44540 10102 45000
rect 10322 44540 10378 45000
rect 10598 44540 10654 45000
rect 10874 44540 10930 45000
rect 11150 44540 11206 45000
rect 11426 44540 11482 45000
rect 11702 44540 11758 45000
rect 11978 44540 12034 45000
rect 12254 44540 12310 45000
rect 12530 44540 12586 45000
rect 12806 44540 12862 45000
rect 13082 44540 13138 45000
rect 13358 44540 13414 45000
rect 13634 44540 13690 45000
rect 13910 44540 13966 45000
rect 14186 44540 14242 45000
rect 14462 44540 14518 45000
rect 14738 44540 14794 45000
rect 15014 44540 15070 45000
rect 15290 44540 15346 45000
rect 15566 44540 15622 45000
rect 15842 44540 15898 45000
rect 16118 44540 16174 45000
rect 16394 44540 16450 45000
rect 16670 44540 16726 45000
rect 16946 44540 17002 45000
rect 17222 44540 17278 45000
rect 17498 44540 17554 45000
rect 17774 44540 17830 45000
rect 18050 44540 18106 45000
rect 18326 44540 18382 45000
rect 18602 44540 18658 45000
rect 18878 44540 18934 45000
rect 19154 44540 19210 45000
rect 19430 44540 19486 45000
rect 19706 44540 19762 45000
rect 19982 44540 20038 45000
rect 20258 44540 20314 45000
rect 20534 44540 20590 45000
rect 20810 44540 20866 45000
rect 21086 44540 21142 45000
rect 21362 44540 21418 45000
rect 21638 44540 21694 45000
rect 21914 44540 21970 45000
rect 22190 44540 22246 45000
rect 22466 44540 22522 45000
rect 22742 44540 22798 45000
rect 23018 44540 23074 45000
rect 23294 44540 23350 45000
rect 23570 44540 23626 45000
rect 23846 44540 23902 45000
rect 24122 44540 24178 45000
rect 24398 44540 24454 45000
rect 24674 44540 24730 45000
rect 24950 44540 25006 45000
rect 25226 44540 25282 45000
rect 25502 44540 25558 45000
rect 25778 44540 25834 45000
rect 26054 44540 26110 45000
rect 26330 44540 26386 45000
rect 26606 44540 26662 45000
rect 26882 44540 26938 45000
rect 27158 44540 27214 45000
rect 27434 44540 27490 45000
rect 27710 44540 27766 45000
rect 27986 44540 28042 45000
rect 28262 44540 28318 45000
rect 28538 44540 28594 45000
rect 28814 44540 28870 45000
rect 29090 44540 29146 45000
rect 29366 44540 29422 45000
rect 29642 44540 29698 45000
rect 29918 44540 29974 45000
rect 30194 44540 30250 45000
rect 30470 44540 30526 45000
rect 30746 44540 30802 45000
rect 31022 44540 31078 45000
rect 31298 44540 31354 45000
rect 31574 44540 31630 45000
rect 31850 44540 31906 45000
rect 32126 44540 32182 45000
rect 32402 44540 32458 45000
rect 32678 44540 32734 45000
rect 32954 44540 33010 45000
rect 33230 44540 33286 45000
rect 33506 44540 33562 45000
rect 33782 44540 33838 45000
rect 34058 44540 34114 45000
rect 34334 44540 34390 45000
rect 34610 44540 34666 45000
rect 34886 44540 34942 45000
rect 35162 44540 35218 45000
rect 35438 44540 35494 45000
rect 35714 44540 35770 45000
rect 35990 44540 36046 45000
rect 36266 44540 36322 45000
rect 36542 44540 36598 45000
rect 36818 44540 36874 45000
rect 37094 44540 37150 45000
rect 37370 44540 37426 45000
rect 37646 44540 37702 45000
rect 37922 44540 37978 45000
rect 38198 44540 38254 45000
rect 38474 44540 38530 45000
rect 38750 44540 38806 45000
rect 39026 44540 39082 45000
rect 39302 44540 39358 45000
rect 39578 44540 39634 45000
rect 5078 -300 5134 160
rect 5354 -300 5410 160
rect 5630 -300 5686 160
rect 5906 -300 5962 160
rect 6182 -300 6238 160
rect 6458 -300 6514 160
rect 6734 -300 6790 160
rect 7010 -300 7066 160
rect 7286 -300 7342 160
rect 7562 -300 7618 160
rect 7838 -300 7894 160
rect 8114 -300 8170 160
rect 8390 -300 8446 160
rect 8666 -300 8722 160
rect 8942 -300 8998 160
rect 9218 -300 9274 160
rect 9494 -300 9550 160
rect 9770 -300 9826 160
rect 10046 -300 10102 160
rect 10322 -300 10378 160
rect 10598 -300 10654 160
rect 10874 -300 10930 160
rect 11150 -300 11206 160
rect 11426 -300 11482 160
rect 11702 -300 11758 160
rect 11978 -300 12034 160
rect 12254 -300 12310 160
rect 12530 -300 12586 160
rect 12806 -300 12862 160
rect 13082 -300 13138 160
rect 13358 -300 13414 160
rect 13634 -300 13690 160
rect 13910 -300 13966 160
rect 14186 -300 14242 160
rect 14462 -300 14518 160
rect 14738 -300 14794 160
rect 15014 -300 15070 160
rect 15290 -300 15346 160
rect 15566 -300 15622 160
rect 15842 -300 15898 160
rect 16118 -300 16174 160
rect 16394 -300 16450 160
rect 16670 -300 16726 160
rect 16946 -300 17002 160
rect 17222 -300 17278 160
rect 17498 -300 17554 160
rect 17774 -300 17830 160
rect 18050 -300 18106 160
rect 18326 -300 18382 160
rect 18602 -300 18658 160
rect 18878 -300 18934 160
rect 19154 -300 19210 160
rect 19430 -300 19486 160
rect 19706 -300 19762 160
rect 19982 -300 20038 160
rect 20258 -300 20314 160
rect 20534 -300 20590 160
rect 20810 -300 20866 160
rect 21086 -300 21142 160
rect 21362 -300 21418 160
rect 21638 -300 21694 160
rect 21914 -300 21970 160
rect 22190 -300 22246 160
rect 22466 -300 22522 160
rect 22742 -300 22798 160
rect 23018 -300 23074 160
rect 23294 -300 23350 160
rect 23570 -300 23626 160
rect 23846 -300 23902 160
rect 24122 -300 24178 160
rect 24398 -300 24454 160
rect 24674 -300 24730 160
rect 24950 -300 25006 160
rect 25226 -300 25282 160
rect 25502 -300 25558 160
rect 25778 -300 25834 160
rect 26054 -300 26110 160
rect 26330 -300 26386 160
rect 26606 -300 26662 160
rect 26882 -300 26938 160
rect 27158 -300 27214 160
rect 27434 -300 27490 160
rect 27710 -300 27766 160
rect 27986 -300 28042 160
rect 28262 -300 28318 160
rect 28538 -300 28594 160
rect 28814 -300 28870 160
rect 29090 -300 29146 160
rect 29366 -300 29422 160
rect 29642 -300 29698 160
rect 29918 -300 29974 160
rect 30194 -300 30250 160
rect 30470 -300 30526 160
rect 30746 -300 30802 160
rect 31022 -300 31078 160
rect 31298 -300 31354 160
rect 31574 -300 31630 160
rect 31850 -300 31906 160
rect 32126 -300 32182 160
rect 32402 -300 32458 160
rect 32678 -300 32734 160
rect 32954 -300 33010 160
rect 33230 -300 33286 160
rect 33506 -300 33562 160
rect 33782 -300 33838 160
rect 34058 -300 34114 160
rect 34334 -300 34390 160
rect 34610 -300 34666 160
rect 34886 -300 34942 160
rect 35162 -300 35218 160
rect 35438 -300 35494 160
rect 35714 -300 35770 160
rect 35990 -300 36046 160
rect 36266 -300 36322 160
rect 36542 -300 36598 160
rect 36818 -300 36874 160
rect 37094 -300 37150 160
rect 37370 -300 37426 160
rect 37646 -300 37702 160
rect 37922 -300 37978 160
rect 38198 -300 38254 160
rect 38474 -300 38530 160
rect 38750 -300 38806 160
rect 39026 -300 39082 160
rect 39302 -300 39358 160
rect 39578 -300 39634 160
<< obsm2 >>
rect 20 44484 5022 44606
rect 5190 44484 5298 44606
rect 5466 44484 5574 44606
rect 5742 44484 5850 44606
rect 6018 44484 6126 44606
rect 6294 44484 6402 44606
rect 6570 44484 6678 44606
rect 6846 44484 6954 44606
rect 7122 44484 7230 44606
rect 7398 44484 7506 44606
rect 7674 44484 7782 44606
rect 7950 44484 8058 44606
rect 8226 44484 8334 44606
rect 8502 44484 8610 44606
rect 8778 44484 8886 44606
rect 9054 44484 9162 44606
rect 9330 44484 9438 44606
rect 9606 44484 9714 44606
rect 9882 44484 9990 44606
rect 10158 44484 10266 44606
rect 10434 44484 10542 44606
rect 10710 44484 10818 44606
rect 10986 44484 11094 44606
rect 11262 44484 11370 44606
rect 11538 44484 11646 44606
rect 11814 44484 11922 44606
rect 12090 44484 12198 44606
rect 12366 44484 12474 44606
rect 12642 44484 12750 44606
rect 12918 44484 13026 44606
rect 13194 44484 13302 44606
rect 13470 44484 13578 44606
rect 13746 44484 13854 44606
rect 14022 44484 14130 44606
rect 14298 44484 14406 44606
rect 14574 44484 14682 44606
rect 14850 44484 14958 44606
rect 15126 44484 15234 44606
rect 15402 44484 15510 44606
rect 15678 44484 15786 44606
rect 15954 44484 16062 44606
rect 16230 44484 16338 44606
rect 16506 44484 16614 44606
rect 16782 44484 16890 44606
rect 17058 44484 17166 44606
rect 17334 44484 17442 44606
rect 17610 44484 17718 44606
rect 17886 44484 17994 44606
rect 18162 44484 18270 44606
rect 18438 44484 18546 44606
rect 18714 44484 18822 44606
rect 18990 44484 19098 44606
rect 19266 44484 19374 44606
rect 19542 44484 19650 44606
rect 19818 44484 19926 44606
rect 20094 44484 20202 44606
rect 20370 44484 20478 44606
rect 20646 44484 20754 44606
rect 20922 44484 21030 44606
rect 21198 44484 21306 44606
rect 21474 44484 21582 44606
rect 21750 44484 21858 44606
rect 22026 44484 22134 44606
rect 22302 44484 22410 44606
rect 22578 44484 22686 44606
rect 22854 44484 22962 44606
rect 23130 44484 23238 44606
rect 23406 44484 23514 44606
rect 23682 44484 23790 44606
rect 23958 44484 24066 44606
rect 24234 44484 24342 44606
rect 24510 44484 24618 44606
rect 24786 44484 24894 44606
rect 25062 44484 25170 44606
rect 25338 44484 25446 44606
rect 25614 44484 25722 44606
rect 25890 44484 25998 44606
rect 26166 44484 26274 44606
rect 26442 44484 26550 44606
rect 26718 44484 26826 44606
rect 26994 44484 27102 44606
rect 27270 44484 27378 44606
rect 27546 44484 27654 44606
rect 27822 44484 27930 44606
rect 28098 44484 28206 44606
rect 28374 44484 28482 44606
rect 28650 44484 28758 44606
rect 28926 44484 29034 44606
rect 29202 44484 29310 44606
rect 29478 44484 29586 44606
rect 29754 44484 29862 44606
rect 30030 44484 30138 44606
rect 30306 44484 30414 44606
rect 30582 44484 30690 44606
rect 30858 44484 30966 44606
rect 31134 44484 31242 44606
rect 31410 44484 31518 44606
rect 31686 44484 31794 44606
rect 31962 44484 32070 44606
rect 32238 44484 32346 44606
rect 32514 44484 32622 44606
rect 32790 44484 32898 44606
rect 33066 44484 33174 44606
rect 33342 44484 33450 44606
rect 33618 44484 33726 44606
rect 33894 44484 34002 44606
rect 34170 44484 34278 44606
rect 34446 44484 34554 44606
rect 34722 44484 34830 44606
rect 34998 44484 35106 44606
rect 35274 44484 35382 44606
rect 35550 44484 35658 44606
rect 35826 44484 35934 44606
rect 36102 44484 36210 44606
rect 36378 44484 36486 44606
rect 36654 44484 36762 44606
rect 36930 44484 37038 44606
rect 37206 44484 37314 44606
rect 37482 44484 37590 44606
rect 37758 44484 37866 44606
rect 38034 44484 38142 44606
rect 38310 44484 38418 44606
rect 38586 44484 38694 44606
rect 38862 44484 38970 44606
rect 39138 44484 39246 44606
rect 39414 44484 39522 44606
rect 39690 44484 44692 44606
rect 20 216 44692 44484
rect 20 54 5022 216
rect 5190 54 5298 216
rect 5466 54 5574 216
rect 5742 54 5850 216
rect 6018 54 6126 216
rect 6294 54 6402 216
rect 6570 54 6678 216
rect 6846 54 6954 216
rect 7122 54 7230 216
rect 7398 54 7506 216
rect 7674 54 7782 216
rect 7950 54 8058 216
rect 8226 54 8334 216
rect 8502 54 8610 216
rect 8778 54 8886 216
rect 9054 54 9162 216
rect 9330 54 9438 216
rect 9606 54 9714 216
rect 9882 54 9990 216
rect 10158 54 10266 216
rect 10434 54 10542 216
rect 10710 54 10818 216
rect 10986 54 11094 216
rect 11262 54 11370 216
rect 11538 54 11646 216
rect 11814 54 11922 216
rect 12090 54 12198 216
rect 12366 54 12474 216
rect 12642 54 12750 216
rect 12918 54 13026 216
rect 13194 54 13302 216
rect 13470 54 13578 216
rect 13746 54 13854 216
rect 14022 54 14130 216
rect 14298 54 14406 216
rect 14574 54 14682 216
rect 14850 54 14958 216
rect 15126 54 15234 216
rect 15402 54 15510 216
rect 15678 54 15786 216
rect 15954 54 16062 216
rect 16230 54 16338 216
rect 16506 54 16614 216
rect 16782 54 16890 216
rect 17058 54 17166 216
rect 17334 54 17442 216
rect 17610 54 17718 216
rect 17886 54 17994 216
rect 18162 54 18270 216
rect 18438 54 18546 216
rect 18714 54 18822 216
rect 18990 54 19098 216
rect 19266 54 19374 216
rect 19542 54 19650 216
rect 19818 54 19926 216
rect 20094 54 20202 216
rect 20370 54 20478 216
rect 20646 54 20754 216
rect 20922 54 21030 216
rect 21198 54 21306 216
rect 21474 54 21582 216
rect 21750 54 21858 216
rect 22026 54 22134 216
rect 22302 54 22410 216
rect 22578 54 22686 216
rect 22854 54 22962 216
rect 23130 54 23238 216
rect 23406 54 23514 216
rect 23682 54 23790 216
rect 23958 54 24066 216
rect 24234 54 24342 216
rect 24510 54 24618 216
rect 24786 54 24894 216
rect 25062 54 25170 216
rect 25338 54 25446 216
rect 25614 54 25722 216
rect 25890 54 25998 216
rect 26166 54 26274 216
rect 26442 54 26550 216
rect 26718 54 26826 216
rect 26994 54 27102 216
rect 27270 54 27378 216
rect 27546 54 27654 216
rect 27822 54 27930 216
rect 28098 54 28206 216
rect 28374 54 28482 216
rect 28650 54 28758 216
rect 28926 54 29034 216
rect 29202 54 29310 216
rect 29478 54 29586 216
rect 29754 54 29862 216
rect 30030 54 30138 216
rect 30306 54 30414 216
rect 30582 54 30690 216
rect 30858 54 30966 216
rect 31134 54 31242 216
rect 31410 54 31518 216
rect 31686 54 31794 216
rect 31962 54 32070 216
rect 32238 54 32346 216
rect 32514 54 32622 216
rect 32790 54 32898 216
rect 33066 54 33174 216
rect 33342 54 33450 216
rect 33618 54 33726 216
rect 33894 54 34002 216
rect 34170 54 34278 216
rect 34446 54 34554 216
rect 34722 54 34830 216
rect 34998 54 35106 216
rect 35274 54 35382 216
rect 35550 54 35658 216
rect 35826 54 35934 216
rect 36102 54 36210 216
rect 36378 54 36486 216
rect 36654 54 36762 216
rect 36930 54 37038 216
rect 37206 54 37314 216
rect 37482 54 37590 216
rect 37758 54 37866 216
rect 38034 54 38142 216
rect 38310 54 38418 216
rect 38586 54 38694 216
rect 38862 54 38970 216
rect 39138 54 39246 216
rect 39414 54 39522 216
rect 39690 54 44692 216
<< metal3 >>
rect -300 39448 160 39568
rect -300 39176 160 39296
rect -300 38904 160 39024
rect -300 38632 160 38752
rect -300 38360 160 38480
rect -300 38088 160 38208
rect -300 37816 160 37936
rect -300 37544 160 37664
rect -300 37272 160 37392
rect -300 37000 160 37120
rect -300 36728 160 36848
rect -300 36456 160 36576
rect -300 36184 160 36304
rect -300 35912 160 36032
rect -300 35640 160 35760
rect -300 35368 160 35488
rect -300 35096 160 35216
rect -300 34824 160 34944
rect -300 34552 160 34672
rect -300 34280 160 34400
rect -300 34008 160 34128
rect -300 33736 160 33856
rect -300 33464 160 33584
rect -300 33192 160 33312
rect -300 32920 160 33040
rect -300 32648 160 32768
rect -300 32376 160 32496
rect -300 32104 160 32224
rect -300 31832 160 31952
rect -300 31560 160 31680
rect -300 31288 160 31408
rect -300 31016 160 31136
rect -300 30744 160 30864
rect -300 30472 160 30592
rect -300 30200 160 30320
rect -300 29928 160 30048
rect -300 29656 160 29776
rect -300 29384 160 29504
rect -300 29112 160 29232
rect -300 28840 160 28960
rect -300 28568 160 28688
rect -300 28296 160 28416
rect -300 28024 160 28144
rect -300 27752 160 27872
rect -300 27480 160 27600
rect -300 27208 160 27328
rect -300 26936 160 27056
rect -300 26664 160 26784
rect -300 26392 160 26512
rect -300 26120 160 26240
rect -300 25848 160 25968
rect -300 25576 160 25696
rect -300 25304 160 25424
rect -300 25032 160 25152
rect -300 24760 160 24880
rect -300 24488 160 24608
rect -300 24216 160 24336
rect -300 23944 160 24064
rect -300 23672 160 23792
rect -300 23400 160 23520
rect -300 23128 160 23248
rect -300 22856 160 22976
rect -300 22584 160 22704
rect -300 22312 160 22432
rect -300 22040 160 22160
rect -300 21768 160 21888
rect -300 21496 160 21616
rect -300 21224 160 21344
rect -300 20952 160 21072
rect -300 20680 160 20800
rect -300 20408 160 20528
rect -300 20136 160 20256
rect -300 19864 160 19984
rect -300 19592 160 19712
rect -300 19320 160 19440
rect -300 19048 160 19168
rect -300 18776 160 18896
rect -300 18504 160 18624
rect -300 18232 160 18352
rect -300 17960 160 18080
rect -300 17688 160 17808
rect -300 17416 160 17536
rect -300 17144 160 17264
rect -300 16872 160 16992
rect -300 16600 160 16720
rect -300 16328 160 16448
rect -300 16056 160 16176
rect -300 15784 160 15904
rect -300 15512 160 15632
rect -300 15240 160 15360
rect -300 14968 160 15088
rect -300 14696 160 14816
rect -300 14424 160 14544
rect -300 14152 160 14272
rect -300 13880 160 14000
rect -300 13608 160 13728
rect -300 13336 160 13456
rect -300 13064 160 13184
rect -300 12792 160 12912
rect -300 12520 160 12640
rect -300 12248 160 12368
rect -300 11976 160 12096
rect -300 11704 160 11824
rect -300 11432 160 11552
rect -300 11160 160 11280
rect -300 10888 160 11008
rect -300 10616 160 10736
rect -300 10344 160 10464
rect -300 10072 160 10192
rect -300 9800 160 9920
rect -300 9528 160 9648
rect -300 9256 160 9376
rect -300 8984 160 9104
rect -300 8712 160 8832
rect -300 8440 160 8560
rect -300 8168 160 8288
rect -300 7896 160 8016
rect -300 7624 160 7744
rect -300 7352 160 7472
rect -300 7080 160 7200
rect -300 6808 160 6928
rect -300 6536 160 6656
rect -300 6264 160 6384
rect -300 5992 160 6112
rect -300 5720 160 5840
rect -300 5448 160 5568
rect -300 5176 160 5296
rect -300 4904 160 5024
rect 44540 39448 45000 39568
rect 44540 39176 45000 39296
rect 44540 38904 45000 39024
rect 44540 38632 45000 38752
rect 44540 38360 45000 38480
rect 44540 38088 45000 38208
rect 44540 37816 45000 37936
rect 44540 37544 45000 37664
rect 44540 37272 45000 37392
rect 44540 37000 45000 37120
rect 44540 36728 45000 36848
rect 44540 36456 45000 36576
rect 44540 36184 45000 36304
rect 44540 35912 45000 36032
rect 44540 35640 45000 35760
rect 44540 35368 45000 35488
rect 44540 35096 45000 35216
rect 44540 34824 45000 34944
rect 44540 34552 45000 34672
rect 44540 34280 45000 34400
rect 44540 34008 45000 34128
rect 44540 33736 45000 33856
rect 44540 33464 45000 33584
rect 44540 33192 45000 33312
rect 44540 32920 45000 33040
rect 44540 32648 45000 32768
rect 44540 32376 45000 32496
rect 44540 32104 45000 32224
rect 44540 31832 45000 31952
rect 44540 31560 45000 31680
rect 44540 31288 45000 31408
rect 44540 31016 45000 31136
rect 44540 30744 45000 30864
rect 44540 30472 45000 30592
rect 44540 30200 45000 30320
rect 44540 29928 45000 30048
rect 44540 29656 45000 29776
rect 44540 29384 45000 29504
rect 44540 29112 45000 29232
rect 44540 28840 45000 28960
rect 44540 28568 45000 28688
rect 44540 28296 45000 28416
rect 44540 28024 45000 28144
rect 44540 27752 45000 27872
rect 44540 27480 45000 27600
rect 44540 27208 45000 27328
rect 44540 26936 45000 27056
rect 44540 26664 45000 26784
rect 44540 26392 45000 26512
rect 44540 26120 45000 26240
rect 44540 25848 45000 25968
rect 44540 25576 45000 25696
rect 44540 25304 45000 25424
rect 44540 25032 45000 25152
rect 44540 24760 45000 24880
rect 44540 24488 45000 24608
rect 44540 24216 45000 24336
rect 44540 23944 45000 24064
rect 44540 23672 45000 23792
rect 44540 23400 45000 23520
rect 44540 23128 45000 23248
rect 44540 22856 45000 22976
rect 44540 22584 45000 22704
rect 44540 22312 45000 22432
rect 44540 22040 45000 22160
rect 44540 21768 45000 21888
rect 44540 21496 45000 21616
rect 44540 21224 45000 21344
rect 44540 20952 45000 21072
rect 44540 20680 45000 20800
rect 44540 20408 45000 20528
rect 44540 20136 45000 20256
rect 44540 19864 45000 19984
rect 44540 19592 45000 19712
rect 44540 19320 45000 19440
rect 44540 19048 45000 19168
rect 44540 18776 45000 18896
rect 44540 18504 45000 18624
rect 44540 18232 45000 18352
rect 44540 17960 45000 18080
rect 44540 17688 45000 17808
rect 44540 17416 45000 17536
rect 44540 17144 45000 17264
rect 44540 16872 45000 16992
rect 44540 16600 45000 16720
rect 44540 16328 45000 16448
rect 44540 16056 45000 16176
rect 44540 15784 45000 15904
rect 44540 15512 45000 15632
rect 44540 15240 45000 15360
rect 44540 14968 45000 15088
rect 44540 14696 45000 14816
rect 44540 14424 45000 14544
rect 44540 14152 45000 14272
rect 44540 13880 45000 14000
rect 44540 13608 45000 13728
rect 44540 13336 45000 13456
rect 44540 13064 45000 13184
rect 44540 12792 45000 12912
rect 44540 12520 45000 12640
rect 44540 12248 45000 12368
rect 44540 11976 45000 12096
rect 44540 11704 45000 11824
rect 44540 11432 45000 11552
rect 44540 11160 45000 11280
rect 44540 10888 45000 11008
rect 44540 10616 45000 10736
rect 44540 10344 45000 10464
rect 44540 10072 45000 10192
rect 44540 9800 45000 9920
rect 44540 9528 45000 9648
rect 44540 9256 45000 9376
rect 44540 8984 45000 9104
rect 44540 8712 45000 8832
rect 44540 8440 45000 8560
rect 44540 8168 45000 8288
rect 44540 7896 45000 8016
rect 44540 7624 45000 7744
rect 44540 7352 45000 7472
rect 44540 7080 45000 7200
rect 44540 6808 45000 6928
rect 44540 6536 45000 6656
rect 44540 6264 45000 6384
rect 44540 5992 45000 6112
rect 44540 5720 45000 5840
rect 44540 5448 45000 5568
rect 44540 5176 45000 5296
rect 44540 4904 45000 5024
<< obsm3 >>
rect 160 39648 44607 44437
rect 240 4824 44460 39648
rect 160 36 44607 4824
<< metal4 >>
rect 3564 1040 3884 43568
rect 11064 1040 11384 43568
rect 18564 1040 18884 43568
rect 26064 1040 26384 43568
rect 33564 1040 33884 43568
rect 41064 1040 41384 43568
<< obsm4 >>
rect 243 43648 44101 44437
rect 243 960 3484 43648
rect 3964 960 10984 43648
rect 11464 960 18484 43648
rect 18964 960 25984 43648
rect 26464 960 33484 43648
rect 33964 960 40984 43648
rect 41464 960 44101 43648
rect 243 35 44101 960
<< labels >>
rlabel metal2 s 34058 -300 34114 160 8 Ci
port 1 nsew signal input
rlabel metal2 s 34058 44540 34114 45000 6 Co
port 2 nsew signal output
rlabel metal3 s 44540 17960 45000 18080 6 E1BEG[0]
port 3 nsew signal output
rlabel metal3 s 44540 18232 45000 18352 6 E1BEG[1]
port 4 nsew signal output
rlabel metal3 s 44540 18504 45000 18624 6 E1BEG[2]
port 5 nsew signal output
rlabel metal3 s 44540 18776 45000 18896 6 E1BEG[3]
port 6 nsew signal output
rlabel metal3 s -300 17960 160 18080 4 E1END[0]
port 7 nsew signal input
rlabel metal3 s -300 18232 160 18352 4 E1END[1]
port 8 nsew signal input
rlabel metal3 s -300 18504 160 18624 4 E1END[2]
port 9 nsew signal input
rlabel metal3 s -300 18776 160 18896 4 E1END[3]
port 10 nsew signal input
rlabel metal3 s 44540 19048 45000 19168 6 E2BEG[0]
port 11 nsew signal output
rlabel metal3 s 44540 19320 45000 19440 6 E2BEG[1]
port 12 nsew signal output
rlabel metal3 s 44540 19592 45000 19712 6 E2BEG[2]
port 13 nsew signal output
rlabel metal3 s 44540 19864 45000 19984 6 E2BEG[3]
port 14 nsew signal output
rlabel metal3 s 44540 20136 45000 20256 6 E2BEG[4]
port 15 nsew signal output
rlabel metal3 s 44540 20408 45000 20528 6 E2BEG[5]
port 16 nsew signal output
rlabel metal3 s 44540 20680 45000 20800 6 E2BEG[6]
port 17 nsew signal output
rlabel metal3 s 44540 20952 45000 21072 6 E2BEG[7]
port 18 nsew signal output
rlabel metal3 s 44540 21224 45000 21344 6 E2BEGb[0]
port 19 nsew signal output
rlabel metal3 s 44540 21496 45000 21616 6 E2BEGb[1]
port 20 nsew signal output
rlabel metal3 s 44540 21768 45000 21888 6 E2BEGb[2]
port 21 nsew signal output
rlabel metal3 s 44540 22040 45000 22160 6 E2BEGb[3]
port 22 nsew signal output
rlabel metal3 s 44540 22312 45000 22432 6 E2BEGb[4]
port 23 nsew signal output
rlabel metal3 s 44540 22584 45000 22704 6 E2BEGb[5]
port 24 nsew signal output
rlabel metal3 s 44540 22856 45000 22976 6 E2BEGb[6]
port 25 nsew signal output
rlabel metal3 s 44540 23128 45000 23248 6 E2BEGb[7]
port 26 nsew signal output
rlabel metal3 s -300 21224 160 21344 4 E2END[0]
port 27 nsew signal input
rlabel metal3 s -300 21496 160 21616 4 E2END[1]
port 28 nsew signal input
rlabel metal3 s -300 21768 160 21888 4 E2END[2]
port 29 nsew signal input
rlabel metal3 s -300 22040 160 22160 4 E2END[3]
port 30 nsew signal input
rlabel metal3 s -300 22312 160 22432 4 E2END[4]
port 31 nsew signal input
rlabel metal3 s -300 22584 160 22704 4 E2END[5]
port 32 nsew signal input
rlabel metal3 s -300 22856 160 22976 4 E2END[6]
port 33 nsew signal input
rlabel metal3 s -300 23128 160 23248 4 E2END[7]
port 34 nsew signal input
rlabel metal3 s -300 19048 160 19168 4 E2MID[0]
port 35 nsew signal input
rlabel metal3 s -300 19320 160 19440 4 E2MID[1]
port 36 nsew signal input
rlabel metal3 s -300 19592 160 19712 4 E2MID[2]
port 37 nsew signal input
rlabel metal3 s -300 19864 160 19984 4 E2MID[3]
port 38 nsew signal input
rlabel metal3 s -300 20136 160 20256 4 E2MID[4]
port 39 nsew signal input
rlabel metal3 s -300 20408 160 20528 4 E2MID[5]
port 40 nsew signal input
rlabel metal3 s -300 20680 160 20800 4 E2MID[6]
port 41 nsew signal input
rlabel metal3 s -300 20952 160 21072 4 E2MID[7]
port 42 nsew signal input
rlabel metal3 s 44540 27752 45000 27872 6 E6BEG[0]
port 43 nsew signal output
rlabel metal3 s 44540 30472 45000 30592 6 E6BEG[10]
port 44 nsew signal output
rlabel metal3 s 44540 30744 45000 30864 6 E6BEG[11]
port 45 nsew signal output
rlabel metal3 s 44540 28024 45000 28144 6 E6BEG[1]
port 46 nsew signal output
rlabel metal3 s 44540 28296 45000 28416 6 E6BEG[2]
port 47 nsew signal output
rlabel metal3 s 44540 28568 45000 28688 6 E6BEG[3]
port 48 nsew signal output
rlabel metal3 s 44540 28840 45000 28960 6 E6BEG[4]
port 49 nsew signal output
rlabel metal3 s 44540 29112 45000 29232 6 E6BEG[5]
port 50 nsew signal output
rlabel metal3 s 44540 29384 45000 29504 6 E6BEG[6]
port 51 nsew signal output
rlabel metal3 s 44540 29656 45000 29776 6 E6BEG[7]
port 52 nsew signal output
rlabel metal3 s 44540 29928 45000 30048 6 E6BEG[8]
port 53 nsew signal output
rlabel metal3 s 44540 30200 45000 30320 6 E6BEG[9]
port 54 nsew signal output
rlabel metal3 s -300 27752 160 27872 4 E6END[0]
port 55 nsew signal input
rlabel metal3 s -300 30472 160 30592 4 E6END[10]
port 56 nsew signal input
rlabel metal3 s -300 30744 160 30864 4 E6END[11]
port 57 nsew signal input
rlabel metal3 s -300 28024 160 28144 4 E6END[1]
port 58 nsew signal input
rlabel metal3 s -300 28296 160 28416 4 E6END[2]
port 59 nsew signal input
rlabel metal3 s -300 28568 160 28688 4 E6END[3]
port 60 nsew signal input
rlabel metal3 s -300 28840 160 28960 4 E6END[4]
port 61 nsew signal input
rlabel metal3 s -300 29112 160 29232 4 E6END[5]
port 62 nsew signal input
rlabel metal3 s -300 29384 160 29504 4 E6END[6]
port 63 nsew signal input
rlabel metal3 s -300 29656 160 29776 4 E6END[7]
port 64 nsew signal input
rlabel metal3 s -300 29928 160 30048 4 E6END[8]
port 65 nsew signal input
rlabel metal3 s -300 30200 160 30320 4 E6END[9]
port 66 nsew signal input
rlabel metal3 s 44540 23400 45000 23520 6 EE4BEG[0]
port 67 nsew signal output
rlabel metal3 s 44540 26120 45000 26240 6 EE4BEG[10]
port 68 nsew signal output
rlabel metal3 s 44540 26392 45000 26512 6 EE4BEG[11]
port 69 nsew signal output
rlabel metal3 s 44540 26664 45000 26784 6 EE4BEG[12]
port 70 nsew signal output
rlabel metal3 s 44540 26936 45000 27056 6 EE4BEG[13]
port 71 nsew signal output
rlabel metal3 s 44540 27208 45000 27328 6 EE4BEG[14]
port 72 nsew signal output
rlabel metal3 s 44540 27480 45000 27600 6 EE4BEG[15]
port 73 nsew signal output
rlabel metal3 s 44540 23672 45000 23792 6 EE4BEG[1]
port 74 nsew signal output
rlabel metal3 s 44540 23944 45000 24064 6 EE4BEG[2]
port 75 nsew signal output
rlabel metal3 s 44540 24216 45000 24336 6 EE4BEG[3]
port 76 nsew signal output
rlabel metal3 s 44540 24488 45000 24608 6 EE4BEG[4]
port 77 nsew signal output
rlabel metal3 s 44540 24760 45000 24880 6 EE4BEG[5]
port 78 nsew signal output
rlabel metal3 s 44540 25032 45000 25152 6 EE4BEG[6]
port 79 nsew signal output
rlabel metal3 s 44540 25304 45000 25424 6 EE4BEG[7]
port 80 nsew signal output
rlabel metal3 s 44540 25576 45000 25696 6 EE4BEG[8]
port 81 nsew signal output
rlabel metal3 s 44540 25848 45000 25968 6 EE4BEG[9]
port 82 nsew signal output
rlabel metal3 s -300 23400 160 23520 4 EE4END[0]
port 83 nsew signal input
rlabel metal3 s -300 26120 160 26240 4 EE4END[10]
port 84 nsew signal input
rlabel metal3 s -300 26392 160 26512 4 EE4END[11]
port 85 nsew signal input
rlabel metal3 s -300 26664 160 26784 4 EE4END[12]
port 86 nsew signal input
rlabel metal3 s -300 26936 160 27056 4 EE4END[13]
port 87 nsew signal input
rlabel metal3 s -300 27208 160 27328 4 EE4END[14]
port 88 nsew signal input
rlabel metal3 s -300 27480 160 27600 4 EE4END[15]
port 89 nsew signal input
rlabel metal3 s -300 23672 160 23792 4 EE4END[1]
port 90 nsew signal input
rlabel metal3 s -300 23944 160 24064 4 EE4END[2]
port 91 nsew signal input
rlabel metal3 s -300 24216 160 24336 4 EE4END[3]
port 92 nsew signal input
rlabel metal3 s -300 24488 160 24608 4 EE4END[4]
port 93 nsew signal input
rlabel metal3 s -300 24760 160 24880 4 EE4END[5]
port 94 nsew signal input
rlabel metal3 s -300 25032 160 25152 4 EE4END[6]
port 95 nsew signal input
rlabel metal3 s -300 25304 160 25424 4 EE4END[7]
port 96 nsew signal input
rlabel metal3 s -300 25576 160 25696 4 EE4END[8]
port 97 nsew signal input
rlabel metal3 s -300 25848 160 25968 4 EE4END[9]
port 98 nsew signal input
rlabel metal3 s -300 31016 160 31136 4 FrameData[0]
port 99 nsew signal input
rlabel metal3 s -300 33736 160 33856 4 FrameData[10]
port 100 nsew signal input
rlabel metal3 s -300 34008 160 34128 4 FrameData[11]
port 101 nsew signal input
rlabel metal3 s -300 34280 160 34400 4 FrameData[12]
port 102 nsew signal input
rlabel metal3 s -300 34552 160 34672 4 FrameData[13]
port 103 nsew signal input
rlabel metal3 s -300 34824 160 34944 4 FrameData[14]
port 104 nsew signal input
rlabel metal3 s -300 35096 160 35216 4 FrameData[15]
port 105 nsew signal input
rlabel metal3 s -300 35368 160 35488 4 FrameData[16]
port 106 nsew signal input
rlabel metal3 s -300 35640 160 35760 4 FrameData[17]
port 107 nsew signal input
rlabel metal3 s -300 35912 160 36032 4 FrameData[18]
port 108 nsew signal input
rlabel metal3 s -300 36184 160 36304 4 FrameData[19]
port 109 nsew signal input
rlabel metal3 s -300 31288 160 31408 4 FrameData[1]
port 110 nsew signal input
rlabel metal3 s -300 36456 160 36576 4 FrameData[20]
port 111 nsew signal input
rlabel metal3 s -300 36728 160 36848 4 FrameData[21]
port 112 nsew signal input
rlabel metal3 s -300 37000 160 37120 4 FrameData[22]
port 113 nsew signal input
rlabel metal3 s -300 37272 160 37392 4 FrameData[23]
port 114 nsew signal input
rlabel metal3 s -300 37544 160 37664 4 FrameData[24]
port 115 nsew signal input
rlabel metal3 s -300 37816 160 37936 4 FrameData[25]
port 116 nsew signal input
rlabel metal3 s -300 38088 160 38208 4 FrameData[26]
port 117 nsew signal input
rlabel metal3 s -300 38360 160 38480 4 FrameData[27]
port 118 nsew signal input
rlabel metal3 s -300 38632 160 38752 4 FrameData[28]
port 119 nsew signal input
rlabel metal3 s -300 38904 160 39024 4 FrameData[29]
port 120 nsew signal input
rlabel metal3 s -300 31560 160 31680 4 FrameData[2]
port 121 nsew signal input
rlabel metal3 s -300 39176 160 39296 4 FrameData[30]
port 122 nsew signal input
rlabel metal3 s -300 39448 160 39568 4 FrameData[31]
port 123 nsew signal input
rlabel metal3 s -300 31832 160 31952 4 FrameData[3]
port 124 nsew signal input
rlabel metal3 s -300 32104 160 32224 4 FrameData[4]
port 125 nsew signal input
rlabel metal3 s -300 32376 160 32496 4 FrameData[5]
port 126 nsew signal input
rlabel metal3 s -300 32648 160 32768 4 FrameData[6]
port 127 nsew signal input
rlabel metal3 s -300 32920 160 33040 4 FrameData[7]
port 128 nsew signal input
rlabel metal3 s -300 33192 160 33312 4 FrameData[8]
port 129 nsew signal input
rlabel metal3 s -300 33464 160 33584 4 FrameData[9]
port 130 nsew signal input
rlabel metal3 s 44540 31016 45000 31136 6 FrameData_O[0]
port 131 nsew signal output
rlabel metal3 s 44540 33736 45000 33856 6 FrameData_O[10]
port 132 nsew signal output
rlabel metal3 s 44540 34008 45000 34128 6 FrameData_O[11]
port 133 nsew signal output
rlabel metal3 s 44540 34280 45000 34400 6 FrameData_O[12]
port 134 nsew signal output
rlabel metal3 s 44540 34552 45000 34672 6 FrameData_O[13]
port 135 nsew signal output
rlabel metal3 s 44540 34824 45000 34944 6 FrameData_O[14]
port 136 nsew signal output
rlabel metal3 s 44540 35096 45000 35216 6 FrameData_O[15]
port 137 nsew signal output
rlabel metal3 s 44540 35368 45000 35488 6 FrameData_O[16]
port 138 nsew signal output
rlabel metal3 s 44540 35640 45000 35760 6 FrameData_O[17]
port 139 nsew signal output
rlabel metal3 s 44540 35912 45000 36032 6 FrameData_O[18]
port 140 nsew signal output
rlabel metal3 s 44540 36184 45000 36304 6 FrameData_O[19]
port 141 nsew signal output
rlabel metal3 s 44540 31288 45000 31408 6 FrameData_O[1]
port 142 nsew signal output
rlabel metal3 s 44540 36456 45000 36576 6 FrameData_O[20]
port 143 nsew signal output
rlabel metal3 s 44540 36728 45000 36848 6 FrameData_O[21]
port 144 nsew signal output
rlabel metal3 s 44540 37000 45000 37120 6 FrameData_O[22]
port 145 nsew signal output
rlabel metal3 s 44540 37272 45000 37392 6 FrameData_O[23]
port 146 nsew signal output
rlabel metal3 s 44540 37544 45000 37664 6 FrameData_O[24]
port 147 nsew signal output
rlabel metal3 s 44540 37816 45000 37936 6 FrameData_O[25]
port 148 nsew signal output
rlabel metal3 s 44540 38088 45000 38208 6 FrameData_O[26]
port 149 nsew signal output
rlabel metal3 s 44540 38360 45000 38480 6 FrameData_O[27]
port 150 nsew signal output
rlabel metal3 s 44540 38632 45000 38752 6 FrameData_O[28]
port 151 nsew signal output
rlabel metal3 s 44540 38904 45000 39024 6 FrameData_O[29]
port 152 nsew signal output
rlabel metal3 s 44540 31560 45000 31680 6 FrameData_O[2]
port 153 nsew signal output
rlabel metal3 s 44540 39176 45000 39296 6 FrameData_O[30]
port 154 nsew signal output
rlabel metal3 s 44540 39448 45000 39568 6 FrameData_O[31]
port 155 nsew signal output
rlabel metal3 s 44540 31832 45000 31952 6 FrameData_O[3]
port 156 nsew signal output
rlabel metal3 s 44540 32104 45000 32224 6 FrameData_O[4]
port 157 nsew signal output
rlabel metal3 s 44540 32376 45000 32496 6 FrameData_O[5]
port 158 nsew signal output
rlabel metal3 s 44540 32648 45000 32768 6 FrameData_O[6]
port 159 nsew signal output
rlabel metal3 s 44540 32920 45000 33040 6 FrameData_O[7]
port 160 nsew signal output
rlabel metal3 s 44540 33192 45000 33312 6 FrameData_O[8]
port 161 nsew signal output
rlabel metal3 s 44540 33464 45000 33584 6 FrameData_O[9]
port 162 nsew signal output
rlabel metal2 s 34334 -300 34390 160 8 FrameStrobe[0]
port 163 nsew signal input
rlabel metal2 s 37094 -300 37150 160 8 FrameStrobe[10]
port 164 nsew signal input
rlabel metal2 s 37370 -300 37426 160 8 FrameStrobe[11]
port 165 nsew signal input
rlabel metal2 s 37646 -300 37702 160 8 FrameStrobe[12]
port 166 nsew signal input
rlabel metal2 s 37922 -300 37978 160 8 FrameStrobe[13]
port 167 nsew signal input
rlabel metal2 s 38198 -300 38254 160 8 FrameStrobe[14]
port 168 nsew signal input
rlabel metal2 s 38474 -300 38530 160 8 FrameStrobe[15]
port 169 nsew signal input
rlabel metal2 s 38750 -300 38806 160 8 FrameStrobe[16]
port 170 nsew signal input
rlabel metal2 s 39026 -300 39082 160 8 FrameStrobe[17]
port 171 nsew signal input
rlabel metal2 s 39302 -300 39358 160 8 FrameStrobe[18]
port 172 nsew signal input
rlabel metal2 s 39578 -300 39634 160 8 FrameStrobe[19]
port 173 nsew signal input
rlabel metal2 s 34610 -300 34666 160 8 FrameStrobe[1]
port 174 nsew signal input
rlabel metal2 s 34886 -300 34942 160 8 FrameStrobe[2]
port 175 nsew signal input
rlabel metal2 s 35162 -300 35218 160 8 FrameStrobe[3]
port 176 nsew signal input
rlabel metal2 s 35438 -300 35494 160 8 FrameStrobe[4]
port 177 nsew signal input
rlabel metal2 s 35714 -300 35770 160 8 FrameStrobe[5]
port 178 nsew signal input
rlabel metal2 s 35990 -300 36046 160 8 FrameStrobe[6]
port 179 nsew signal input
rlabel metal2 s 36266 -300 36322 160 8 FrameStrobe[7]
port 180 nsew signal input
rlabel metal2 s 36542 -300 36598 160 8 FrameStrobe[8]
port 181 nsew signal input
rlabel metal2 s 36818 -300 36874 160 8 FrameStrobe[9]
port 182 nsew signal input
rlabel metal2 s 34334 44540 34390 45000 6 FrameStrobe_O[0]
port 183 nsew signal output
rlabel metal2 s 37094 44540 37150 45000 6 FrameStrobe_O[10]
port 184 nsew signal output
rlabel metal2 s 37370 44540 37426 45000 6 FrameStrobe_O[11]
port 185 nsew signal output
rlabel metal2 s 37646 44540 37702 45000 6 FrameStrobe_O[12]
port 186 nsew signal output
rlabel metal2 s 37922 44540 37978 45000 6 FrameStrobe_O[13]
port 187 nsew signal output
rlabel metal2 s 38198 44540 38254 45000 6 FrameStrobe_O[14]
port 188 nsew signal output
rlabel metal2 s 38474 44540 38530 45000 6 FrameStrobe_O[15]
port 189 nsew signal output
rlabel metal2 s 38750 44540 38806 45000 6 FrameStrobe_O[16]
port 190 nsew signal output
rlabel metal2 s 39026 44540 39082 45000 6 FrameStrobe_O[17]
port 191 nsew signal output
rlabel metal2 s 39302 44540 39358 45000 6 FrameStrobe_O[18]
port 192 nsew signal output
rlabel metal2 s 39578 44540 39634 45000 6 FrameStrobe_O[19]
port 193 nsew signal output
rlabel metal2 s 34610 44540 34666 45000 6 FrameStrobe_O[1]
port 194 nsew signal output
rlabel metal2 s 34886 44540 34942 45000 6 FrameStrobe_O[2]
port 195 nsew signal output
rlabel metal2 s 35162 44540 35218 45000 6 FrameStrobe_O[3]
port 196 nsew signal output
rlabel metal2 s 35438 44540 35494 45000 6 FrameStrobe_O[4]
port 197 nsew signal output
rlabel metal2 s 35714 44540 35770 45000 6 FrameStrobe_O[5]
port 198 nsew signal output
rlabel metal2 s 35990 44540 36046 45000 6 FrameStrobe_O[6]
port 199 nsew signal output
rlabel metal2 s 36266 44540 36322 45000 6 FrameStrobe_O[7]
port 200 nsew signal output
rlabel metal2 s 36542 44540 36598 45000 6 FrameStrobe_O[8]
port 201 nsew signal output
rlabel metal2 s 36818 44540 36874 45000 6 FrameStrobe_O[9]
port 202 nsew signal output
rlabel metal2 s 5078 44540 5134 45000 6 N1BEG[0]
port 203 nsew signal output
rlabel metal2 s 5354 44540 5410 45000 6 N1BEG[1]
port 204 nsew signal output
rlabel metal2 s 5630 44540 5686 45000 6 N1BEG[2]
port 205 nsew signal output
rlabel metal2 s 5906 44540 5962 45000 6 N1BEG[3]
port 206 nsew signal output
rlabel metal2 s 5078 -300 5134 160 8 N1END[0]
port 207 nsew signal input
rlabel metal2 s 5354 -300 5410 160 8 N1END[1]
port 208 nsew signal input
rlabel metal2 s 5630 -300 5686 160 8 N1END[2]
port 209 nsew signal input
rlabel metal2 s 5906 -300 5962 160 8 N1END[3]
port 210 nsew signal input
rlabel metal2 s 6182 44540 6238 45000 6 N2BEG[0]
port 211 nsew signal output
rlabel metal2 s 6458 44540 6514 45000 6 N2BEG[1]
port 212 nsew signal output
rlabel metal2 s 6734 44540 6790 45000 6 N2BEG[2]
port 213 nsew signal output
rlabel metal2 s 7010 44540 7066 45000 6 N2BEG[3]
port 214 nsew signal output
rlabel metal2 s 7286 44540 7342 45000 6 N2BEG[4]
port 215 nsew signal output
rlabel metal2 s 7562 44540 7618 45000 6 N2BEG[5]
port 216 nsew signal output
rlabel metal2 s 7838 44540 7894 45000 6 N2BEG[6]
port 217 nsew signal output
rlabel metal2 s 8114 44540 8170 45000 6 N2BEG[7]
port 218 nsew signal output
rlabel metal2 s 8390 44540 8446 45000 6 N2BEGb[0]
port 219 nsew signal output
rlabel metal2 s 8666 44540 8722 45000 6 N2BEGb[1]
port 220 nsew signal output
rlabel metal2 s 8942 44540 8998 45000 6 N2BEGb[2]
port 221 nsew signal output
rlabel metal2 s 9218 44540 9274 45000 6 N2BEGb[3]
port 222 nsew signal output
rlabel metal2 s 9494 44540 9550 45000 6 N2BEGb[4]
port 223 nsew signal output
rlabel metal2 s 9770 44540 9826 45000 6 N2BEGb[5]
port 224 nsew signal output
rlabel metal2 s 10046 44540 10102 45000 6 N2BEGb[6]
port 225 nsew signal output
rlabel metal2 s 10322 44540 10378 45000 6 N2BEGb[7]
port 226 nsew signal output
rlabel metal2 s 8390 -300 8446 160 8 N2END[0]
port 227 nsew signal input
rlabel metal2 s 8666 -300 8722 160 8 N2END[1]
port 228 nsew signal input
rlabel metal2 s 8942 -300 8998 160 8 N2END[2]
port 229 nsew signal input
rlabel metal2 s 9218 -300 9274 160 8 N2END[3]
port 230 nsew signal input
rlabel metal2 s 9494 -300 9550 160 8 N2END[4]
port 231 nsew signal input
rlabel metal2 s 9770 -300 9826 160 8 N2END[5]
port 232 nsew signal input
rlabel metal2 s 10046 -300 10102 160 8 N2END[6]
port 233 nsew signal input
rlabel metal2 s 10322 -300 10378 160 8 N2END[7]
port 234 nsew signal input
rlabel metal2 s 6182 -300 6238 160 8 N2MID[0]
port 235 nsew signal input
rlabel metal2 s 6458 -300 6514 160 8 N2MID[1]
port 236 nsew signal input
rlabel metal2 s 6734 -300 6790 160 8 N2MID[2]
port 237 nsew signal input
rlabel metal2 s 7010 -300 7066 160 8 N2MID[3]
port 238 nsew signal input
rlabel metal2 s 7286 -300 7342 160 8 N2MID[4]
port 239 nsew signal input
rlabel metal2 s 7562 -300 7618 160 8 N2MID[5]
port 240 nsew signal input
rlabel metal2 s 7838 -300 7894 160 8 N2MID[6]
port 241 nsew signal input
rlabel metal2 s 8114 -300 8170 160 8 N2MID[7]
port 242 nsew signal input
rlabel metal2 s 10598 44540 10654 45000 6 N4BEG[0]
port 243 nsew signal output
rlabel metal2 s 13358 44540 13414 45000 6 N4BEG[10]
port 244 nsew signal output
rlabel metal2 s 13634 44540 13690 45000 6 N4BEG[11]
port 245 nsew signal output
rlabel metal2 s 13910 44540 13966 45000 6 N4BEG[12]
port 246 nsew signal output
rlabel metal2 s 14186 44540 14242 45000 6 N4BEG[13]
port 247 nsew signal output
rlabel metal2 s 14462 44540 14518 45000 6 N4BEG[14]
port 248 nsew signal output
rlabel metal2 s 14738 44540 14794 45000 6 N4BEG[15]
port 249 nsew signal output
rlabel metal2 s 10874 44540 10930 45000 6 N4BEG[1]
port 250 nsew signal output
rlabel metal2 s 11150 44540 11206 45000 6 N4BEG[2]
port 251 nsew signal output
rlabel metal2 s 11426 44540 11482 45000 6 N4BEG[3]
port 252 nsew signal output
rlabel metal2 s 11702 44540 11758 45000 6 N4BEG[4]
port 253 nsew signal output
rlabel metal2 s 11978 44540 12034 45000 6 N4BEG[5]
port 254 nsew signal output
rlabel metal2 s 12254 44540 12310 45000 6 N4BEG[6]
port 255 nsew signal output
rlabel metal2 s 12530 44540 12586 45000 6 N4BEG[7]
port 256 nsew signal output
rlabel metal2 s 12806 44540 12862 45000 6 N4BEG[8]
port 257 nsew signal output
rlabel metal2 s 13082 44540 13138 45000 6 N4BEG[9]
port 258 nsew signal output
rlabel metal2 s 10598 -300 10654 160 8 N4END[0]
port 259 nsew signal input
rlabel metal2 s 13358 -300 13414 160 8 N4END[10]
port 260 nsew signal input
rlabel metal2 s 13634 -300 13690 160 8 N4END[11]
port 261 nsew signal input
rlabel metal2 s 13910 -300 13966 160 8 N4END[12]
port 262 nsew signal input
rlabel metal2 s 14186 -300 14242 160 8 N4END[13]
port 263 nsew signal input
rlabel metal2 s 14462 -300 14518 160 8 N4END[14]
port 264 nsew signal input
rlabel metal2 s 14738 -300 14794 160 8 N4END[15]
port 265 nsew signal input
rlabel metal2 s 10874 -300 10930 160 8 N4END[1]
port 266 nsew signal input
rlabel metal2 s 11150 -300 11206 160 8 N4END[2]
port 267 nsew signal input
rlabel metal2 s 11426 -300 11482 160 8 N4END[3]
port 268 nsew signal input
rlabel metal2 s 11702 -300 11758 160 8 N4END[4]
port 269 nsew signal input
rlabel metal2 s 11978 -300 12034 160 8 N4END[5]
port 270 nsew signal input
rlabel metal2 s 12254 -300 12310 160 8 N4END[6]
port 271 nsew signal input
rlabel metal2 s 12530 -300 12586 160 8 N4END[7]
port 272 nsew signal input
rlabel metal2 s 12806 -300 12862 160 8 N4END[8]
port 273 nsew signal input
rlabel metal2 s 13082 -300 13138 160 8 N4END[9]
port 274 nsew signal input
rlabel metal2 s 15014 44540 15070 45000 6 NN4BEG[0]
port 275 nsew signal output
rlabel metal2 s 17774 44540 17830 45000 6 NN4BEG[10]
port 276 nsew signal output
rlabel metal2 s 18050 44540 18106 45000 6 NN4BEG[11]
port 277 nsew signal output
rlabel metal2 s 18326 44540 18382 45000 6 NN4BEG[12]
port 278 nsew signal output
rlabel metal2 s 18602 44540 18658 45000 6 NN4BEG[13]
port 279 nsew signal output
rlabel metal2 s 18878 44540 18934 45000 6 NN4BEG[14]
port 280 nsew signal output
rlabel metal2 s 19154 44540 19210 45000 6 NN4BEG[15]
port 281 nsew signal output
rlabel metal2 s 15290 44540 15346 45000 6 NN4BEG[1]
port 282 nsew signal output
rlabel metal2 s 15566 44540 15622 45000 6 NN4BEG[2]
port 283 nsew signal output
rlabel metal2 s 15842 44540 15898 45000 6 NN4BEG[3]
port 284 nsew signal output
rlabel metal2 s 16118 44540 16174 45000 6 NN4BEG[4]
port 285 nsew signal output
rlabel metal2 s 16394 44540 16450 45000 6 NN4BEG[5]
port 286 nsew signal output
rlabel metal2 s 16670 44540 16726 45000 6 NN4BEG[6]
port 287 nsew signal output
rlabel metal2 s 16946 44540 17002 45000 6 NN4BEG[7]
port 288 nsew signal output
rlabel metal2 s 17222 44540 17278 45000 6 NN4BEG[8]
port 289 nsew signal output
rlabel metal2 s 17498 44540 17554 45000 6 NN4BEG[9]
port 290 nsew signal output
rlabel metal2 s 15014 -300 15070 160 8 NN4END[0]
port 291 nsew signal input
rlabel metal2 s 17774 -300 17830 160 8 NN4END[10]
port 292 nsew signal input
rlabel metal2 s 18050 -300 18106 160 8 NN4END[11]
port 293 nsew signal input
rlabel metal2 s 18326 -300 18382 160 8 NN4END[12]
port 294 nsew signal input
rlabel metal2 s 18602 -300 18658 160 8 NN4END[13]
port 295 nsew signal input
rlabel metal2 s 18878 -300 18934 160 8 NN4END[14]
port 296 nsew signal input
rlabel metal2 s 19154 -300 19210 160 8 NN4END[15]
port 297 nsew signal input
rlabel metal2 s 15290 -300 15346 160 8 NN4END[1]
port 298 nsew signal input
rlabel metal2 s 15566 -300 15622 160 8 NN4END[2]
port 299 nsew signal input
rlabel metal2 s 15842 -300 15898 160 8 NN4END[3]
port 300 nsew signal input
rlabel metal2 s 16118 -300 16174 160 8 NN4END[4]
port 301 nsew signal input
rlabel metal2 s 16394 -300 16450 160 8 NN4END[5]
port 302 nsew signal input
rlabel metal2 s 16670 -300 16726 160 8 NN4END[6]
port 303 nsew signal input
rlabel metal2 s 16946 -300 17002 160 8 NN4END[7]
port 304 nsew signal input
rlabel metal2 s 17222 -300 17278 160 8 NN4END[8]
port 305 nsew signal input
rlabel metal2 s 17498 -300 17554 160 8 NN4END[9]
port 306 nsew signal input
rlabel metal2 s 19430 -300 19486 160 8 S1BEG[0]
port 307 nsew signal output
rlabel metal2 s 19706 -300 19762 160 8 S1BEG[1]
port 308 nsew signal output
rlabel metal2 s 19982 -300 20038 160 8 S1BEG[2]
port 309 nsew signal output
rlabel metal2 s 20258 -300 20314 160 8 S1BEG[3]
port 310 nsew signal output
rlabel metal2 s 19430 44540 19486 45000 6 S1END[0]
port 311 nsew signal input
rlabel metal2 s 19706 44540 19762 45000 6 S1END[1]
port 312 nsew signal input
rlabel metal2 s 19982 44540 20038 45000 6 S1END[2]
port 313 nsew signal input
rlabel metal2 s 20258 44540 20314 45000 6 S1END[3]
port 314 nsew signal input
rlabel metal2 s 22742 -300 22798 160 8 S2BEG[0]
port 315 nsew signal output
rlabel metal2 s 23018 -300 23074 160 8 S2BEG[1]
port 316 nsew signal output
rlabel metal2 s 23294 -300 23350 160 8 S2BEG[2]
port 317 nsew signal output
rlabel metal2 s 23570 -300 23626 160 8 S2BEG[3]
port 318 nsew signal output
rlabel metal2 s 23846 -300 23902 160 8 S2BEG[4]
port 319 nsew signal output
rlabel metal2 s 24122 -300 24178 160 8 S2BEG[5]
port 320 nsew signal output
rlabel metal2 s 24398 -300 24454 160 8 S2BEG[6]
port 321 nsew signal output
rlabel metal2 s 24674 -300 24730 160 8 S2BEG[7]
port 322 nsew signal output
rlabel metal2 s 20534 -300 20590 160 8 S2BEGb[0]
port 323 nsew signal output
rlabel metal2 s 20810 -300 20866 160 8 S2BEGb[1]
port 324 nsew signal output
rlabel metal2 s 21086 -300 21142 160 8 S2BEGb[2]
port 325 nsew signal output
rlabel metal2 s 21362 -300 21418 160 8 S2BEGb[3]
port 326 nsew signal output
rlabel metal2 s 21638 -300 21694 160 8 S2BEGb[4]
port 327 nsew signal output
rlabel metal2 s 21914 -300 21970 160 8 S2BEGb[5]
port 328 nsew signal output
rlabel metal2 s 22190 -300 22246 160 8 S2BEGb[6]
port 329 nsew signal output
rlabel metal2 s 22466 -300 22522 160 8 S2BEGb[7]
port 330 nsew signal output
rlabel metal2 s 20534 44540 20590 45000 6 S2END[0]
port 331 nsew signal input
rlabel metal2 s 20810 44540 20866 45000 6 S2END[1]
port 332 nsew signal input
rlabel metal2 s 21086 44540 21142 45000 6 S2END[2]
port 333 nsew signal input
rlabel metal2 s 21362 44540 21418 45000 6 S2END[3]
port 334 nsew signal input
rlabel metal2 s 21638 44540 21694 45000 6 S2END[4]
port 335 nsew signal input
rlabel metal2 s 21914 44540 21970 45000 6 S2END[5]
port 336 nsew signal input
rlabel metal2 s 22190 44540 22246 45000 6 S2END[6]
port 337 nsew signal input
rlabel metal2 s 22466 44540 22522 45000 6 S2END[7]
port 338 nsew signal input
rlabel metal2 s 22742 44540 22798 45000 6 S2MID[0]
port 339 nsew signal input
rlabel metal2 s 23018 44540 23074 45000 6 S2MID[1]
port 340 nsew signal input
rlabel metal2 s 23294 44540 23350 45000 6 S2MID[2]
port 341 nsew signal input
rlabel metal2 s 23570 44540 23626 45000 6 S2MID[3]
port 342 nsew signal input
rlabel metal2 s 23846 44540 23902 45000 6 S2MID[4]
port 343 nsew signal input
rlabel metal2 s 24122 44540 24178 45000 6 S2MID[5]
port 344 nsew signal input
rlabel metal2 s 24398 44540 24454 45000 6 S2MID[6]
port 345 nsew signal input
rlabel metal2 s 24674 44540 24730 45000 6 S2MID[7]
port 346 nsew signal input
rlabel metal2 s 24950 -300 25006 160 8 S4BEG[0]
port 347 nsew signal output
rlabel metal2 s 27710 -300 27766 160 8 S4BEG[10]
port 348 nsew signal output
rlabel metal2 s 27986 -300 28042 160 8 S4BEG[11]
port 349 nsew signal output
rlabel metal2 s 28262 -300 28318 160 8 S4BEG[12]
port 350 nsew signal output
rlabel metal2 s 28538 -300 28594 160 8 S4BEG[13]
port 351 nsew signal output
rlabel metal2 s 28814 -300 28870 160 8 S4BEG[14]
port 352 nsew signal output
rlabel metal2 s 29090 -300 29146 160 8 S4BEG[15]
port 353 nsew signal output
rlabel metal2 s 25226 -300 25282 160 8 S4BEG[1]
port 354 nsew signal output
rlabel metal2 s 25502 -300 25558 160 8 S4BEG[2]
port 355 nsew signal output
rlabel metal2 s 25778 -300 25834 160 8 S4BEG[3]
port 356 nsew signal output
rlabel metal2 s 26054 -300 26110 160 8 S4BEG[4]
port 357 nsew signal output
rlabel metal2 s 26330 -300 26386 160 8 S4BEG[5]
port 358 nsew signal output
rlabel metal2 s 26606 -300 26662 160 8 S4BEG[6]
port 359 nsew signal output
rlabel metal2 s 26882 -300 26938 160 8 S4BEG[7]
port 360 nsew signal output
rlabel metal2 s 27158 -300 27214 160 8 S4BEG[8]
port 361 nsew signal output
rlabel metal2 s 27434 -300 27490 160 8 S4BEG[9]
port 362 nsew signal output
rlabel metal2 s 24950 44540 25006 45000 6 S4END[0]
port 363 nsew signal input
rlabel metal2 s 27710 44540 27766 45000 6 S4END[10]
port 364 nsew signal input
rlabel metal2 s 27986 44540 28042 45000 6 S4END[11]
port 365 nsew signal input
rlabel metal2 s 28262 44540 28318 45000 6 S4END[12]
port 366 nsew signal input
rlabel metal2 s 28538 44540 28594 45000 6 S4END[13]
port 367 nsew signal input
rlabel metal2 s 28814 44540 28870 45000 6 S4END[14]
port 368 nsew signal input
rlabel metal2 s 29090 44540 29146 45000 6 S4END[15]
port 369 nsew signal input
rlabel metal2 s 25226 44540 25282 45000 6 S4END[1]
port 370 nsew signal input
rlabel metal2 s 25502 44540 25558 45000 6 S4END[2]
port 371 nsew signal input
rlabel metal2 s 25778 44540 25834 45000 6 S4END[3]
port 372 nsew signal input
rlabel metal2 s 26054 44540 26110 45000 6 S4END[4]
port 373 nsew signal input
rlabel metal2 s 26330 44540 26386 45000 6 S4END[5]
port 374 nsew signal input
rlabel metal2 s 26606 44540 26662 45000 6 S4END[6]
port 375 nsew signal input
rlabel metal2 s 26882 44540 26938 45000 6 S4END[7]
port 376 nsew signal input
rlabel metal2 s 27158 44540 27214 45000 6 S4END[8]
port 377 nsew signal input
rlabel metal2 s 27434 44540 27490 45000 6 S4END[9]
port 378 nsew signal input
rlabel metal2 s 29366 -300 29422 160 8 SS4BEG[0]
port 379 nsew signal output
rlabel metal2 s 32126 -300 32182 160 8 SS4BEG[10]
port 380 nsew signal output
rlabel metal2 s 32402 -300 32458 160 8 SS4BEG[11]
port 381 nsew signal output
rlabel metal2 s 32678 -300 32734 160 8 SS4BEG[12]
port 382 nsew signal output
rlabel metal2 s 32954 -300 33010 160 8 SS4BEG[13]
port 383 nsew signal output
rlabel metal2 s 33230 -300 33286 160 8 SS4BEG[14]
port 384 nsew signal output
rlabel metal2 s 33506 -300 33562 160 8 SS4BEG[15]
port 385 nsew signal output
rlabel metal2 s 29642 -300 29698 160 8 SS4BEG[1]
port 386 nsew signal output
rlabel metal2 s 29918 -300 29974 160 8 SS4BEG[2]
port 387 nsew signal output
rlabel metal2 s 30194 -300 30250 160 8 SS4BEG[3]
port 388 nsew signal output
rlabel metal2 s 30470 -300 30526 160 8 SS4BEG[4]
port 389 nsew signal output
rlabel metal2 s 30746 -300 30802 160 8 SS4BEG[5]
port 390 nsew signal output
rlabel metal2 s 31022 -300 31078 160 8 SS4BEG[6]
port 391 nsew signal output
rlabel metal2 s 31298 -300 31354 160 8 SS4BEG[7]
port 392 nsew signal output
rlabel metal2 s 31574 -300 31630 160 8 SS4BEG[8]
port 393 nsew signal output
rlabel metal2 s 31850 -300 31906 160 8 SS4BEG[9]
port 394 nsew signal output
rlabel metal2 s 29366 44540 29422 45000 6 SS4END[0]
port 395 nsew signal input
rlabel metal2 s 32126 44540 32182 45000 6 SS4END[10]
port 396 nsew signal input
rlabel metal2 s 32402 44540 32458 45000 6 SS4END[11]
port 397 nsew signal input
rlabel metal2 s 32678 44540 32734 45000 6 SS4END[12]
port 398 nsew signal input
rlabel metal2 s 32954 44540 33010 45000 6 SS4END[13]
port 399 nsew signal input
rlabel metal2 s 33230 44540 33286 45000 6 SS4END[14]
port 400 nsew signal input
rlabel metal2 s 33506 44540 33562 45000 6 SS4END[15]
port 401 nsew signal input
rlabel metal2 s 29642 44540 29698 45000 6 SS4END[1]
port 402 nsew signal input
rlabel metal2 s 29918 44540 29974 45000 6 SS4END[2]
port 403 nsew signal input
rlabel metal2 s 30194 44540 30250 45000 6 SS4END[3]
port 404 nsew signal input
rlabel metal2 s 30470 44540 30526 45000 6 SS4END[4]
port 405 nsew signal input
rlabel metal2 s 30746 44540 30802 45000 6 SS4END[5]
port 406 nsew signal input
rlabel metal2 s 31022 44540 31078 45000 6 SS4END[6]
port 407 nsew signal input
rlabel metal2 s 31298 44540 31354 45000 6 SS4END[7]
port 408 nsew signal input
rlabel metal2 s 31574 44540 31630 45000 6 SS4END[8]
port 409 nsew signal input
rlabel metal2 s 31850 44540 31906 45000 6 SS4END[9]
port 410 nsew signal input
rlabel metal2 s 33782 -300 33838 160 8 UserCLK
port 411 nsew signal input
rlabel metal2 s 33782 44540 33838 45000 6 UserCLKo
port 412 nsew signal output
rlabel metal3 s -300 4904 160 5024 4 W1BEG[0]
port 413 nsew signal output
rlabel metal3 s -300 5176 160 5296 4 W1BEG[1]
port 414 nsew signal output
rlabel metal3 s -300 5448 160 5568 4 W1BEG[2]
port 415 nsew signal output
rlabel metal3 s -300 5720 160 5840 4 W1BEG[3]
port 416 nsew signal output
rlabel metal3 s 44540 4904 45000 5024 6 W1END[0]
port 417 nsew signal input
rlabel metal3 s 44540 5176 45000 5296 6 W1END[1]
port 418 nsew signal input
rlabel metal3 s 44540 5448 45000 5568 6 W1END[2]
port 419 nsew signal input
rlabel metal3 s 44540 5720 45000 5840 6 W1END[3]
port 420 nsew signal input
rlabel metal3 s -300 5992 160 6112 4 W2BEG[0]
port 421 nsew signal output
rlabel metal3 s -300 6264 160 6384 4 W2BEG[1]
port 422 nsew signal output
rlabel metal3 s -300 6536 160 6656 4 W2BEG[2]
port 423 nsew signal output
rlabel metal3 s -300 6808 160 6928 4 W2BEG[3]
port 424 nsew signal output
rlabel metal3 s -300 7080 160 7200 4 W2BEG[4]
port 425 nsew signal output
rlabel metal3 s -300 7352 160 7472 4 W2BEG[5]
port 426 nsew signal output
rlabel metal3 s -300 7624 160 7744 4 W2BEG[6]
port 427 nsew signal output
rlabel metal3 s -300 7896 160 8016 4 W2BEG[7]
port 428 nsew signal output
rlabel metal3 s -300 8168 160 8288 4 W2BEGb[0]
port 429 nsew signal output
rlabel metal3 s -300 8440 160 8560 4 W2BEGb[1]
port 430 nsew signal output
rlabel metal3 s -300 8712 160 8832 4 W2BEGb[2]
port 431 nsew signal output
rlabel metal3 s -300 8984 160 9104 4 W2BEGb[3]
port 432 nsew signal output
rlabel metal3 s -300 9256 160 9376 4 W2BEGb[4]
port 433 nsew signal output
rlabel metal3 s -300 9528 160 9648 4 W2BEGb[5]
port 434 nsew signal output
rlabel metal3 s -300 9800 160 9920 4 W2BEGb[6]
port 435 nsew signal output
rlabel metal3 s -300 10072 160 10192 4 W2BEGb[7]
port 436 nsew signal output
rlabel metal3 s 44540 8168 45000 8288 6 W2END[0]
port 437 nsew signal input
rlabel metal3 s 44540 8440 45000 8560 6 W2END[1]
port 438 nsew signal input
rlabel metal3 s 44540 8712 45000 8832 6 W2END[2]
port 439 nsew signal input
rlabel metal3 s 44540 8984 45000 9104 6 W2END[3]
port 440 nsew signal input
rlabel metal3 s 44540 9256 45000 9376 6 W2END[4]
port 441 nsew signal input
rlabel metal3 s 44540 9528 45000 9648 6 W2END[5]
port 442 nsew signal input
rlabel metal3 s 44540 9800 45000 9920 6 W2END[6]
port 443 nsew signal input
rlabel metal3 s 44540 10072 45000 10192 6 W2END[7]
port 444 nsew signal input
rlabel metal3 s 44540 5992 45000 6112 6 W2MID[0]
port 445 nsew signal input
rlabel metal3 s 44540 6264 45000 6384 6 W2MID[1]
port 446 nsew signal input
rlabel metal3 s 44540 6536 45000 6656 6 W2MID[2]
port 447 nsew signal input
rlabel metal3 s 44540 6808 45000 6928 6 W2MID[3]
port 448 nsew signal input
rlabel metal3 s 44540 7080 45000 7200 6 W2MID[4]
port 449 nsew signal input
rlabel metal3 s 44540 7352 45000 7472 6 W2MID[5]
port 450 nsew signal input
rlabel metal3 s 44540 7624 45000 7744 6 W2MID[6]
port 451 nsew signal input
rlabel metal3 s 44540 7896 45000 8016 6 W2MID[7]
port 452 nsew signal input
rlabel metal3 s -300 14696 160 14816 4 W6BEG[0]
port 453 nsew signal output
rlabel metal3 s -300 17416 160 17536 4 W6BEG[10]
port 454 nsew signal output
rlabel metal3 s -300 17688 160 17808 4 W6BEG[11]
port 455 nsew signal output
rlabel metal3 s -300 14968 160 15088 4 W6BEG[1]
port 456 nsew signal output
rlabel metal3 s -300 15240 160 15360 4 W6BEG[2]
port 457 nsew signal output
rlabel metal3 s -300 15512 160 15632 4 W6BEG[3]
port 458 nsew signal output
rlabel metal3 s -300 15784 160 15904 4 W6BEG[4]
port 459 nsew signal output
rlabel metal3 s -300 16056 160 16176 4 W6BEG[5]
port 460 nsew signal output
rlabel metal3 s -300 16328 160 16448 4 W6BEG[6]
port 461 nsew signal output
rlabel metal3 s -300 16600 160 16720 4 W6BEG[7]
port 462 nsew signal output
rlabel metal3 s -300 16872 160 16992 4 W6BEG[8]
port 463 nsew signal output
rlabel metal3 s -300 17144 160 17264 4 W6BEG[9]
port 464 nsew signal output
rlabel metal3 s 44540 14696 45000 14816 6 W6END[0]
port 465 nsew signal input
rlabel metal3 s 44540 17416 45000 17536 6 W6END[10]
port 466 nsew signal input
rlabel metal3 s 44540 17688 45000 17808 6 W6END[11]
port 467 nsew signal input
rlabel metal3 s 44540 14968 45000 15088 6 W6END[1]
port 468 nsew signal input
rlabel metal3 s 44540 15240 45000 15360 6 W6END[2]
port 469 nsew signal input
rlabel metal3 s 44540 15512 45000 15632 6 W6END[3]
port 470 nsew signal input
rlabel metal3 s 44540 15784 45000 15904 6 W6END[4]
port 471 nsew signal input
rlabel metal3 s 44540 16056 45000 16176 6 W6END[5]
port 472 nsew signal input
rlabel metal3 s 44540 16328 45000 16448 6 W6END[6]
port 473 nsew signal input
rlabel metal3 s 44540 16600 45000 16720 6 W6END[7]
port 474 nsew signal input
rlabel metal3 s 44540 16872 45000 16992 6 W6END[8]
port 475 nsew signal input
rlabel metal3 s 44540 17144 45000 17264 6 W6END[9]
port 476 nsew signal input
rlabel metal3 s -300 10344 160 10464 4 WW4BEG[0]
port 477 nsew signal output
rlabel metal3 s -300 13064 160 13184 4 WW4BEG[10]
port 478 nsew signal output
rlabel metal3 s -300 13336 160 13456 4 WW4BEG[11]
port 479 nsew signal output
rlabel metal3 s -300 13608 160 13728 4 WW4BEG[12]
port 480 nsew signal output
rlabel metal3 s -300 13880 160 14000 4 WW4BEG[13]
port 481 nsew signal output
rlabel metal3 s -300 14152 160 14272 4 WW4BEG[14]
port 482 nsew signal output
rlabel metal3 s -300 14424 160 14544 4 WW4BEG[15]
port 483 nsew signal output
rlabel metal3 s -300 10616 160 10736 4 WW4BEG[1]
port 484 nsew signal output
rlabel metal3 s -300 10888 160 11008 4 WW4BEG[2]
port 485 nsew signal output
rlabel metal3 s -300 11160 160 11280 4 WW4BEG[3]
port 486 nsew signal output
rlabel metal3 s -300 11432 160 11552 4 WW4BEG[4]
port 487 nsew signal output
rlabel metal3 s -300 11704 160 11824 4 WW4BEG[5]
port 488 nsew signal output
rlabel metal3 s -300 11976 160 12096 4 WW4BEG[6]
port 489 nsew signal output
rlabel metal3 s -300 12248 160 12368 4 WW4BEG[7]
port 490 nsew signal output
rlabel metal3 s -300 12520 160 12640 4 WW4BEG[8]
port 491 nsew signal output
rlabel metal3 s -300 12792 160 12912 4 WW4BEG[9]
port 492 nsew signal output
rlabel metal3 s 44540 10344 45000 10464 6 WW4END[0]
port 493 nsew signal input
rlabel metal3 s 44540 13064 45000 13184 6 WW4END[10]
port 494 nsew signal input
rlabel metal3 s 44540 13336 45000 13456 6 WW4END[11]
port 495 nsew signal input
rlabel metal3 s 44540 13608 45000 13728 6 WW4END[12]
port 496 nsew signal input
rlabel metal3 s 44540 13880 45000 14000 6 WW4END[13]
port 497 nsew signal input
rlabel metal3 s 44540 14152 45000 14272 6 WW4END[14]
port 498 nsew signal input
rlabel metal3 s 44540 14424 45000 14544 6 WW4END[15]
port 499 nsew signal input
rlabel metal3 s 44540 10616 45000 10736 6 WW4END[1]
port 500 nsew signal input
rlabel metal3 s 44540 10888 45000 11008 6 WW4END[2]
port 501 nsew signal input
rlabel metal3 s 44540 11160 45000 11280 6 WW4END[3]
port 502 nsew signal input
rlabel metal3 s 44540 11432 45000 11552 6 WW4END[4]
port 503 nsew signal input
rlabel metal3 s 44540 11704 45000 11824 6 WW4END[5]
port 504 nsew signal input
rlabel metal3 s 44540 11976 45000 12096 6 WW4END[6]
port 505 nsew signal input
rlabel metal3 s 44540 12248 45000 12368 6 WW4END[7]
port 506 nsew signal input
rlabel metal3 s 44540 12520 45000 12640 6 WW4END[8]
port 507 nsew signal input
rlabel metal3 s 44540 12792 45000 12912 6 WW4END[9]
port 508 nsew signal input
rlabel metal4 s 3564 1040 3884 43568 6 vccd1
port 509 nsew power bidirectional
rlabel metal4 s 18564 1040 18884 43568 6 vccd1
port 509 nsew power bidirectional
rlabel metal4 s 33564 1040 33884 43568 6 vccd1
port 509 nsew power bidirectional
rlabel metal4 s 11064 1040 11384 43568 6 vssd1
port 510 nsew ground bidirectional
rlabel metal4 s 26064 1040 26384 43568 6 vssd1
port 510 nsew ground bidirectional
rlabel metal4 s 41064 1040 41384 43568 6 vssd1
port 510 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 44700 44700
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9775556
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/LUT4AB/runs/24_12_07_21_53/results/signoff/LUT4AB.magic.gds
string GDS_START 214348
<< end >>

