VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbyte_1rw1r_32x256_8
   CLASS BLOCK ;
   SIZE 492.56 BY 399.67 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.0 0.0 108.38 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.84 0.0 114.22 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.68 0.0 120.06 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.52 0.0 125.9 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  131.36 0.0 131.74 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  137.2 0.0 137.58 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.04 0.0 143.42 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.88 0.0 149.26 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.72 0.0 155.1 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  160.56 0.0 160.94 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  166.4 0.0 166.78 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.24 0.0 172.62 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.08 0.0 178.46 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  183.92 0.0 184.3 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.76 0.0 190.14 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.6 0.0 195.98 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.44 0.0 201.82 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.28 0.0 207.66 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  213.12 0.0 213.5 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  218.96 0.0 219.34 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.8 0.0 225.18 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.64 0.0 231.02 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  236.48 0.0 236.86 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  242.32 0.0 242.7 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.16 0.0 248.54 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  254.0 0.0 254.38 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.84 0.0 260.22 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.68 0.0 266.06 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  271.52 0.0 271.9 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  277.36 0.0 277.74 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  283.2 0.0 283.58 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  289.04 0.0 289.42 0.38 ;
      END
   END din0[31]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  78.8 0.0 79.18 0.38 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 129.77 0.38 130.15 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 138.27 0.38 138.65 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 143.185 0.38 143.565 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 153.075 0.38 153.455 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 158.05 0.38 158.43 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 166.55 0.38 166.93 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 172.19 0.38 172.57 ;
      END
   END addr0[7]
   PIN addr1[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  408.92 399.29 409.3 399.67 ;
      END
   END addr1[0]
   PIN addr1[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  492.18 84.385 492.56 84.765 ;
      END
   END addr1[1]
   PIN addr1[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  492.18 75.985 492.56 76.365 ;
      END
   END addr1[2]
   PIN addr1[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  492.18 70.49 492.56 70.87 ;
      END
   END addr1[3]
   PIN addr1[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  427.98 0.0 428.36 0.38 ;
      END
   END addr1[4]
   PIN addr1[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  425.005 0.0 425.385 0.38 ;
      END
   END addr1[5]
   PIN addr1[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  425.695 0.0 426.075 0.38 ;
      END
   END addr1[6]
   PIN addr1[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  426.44 0.0 426.82 0.38 ;
      END
   END addr1[7]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 28.89 0.38 29.27 ;
      END
   END csb0
   PIN csb1
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  492.18 384.42 492.56 384.8 ;
      END
   END csb1
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 37.39 0.38 37.77 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.1 0.0 31.48 0.38 ;
      END
   END clk0
   PIN clk1
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  461.92 399.29 462.3 399.67 ;
      END
   END clk1
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  84.64 0.0 85.02 0.38 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  90.48 0.0 90.86 0.38 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  96.32 0.0 96.7 0.38 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.16 0.0 102.54 0.38 ;
      END
   END wmask0[3]
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  146.04 0.0 146.42 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  152.86 0.0 153.24 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  158.755 0.0 159.135 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.405 0.0 167.785 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.93 0.0 173.31 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.77 0.0 179.15 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.745 0.0 185.125 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  190.985 0.0 191.365 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.605 0.0 198.985 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.465 0.0 203.845 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.705 0.0 210.085 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.945 0.0 216.325 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.185 0.0 222.565 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.425 0.0 228.805 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  234.665 0.0 235.045 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  240.515 0.0 240.895 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  245.88 0.0 246.26 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  252.195 0.0 252.575 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  261.005 0.0 261.385 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  266.37 0.0 266.75 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.21 0.0 272.59 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.345 0.0 278.725 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.585 0.0 284.965 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  290.825 0.0 291.205 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  298.445 0.0 298.825 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.305 0.0 303.685 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.545 0.0 309.925 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  315.785 0.0 316.165 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  322.025 0.0 322.405 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.265 0.0 328.645 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  334.505 0.0 334.885 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  340.745 0.0 341.125 0.38 ;
      END
   END dout0[31]
   PIN dout1[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  147.365 399.29 147.745 399.67 ;
      END
   END dout1[0]
   PIN dout1[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  153.605 399.29 153.985 399.67 ;
      END
   END dout1[1]
   PIN dout1[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  159.845 399.29 160.225 399.67 ;
      END
   END dout1[2]
   PIN dout1[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  166.085 399.29 166.465 399.67 ;
      END
   END dout1[3]
   PIN dout1[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.325 399.29 172.705 399.67 ;
      END
   END dout1[4]
   PIN dout1[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.565 399.29 178.945 399.67 ;
      END
   END dout1[5]
   PIN dout1[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.805 399.29 185.185 399.67 ;
      END
   END dout1[6]
   PIN dout1[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  191.045 399.29 191.425 399.67 ;
      END
   END dout1[7]
   PIN dout1[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.285 399.29 197.665 399.67 ;
      END
   END dout1[8]
   PIN dout1[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.525 399.29 203.905 399.67 ;
      END
   END dout1[9]
   PIN dout1[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  209.765 399.29 210.145 399.67 ;
      END
   END dout1[10]
   PIN dout1[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  216.005 399.29 216.385 399.67 ;
      END
   END dout1[11]
   PIN dout1[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.245 399.29 222.625 399.67 ;
      END
   END dout1[12]
   PIN dout1[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  228.485 399.29 228.865 399.67 ;
      END
   END dout1[13]
   PIN dout1[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  234.725 399.29 235.105 399.67 ;
      END
   END dout1[14]
   PIN dout1[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  240.965 399.29 241.345 399.67 ;
      END
   END dout1[15]
   PIN dout1[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  247.205 399.29 247.585 399.67 ;
      END
   END dout1[16]
   PIN dout1[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  253.445 399.29 253.825 399.67 ;
      END
   END dout1[17]
   PIN dout1[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  259.685 399.29 260.065 399.67 ;
      END
   END dout1[18]
   PIN dout1[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.925 399.29 266.305 399.67 ;
      END
   END dout1[19]
   PIN dout1[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  272.165 399.29 272.545 399.67 ;
      END
   END dout1[20]
   PIN dout1[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  278.405 399.29 278.785 399.67 ;
      END
   END dout1[21]
   PIN dout1[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  284.645 399.29 285.025 399.67 ;
      END
   END dout1[22]
   PIN dout1[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  290.885 399.29 291.265 399.67 ;
      END
   END dout1[23]
   PIN dout1[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  297.125 399.29 297.505 399.67 ;
      END
   END dout1[24]
   PIN dout1[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  303.365 399.29 303.745 399.67 ;
      END
   END dout1[25]
   PIN dout1[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  309.605 399.29 309.985 399.67 ;
      END
   END dout1[26]
   PIN dout1[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  315.845 399.29 316.225 399.67 ;
      END
   END dout1[27]
   PIN dout1[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  322.085 399.29 322.465 399.67 ;
      END
   END dout1[28]
   PIN dout1[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  328.325 399.29 328.705 399.67 ;
      END
   END dout1[29]
   PIN dout1[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  334.565 399.29 334.945 399.67 ;
      END
   END dout1[30]
   PIN dout1[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  340.805 399.29 341.185 399.67 ;
      END
   END dout1[31]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  490.82 0.0 492.56 399.67 ;
         LAYER met3 ;
         RECT  0.0 0.0 492.56 1.74 ;
         LAYER met3 ;
         RECT  0.0 397.93 492.56 399.67 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 399.67 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  3.48 3.48 5.22 396.19 ;
         LAYER met3 ;
         RECT  3.48 3.48 489.08 5.22 ;
         LAYER met3 ;
         RECT  3.48 394.45 489.08 396.19 ;
         LAYER met4 ;
         RECT  487.34 3.48 489.08 396.19 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 491.94 399.05 ;
   LAYER  met2 ;
      RECT  0.62 0.62 491.94 399.05 ;
   LAYER  met3 ;
      RECT  0.98 129.17 491.94 130.75 ;
      RECT  0.62 130.75 0.98 137.67 ;
      RECT  0.62 139.25 0.98 142.585 ;
      RECT  0.62 144.165 0.98 152.475 ;
      RECT  0.62 154.055 0.98 157.45 ;
      RECT  0.62 159.03 0.98 165.95 ;
      RECT  0.62 167.53 0.98 171.59 ;
      RECT  0.98 83.785 491.58 85.365 ;
      RECT  0.98 85.365 491.58 129.17 ;
      RECT  491.58 85.365 491.94 129.17 ;
      RECT  491.58 76.965 491.94 83.785 ;
      RECT  491.58 71.47 491.94 75.385 ;
      RECT  0.98 130.75 491.58 383.82 ;
      RECT  0.98 383.82 491.58 385.4 ;
      RECT  491.58 130.75 491.94 383.82 ;
      RECT  0.62 29.87 0.98 36.79 ;
      RECT  0.62 38.37 0.98 129.17 ;
      RECT  491.58 2.34 491.94 69.89 ;
      RECT  0.62 2.34 0.98 28.29 ;
      RECT  0.62 173.17 0.98 397.33 ;
      RECT  491.58 385.4 491.94 397.33 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 83.785 ;
      RECT  2.88 2.34 489.68 2.88 ;
      RECT  2.88 5.82 489.68 83.785 ;
      RECT  489.68 2.34 491.58 2.88 ;
      RECT  489.68 2.88 491.58 5.82 ;
      RECT  489.68 5.82 491.58 83.785 ;
      RECT  0.98 385.4 2.88 393.85 ;
      RECT  0.98 393.85 2.88 396.79 ;
      RECT  0.98 396.79 2.88 397.33 ;
      RECT  2.88 385.4 489.68 393.85 ;
      RECT  2.88 396.79 489.68 397.33 ;
      RECT  489.68 385.4 491.58 393.85 ;
      RECT  489.68 393.85 491.58 396.79 ;
      RECT  489.68 396.79 491.58 397.33 ;
   LAYER  met4 ;
      RECT  107.4 0.98 108.98 399.05 ;
      RECT  108.98 0.62 113.24 0.98 ;
      RECT  114.82 0.62 119.08 0.98 ;
      RECT  120.66 0.62 124.92 0.98 ;
      RECT  126.5 0.62 130.76 0.98 ;
      RECT  132.34 0.62 136.6 0.98 ;
      RECT  138.18 0.62 142.44 0.98 ;
      RECT  161.54 0.62 165.8 0.98 ;
      RECT  254.98 0.62 259.24 0.98 ;
      RECT  108.98 0.98 408.32 398.69 ;
      RECT  408.32 0.98 409.9 398.69 ;
      RECT  32.08 0.62 78.2 0.98 ;
      RECT  409.9 398.69 461.32 399.05 ;
      RECT  79.78 0.62 84.04 0.98 ;
      RECT  85.62 0.62 89.88 0.98 ;
      RECT  91.46 0.62 95.72 0.98 ;
      RECT  97.3 0.62 101.56 0.98 ;
      RECT  103.14 0.62 107.4 0.98 ;
      RECT  144.02 0.62 145.44 0.98 ;
      RECT  147.02 0.62 148.28 0.98 ;
      RECT  149.86 0.62 152.26 0.98 ;
      RECT  153.84 0.62 154.12 0.98 ;
      RECT  155.7 0.62 158.155 0.98 ;
      RECT  159.735 0.62 159.96 0.98 ;
      RECT  168.385 0.62 171.64 0.98 ;
      RECT  173.91 0.62 177.48 0.98 ;
      RECT  179.75 0.62 183.32 0.98 ;
      RECT  185.725 0.62 189.16 0.98 ;
      RECT  191.965 0.62 195.0 0.98 ;
      RECT  196.58 0.62 198.005 0.98 ;
      RECT  199.585 0.62 200.84 0.98 ;
      RECT  202.42 0.62 202.865 0.98 ;
      RECT  204.445 0.62 206.68 0.98 ;
      RECT  208.26 0.62 209.105 0.98 ;
      RECT  210.685 0.62 212.52 0.98 ;
      RECT  214.1 0.62 215.345 0.98 ;
      RECT  216.925 0.62 218.36 0.98 ;
      RECT  219.94 0.62 221.585 0.98 ;
      RECT  223.165 0.62 224.2 0.98 ;
      RECT  225.78 0.62 227.825 0.98 ;
      RECT  229.405 0.62 230.04 0.98 ;
      RECT  231.62 0.62 234.065 0.98 ;
      RECT  235.645 0.62 235.88 0.98 ;
      RECT  237.46 0.62 239.915 0.98 ;
      RECT  241.495 0.62 241.72 0.98 ;
      RECT  243.3 0.62 245.28 0.98 ;
      RECT  246.86 0.62 247.56 0.98 ;
      RECT  249.14 0.62 251.595 0.98 ;
      RECT  253.175 0.62 253.4 0.98 ;
      RECT  261.985 0.62 265.08 0.98 ;
      RECT  267.35 0.62 270.92 0.98 ;
      RECT  273.19 0.62 276.76 0.98 ;
      RECT  279.325 0.62 282.6 0.98 ;
      RECT  285.565 0.62 288.44 0.98 ;
      RECT  290.02 0.62 290.225 0.98 ;
      RECT  291.805 0.62 297.845 0.98 ;
      RECT  299.425 0.62 302.705 0.98 ;
      RECT  304.285 0.62 308.945 0.98 ;
      RECT  310.525 0.62 315.185 0.98 ;
      RECT  316.765 0.62 321.425 0.98 ;
      RECT  323.005 0.62 327.665 0.98 ;
      RECT  329.245 0.62 333.905 0.98 ;
      RECT  335.485 0.62 340.145 0.98 ;
      RECT  341.725 0.62 424.405 0.98 ;
      RECT  108.98 398.69 146.765 399.05 ;
      RECT  148.345 398.69 153.005 399.05 ;
      RECT  154.585 398.69 159.245 399.05 ;
      RECT  160.825 398.69 165.485 399.05 ;
      RECT  167.065 398.69 171.725 399.05 ;
      RECT  173.305 398.69 177.965 399.05 ;
      RECT  179.545 398.69 184.205 399.05 ;
      RECT  185.785 398.69 190.445 399.05 ;
      RECT  192.025 398.69 196.685 399.05 ;
      RECT  198.265 398.69 202.925 399.05 ;
      RECT  204.505 398.69 209.165 399.05 ;
      RECT  210.745 398.69 215.405 399.05 ;
      RECT  216.985 398.69 221.645 399.05 ;
      RECT  223.225 398.69 227.885 399.05 ;
      RECT  229.465 398.69 234.125 399.05 ;
      RECT  235.705 398.69 240.365 399.05 ;
      RECT  241.945 398.69 246.605 399.05 ;
      RECT  248.185 398.69 252.845 399.05 ;
      RECT  254.425 398.69 259.085 399.05 ;
      RECT  260.665 398.69 265.325 399.05 ;
      RECT  266.905 398.69 271.565 399.05 ;
      RECT  273.145 398.69 277.805 399.05 ;
      RECT  279.385 398.69 284.045 399.05 ;
      RECT  285.625 398.69 290.285 399.05 ;
      RECT  291.865 398.69 296.525 399.05 ;
      RECT  298.105 398.69 302.765 399.05 ;
      RECT  304.345 398.69 309.005 399.05 ;
      RECT  310.585 398.69 315.245 399.05 ;
      RECT  316.825 398.69 321.485 399.05 ;
      RECT  323.065 398.69 327.725 399.05 ;
      RECT  329.305 398.69 333.965 399.05 ;
      RECT  335.545 398.69 340.205 399.05 ;
      RECT  341.785 398.69 408.32 399.05 ;
      RECT  428.96 0.62 490.22 0.98 ;
      RECT  462.9 398.69 490.22 399.05 ;
      RECT  2.34 0.62 30.5 0.98 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 396.79 ;
      RECT  2.34 396.79 2.88 399.05 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 396.79 5.82 399.05 ;
      RECT  5.82 0.98 107.4 2.88 ;
      RECT  5.82 2.88 107.4 396.79 ;
      RECT  5.82 396.79 107.4 399.05 ;
      RECT  409.9 0.98 486.74 2.88 ;
      RECT  409.9 2.88 486.74 396.79 ;
      RECT  409.9 396.79 486.74 398.69 ;
      RECT  486.74 0.98 489.68 2.88 ;
      RECT  486.74 396.79 489.68 398.69 ;
      RECT  489.68 0.98 490.22 2.88 ;
      RECT  489.68 2.88 490.22 396.79 ;
      RECT  489.68 396.79 490.22 398.69 ;
   END
END    sky130_sram_1kbyte_1rw1r_32x256_8
END    LIBRARY
