magic
tech sky130A
magscale 1 2
timestamp 1733618678
<< viali >>
rect 3893 8585 3927 8619
rect 5641 8585 5675 8619
rect 8033 8585 8067 8619
rect 10241 8585 10275 8619
rect 14657 8585 14691 8619
rect 19441 8585 19475 8619
rect 21281 8585 21315 8619
rect 25697 8585 25731 8619
rect 27721 8585 27755 8619
rect 30113 8585 30147 8619
rect 32321 8585 32355 8619
rect 34897 8585 34931 8619
rect 36737 8585 36771 8619
rect 38761 8585 38795 8619
rect 41153 8585 41187 8619
rect 43361 8585 43395 8619
rect 44741 8585 44775 8619
rect 1409 8517 1443 8551
rect 1777 8517 1811 8551
rect 12173 8517 12207 8551
rect 12541 8517 12575 8551
rect 16681 8517 16715 8551
rect 23213 8517 23247 8551
rect 4077 8449 4111 8483
rect 5917 8449 5951 8483
rect 8217 8449 8251 8483
rect 10425 8449 10459 8483
rect 14841 8449 14875 8483
rect 17049 8449 17083 8483
rect 19349 8449 19383 8483
rect 21465 8449 21499 8483
rect 23581 8449 23615 8483
rect 25881 8449 25915 8483
rect 27997 8449 28031 8483
rect 30297 8449 30331 8483
rect 32505 8449 32539 8483
rect 34805 8449 34839 8483
rect 36921 8449 36955 8483
rect 39037 8449 39071 8483
rect 41337 8449 41371 8483
rect 43545 8449 43579 8483
rect 44557 8449 44591 8483
rect 22937 3145 22971 3179
rect 21833 3009 21867 3043
rect 22385 3009 22419 3043
rect 22753 3009 22787 3043
rect 23397 3009 23431 3043
rect 22017 2805 22051 2839
rect 22569 2805 22603 2839
rect 23213 2805 23247 2839
rect 17049 2601 17083 2635
rect 19349 2601 19383 2635
rect 20637 2601 20671 2635
rect 21557 2601 21591 2635
rect 22385 2601 22419 2635
rect 22937 2601 22971 2635
rect 23305 2601 23339 2635
rect 24409 2601 24443 2635
rect 25973 2601 26007 2635
rect 28181 2601 28215 2635
rect 29193 2601 29227 2635
rect 30389 2601 30423 2635
rect 32597 2601 32631 2635
rect 34805 2601 34839 2635
rect 37013 2601 37047 2635
rect 39129 2601 39163 2635
rect 41337 2601 41371 2635
rect 43821 2601 43855 2635
rect 44557 2601 44591 2635
rect 22845 2533 22879 2567
rect 23949 2533 23983 2567
rect 27997 2533 28031 2567
rect 17233 2397 17267 2431
rect 18797 2397 18831 2431
rect 19533 2397 19567 2431
rect 19625 2397 19659 2431
rect 19901 2397 19935 2431
rect 20361 2397 20395 2431
rect 20821 2397 20855 2431
rect 21281 2397 21315 2431
rect 21741 2397 21775 2431
rect 21833 2397 21867 2431
rect 22109 2397 22143 2431
rect 22569 2397 22603 2431
rect 22661 2397 22695 2431
rect 23129 2397 23163 2431
rect 23489 2397 23523 2431
rect 24133 2397 24167 2431
rect 24593 2397 24627 2431
rect 26157 2397 26191 2431
rect 27813 2397 27847 2431
rect 28365 2397 28399 2431
rect 29377 2397 29411 2431
rect 30573 2397 30607 2431
rect 30665 2397 30699 2431
rect 30941 2397 30975 2431
rect 31217 2397 31251 2431
rect 32781 2397 32815 2431
rect 34989 2397 35023 2431
rect 37197 2397 37231 2431
rect 39313 2397 39347 2431
rect 41521 2397 41555 2431
rect 44005 2397 44039 2431
rect 44373 2397 44407 2431
rect 44833 2397 44867 2431
rect 45201 2397 45235 2431
rect 23765 2329 23799 2363
rect 18981 2261 19015 2295
rect 19809 2261 19843 2295
rect 20085 2261 20119 2295
rect 20545 2261 20579 2295
rect 21097 2261 21131 2295
rect 22017 2261 22051 2295
rect 22293 2261 22327 2295
rect 23673 2261 23707 2295
rect 30849 2261 30883 2295
rect 31125 2261 31159 2295
rect 31401 2261 31435 2295
rect 44649 2261 44683 2295
rect 45017 2261 45051 2295
rect 3341 2057 3375 2091
rect 15393 2057 15427 2091
rect 16221 2057 16255 2091
rect 16497 2057 16531 2091
rect 17049 2057 17083 2091
rect 17601 2057 17635 2091
rect 18153 2057 18187 2091
rect 18705 2057 18739 2091
rect 19257 2057 19291 2091
rect 20085 2057 20119 2091
rect 20913 2057 20947 2091
rect 23489 2057 23523 2091
rect 24041 2057 24075 2091
rect 24961 2057 24995 2091
rect 27261 2057 27295 2091
rect 28273 2057 28307 2091
rect 31861 2057 31895 2091
rect 32137 2057 32171 2091
rect 33241 2057 33275 2091
rect 35173 2057 35207 2091
rect 37381 2057 37415 2091
rect 39681 2057 39715 2091
rect 40141 2057 40175 2091
rect 40417 2057 40451 2091
rect 40693 2057 40727 2091
rect 41797 2057 41831 2091
rect 44373 2057 44407 2091
rect 22017 1989 22051 2023
rect 31217 1989 31251 2023
rect 36369 1989 36403 2023
rect 1409 1921 1443 1955
rect 1685 1921 1719 1955
rect 2329 1921 2363 1955
rect 3157 1921 3191 1955
rect 15025 1921 15059 1955
rect 15485 1921 15519 1955
rect 15761 1921 15795 1955
rect 16037 1921 16071 1955
rect 16313 1921 16347 1955
rect 16865 1921 16899 1955
rect 17141 1921 17175 1955
rect 17417 1921 17451 1955
rect 17693 1921 17727 1955
rect 17969 1921 18003 1955
rect 18245 1921 18279 1955
rect 18521 1921 18555 1955
rect 18797 1921 18831 1955
rect 19073 1921 19107 1955
rect 19341 1925 19375 1959
rect 19625 1921 19659 1955
rect 19901 1921 19935 1955
rect 20177 1921 20211 1955
rect 20453 1921 20487 1955
rect 20729 1921 20763 1955
rect 21005 1921 21039 1955
rect 21465 1921 21499 1955
rect 22477 1921 22511 1955
rect 23029 1921 23063 1955
rect 23305 1921 23339 1955
rect 23581 1921 23615 1955
rect 24225 1921 24259 1955
rect 24317 1921 24351 1955
rect 24685 1921 24719 1955
rect 25145 1921 25179 1955
rect 25237 1921 25271 1955
rect 25513 1921 25547 1955
rect 25973 1921 26007 1955
rect 26341 1921 26375 1955
rect 26617 1921 26651 1955
rect 26985 1921 27019 1955
rect 27421 1921 27455 1955
rect 27537 1921 27571 1955
rect 27813 1921 27847 1955
rect 28089 1921 28123 1955
rect 28457 1921 28491 1955
rect 28825 1921 28859 1955
rect 29101 1921 29135 1955
rect 29377 1921 29411 1955
rect 29653 1921 29687 1955
rect 29929 1921 29963 1955
rect 30297 1921 30331 1955
rect 30573 1921 30607 1955
rect 30849 1921 30883 1955
rect 31677 1921 31711 1955
rect 32321 1921 32355 1955
rect 32873 1921 32907 1955
rect 33425 1921 33459 1955
rect 33793 1921 33827 1955
rect 34253 1921 34287 1955
rect 35357 1921 35391 1955
rect 35449 1921 35483 1955
rect 37565 1921 37599 1955
rect 38025 1921 38059 1955
rect 38393 1921 38427 1955
rect 39865 1921 39899 1955
rect 40325 1921 40359 1955
rect 40601 1921 40635 1955
rect 40877 1921 40911 1955
rect 41981 1921 42015 1955
rect 44557 1921 44591 1955
rect 44833 1921 44867 1955
rect 45201 1921 45235 1955
rect 2053 1853 2087 1887
rect 1869 1785 1903 1819
rect 17325 1785 17359 1819
rect 18981 1785 19015 1819
rect 19533 1785 19567 1819
rect 20637 1785 20671 1819
rect 21649 1785 21683 1819
rect 23213 1785 23247 1819
rect 25421 1785 25455 1819
rect 44649 1785 44683 1819
rect 45017 1785 45051 1819
rect 1593 1717 1627 1751
rect 15209 1717 15243 1751
rect 15945 1717 15979 1751
rect 17877 1717 17911 1751
rect 18429 1717 18463 1751
rect 19809 1717 19843 1751
rect 20361 1717 20395 1751
rect 21189 1717 21223 1751
rect 22109 1717 22143 1751
rect 22661 1717 22695 1751
rect 23765 1717 23799 1751
rect 24501 1717 24535 1751
rect 24869 1717 24903 1751
rect 25697 1717 25731 1751
rect 26157 1717 26191 1751
rect 26525 1717 26559 1751
rect 26801 1717 26835 1751
rect 27169 1717 27203 1751
rect 27721 1717 27755 1751
rect 27997 1717 28031 1751
rect 28641 1717 28675 1751
rect 29009 1717 29043 1751
rect 29285 1717 29319 1751
rect 29561 1717 29595 1751
rect 29837 1717 29871 1751
rect 30113 1717 30147 1751
rect 30481 1717 30515 1751
rect 30757 1717 30791 1751
rect 31033 1717 31067 1751
rect 31309 1717 31343 1751
rect 33057 1717 33091 1751
rect 33885 1717 33919 1751
rect 34437 1717 34471 1751
rect 35633 1717 35667 1751
rect 36461 1717 36495 1751
rect 38209 1717 38243 1751
rect 38577 1717 38611 1751
rect 14565 1513 14599 1547
rect 15117 1513 15151 1547
rect 15393 1513 15427 1547
rect 16497 1513 16531 1547
rect 16957 1513 16991 1547
rect 17325 1513 17359 1547
rect 18061 1513 18095 1547
rect 18337 1513 18371 1547
rect 18613 1513 18647 1547
rect 18889 1513 18923 1547
rect 25053 1513 25087 1547
rect 27905 1513 27939 1547
rect 29745 1513 29779 1547
rect 31033 1513 31067 1547
rect 32321 1513 32355 1547
rect 33425 1513 33459 1547
rect 33977 1513 34011 1547
rect 34897 1513 34931 1547
rect 35449 1513 35483 1547
rect 36001 1513 36035 1547
rect 36553 1513 36587 1547
rect 38025 1513 38059 1547
rect 39129 1513 39163 1547
rect 40417 1513 40451 1547
rect 42441 1513 42475 1547
rect 44649 1513 44683 1547
rect 1869 1445 1903 1479
rect 14289 1445 14323 1479
rect 15669 1445 15703 1479
rect 17601 1445 17635 1479
rect 38669 1445 38703 1479
rect 40141 1445 40175 1479
rect 43545 1445 43579 1479
rect 43821 1445 43855 1479
rect 44373 1445 44407 1479
rect 45017 1445 45051 1479
rect 22477 1377 22511 1411
rect 23581 1377 23615 1411
rect 26433 1377 26467 1411
rect 28917 1377 28951 1411
rect 31769 1377 31803 1411
rect 37657 1377 37691 1411
rect 1409 1309 1443 1343
rect 1685 1309 1719 1343
rect 2145 1309 2179 1343
rect 2421 1309 2455 1343
rect 2697 1309 2731 1343
rect 3433 1309 3467 1343
rect 3893 1309 3927 1343
rect 4261 1309 4295 1343
rect 4629 1309 4663 1343
rect 4997 1309 5031 1343
rect 5365 1309 5399 1343
rect 5733 1309 5767 1343
rect 6009 1309 6043 1343
rect 6469 1309 6503 1343
rect 6837 1309 6871 1343
rect 7205 1309 7239 1343
rect 7573 1309 7607 1343
rect 7941 1309 7975 1343
rect 8309 1309 8343 1343
rect 8585 1309 8619 1343
rect 9045 1309 9079 1343
rect 9413 1309 9447 1343
rect 9781 1309 9815 1343
rect 10149 1309 10183 1343
rect 10517 1309 10551 1343
rect 10885 1309 10919 1343
rect 11161 1309 11195 1343
rect 11621 1309 11655 1343
rect 11989 1309 12023 1343
rect 12357 1309 12391 1343
rect 12633 1309 12667 1343
rect 12909 1309 12943 1343
rect 13185 1309 13219 1343
rect 13461 1309 13495 1343
rect 13737 1309 13771 1343
rect 14105 1309 14139 1343
rect 14381 1309 14415 1343
rect 14657 1309 14691 1343
rect 14933 1309 14967 1343
rect 15209 1309 15243 1343
rect 15485 1309 15519 1343
rect 15761 1309 15795 1343
rect 16037 1309 16071 1343
rect 16313 1309 16347 1343
rect 16773 1309 16807 1343
rect 17049 1309 17083 1343
rect 17509 1309 17543 1343
rect 17785 1309 17819 1343
rect 18245 1309 18279 1343
rect 18521 1309 18555 1343
rect 18797 1309 18831 1343
rect 19073 1309 19107 1343
rect 19257 1309 19291 1343
rect 19533 1309 19567 1343
rect 19901 1309 19935 1343
rect 20269 1309 20303 1343
rect 21373 1309 21407 1343
rect 21833 1309 21867 1343
rect 22845 1309 22879 1343
rect 23949 1309 23983 1343
rect 24501 1309 24535 1343
rect 25421 1309 25455 1343
rect 25789 1309 25823 1343
rect 26709 1309 26743 1343
rect 26985 1309 27019 1343
rect 27353 1309 27387 1343
rect 27813 1309 27847 1343
rect 28273 1309 28307 1343
rect 29193 1309 29227 1343
rect 29653 1309 29687 1343
rect 30665 1309 30699 1343
rect 30941 1309 30975 1343
rect 31493 1309 31527 1343
rect 32229 1309 32263 1343
rect 32689 1309 32723 1343
rect 35909 1309 35943 1343
rect 39681 1309 39715 1343
rect 40601 1309 40635 1343
rect 40877 1309 40911 1343
rect 41153 1309 41187 1343
rect 41981 1309 42015 1343
rect 42257 1309 42291 1343
rect 42625 1309 42659 1343
rect 42901 1309 42935 1343
rect 43177 1309 43211 1343
rect 43453 1309 43487 1343
rect 43729 1309 43763 1343
rect 44005 1309 44039 1343
rect 44281 1309 44315 1343
rect 44557 1309 44591 1343
rect 44833 1309 44867 1343
rect 45201 1309 45235 1343
rect 20729 1241 20763 1275
rect 22201 1241 22235 1275
rect 23305 1241 23339 1275
rect 24961 1241 24995 1275
rect 30297 1241 30331 1275
rect 33333 1241 33367 1275
rect 33885 1241 33919 1275
rect 34805 1241 34839 1275
rect 35357 1241 35391 1275
rect 36461 1241 36495 1275
rect 37381 1241 37415 1275
rect 37933 1241 37967 1275
rect 38485 1241 38519 1275
rect 39037 1241 39071 1275
rect 39957 1241 39991 1275
rect 1593 1173 1627 1207
rect 2329 1173 2363 1207
rect 3617 1173 3651 1207
rect 4077 1173 4111 1207
rect 4445 1173 4479 1207
rect 4813 1173 4847 1207
rect 5181 1173 5215 1207
rect 5549 1173 5583 1207
rect 5917 1173 5951 1207
rect 6193 1173 6227 1207
rect 6653 1173 6687 1207
rect 7021 1173 7055 1207
rect 7389 1173 7423 1207
rect 7757 1173 7791 1207
rect 8125 1173 8159 1207
rect 8493 1173 8527 1207
rect 8769 1173 8803 1207
rect 9229 1173 9263 1207
rect 9597 1173 9631 1207
rect 9965 1173 9999 1207
rect 10333 1173 10367 1207
rect 10701 1173 10735 1207
rect 11069 1173 11103 1207
rect 11345 1173 11379 1207
rect 11805 1173 11839 1207
rect 12173 1173 12207 1207
rect 12541 1173 12575 1207
rect 12817 1173 12851 1207
rect 13093 1173 13127 1207
rect 13369 1173 13403 1207
rect 13645 1173 13679 1207
rect 13921 1173 13955 1207
rect 14841 1173 14875 1207
rect 15945 1173 15979 1207
rect 16221 1173 16255 1207
rect 17233 1173 17267 1207
rect 19441 1173 19475 1207
rect 19717 1173 19751 1207
rect 20085 1173 20119 1207
rect 20453 1173 20487 1207
rect 20821 1173 20855 1207
rect 21557 1173 21591 1207
rect 22017 1173 22051 1207
rect 23029 1173 23063 1207
rect 24133 1173 24167 1207
rect 24685 1173 24719 1207
rect 25605 1173 25639 1207
rect 25973 1173 26007 1207
rect 27169 1173 27203 1207
rect 27537 1173 27571 1207
rect 28457 1173 28491 1207
rect 32873 1173 32907 1207
rect 39497 1173 39531 1207
rect 41797 1173 41831 1207
rect 42073 1173 42107 1207
rect 42717 1173 42751 1207
rect 42993 1173 43027 1207
rect 43269 1173 43303 1207
rect 44097 1173 44131 1207
<< metal1 >>
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 22370 8956 22376 8968
rect 17368 8928 22376 8956
rect 17368 8916 17374 8928
rect 22370 8916 22376 8928
rect 22428 8916 22434 8968
rect 8202 8848 8208 8900
rect 8260 8888 8266 8900
rect 22922 8888 22928 8900
rect 8260 8860 22928 8888
rect 8260 8848 8266 8860
rect 22922 8848 22928 8860
rect 22980 8848 22986 8900
rect 4062 8780 4068 8832
rect 4120 8820 4126 8832
rect 23658 8820 23664 8832
rect 4120 8792 23664 8820
rect 4120 8780 4126 8792
rect 23658 8780 23664 8792
rect 23716 8780 23722 8832
rect 1104 8730 45696 8752
rect 1104 8678 12058 8730
rect 12110 8678 12122 8730
rect 12174 8678 12186 8730
rect 12238 8678 12250 8730
rect 12302 8678 12314 8730
rect 12366 8678 23166 8730
rect 23218 8678 23230 8730
rect 23282 8678 23294 8730
rect 23346 8678 23358 8730
rect 23410 8678 23422 8730
rect 23474 8678 34274 8730
rect 34326 8678 34338 8730
rect 34390 8678 34402 8730
rect 34454 8678 34466 8730
rect 34518 8678 34530 8730
rect 34582 8678 45382 8730
rect 45434 8678 45446 8730
rect 45498 8678 45510 8730
rect 45562 8678 45574 8730
rect 45626 8678 45638 8730
rect 45690 8678 45696 8730
rect 1104 8656 45696 8678
rect 3418 8576 3424 8628
rect 3476 8616 3482 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3476 8588 3893 8616
rect 3476 8576 3482 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 3881 8579 3939 8585
rect 5626 8576 5632 8628
rect 5684 8576 5690 8628
rect 7834 8576 7840 8628
rect 7892 8616 7898 8628
rect 8021 8619 8079 8625
rect 8021 8616 8033 8619
rect 7892 8588 8033 8616
rect 7892 8576 7898 8588
rect 8021 8585 8033 8588
rect 8067 8585 8079 8619
rect 8021 8579 8079 8585
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10229 8619 10287 8625
rect 10229 8616 10241 8619
rect 10100 8588 10241 8616
rect 10100 8576 10106 8588
rect 10229 8585 10241 8588
rect 10275 8585 10287 8619
rect 10229 8579 10287 8585
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 14516 8588 14657 8616
rect 14516 8576 14522 8588
rect 14645 8585 14657 8588
rect 14691 8585 14703 8619
rect 17310 8616 17316 8628
rect 14645 8579 14703 8585
rect 16592 8588 17316 8616
rect 1394 8508 1400 8560
rect 1452 8508 1458 8560
rect 1765 8551 1823 8557
rect 1765 8517 1777 8551
rect 1811 8548 1823 8551
rect 1811 8520 10548 8548
rect 1811 8517 1823 8520
rect 1765 8511 1823 8517
rect 4062 8440 4068 8492
rect 4120 8440 4126 8492
rect 5905 8483 5963 8489
rect 5905 8449 5917 8483
rect 5951 8480 5963 8483
rect 5951 8452 6914 8480
rect 5951 8449 5963 8452
rect 5905 8443 5963 8449
rect 6886 8344 6914 8452
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8449 10471 8483
rect 10520 8480 10548 8520
rect 12158 8508 12164 8560
rect 12216 8508 12222 8560
rect 12529 8551 12587 8557
rect 12529 8517 12541 8551
rect 12575 8548 12587 8551
rect 16592 8548 16620 8588
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 18932 8588 19441 8616
rect 18932 8576 18938 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 21082 8576 21088 8628
rect 21140 8616 21146 8628
rect 21269 8619 21327 8625
rect 21269 8616 21281 8619
rect 21140 8588 21281 8616
rect 21140 8576 21146 8588
rect 21269 8585 21281 8588
rect 21315 8585 21327 8619
rect 21269 8579 21327 8585
rect 25498 8576 25504 8628
rect 25556 8616 25562 8628
rect 25685 8619 25743 8625
rect 25685 8616 25697 8619
rect 25556 8588 25697 8616
rect 25556 8576 25562 8588
rect 25685 8585 25697 8588
rect 25731 8585 25743 8619
rect 25685 8579 25743 8585
rect 27706 8576 27712 8628
rect 27764 8576 27770 8628
rect 29914 8576 29920 8628
rect 29972 8616 29978 8628
rect 30101 8619 30159 8625
rect 30101 8616 30113 8619
rect 29972 8588 30113 8616
rect 29972 8576 29978 8588
rect 30101 8585 30113 8588
rect 30147 8585 30159 8619
rect 30101 8579 30159 8585
rect 32122 8576 32128 8628
rect 32180 8616 32186 8628
rect 32309 8619 32367 8625
rect 32309 8616 32321 8619
rect 32180 8588 32321 8616
rect 32180 8576 32186 8588
rect 32309 8585 32321 8588
rect 32355 8585 32367 8619
rect 32309 8579 32367 8585
rect 34146 8576 34152 8628
rect 34204 8616 34210 8628
rect 34885 8619 34943 8625
rect 34885 8616 34897 8619
rect 34204 8588 34897 8616
rect 34204 8576 34210 8588
rect 34885 8585 34897 8588
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 36538 8576 36544 8628
rect 36596 8616 36602 8628
rect 36725 8619 36783 8625
rect 36725 8616 36737 8619
rect 36596 8588 36737 8616
rect 36596 8576 36602 8588
rect 36725 8585 36737 8588
rect 36771 8585 36783 8619
rect 36725 8579 36783 8585
rect 38746 8576 38752 8628
rect 38804 8576 38810 8628
rect 40954 8576 40960 8628
rect 41012 8616 41018 8628
rect 41141 8619 41199 8625
rect 41141 8616 41153 8619
rect 41012 8588 41153 8616
rect 41012 8576 41018 8588
rect 41141 8585 41153 8588
rect 41187 8585 41199 8619
rect 41141 8579 41199 8585
rect 43162 8576 43168 8628
rect 43220 8616 43226 8628
rect 43349 8619 43407 8625
rect 43349 8616 43361 8619
rect 43220 8588 43361 8616
rect 43220 8576 43226 8588
rect 43349 8585 43361 8588
rect 43395 8585 43407 8619
rect 43349 8579 43407 8585
rect 44729 8619 44787 8625
rect 44729 8585 44741 8619
rect 44775 8616 44787 8619
rect 45278 8616 45284 8628
rect 44775 8588 45284 8616
rect 44775 8585 44787 8588
rect 44729 8579 44787 8585
rect 45278 8576 45284 8588
rect 45336 8576 45342 8628
rect 12575 8520 16620 8548
rect 12575 8517 12587 8520
rect 12529 8511 12587 8517
rect 16666 8508 16672 8560
rect 16724 8508 16730 8560
rect 20622 8548 20628 8560
rect 16960 8520 20628 8548
rect 13814 8480 13820 8492
rect 10520 8452 13820 8480
rect 10413 8443 10471 8449
rect 10428 8412 10456 8443
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14829 8483 14887 8489
rect 14829 8449 14841 8483
rect 14875 8480 14887 8483
rect 16960 8480 16988 8520
rect 20622 8508 20628 8520
rect 20680 8508 20686 8560
rect 23014 8508 23020 8560
rect 23072 8548 23078 8560
rect 23201 8551 23259 8557
rect 23201 8548 23213 8551
rect 23072 8520 23213 8548
rect 23072 8508 23078 8520
rect 23201 8517 23213 8520
rect 23247 8517 23259 8551
rect 23201 8511 23259 8517
rect 14875 8452 16988 8480
rect 14875 8449 14887 8452
rect 14829 8443 14887 8449
rect 17034 8440 17040 8492
rect 17092 8440 17098 8492
rect 19242 8480 19248 8492
rect 17512 8452 19248 8480
rect 17512 8412 17540 8452
rect 19242 8440 19248 8452
rect 19300 8440 19306 8492
rect 19334 8440 19340 8492
rect 19392 8440 19398 8492
rect 21450 8440 21456 8492
rect 21508 8440 21514 8492
rect 23566 8440 23572 8492
rect 23624 8440 23630 8492
rect 25866 8440 25872 8492
rect 25924 8440 25930 8492
rect 27982 8440 27988 8492
rect 28040 8440 28046 8492
rect 30285 8483 30343 8489
rect 30285 8449 30297 8483
rect 30331 8480 30343 8483
rect 30374 8480 30380 8492
rect 30331 8452 30380 8480
rect 30331 8449 30343 8452
rect 30285 8443 30343 8449
rect 30374 8440 30380 8452
rect 30432 8440 30438 8492
rect 32490 8440 32496 8492
rect 32548 8440 32554 8492
rect 34790 8440 34796 8492
rect 34848 8440 34854 8492
rect 36906 8440 36912 8492
rect 36964 8440 36970 8492
rect 39022 8440 39028 8492
rect 39080 8440 39086 8492
rect 41322 8440 41328 8492
rect 41380 8440 41386 8492
rect 43530 8440 43536 8492
rect 43588 8440 43594 8492
rect 44542 8440 44548 8492
rect 44600 8440 44606 8492
rect 23014 8412 23020 8424
rect 10428 8384 17540 8412
rect 17788 8384 23020 8412
rect 6886 8316 9674 8344
rect 9646 8276 9674 8316
rect 17788 8276 17816 8384
rect 23014 8372 23020 8384
rect 23072 8372 23078 8424
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 24394 8344 24400 8356
rect 19300 8316 24400 8344
rect 19300 8304 19306 8316
rect 24394 8304 24400 8316
rect 24452 8304 24458 8356
rect 9646 8248 17816 8276
rect 1104 8186 45540 8208
rect 1104 8134 6504 8186
rect 6556 8134 6568 8186
rect 6620 8134 6632 8186
rect 6684 8134 6696 8186
rect 6748 8134 6760 8186
rect 6812 8134 17612 8186
rect 17664 8134 17676 8186
rect 17728 8134 17740 8186
rect 17792 8134 17804 8186
rect 17856 8134 17868 8186
rect 17920 8134 28720 8186
rect 28772 8134 28784 8186
rect 28836 8134 28848 8186
rect 28900 8134 28912 8186
rect 28964 8134 28976 8186
rect 29028 8134 39828 8186
rect 39880 8134 39892 8186
rect 39944 8134 39956 8186
rect 40008 8134 40020 8186
rect 40072 8134 40084 8186
rect 40136 8134 45540 8186
rect 1104 8112 45540 8134
rect 1104 7642 45696 7664
rect 1104 7590 12058 7642
rect 12110 7590 12122 7642
rect 12174 7590 12186 7642
rect 12238 7590 12250 7642
rect 12302 7590 12314 7642
rect 12366 7590 23166 7642
rect 23218 7590 23230 7642
rect 23282 7590 23294 7642
rect 23346 7590 23358 7642
rect 23410 7590 23422 7642
rect 23474 7590 34274 7642
rect 34326 7590 34338 7642
rect 34390 7590 34402 7642
rect 34454 7590 34466 7642
rect 34518 7590 34530 7642
rect 34582 7590 45382 7642
rect 45434 7590 45446 7642
rect 45498 7590 45510 7642
rect 45562 7590 45574 7642
rect 45626 7590 45638 7642
rect 45690 7590 45696 7642
rect 1104 7568 45696 7590
rect 1104 7098 45540 7120
rect 1104 7046 6504 7098
rect 6556 7046 6568 7098
rect 6620 7046 6632 7098
rect 6684 7046 6696 7098
rect 6748 7046 6760 7098
rect 6812 7046 17612 7098
rect 17664 7046 17676 7098
rect 17728 7046 17740 7098
rect 17792 7046 17804 7098
rect 17856 7046 17868 7098
rect 17920 7046 28720 7098
rect 28772 7046 28784 7098
rect 28836 7046 28848 7098
rect 28900 7046 28912 7098
rect 28964 7046 28976 7098
rect 29028 7046 39828 7098
rect 39880 7046 39892 7098
rect 39944 7046 39956 7098
rect 40008 7046 40020 7098
rect 40072 7046 40084 7098
rect 40136 7046 45540 7098
rect 1104 7024 45540 7046
rect 1104 6554 45696 6576
rect 1104 6502 12058 6554
rect 12110 6502 12122 6554
rect 12174 6502 12186 6554
rect 12238 6502 12250 6554
rect 12302 6502 12314 6554
rect 12366 6502 23166 6554
rect 23218 6502 23230 6554
rect 23282 6502 23294 6554
rect 23346 6502 23358 6554
rect 23410 6502 23422 6554
rect 23474 6502 34274 6554
rect 34326 6502 34338 6554
rect 34390 6502 34402 6554
rect 34454 6502 34466 6554
rect 34518 6502 34530 6554
rect 34582 6502 45382 6554
rect 45434 6502 45446 6554
rect 45498 6502 45510 6554
rect 45562 6502 45574 6554
rect 45626 6502 45638 6554
rect 45690 6502 45696 6554
rect 1104 6480 45696 6502
rect 1104 6010 45540 6032
rect 1104 5958 6504 6010
rect 6556 5958 6568 6010
rect 6620 5958 6632 6010
rect 6684 5958 6696 6010
rect 6748 5958 6760 6010
rect 6812 5958 17612 6010
rect 17664 5958 17676 6010
rect 17728 5958 17740 6010
rect 17792 5958 17804 6010
rect 17856 5958 17868 6010
rect 17920 5958 28720 6010
rect 28772 5958 28784 6010
rect 28836 5958 28848 6010
rect 28900 5958 28912 6010
rect 28964 5958 28976 6010
rect 29028 5958 39828 6010
rect 39880 5958 39892 6010
rect 39944 5958 39956 6010
rect 40008 5958 40020 6010
rect 40072 5958 40084 6010
rect 40136 5958 45540 6010
rect 1104 5936 45540 5958
rect 1104 5466 45696 5488
rect 1104 5414 12058 5466
rect 12110 5414 12122 5466
rect 12174 5414 12186 5466
rect 12238 5414 12250 5466
rect 12302 5414 12314 5466
rect 12366 5414 23166 5466
rect 23218 5414 23230 5466
rect 23282 5414 23294 5466
rect 23346 5414 23358 5466
rect 23410 5414 23422 5466
rect 23474 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 34530 5466
rect 34582 5414 45382 5466
rect 45434 5414 45446 5466
rect 45498 5414 45510 5466
rect 45562 5414 45574 5466
rect 45626 5414 45638 5466
rect 45690 5414 45696 5466
rect 1104 5392 45696 5414
rect 1104 4922 45540 4944
rect 1104 4870 6504 4922
rect 6556 4870 6568 4922
rect 6620 4870 6632 4922
rect 6684 4870 6696 4922
rect 6748 4870 6760 4922
rect 6812 4870 17612 4922
rect 17664 4870 17676 4922
rect 17728 4870 17740 4922
rect 17792 4870 17804 4922
rect 17856 4870 17868 4922
rect 17920 4870 28720 4922
rect 28772 4870 28784 4922
rect 28836 4870 28848 4922
rect 28900 4870 28912 4922
rect 28964 4870 28976 4922
rect 29028 4870 39828 4922
rect 39880 4870 39892 4922
rect 39944 4870 39956 4922
rect 40008 4870 40020 4922
rect 40072 4870 40084 4922
rect 40136 4870 45540 4922
rect 1104 4848 45540 4870
rect 5534 4496 5540 4548
rect 5592 4536 5598 4548
rect 24302 4536 24308 4548
rect 5592 4508 24308 4536
rect 5592 4496 5598 4508
rect 24302 4496 24308 4508
rect 24360 4496 24366 4548
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 26602 4468 26608 4480
rect 2372 4440 26608 4468
rect 2372 4428 2378 4440
rect 26602 4428 26608 4440
rect 26660 4428 26666 4480
rect 1104 4378 45696 4400
rect 1104 4326 12058 4378
rect 12110 4326 12122 4378
rect 12174 4326 12186 4378
rect 12238 4326 12250 4378
rect 12302 4326 12314 4378
rect 12366 4326 23166 4378
rect 23218 4326 23230 4378
rect 23282 4326 23294 4378
rect 23346 4326 23358 4378
rect 23410 4326 23422 4378
rect 23474 4326 34274 4378
rect 34326 4326 34338 4378
rect 34390 4326 34402 4378
rect 34454 4326 34466 4378
rect 34518 4326 34530 4378
rect 34582 4326 45382 4378
rect 45434 4326 45446 4378
rect 45498 4326 45510 4378
rect 45562 4326 45574 4378
rect 45626 4326 45638 4378
rect 45690 4326 45696 4378
rect 1104 4304 45696 4326
rect 18506 4224 18512 4276
rect 18564 4264 18570 4276
rect 42426 4264 42432 4276
rect 18564 4236 42432 4264
rect 18564 4224 18570 4236
rect 42426 4224 42432 4236
rect 42484 4224 42490 4276
rect 16942 4156 16948 4208
rect 17000 4196 17006 4208
rect 41138 4196 41144 4208
rect 17000 4168 41144 4196
rect 17000 4156 17006 4168
rect 41138 4156 41144 4168
rect 41196 4156 41202 4208
rect 1104 3834 45540 3856
rect 1104 3782 6504 3834
rect 6556 3782 6568 3834
rect 6620 3782 6632 3834
rect 6684 3782 6696 3834
rect 6748 3782 6760 3834
rect 6812 3782 17612 3834
rect 17664 3782 17676 3834
rect 17728 3782 17740 3834
rect 17792 3782 17804 3834
rect 17856 3782 17868 3834
rect 17920 3782 28720 3834
rect 28772 3782 28784 3834
rect 28836 3782 28848 3834
rect 28900 3782 28912 3834
rect 28964 3782 28976 3834
rect 29028 3782 39828 3834
rect 39880 3782 39892 3834
rect 39944 3782 39956 3834
rect 40008 3782 40020 3834
rect 40072 3782 40084 3834
rect 40136 3782 45540 3834
rect 1104 3760 45540 3782
rect 16206 3612 16212 3664
rect 16264 3652 16270 3664
rect 35250 3652 35256 3664
rect 16264 3624 35256 3652
rect 16264 3612 16270 3624
rect 35250 3612 35256 3624
rect 35308 3612 35314 3664
rect 12406 3556 25544 3584
rect 8110 3408 8116 3460
rect 8168 3448 8174 3460
rect 12406 3448 12434 3556
rect 25516 3528 25544 3556
rect 22738 3476 22744 3528
rect 22796 3516 22802 3528
rect 23014 3516 23020 3528
rect 22796 3488 23020 3516
rect 22796 3476 22802 3488
rect 23014 3476 23020 3488
rect 23072 3476 23078 3528
rect 25498 3476 25504 3528
rect 25556 3476 25562 3528
rect 8168 3420 12434 3448
rect 8168 3408 8174 3420
rect 20438 3408 20444 3460
rect 20496 3448 20502 3460
rect 28626 3448 28632 3460
rect 20496 3420 28632 3448
rect 20496 3408 20502 3420
rect 28626 3408 28632 3420
rect 28684 3408 28690 3460
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 25038 3380 25044 3392
rect 17552 3352 25044 3380
rect 17552 3340 17558 3352
rect 25038 3340 25044 3352
rect 25096 3340 25102 3392
rect 1104 3290 45696 3312
rect 1104 3238 12058 3290
rect 12110 3238 12122 3290
rect 12174 3238 12186 3290
rect 12238 3238 12250 3290
rect 12302 3238 12314 3290
rect 12366 3238 23166 3290
rect 23218 3238 23230 3290
rect 23282 3238 23294 3290
rect 23346 3238 23358 3290
rect 23410 3238 23422 3290
rect 23474 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 34530 3290
rect 34582 3238 45382 3290
rect 45434 3238 45446 3290
rect 45498 3238 45510 3290
rect 45562 3238 45574 3290
rect 45626 3238 45638 3290
rect 45690 3238 45696 3290
rect 1104 3216 45696 3238
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 19242 3176 19248 3188
rect 13688 3148 19248 3176
rect 13688 3136 13694 3148
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 22925 3179 22983 3185
rect 22925 3145 22937 3179
rect 22971 3176 22983 3179
rect 39666 3176 39672 3188
rect 22971 3148 39672 3176
rect 22971 3145 22983 3148
rect 22925 3139 22983 3145
rect 39666 3136 39672 3148
rect 39724 3136 39730 3188
rect 12526 3068 12532 3120
rect 12584 3108 12590 3120
rect 29086 3108 29092 3120
rect 12584 3080 29092 3108
rect 12584 3068 12590 3080
rect 29086 3068 29092 3080
rect 29144 3068 29150 3120
rect 8202 3000 8208 3052
rect 8260 3040 8266 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 8260 3012 21833 3040
rect 8260 3000 8266 3012
rect 21821 3009 21833 3012
rect 21867 3009 21879 3043
rect 21821 3003 21879 3009
rect 22373 3043 22431 3049
rect 22373 3009 22385 3043
rect 22419 3009 22431 3043
rect 22373 3003 22431 3009
rect 22741 3043 22799 3049
rect 22741 3009 22753 3043
rect 22787 3009 22799 3043
rect 22741 3003 22799 3009
rect 23385 3043 23443 3049
rect 23385 3009 23397 3043
rect 23431 3040 23443 3043
rect 30098 3040 30104 3052
rect 23431 3012 30104 3040
rect 23431 3009 23443 3012
rect 23385 3003 23443 3009
rect 12986 2932 12992 2984
rect 13044 2972 13050 2984
rect 22388 2972 22416 3003
rect 13044 2944 22416 2972
rect 13044 2932 13050 2944
rect 14090 2864 14096 2916
rect 14148 2904 14154 2916
rect 22756 2904 22784 3003
rect 30098 3000 30104 3012
rect 30156 3000 30162 3052
rect 23474 2904 23480 2916
rect 14148 2876 22784 2904
rect 23124 2876 23480 2904
rect 14148 2864 14154 2876
rect 16850 2796 16856 2848
rect 16908 2836 16914 2848
rect 19426 2836 19432 2848
rect 16908 2808 19432 2836
rect 16908 2796 16914 2808
rect 19426 2796 19432 2808
rect 19484 2796 19490 2848
rect 22005 2839 22063 2845
rect 22005 2805 22017 2839
rect 22051 2836 22063 2839
rect 22278 2836 22284 2848
rect 22051 2808 22284 2836
rect 22051 2805 22063 2808
rect 22005 2799 22063 2805
rect 22278 2796 22284 2808
rect 22336 2796 22342 2848
rect 22557 2839 22615 2845
rect 22557 2805 22569 2839
rect 22603 2836 22615 2839
rect 23124 2836 23152 2876
rect 23474 2864 23480 2876
rect 23532 2864 23538 2916
rect 22603 2808 23152 2836
rect 22603 2805 22615 2808
rect 22557 2799 22615 2805
rect 23198 2796 23204 2848
rect 23256 2796 23262 2848
rect 30282 2796 30288 2848
rect 30340 2836 30346 2848
rect 32858 2836 32864 2848
rect 30340 2808 32864 2836
rect 30340 2796 30346 2808
rect 32858 2796 32864 2808
rect 32916 2796 32922 2848
rect 1104 2746 45540 2768
rect 1104 2694 6504 2746
rect 6556 2694 6568 2746
rect 6620 2694 6632 2746
rect 6684 2694 6696 2746
rect 6748 2694 6760 2746
rect 6812 2694 17612 2746
rect 17664 2694 17676 2746
rect 17728 2694 17740 2746
rect 17792 2694 17804 2746
rect 17856 2694 17868 2746
rect 17920 2694 28720 2746
rect 28772 2694 28784 2746
rect 28836 2694 28848 2746
rect 28900 2694 28912 2746
rect 28964 2694 28976 2746
rect 29028 2694 39828 2746
rect 39880 2694 39892 2746
rect 39944 2694 39956 2746
rect 40008 2694 40020 2746
rect 40072 2694 40084 2746
rect 40136 2694 45540 2746
rect 1104 2672 45540 2694
rect 17034 2592 17040 2644
rect 17092 2592 17098 2644
rect 19337 2635 19395 2641
rect 19337 2601 19349 2635
rect 19383 2632 19395 2635
rect 19518 2632 19524 2644
rect 19383 2604 19524 2632
rect 19383 2601 19395 2604
rect 19337 2595 19395 2601
rect 19518 2592 19524 2604
rect 19576 2592 19582 2644
rect 20622 2592 20628 2644
rect 20680 2592 20686 2644
rect 21450 2592 21456 2644
rect 21508 2632 21514 2644
rect 21545 2635 21603 2641
rect 21545 2632 21557 2635
rect 21508 2604 21557 2632
rect 21508 2592 21514 2604
rect 21545 2601 21557 2604
rect 21591 2601 21603 2635
rect 22002 2632 22008 2644
rect 21545 2595 21603 2601
rect 21652 2604 22008 2632
rect 17052 2536 17448 2564
rect 10962 2456 10968 2508
rect 11020 2496 11026 2508
rect 17052 2496 17080 2536
rect 11020 2468 17080 2496
rect 17420 2496 17448 2536
rect 18138 2524 18144 2576
rect 18196 2564 18202 2576
rect 21652 2564 21680 2604
rect 22002 2592 22008 2604
rect 22060 2592 22066 2644
rect 22370 2592 22376 2644
rect 22428 2592 22434 2644
rect 22738 2592 22744 2644
rect 22796 2632 22802 2644
rect 22925 2635 22983 2641
rect 22925 2632 22937 2635
rect 22796 2604 22937 2632
rect 22796 2592 22802 2604
rect 22925 2601 22937 2604
rect 22971 2601 22983 2635
rect 22925 2595 22983 2601
rect 23014 2592 23020 2644
rect 23072 2632 23078 2644
rect 23293 2635 23351 2641
rect 23293 2632 23305 2635
rect 23072 2604 23305 2632
rect 23072 2592 23078 2604
rect 23293 2601 23305 2604
rect 23339 2601 23351 2635
rect 23293 2595 23351 2601
rect 23400 2604 24072 2632
rect 18196 2536 21680 2564
rect 22833 2567 22891 2573
rect 18196 2524 18202 2536
rect 22833 2533 22845 2567
rect 22879 2564 22891 2567
rect 22879 2536 23060 2564
rect 22879 2533 22891 2536
rect 22833 2527 22891 2533
rect 17420 2468 19748 2496
rect 11020 2456 11026 2468
rect 19720 2440 19748 2468
rect 19794 2456 19800 2508
rect 19852 2496 19858 2508
rect 22186 2496 22192 2508
rect 19852 2468 22192 2496
rect 19852 2456 19858 2468
rect 22186 2456 22192 2468
rect 22244 2456 22250 2508
rect 22738 2496 22744 2508
rect 22480 2468 22744 2496
rect 17218 2388 17224 2440
rect 17276 2388 17282 2440
rect 18782 2388 18788 2440
rect 18840 2388 18846 2440
rect 19150 2388 19156 2440
rect 19208 2428 19214 2440
rect 19521 2431 19579 2437
rect 19521 2428 19533 2431
rect 19208 2400 19533 2428
rect 19208 2388 19214 2400
rect 19521 2397 19533 2400
rect 19567 2397 19579 2431
rect 19521 2391 19579 2397
rect 19610 2388 19616 2440
rect 19668 2388 19674 2440
rect 19702 2388 19708 2440
rect 19760 2388 19766 2440
rect 19886 2388 19892 2440
rect 19944 2388 19950 2440
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2428 20867 2431
rect 21269 2431 21327 2437
rect 20855 2400 21128 2428
rect 20855 2397 20867 2400
rect 20809 2391 20867 2397
rect 11238 2320 11244 2372
rect 11296 2360 11302 2372
rect 18046 2360 18052 2372
rect 11296 2332 18052 2360
rect 11296 2320 11302 2332
rect 18046 2320 18052 2332
rect 18104 2320 18110 2372
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 20364 2360 20392 2391
rect 18380 2332 20392 2360
rect 18380 2320 18386 2332
rect 15286 2252 15292 2304
rect 15344 2292 15350 2304
rect 18874 2292 18880 2304
rect 15344 2264 18880 2292
rect 15344 2252 15350 2264
rect 18874 2252 18880 2264
rect 18932 2252 18938 2304
rect 18966 2252 18972 2304
rect 19024 2252 19030 2304
rect 19797 2295 19855 2301
rect 19797 2261 19809 2295
rect 19843 2292 19855 2295
rect 19978 2292 19984 2304
rect 19843 2264 19984 2292
rect 19843 2261 19855 2264
rect 19797 2255 19855 2261
rect 19978 2252 19984 2264
rect 20036 2252 20042 2304
rect 20073 2295 20131 2301
rect 20073 2261 20085 2295
rect 20119 2292 20131 2295
rect 20162 2292 20168 2304
rect 20119 2264 20168 2292
rect 20119 2261 20131 2264
rect 20073 2255 20131 2261
rect 20162 2252 20168 2264
rect 20220 2252 20226 2304
rect 20533 2295 20591 2301
rect 20533 2261 20545 2295
rect 20579 2292 20591 2295
rect 20990 2292 20996 2304
rect 20579 2264 20996 2292
rect 20579 2261 20591 2264
rect 20533 2255 20591 2261
rect 20990 2252 20996 2264
rect 21048 2252 21054 2304
rect 21100 2301 21128 2400
rect 21269 2397 21281 2431
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 21284 2360 21312 2391
rect 21358 2388 21364 2440
rect 21416 2428 21422 2440
rect 21729 2431 21787 2437
rect 21729 2428 21741 2431
rect 21416 2400 21741 2428
rect 21416 2388 21422 2400
rect 21729 2397 21741 2400
rect 21775 2397 21787 2431
rect 21729 2391 21787 2397
rect 21818 2388 21824 2440
rect 21876 2388 21882 2440
rect 22094 2388 22100 2440
rect 22152 2388 22158 2440
rect 22480 2360 22508 2468
rect 22738 2456 22744 2468
rect 22796 2456 22802 2508
rect 23032 2496 23060 2536
rect 23106 2524 23112 2576
rect 23164 2564 23170 2576
rect 23400 2564 23428 2604
rect 23164 2536 23428 2564
rect 23164 2524 23170 2536
rect 23566 2524 23572 2576
rect 23624 2564 23630 2576
rect 23937 2567 23995 2573
rect 23937 2564 23949 2567
rect 23624 2536 23949 2564
rect 23624 2524 23630 2536
rect 23937 2533 23949 2536
rect 23983 2533 23995 2567
rect 24044 2564 24072 2604
rect 24394 2592 24400 2644
rect 24452 2592 24458 2644
rect 25866 2592 25872 2644
rect 25924 2632 25930 2644
rect 25961 2635 26019 2641
rect 25961 2632 25973 2635
rect 25924 2604 25973 2632
rect 25924 2592 25930 2604
rect 25961 2601 25973 2604
rect 26007 2601 26019 2635
rect 25961 2595 26019 2601
rect 28074 2592 28080 2644
rect 28132 2632 28138 2644
rect 28169 2635 28227 2641
rect 28169 2632 28181 2635
rect 28132 2604 28181 2632
rect 28132 2592 28138 2604
rect 28169 2601 28181 2604
rect 28215 2601 28227 2635
rect 28169 2595 28227 2601
rect 29178 2592 29184 2644
rect 29236 2592 29242 2644
rect 30374 2592 30380 2644
rect 30432 2592 30438 2644
rect 30466 2592 30472 2644
rect 30524 2632 30530 2644
rect 30524 2604 31432 2632
rect 30524 2592 30530 2604
rect 27890 2564 27896 2576
rect 24044 2536 27896 2564
rect 23937 2527 23995 2533
rect 27890 2524 27896 2536
rect 27948 2524 27954 2576
rect 27985 2567 28043 2573
rect 27985 2533 27997 2567
rect 28031 2564 28043 2567
rect 30282 2564 30288 2576
rect 28031 2536 30288 2564
rect 28031 2533 28043 2536
rect 27985 2527 28043 2533
rect 30282 2524 30288 2536
rect 30340 2524 30346 2576
rect 31404 2564 31432 2604
rect 32490 2592 32496 2644
rect 32548 2632 32554 2644
rect 32585 2635 32643 2641
rect 32585 2632 32597 2635
rect 32548 2604 32597 2632
rect 32548 2592 32554 2604
rect 32585 2601 32597 2604
rect 32631 2601 32643 2635
rect 32585 2595 32643 2601
rect 34790 2592 34796 2644
rect 34848 2592 34854 2644
rect 34900 2604 36860 2632
rect 34900 2564 34928 2604
rect 31404 2536 34928 2564
rect 35066 2524 35072 2576
rect 35124 2564 35130 2576
rect 36832 2564 36860 2604
rect 36906 2592 36912 2644
rect 36964 2632 36970 2644
rect 37001 2635 37059 2641
rect 37001 2632 37013 2635
rect 36964 2604 37013 2632
rect 36964 2592 36970 2604
rect 37001 2601 37013 2604
rect 37047 2601 37059 2635
rect 37001 2595 37059 2601
rect 39022 2592 39028 2644
rect 39080 2632 39086 2644
rect 39117 2635 39175 2641
rect 39117 2632 39129 2635
rect 39080 2604 39129 2632
rect 39080 2592 39086 2604
rect 39117 2601 39129 2604
rect 39163 2601 39175 2635
rect 39117 2595 39175 2601
rect 41322 2592 41328 2644
rect 41380 2592 41386 2644
rect 43530 2592 43536 2644
rect 43588 2632 43594 2644
rect 43809 2635 43867 2641
rect 43809 2632 43821 2635
rect 43588 2604 43821 2632
rect 43588 2592 43594 2604
rect 43809 2601 43821 2604
rect 43855 2601 43867 2635
rect 43809 2595 43867 2601
rect 44542 2592 44548 2644
rect 44600 2592 44606 2644
rect 40402 2564 40408 2576
rect 35124 2536 36768 2564
rect 36832 2536 40408 2564
rect 35124 2524 35130 2536
rect 23032 2468 23520 2496
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2397 22615 2431
rect 22557 2391 22615 2397
rect 21284 2332 22508 2360
rect 21085 2295 21143 2301
rect 21085 2261 21097 2295
rect 21131 2261 21143 2295
rect 21085 2255 21143 2261
rect 22005 2295 22063 2301
rect 22005 2261 22017 2295
rect 22051 2292 22063 2295
rect 22186 2292 22192 2304
rect 22051 2264 22192 2292
rect 22051 2261 22063 2264
rect 22005 2255 22063 2261
rect 22186 2252 22192 2264
rect 22244 2252 22250 2304
rect 22278 2252 22284 2304
rect 22336 2252 22342 2304
rect 22572 2292 22600 2391
rect 22646 2388 22652 2440
rect 22704 2388 22710 2440
rect 23106 2388 23112 2440
rect 23164 2437 23170 2440
rect 23492 2437 23520 2468
rect 25774 2456 25780 2508
rect 25832 2496 25838 2508
rect 30466 2496 30472 2508
rect 25832 2468 30472 2496
rect 25832 2456 25838 2468
rect 30466 2456 30472 2468
rect 30524 2456 30530 2508
rect 32122 2496 32128 2508
rect 30576 2468 32128 2496
rect 23164 2391 23175 2437
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23842 2428 23848 2440
rect 23477 2391 23535 2397
rect 23676 2400 23848 2428
rect 23164 2388 23170 2391
rect 23198 2292 23204 2304
rect 22572 2264 23204 2292
rect 23198 2252 23204 2264
rect 23256 2252 23262 2304
rect 23676 2301 23704 2400
rect 23842 2388 23848 2400
rect 23900 2388 23906 2440
rect 24118 2388 24124 2440
rect 24176 2388 24182 2440
rect 24578 2388 24584 2440
rect 24636 2388 24642 2440
rect 26142 2388 26148 2440
rect 26200 2388 26206 2440
rect 27798 2388 27804 2440
rect 27856 2388 27862 2440
rect 28353 2431 28411 2437
rect 28353 2397 28365 2431
rect 28399 2428 28411 2431
rect 29178 2428 29184 2440
rect 28399 2400 29184 2428
rect 28399 2397 28411 2400
rect 28353 2391 28411 2397
rect 29178 2388 29184 2400
rect 29236 2388 29242 2440
rect 30576 2437 30604 2468
rect 32122 2456 32128 2468
rect 32180 2456 32186 2508
rect 36630 2496 36636 2508
rect 32324 2468 36636 2496
rect 32324 2440 32352 2468
rect 36630 2456 36636 2468
rect 36688 2456 36694 2508
rect 36740 2496 36768 2536
rect 40402 2524 40408 2536
rect 40460 2524 40466 2576
rect 40678 2496 40684 2508
rect 36740 2468 40684 2496
rect 40678 2456 40684 2468
rect 40736 2456 40742 2508
rect 29365 2431 29423 2437
rect 29365 2397 29377 2431
rect 29411 2397 29423 2431
rect 29365 2391 29423 2397
rect 30561 2431 30619 2437
rect 30561 2397 30573 2431
rect 30607 2397 30619 2431
rect 30561 2391 30619 2397
rect 23750 2320 23756 2372
rect 23808 2320 23814 2372
rect 24210 2320 24216 2372
rect 24268 2360 24274 2372
rect 29270 2360 29276 2372
rect 24268 2332 29276 2360
rect 24268 2320 24274 2332
rect 29270 2320 29276 2332
rect 29328 2320 29334 2372
rect 29380 2360 29408 2391
rect 30650 2388 30656 2440
rect 30708 2388 30714 2440
rect 30926 2388 30932 2440
rect 30984 2388 30990 2440
rect 31202 2388 31208 2440
rect 31260 2388 31266 2440
rect 32306 2388 32312 2440
rect 32364 2388 32370 2440
rect 32766 2388 32772 2440
rect 32824 2388 32830 2440
rect 34974 2388 34980 2440
rect 35032 2388 35038 2440
rect 37182 2388 37188 2440
rect 37240 2388 37246 2440
rect 39298 2388 39304 2440
rect 39356 2388 39362 2440
rect 41506 2388 41512 2440
rect 41564 2388 41570 2440
rect 43990 2388 43996 2440
rect 44048 2388 44054 2440
rect 44358 2388 44364 2440
rect 44416 2388 44422 2440
rect 44821 2431 44879 2437
rect 44821 2397 44833 2431
rect 44867 2428 44879 2431
rect 45094 2428 45100 2440
rect 44867 2400 45100 2428
rect 44867 2397 44879 2400
rect 44821 2391 44879 2397
rect 45094 2388 45100 2400
rect 45152 2388 45158 2440
rect 45189 2431 45247 2437
rect 45189 2397 45201 2431
rect 45235 2428 45247 2431
rect 46106 2428 46112 2440
rect 45235 2400 46112 2428
rect 45235 2397 45247 2400
rect 45189 2391 45247 2397
rect 46106 2388 46112 2400
rect 46164 2388 46170 2440
rect 43530 2360 43536 2372
rect 29380 2332 43536 2360
rect 43530 2320 43536 2332
rect 43588 2320 43594 2372
rect 23661 2295 23719 2301
rect 23661 2261 23673 2295
rect 23707 2261 23719 2295
rect 23661 2255 23719 2261
rect 24026 2252 24032 2304
rect 24084 2292 24090 2304
rect 30558 2292 30564 2304
rect 24084 2264 30564 2292
rect 24084 2252 24090 2264
rect 30558 2252 30564 2264
rect 30616 2252 30622 2304
rect 30834 2252 30840 2304
rect 30892 2252 30898 2304
rect 31110 2252 31116 2304
rect 31168 2252 31174 2304
rect 31389 2295 31447 2301
rect 31389 2261 31401 2295
rect 31435 2292 31447 2295
rect 31938 2292 31944 2304
rect 31435 2264 31944 2292
rect 31435 2261 31447 2264
rect 31389 2255 31447 2261
rect 31938 2252 31944 2264
rect 31996 2252 32002 2304
rect 32030 2252 32036 2304
rect 32088 2292 32094 2304
rect 35066 2292 35072 2304
rect 32088 2264 35072 2292
rect 32088 2252 32094 2264
rect 35066 2252 35072 2264
rect 35124 2252 35130 2304
rect 35342 2252 35348 2304
rect 35400 2292 35406 2304
rect 44174 2292 44180 2304
rect 35400 2264 44180 2292
rect 35400 2252 35406 2264
rect 44174 2252 44180 2264
rect 44232 2252 44238 2304
rect 44634 2252 44640 2304
rect 44692 2252 44698 2304
rect 45002 2252 45008 2304
rect 45060 2252 45066 2304
rect 1104 2202 45696 2224
rect 1104 2150 12058 2202
rect 12110 2150 12122 2202
rect 12174 2150 12186 2202
rect 12238 2150 12250 2202
rect 12302 2150 12314 2202
rect 12366 2150 23166 2202
rect 23218 2150 23230 2202
rect 23282 2150 23294 2202
rect 23346 2150 23358 2202
rect 23410 2150 23422 2202
rect 23474 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 34530 2202
rect 34582 2150 45382 2202
rect 45434 2150 45446 2202
rect 45498 2150 45510 2202
rect 45562 2150 45574 2202
rect 45626 2150 45638 2202
rect 45690 2150 45696 2202
rect 1104 2128 45696 2150
rect 3329 2091 3387 2097
rect 3329 2057 3341 2091
rect 3375 2057 3387 2091
rect 3329 2051 3387 2057
rect 474 1912 480 1964
rect 532 1952 538 1964
rect 1397 1955 1455 1961
rect 1397 1952 1409 1955
rect 532 1924 1409 1952
rect 532 1912 538 1924
rect 1397 1921 1409 1924
rect 1443 1921 1455 1955
rect 1397 1915 1455 1921
rect 1673 1955 1731 1961
rect 1673 1921 1685 1955
rect 1719 1921 1731 1955
rect 1673 1915 1731 1921
rect 842 1844 848 1896
rect 900 1884 906 1896
rect 1688 1884 1716 1915
rect 2314 1912 2320 1964
rect 2372 1912 2378 1964
rect 3142 1912 3148 1964
rect 3200 1912 3206 1964
rect 900 1856 1716 1884
rect 900 1844 906 1856
rect 2038 1844 2044 1896
rect 2096 1844 2102 1896
rect 3344 1884 3372 2051
rect 13814 2048 13820 2100
rect 13872 2088 13878 2100
rect 15381 2091 15439 2097
rect 15381 2088 15393 2091
rect 13872 2060 15393 2088
rect 13872 2048 13878 2060
rect 15381 2057 15393 2060
rect 15427 2057 15439 2091
rect 15381 2051 15439 2057
rect 15856 2060 16068 2088
rect 7558 1980 7564 2032
rect 7616 2020 7622 2032
rect 15856 2020 15884 2060
rect 7616 1992 15884 2020
rect 16040 2020 16068 2060
rect 16206 2048 16212 2100
rect 16264 2048 16270 2100
rect 16482 2048 16488 2100
rect 16540 2048 16546 2100
rect 17037 2091 17095 2097
rect 17037 2057 17049 2091
rect 17083 2088 17095 2091
rect 17126 2088 17132 2100
rect 17083 2060 17132 2088
rect 17083 2057 17095 2060
rect 17037 2051 17095 2057
rect 17126 2048 17132 2060
rect 17184 2048 17190 2100
rect 17494 2048 17500 2100
rect 17552 2088 17558 2100
rect 17589 2091 17647 2097
rect 17589 2088 17601 2091
rect 17552 2060 17601 2088
rect 17552 2048 17558 2060
rect 17589 2057 17601 2060
rect 17635 2057 17647 2091
rect 17589 2051 17647 2057
rect 18138 2048 18144 2100
rect 18196 2048 18202 2100
rect 18693 2091 18751 2097
rect 18693 2057 18705 2091
rect 18739 2088 18751 2091
rect 19150 2088 19156 2100
rect 18739 2060 19156 2088
rect 18739 2057 18751 2060
rect 18693 2051 18751 2057
rect 19150 2048 19156 2060
rect 19208 2048 19214 2100
rect 19242 2048 19248 2100
rect 19300 2048 19306 2100
rect 19794 2048 19800 2100
rect 19852 2048 19858 2100
rect 20073 2091 20131 2097
rect 20073 2057 20085 2091
rect 20119 2088 20131 2091
rect 20806 2088 20812 2100
rect 20119 2060 20812 2088
rect 20119 2057 20131 2060
rect 20073 2051 20131 2057
rect 20806 2048 20812 2060
rect 20864 2048 20870 2100
rect 20898 2048 20904 2100
rect 20956 2048 20962 2100
rect 20990 2048 20996 2100
rect 21048 2088 21054 2100
rect 23106 2088 23112 2100
rect 21048 2060 22048 2088
rect 21048 2048 21054 2060
rect 17862 2020 17868 2032
rect 16040 1992 17868 2020
rect 7616 1980 7622 1992
rect 17862 1980 17868 1992
rect 17920 1980 17926 2032
rect 18046 1980 18052 2032
rect 18104 2020 18110 2032
rect 19812 2020 19840 2048
rect 22020 2029 22048 2060
rect 22204 2060 23112 2088
rect 22204 2032 22232 2060
rect 23106 2048 23112 2060
rect 23164 2048 23170 2100
rect 23477 2091 23535 2097
rect 23477 2057 23489 2091
rect 23523 2057 23535 2091
rect 23477 2051 23535 2057
rect 18104 1992 19196 2020
rect 18104 1980 18110 1992
rect 15010 1912 15016 1964
rect 15068 1912 15074 1964
rect 15473 1955 15531 1961
rect 15473 1921 15485 1955
rect 15519 1952 15531 1955
rect 15654 1952 15660 1964
rect 15519 1924 15660 1952
rect 15519 1921 15531 1924
rect 15473 1915 15531 1921
rect 15654 1912 15660 1924
rect 15712 1912 15718 1964
rect 15749 1955 15807 1961
rect 15749 1921 15761 1955
rect 15795 1921 15807 1955
rect 15749 1915 15807 1921
rect 14826 1884 14832 1896
rect 3344 1856 14832 1884
rect 14826 1844 14832 1856
rect 14884 1844 14890 1896
rect 15102 1844 15108 1896
rect 15160 1884 15166 1896
rect 15764 1884 15792 1915
rect 16022 1912 16028 1964
rect 16080 1912 16086 1964
rect 16298 1912 16304 1964
rect 16356 1912 16362 1964
rect 16482 1912 16488 1964
rect 16540 1952 16546 1964
rect 16853 1955 16911 1961
rect 16853 1952 16865 1955
rect 16540 1924 16865 1952
rect 16540 1912 16546 1924
rect 16853 1921 16865 1924
rect 16899 1921 16911 1955
rect 16853 1915 16911 1921
rect 17126 1912 17132 1964
rect 17184 1912 17190 1964
rect 17402 1912 17408 1964
rect 17460 1912 17466 1964
rect 17494 1912 17500 1964
rect 17552 1952 17558 1964
rect 17681 1955 17739 1961
rect 17681 1952 17693 1955
rect 17552 1924 17693 1952
rect 17552 1912 17558 1924
rect 17681 1921 17693 1924
rect 17727 1921 17739 1955
rect 17681 1915 17739 1921
rect 17957 1955 18015 1961
rect 17957 1921 17969 1955
rect 18003 1952 18015 1955
rect 18138 1952 18144 1964
rect 18003 1924 18144 1952
rect 18003 1921 18015 1924
rect 17957 1915 18015 1921
rect 18138 1912 18144 1924
rect 18196 1912 18202 1964
rect 18233 1955 18291 1961
rect 18233 1921 18245 1955
rect 18279 1952 18291 1955
rect 18414 1952 18420 1964
rect 18279 1924 18420 1952
rect 18279 1921 18291 1924
rect 18233 1915 18291 1921
rect 18414 1912 18420 1924
rect 18472 1912 18478 1964
rect 18506 1912 18512 1964
rect 18564 1912 18570 1964
rect 18690 1912 18696 1964
rect 18748 1912 18754 1964
rect 18782 1912 18788 1964
rect 18840 1912 18846 1964
rect 18874 1912 18880 1964
rect 18932 1952 18938 1964
rect 19061 1955 19119 1961
rect 19061 1952 19073 1955
rect 18932 1924 19073 1952
rect 18932 1912 18938 1924
rect 19061 1921 19073 1924
rect 19107 1921 19119 1955
rect 19168 1952 19196 1992
rect 19444 1992 19840 2020
rect 22005 2023 22063 2029
rect 19329 1959 19387 1965
rect 19329 1956 19341 1959
rect 19260 1952 19341 1956
rect 19168 1928 19341 1952
rect 19168 1924 19288 1928
rect 19329 1925 19341 1928
rect 19375 1925 19387 1959
rect 19061 1915 19119 1921
rect 19329 1919 19387 1925
rect 18708 1884 18736 1912
rect 19444 1884 19472 1992
rect 22005 1989 22017 2023
rect 22051 1989 22063 2023
rect 22005 1983 22063 1989
rect 22186 1980 22192 2032
rect 22244 1980 22250 2032
rect 23492 2020 23520 2051
rect 23750 2048 23756 2100
rect 23808 2088 23814 2100
rect 24029 2091 24087 2097
rect 24029 2088 24041 2091
rect 23808 2060 24041 2088
rect 23808 2048 23814 2060
rect 24029 2057 24041 2060
rect 24075 2057 24087 2091
rect 24029 2051 24087 2057
rect 24118 2048 24124 2100
rect 24176 2088 24182 2100
rect 24949 2091 25007 2097
rect 24949 2088 24961 2091
rect 24176 2060 24961 2088
rect 24176 2048 24182 2060
rect 24949 2057 24961 2060
rect 24995 2057 25007 2091
rect 24949 2051 25007 2057
rect 26142 2048 26148 2100
rect 26200 2088 26206 2100
rect 27249 2091 27307 2097
rect 27249 2088 27261 2091
rect 26200 2060 27261 2088
rect 26200 2048 26206 2060
rect 27249 2057 27261 2060
rect 27295 2057 27307 2091
rect 27249 2051 27307 2057
rect 28261 2091 28319 2097
rect 28261 2057 28273 2091
rect 28307 2088 28319 2091
rect 28307 2060 28396 2088
rect 28307 2057 28319 2060
rect 28261 2051 28319 2057
rect 24578 2020 24584 2032
rect 23492 1992 24584 2020
rect 24578 1980 24584 1992
rect 24636 1980 24642 2032
rect 24854 1980 24860 2032
rect 24912 2020 24918 2032
rect 24912 1992 25268 2020
rect 24912 1980 24918 1992
rect 19518 1912 19524 1964
rect 19576 1952 19582 1964
rect 19613 1955 19671 1961
rect 19613 1952 19625 1955
rect 19576 1924 19625 1952
rect 19576 1912 19582 1924
rect 19613 1921 19625 1924
rect 19659 1921 19671 1955
rect 19613 1915 19671 1921
rect 19702 1912 19708 1964
rect 19760 1952 19766 1964
rect 19889 1955 19947 1961
rect 19889 1952 19901 1955
rect 19760 1924 19901 1952
rect 19760 1912 19766 1924
rect 19889 1921 19901 1924
rect 19935 1921 19947 1955
rect 19889 1915 19947 1921
rect 20165 1955 20223 1961
rect 20165 1921 20177 1955
rect 20211 1952 20223 1955
rect 20254 1952 20260 1964
rect 20211 1924 20260 1952
rect 20211 1921 20223 1924
rect 20165 1915 20223 1921
rect 20254 1912 20260 1924
rect 20312 1912 20318 1964
rect 20438 1912 20444 1964
rect 20496 1912 20502 1964
rect 20714 1912 20720 1964
rect 20772 1912 20778 1964
rect 20993 1955 21051 1961
rect 20993 1952 21005 1955
rect 20916 1924 21005 1952
rect 20916 1884 20944 1924
rect 20993 1921 21005 1924
rect 21039 1921 21051 1955
rect 20993 1915 21051 1921
rect 21453 1955 21511 1961
rect 21453 1921 21465 1955
rect 21499 1952 21511 1955
rect 21542 1952 21548 1964
rect 21499 1924 21548 1952
rect 21499 1921 21511 1924
rect 21453 1915 21511 1921
rect 21542 1912 21548 1924
rect 21600 1912 21606 1964
rect 22462 1912 22468 1964
rect 22520 1912 22526 1964
rect 22554 1912 22560 1964
rect 22612 1952 22618 1964
rect 23017 1955 23075 1961
rect 23017 1952 23029 1955
rect 22612 1924 23029 1952
rect 22612 1912 22618 1924
rect 23017 1921 23029 1924
rect 23063 1921 23075 1955
rect 23017 1915 23075 1921
rect 23293 1955 23351 1961
rect 23293 1921 23305 1955
rect 23339 1921 23351 1955
rect 23293 1915 23351 1921
rect 15160 1856 15792 1884
rect 17236 1856 18736 1884
rect 18892 1856 19472 1884
rect 19536 1856 20944 1884
rect 23308 1884 23336 1915
rect 23566 1912 23572 1964
rect 23624 1912 23630 1964
rect 24213 1955 24271 1961
rect 24213 1921 24225 1955
rect 24259 1921 24271 1955
rect 24213 1915 24271 1921
rect 24026 1884 24032 1896
rect 23308 1856 24032 1884
rect 15160 1844 15166 1856
rect 1857 1819 1915 1825
rect 1857 1785 1869 1819
rect 1903 1816 1915 1819
rect 16850 1816 16856 1828
rect 1903 1788 16856 1816
rect 1903 1785 1915 1788
rect 1857 1779 1915 1785
rect 16850 1776 16856 1788
rect 16908 1776 16914 1828
rect 1578 1708 1584 1760
rect 1636 1708 1642 1760
rect 15194 1708 15200 1760
rect 15252 1708 15258 1760
rect 15933 1751 15991 1757
rect 15933 1717 15945 1751
rect 15979 1748 15991 1751
rect 17236 1748 17264 1856
rect 17313 1819 17371 1825
rect 17313 1785 17325 1819
rect 17359 1816 17371 1819
rect 18892 1816 18920 1856
rect 19536 1825 19564 1856
rect 24026 1844 24032 1856
rect 24084 1844 24090 1896
rect 24228 1884 24256 1915
rect 24302 1912 24308 1964
rect 24360 1912 24366 1964
rect 24670 1912 24676 1964
rect 24728 1912 24734 1964
rect 25130 1912 25136 1964
rect 25188 1912 25194 1964
rect 25240 1961 25268 1992
rect 25332 1992 28028 2020
rect 25225 1955 25283 1961
rect 25225 1921 25237 1955
rect 25271 1921 25283 1955
rect 25225 1915 25283 1921
rect 25332 1884 25360 1992
rect 25498 1912 25504 1964
rect 25556 1912 25562 1964
rect 25961 1955 26019 1961
rect 25961 1921 25973 1955
rect 26007 1921 26019 1955
rect 25961 1915 26019 1921
rect 25976 1884 26004 1915
rect 26326 1912 26332 1964
rect 26384 1912 26390 1964
rect 26602 1912 26608 1964
rect 26660 1912 26666 1964
rect 26694 1912 26700 1964
rect 26752 1952 26758 1964
rect 26973 1955 27031 1961
rect 26973 1952 26985 1955
rect 26752 1924 26985 1952
rect 26752 1912 26758 1924
rect 26973 1921 26985 1924
rect 27019 1921 27031 1955
rect 26973 1915 27031 1921
rect 27062 1912 27068 1964
rect 27120 1952 27126 1964
rect 27409 1955 27467 1961
rect 27409 1952 27421 1955
rect 27120 1924 27421 1952
rect 27120 1912 27126 1924
rect 27409 1921 27421 1924
rect 27455 1921 27467 1955
rect 27409 1915 27467 1921
rect 27525 1955 27583 1961
rect 27525 1921 27537 1955
rect 27571 1921 27583 1955
rect 27525 1915 27583 1921
rect 27540 1884 27568 1915
rect 27614 1912 27620 1964
rect 27672 1952 27678 1964
rect 27801 1955 27859 1961
rect 27801 1952 27813 1955
rect 27672 1924 27813 1952
rect 27672 1912 27678 1924
rect 27801 1921 27813 1924
rect 27847 1921 27859 1955
rect 27801 1915 27859 1921
rect 24228 1856 25360 1884
rect 25424 1856 26004 1884
rect 26068 1856 27568 1884
rect 28000 1884 28028 1992
rect 28077 1955 28135 1961
rect 28077 1921 28089 1955
rect 28123 1952 28135 1955
rect 28166 1952 28172 1964
rect 28123 1924 28172 1952
rect 28123 1921 28135 1924
rect 28077 1915 28135 1921
rect 28166 1912 28172 1924
rect 28224 1912 28230 1964
rect 28368 1952 28396 2060
rect 28442 2048 28448 2100
rect 28500 2088 28506 2100
rect 28500 2060 30328 2088
rect 28500 2048 28506 2060
rect 28736 1992 28948 2020
rect 28445 1955 28503 1961
rect 28445 1952 28457 1955
rect 28368 1924 28457 1952
rect 28445 1921 28457 1924
rect 28491 1921 28503 1955
rect 28445 1915 28503 1921
rect 28736 1884 28764 1992
rect 28813 1955 28871 1961
rect 28813 1921 28825 1955
rect 28859 1921 28871 1955
rect 28813 1915 28871 1921
rect 28000 1856 28764 1884
rect 17359 1788 18920 1816
rect 18969 1819 19027 1825
rect 17359 1785 17371 1788
rect 17313 1779 17371 1785
rect 18969 1785 18981 1819
rect 19015 1785 19027 1819
rect 18969 1779 19027 1785
rect 19521 1819 19579 1825
rect 19521 1785 19533 1819
rect 19567 1785 19579 1819
rect 19521 1779 19579 1785
rect 20625 1819 20683 1825
rect 20625 1785 20637 1819
rect 20671 1816 20683 1819
rect 20990 1816 20996 1828
rect 20671 1788 20996 1816
rect 20671 1785 20683 1788
rect 20625 1779 20683 1785
rect 15979 1720 17264 1748
rect 17865 1751 17923 1757
rect 15979 1717 15991 1720
rect 15933 1711 15991 1717
rect 17865 1717 17877 1751
rect 17911 1748 17923 1751
rect 18046 1748 18052 1760
rect 17911 1720 18052 1748
rect 17911 1717 17923 1720
rect 17865 1711 17923 1717
rect 18046 1708 18052 1720
rect 18104 1708 18110 1760
rect 18417 1751 18475 1757
rect 18417 1717 18429 1751
rect 18463 1748 18475 1751
rect 18690 1748 18696 1760
rect 18463 1720 18696 1748
rect 18463 1717 18475 1720
rect 18417 1711 18475 1717
rect 18690 1708 18696 1720
rect 18748 1708 18754 1760
rect 18984 1748 19012 1779
rect 20990 1776 20996 1788
rect 21048 1776 21054 1828
rect 21637 1819 21695 1825
rect 21637 1785 21649 1819
rect 21683 1785 21695 1819
rect 23014 1816 23020 1828
rect 21637 1779 21695 1785
rect 22020 1788 23020 1816
rect 19702 1748 19708 1760
rect 18984 1720 19708 1748
rect 19702 1708 19708 1720
rect 19760 1708 19766 1760
rect 19794 1708 19800 1760
rect 19852 1708 19858 1760
rect 20346 1708 20352 1760
rect 20404 1708 20410 1760
rect 21174 1708 21180 1760
rect 21232 1708 21238 1760
rect 21652 1748 21680 1779
rect 22020 1748 22048 1788
rect 23014 1776 23020 1788
rect 23072 1776 23078 1828
rect 23201 1819 23259 1825
rect 23201 1785 23213 1819
rect 23247 1816 23259 1819
rect 24946 1816 24952 1828
rect 23247 1788 24952 1816
rect 23247 1785 23259 1788
rect 23201 1779 23259 1785
rect 24946 1776 24952 1788
rect 25004 1776 25010 1828
rect 25424 1825 25452 1856
rect 25409 1819 25467 1825
rect 25409 1785 25421 1819
rect 25455 1785 25467 1819
rect 25409 1779 25467 1785
rect 25774 1776 25780 1828
rect 25832 1816 25838 1828
rect 26068 1816 26096 1856
rect 28828 1816 28856 1915
rect 28920 1884 28948 1992
rect 29086 1912 29092 1964
rect 29144 1912 29150 1964
rect 29362 1912 29368 1964
rect 29420 1912 29426 1964
rect 29638 1912 29644 1964
rect 29696 1912 29702 1964
rect 29822 1912 29828 1964
rect 29880 1952 29886 1964
rect 30300 1961 30328 2060
rect 30834 2048 30840 2100
rect 30892 2088 30898 2100
rect 30892 2060 31064 2088
rect 30892 2048 30898 2060
rect 29917 1955 29975 1961
rect 29917 1952 29929 1955
rect 29880 1924 29929 1952
rect 29880 1912 29886 1924
rect 29917 1921 29929 1924
rect 29963 1921 29975 1955
rect 29917 1915 29975 1921
rect 30285 1955 30343 1961
rect 30285 1921 30297 1955
rect 30331 1921 30343 1955
rect 30285 1915 30343 1921
rect 30558 1912 30564 1964
rect 30616 1912 30622 1964
rect 30834 1912 30840 1964
rect 30892 1912 30898 1964
rect 31036 1952 31064 2060
rect 31110 2048 31116 2100
rect 31168 2048 31174 2100
rect 31846 2048 31852 2100
rect 31904 2048 31910 2100
rect 32122 2048 32128 2100
rect 32180 2048 32186 2100
rect 32766 2048 32772 2100
rect 32824 2088 32830 2100
rect 33229 2091 33287 2097
rect 33229 2088 33241 2091
rect 32824 2060 33241 2088
rect 32824 2048 32830 2060
rect 33229 2057 33241 2060
rect 33275 2057 33287 2091
rect 33229 2051 33287 2057
rect 34974 2048 34980 2100
rect 35032 2088 35038 2100
rect 35161 2091 35219 2097
rect 35161 2088 35173 2091
rect 35032 2060 35173 2088
rect 35032 2048 35038 2060
rect 35161 2057 35173 2060
rect 35207 2057 35219 2091
rect 35161 2051 35219 2057
rect 35250 2048 35256 2100
rect 35308 2088 35314 2100
rect 35308 2060 36400 2088
rect 35308 2048 35314 2060
rect 31128 2020 31156 2048
rect 31205 2023 31263 2029
rect 31205 2020 31217 2023
rect 31128 1992 31217 2020
rect 31205 1989 31217 1992
rect 31251 1989 31263 2023
rect 36262 2020 36268 2032
rect 31205 1983 31263 1989
rect 33428 1992 36268 2020
rect 31665 1955 31723 1961
rect 31665 1952 31677 1955
rect 31036 1924 31677 1952
rect 31665 1921 31677 1924
rect 31711 1921 31723 1955
rect 31665 1915 31723 1921
rect 32306 1912 32312 1964
rect 32364 1912 32370 1964
rect 32858 1912 32864 1964
rect 32916 1912 32922 1964
rect 33428 1961 33456 1992
rect 36262 1980 36268 1992
rect 36320 1980 36326 2032
rect 36372 2029 36400 2060
rect 36630 2048 36636 2100
rect 36688 2048 36694 2100
rect 37182 2048 37188 2100
rect 37240 2088 37246 2100
rect 37369 2091 37427 2097
rect 37369 2088 37381 2091
rect 37240 2060 37381 2088
rect 37240 2048 37246 2060
rect 37369 2057 37381 2060
rect 37415 2057 37427 2091
rect 37369 2051 37427 2057
rect 39298 2048 39304 2100
rect 39356 2088 39362 2100
rect 39669 2091 39727 2097
rect 39669 2088 39681 2091
rect 39356 2060 39681 2088
rect 39356 2048 39362 2060
rect 39669 2057 39681 2060
rect 39715 2057 39727 2091
rect 39669 2051 39727 2057
rect 40126 2048 40132 2100
rect 40184 2048 40190 2100
rect 40402 2048 40408 2100
rect 40460 2048 40466 2100
rect 40678 2048 40684 2100
rect 40736 2048 40742 2100
rect 41506 2048 41512 2100
rect 41564 2088 41570 2100
rect 41785 2091 41843 2097
rect 41785 2088 41797 2091
rect 41564 2060 41797 2088
rect 41564 2048 41570 2060
rect 41785 2057 41797 2060
rect 41831 2057 41843 2091
rect 41785 2051 41843 2057
rect 43990 2048 43996 2100
rect 44048 2088 44054 2100
rect 44361 2091 44419 2097
rect 44361 2088 44373 2091
rect 44048 2060 44373 2088
rect 44048 2048 44054 2060
rect 44361 2057 44373 2060
rect 44407 2057 44419 2091
rect 44361 2051 44419 2057
rect 44634 2048 44640 2100
rect 44692 2048 44698 2100
rect 45002 2048 45008 2100
rect 45060 2048 45066 2100
rect 36357 2023 36415 2029
rect 36357 1989 36369 2023
rect 36403 1989 36415 2023
rect 36648 2020 36676 2048
rect 44652 2020 44680 2048
rect 36648 1992 39528 2020
rect 36357 1983 36415 1989
rect 33413 1955 33471 1961
rect 33413 1921 33425 1955
rect 33459 1921 33471 1955
rect 33413 1915 33471 1921
rect 33502 1912 33508 1964
rect 33560 1952 33566 1964
rect 33781 1955 33839 1961
rect 33781 1952 33793 1955
rect 33560 1924 33793 1952
rect 33560 1912 33566 1924
rect 33781 1921 33793 1924
rect 33827 1921 33839 1955
rect 33781 1915 33839 1921
rect 34054 1912 34060 1964
rect 34112 1952 34118 1964
rect 34241 1955 34299 1961
rect 34241 1952 34253 1955
rect 34112 1924 34253 1952
rect 34112 1912 34118 1924
rect 34241 1921 34253 1924
rect 34287 1921 34299 1955
rect 34241 1915 34299 1921
rect 34348 1924 35296 1952
rect 34348 1884 34376 1924
rect 28920 1856 34376 1884
rect 35268 1884 35296 1924
rect 35342 1912 35348 1964
rect 35400 1912 35406 1964
rect 35434 1912 35440 1964
rect 35492 1912 35498 1964
rect 37553 1955 37611 1961
rect 37553 1921 37565 1955
rect 37599 1952 37611 1955
rect 37918 1952 37924 1964
rect 37599 1924 37924 1952
rect 37599 1921 37611 1924
rect 37553 1915 37611 1921
rect 37918 1912 37924 1924
rect 37976 1912 37982 1964
rect 38010 1912 38016 1964
rect 38068 1912 38074 1964
rect 38378 1912 38384 1964
rect 38436 1912 38442 1964
rect 39206 1884 39212 1896
rect 35268 1856 39212 1884
rect 39206 1844 39212 1856
rect 39264 1844 39270 1896
rect 25832 1788 26096 1816
rect 27540 1788 28856 1816
rect 25832 1776 25838 1788
rect 21652 1720 22048 1748
rect 22094 1708 22100 1760
rect 22152 1708 22158 1760
rect 22646 1708 22652 1760
rect 22704 1708 22710 1760
rect 23750 1708 23756 1760
rect 23808 1708 23814 1760
rect 24486 1708 24492 1760
rect 24544 1708 24550 1760
rect 24854 1708 24860 1760
rect 24912 1708 24918 1760
rect 25685 1751 25743 1757
rect 25685 1717 25697 1751
rect 25731 1748 25743 1751
rect 26050 1748 26056 1760
rect 25731 1720 26056 1748
rect 25731 1717 25743 1720
rect 25685 1711 25743 1717
rect 26050 1708 26056 1720
rect 26108 1708 26114 1760
rect 26142 1708 26148 1760
rect 26200 1708 26206 1760
rect 26510 1708 26516 1760
rect 26568 1708 26574 1760
rect 26786 1708 26792 1760
rect 26844 1708 26850 1760
rect 27154 1708 27160 1760
rect 27212 1708 27218 1760
rect 27246 1708 27252 1760
rect 27304 1748 27310 1760
rect 27540 1748 27568 1788
rect 29086 1776 29092 1828
rect 29144 1816 29150 1828
rect 29144 1788 30144 1816
rect 29144 1776 29150 1788
rect 27304 1720 27568 1748
rect 27304 1708 27310 1720
rect 27706 1708 27712 1760
rect 27764 1708 27770 1760
rect 27982 1708 27988 1760
rect 28040 1708 28046 1760
rect 28074 1708 28080 1760
rect 28132 1748 28138 1760
rect 28629 1751 28687 1757
rect 28629 1748 28641 1751
rect 28132 1720 28641 1748
rect 28132 1708 28138 1720
rect 28629 1717 28641 1720
rect 28675 1717 28687 1751
rect 28629 1711 28687 1717
rect 28997 1751 29055 1757
rect 28997 1717 29009 1751
rect 29043 1748 29055 1751
rect 29178 1748 29184 1760
rect 29043 1720 29184 1748
rect 29043 1717 29055 1720
rect 28997 1711 29055 1717
rect 29178 1708 29184 1720
rect 29236 1708 29242 1760
rect 29270 1708 29276 1760
rect 29328 1708 29334 1760
rect 29546 1708 29552 1760
rect 29604 1708 29610 1760
rect 29822 1708 29828 1760
rect 29880 1708 29886 1760
rect 30116 1757 30144 1788
rect 30834 1776 30840 1828
rect 30892 1816 30898 1828
rect 31846 1816 31852 1828
rect 30892 1788 31852 1816
rect 30892 1776 30898 1788
rect 31846 1776 31852 1788
rect 31904 1776 31910 1828
rect 32324 1788 33180 1816
rect 30101 1751 30159 1757
rect 30101 1717 30113 1751
rect 30147 1717 30159 1751
rect 30101 1711 30159 1717
rect 30466 1708 30472 1760
rect 30524 1708 30530 1760
rect 30742 1708 30748 1760
rect 30800 1708 30806 1760
rect 31018 1708 31024 1760
rect 31076 1708 31082 1760
rect 31294 1708 31300 1760
rect 31352 1708 31358 1760
rect 31478 1708 31484 1760
rect 31536 1748 31542 1760
rect 32324 1748 32352 1788
rect 31536 1720 32352 1748
rect 31536 1708 31542 1720
rect 32398 1708 32404 1760
rect 32456 1748 32462 1760
rect 33045 1751 33103 1757
rect 33045 1748 33057 1751
rect 32456 1720 33057 1748
rect 32456 1708 32462 1720
rect 33045 1717 33057 1720
rect 33091 1717 33103 1751
rect 33152 1748 33180 1788
rect 33226 1776 33232 1828
rect 33284 1816 33290 1828
rect 33284 1788 34468 1816
rect 33284 1776 33290 1788
rect 33502 1748 33508 1760
rect 33152 1720 33508 1748
rect 33045 1711 33103 1717
rect 33502 1708 33508 1720
rect 33560 1708 33566 1760
rect 33870 1708 33876 1760
rect 33928 1708 33934 1760
rect 34440 1757 34468 1788
rect 37642 1776 37648 1828
rect 37700 1816 37706 1828
rect 37700 1788 38608 1816
rect 37700 1776 37706 1788
rect 34425 1751 34483 1757
rect 34425 1717 34437 1751
rect 34471 1717 34483 1751
rect 34425 1711 34483 1717
rect 34974 1708 34980 1760
rect 35032 1748 35038 1760
rect 35621 1751 35679 1757
rect 35621 1748 35633 1751
rect 35032 1720 35633 1748
rect 35032 1708 35038 1720
rect 35621 1717 35633 1720
rect 35667 1717 35679 1751
rect 35621 1711 35679 1717
rect 36446 1708 36452 1760
rect 36504 1708 36510 1760
rect 37550 1708 37556 1760
rect 37608 1748 37614 1760
rect 38580 1757 38608 1788
rect 38197 1751 38255 1757
rect 38197 1748 38209 1751
rect 37608 1720 38209 1748
rect 37608 1708 37614 1720
rect 38197 1717 38209 1720
rect 38243 1717 38255 1751
rect 38197 1711 38255 1717
rect 38565 1751 38623 1757
rect 38565 1717 38577 1751
rect 38611 1717 38623 1751
rect 39500 1748 39528 1992
rect 39868 1992 41920 2020
rect 39868 1961 39896 1992
rect 39853 1955 39911 1961
rect 39853 1921 39865 1955
rect 39899 1921 39911 1955
rect 40313 1955 40371 1961
rect 40313 1952 40325 1955
rect 39853 1915 39911 1921
rect 40052 1924 40325 1952
rect 39574 1844 39580 1896
rect 39632 1884 39638 1896
rect 40052 1884 40080 1924
rect 40313 1921 40325 1924
rect 40359 1921 40371 1955
rect 40313 1915 40371 1921
rect 40586 1912 40592 1964
rect 40644 1912 40650 1964
rect 40865 1955 40923 1961
rect 40865 1921 40877 1955
rect 40911 1921 40923 1955
rect 40865 1915 40923 1921
rect 39632 1856 40080 1884
rect 39632 1844 39638 1856
rect 40494 1776 40500 1828
rect 40552 1816 40558 1828
rect 40880 1816 40908 1915
rect 41892 1884 41920 1992
rect 41984 1992 44680 2020
rect 41984 1961 42012 1992
rect 41969 1955 42027 1961
rect 41969 1921 41981 1955
rect 42015 1921 42027 1955
rect 41969 1915 42027 1921
rect 44358 1912 44364 1964
rect 44416 1912 44422 1964
rect 44545 1955 44603 1961
rect 44545 1921 44557 1955
rect 44591 1921 44603 1955
rect 44545 1915 44603 1921
rect 44821 1955 44879 1961
rect 44821 1921 44833 1955
rect 44867 1952 44879 1955
rect 45020 1952 45048 2048
rect 44867 1924 45048 1952
rect 45189 1955 45247 1961
rect 44867 1921 44879 1924
rect 44821 1915 44879 1921
rect 45189 1921 45201 1955
rect 45235 1952 45247 1955
rect 45738 1952 45744 1964
rect 45235 1924 45744 1952
rect 45235 1921 45247 1924
rect 45189 1915 45247 1921
rect 42518 1884 42524 1896
rect 41892 1856 42524 1884
rect 42518 1844 42524 1856
rect 42576 1844 42582 1896
rect 40552 1788 40908 1816
rect 44376 1816 44404 1912
rect 44560 1884 44588 1915
rect 45738 1912 45744 1924
rect 45796 1912 45802 1964
rect 44560 1856 45048 1884
rect 45020 1825 45048 1856
rect 44637 1819 44695 1825
rect 44637 1816 44649 1819
rect 44376 1788 44649 1816
rect 40552 1776 40558 1788
rect 44637 1785 44649 1788
rect 44683 1785 44695 1819
rect 44637 1779 44695 1785
rect 45005 1819 45063 1825
rect 45005 1785 45017 1819
rect 45051 1785 45063 1819
rect 45005 1779 45063 1785
rect 43806 1748 43812 1760
rect 39500 1720 43812 1748
rect 38565 1711 38623 1717
rect 43806 1708 43812 1720
rect 43864 1708 43870 1760
rect 1104 1658 45540 1680
rect 1104 1606 6504 1658
rect 6556 1606 6568 1658
rect 6620 1606 6632 1658
rect 6684 1606 6696 1658
rect 6748 1606 6760 1658
rect 6812 1606 17612 1658
rect 17664 1606 17676 1658
rect 17728 1606 17740 1658
rect 17792 1606 17804 1658
rect 17856 1606 17868 1658
rect 17920 1606 28720 1658
rect 28772 1606 28784 1658
rect 28836 1606 28848 1658
rect 28900 1606 28912 1658
rect 28964 1606 28976 1658
rect 29028 1606 39828 1658
rect 39880 1606 39892 1658
rect 39944 1606 39956 1658
rect 40008 1606 40020 1658
rect 40072 1606 40084 1658
rect 40136 1606 45540 1658
rect 1104 1584 45540 1606
rect 1578 1504 1584 1556
rect 1636 1544 1642 1556
rect 7558 1544 7564 1556
rect 1636 1516 7564 1544
rect 1636 1504 1642 1516
rect 7558 1504 7564 1516
rect 7616 1504 7622 1556
rect 14553 1547 14611 1553
rect 14553 1513 14565 1547
rect 14599 1544 14611 1547
rect 15010 1544 15016 1556
rect 14599 1516 15016 1544
rect 14599 1513 14611 1516
rect 14553 1507 14611 1513
rect 15010 1504 15016 1516
rect 15068 1504 15074 1556
rect 15102 1504 15108 1556
rect 15160 1504 15166 1556
rect 15286 1504 15292 1556
rect 15344 1504 15350 1556
rect 15381 1547 15439 1553
rect 15381 1513 15393 1547
rect 15427 1544 15439 1547
rect 16022 1544 16028 1556
rect 15427 1516 16028 1544
rect 15427 1513 15439 1516
rect 15381 1507 15439 1513
rect 16022 1504 16028 1516
rect 16080 1504 16086 1556
rect 16298 1504 16304 1556
rect 16356 1504 16362 1556
rect 16482 1504 16488 1556
rect 16540 1504 16546 1556
rect 16945 1547 17003 1553
rect 16945 1513 16957 1547
rect 16991 1544 17003 1547
rect 17126 1544 17132 1556
rect 16991 1516 17132 1544
rect 16991 1513 17003 1516
rect 16945 1507 17003 1513
rect 17126 1504 17132 1516
rect 17184 1504 17190 1556
rect 17218 1504 17224 1556
rect 17276 1504 17282 1556
rect 17313 1547 17371 1553
rect 17313 1513 17325 1547
rect 17359 1544 17371 1547
rect 17402 1544 17408 1556
rect 17359 1516 17408 1544
rect 17359 1513 17371 1516
rect 17313 1507 17371 1513
rect 17402 1504 17408 1516
rect 17460 1504 17466 1556
rect 17494 1504 17500 1556
rect 17552 1544 17558 1556
rect 18049 1547 18107 1553
rect 18049 1544 18061 1547
rect 17552 1516 18061 1544
rect 17552 1504 17558 1516
rect 18049 1513 18061 1516
rect 18095 1513 18107 1547
rect 18049 1507 18107 1513
rect 18138 1504 18144 1556
rect 18196 1544 18202 1556
rect 18325 1547 18383 1553
rect 18325 1544 18337 1547
rect 18196 1516 18337 1544
rect 18196 1504 18202 1516
rect 18325 1513 18337 1516
rect 18371 1513 18383 1547
rect 18325 1507 18383 1513
rect 18414 1504 18420 1556
rect 18472 1544 18478 1556
rect 18601 1547 18659 1553
rect 18601 1544 18613 1547
rect 18472 1516 18613 1544
rect 18472 1504 18478 1516
rect 18601 1513 18613 1516
rect 18647 1513 18659 1547
rect 18601 1507 18659 1513
rect 18690 1504 18696 1556
rect 18748 1504 18754 1556
rect 18782 1504 18788 1556
rect 18840 1544 18846 1556
rect 18877 1547 18935 1553
rect 18877 1544 18889 1547
rect 18840 1516 18889 1544
rect 18840 1504 18846 1516
rect 18877 1513 18889 1516
rect 18923 1513 18935 1547
rect 18877 1507 18935 1513
rect 20272 1516 24716 1544
rect 1854 1436 1860 1488
rect 1912 1436 1918 1488
rect 14277 1479 14335 1485
rect 14277 1445 14289 1479
rect 14323 1476 14335 1479
rect 15304 1476 15332 1504
rect 14323 1448 15332 1476
rect 15657 1479 15715 1485
rect 14323 1445 14335 1448
rect 14277 1439 14335 1445
rect 15657 1445 15669 1479
rect 15703 1476 15715 1479
rect 16316 1476 16344 1504
rect 15703 1448 16344 1476
rect 17236 1476 17264 1504
rect 17589 1479 17647 1485
rect 17589 1476 17601 1479
rect 17236 1448 17601 1476
rect 15703 1445 15715 1448
rect 15657 1439 15715 1445
rect 17589 1445 17601 1448
rect 17635 1445 17647 1479
rect 18708 1476 18736 1504
rect 20272 1476 20300 1516
rect 18708 1448 20300 1476
rect 17589 1439 17647 1445
rect 20898 1436 20904 1488
rect 20956 1476 20962 1488
rect 20956 1448 22048 1476
rect 20956 1436 20962 1448
rect 3344 1380 4016 1408
rect 1210 1300 1216 1352
rect 1268 1340 1274 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 1268 1312 1409 1340
rect 1268 1300 1274 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 1670 1300 1676 1352
rect 1728 1300 1734 1352
rect 2133 1343 2191 1349
rect 2133 1309 2145 1343
rect 2179 1309 2191 1343
rect 2133 1303 2191 1309
rect 2148 1272 2176 1303
rect 2406 1300 2412 1352
rect 2464 1300 2470 1352
rect 2685 1343 2743 1349
rect 2685 1309 2697 1343
rect 2731 1309 2743 1343
rect 3344 1340 3372 1380
rect 2685 1303 2743 1309
rect 3160 1312 3372 1340
rect 2498 1272 2504 1284
rect 2148 1244 2504 1272
rect 2498 1232 2504 1244
rect 2556 1232 2562 1284
rect 2700 1272 2728 1303
rect 3160 1272 3188 1312
rect 3418 1300 3424 1352
rect 3476 1300 3482 1352
rect 3878 1300 3884 1352
rect 3936 1300 3942 1352
rect 3988 1272 4016 1380
rect 8036 1380 8248 1408
rect 4246 1300 4252 1352
rect 4304 1300 4310 1352
rect 4614 1300 4620 1352
rect 4672 1300 4678 1352
rect 4982 1300 4988 1352
rect 5040 1300 5046 1352
rect 5350 1300 5356 1352
rect 5408 1300 5414 1352
rect 5718 1300 5724 1352
rect 5776 1300 5782 1352
rect 5994 1300 6000 1352
rect 6052 1300 6058 1352
rect 6454 1300 6460 1352
rect 6512 1300 6518 1352
rect 6822 1300 6828 1352
rect 6880 1300 6886 1352
rect 7190 1300 7196 1352
rect 7248 1300 7254 1352
rect 7558 1300 7564 1352
rect 7616 1300 7622 1352
rect 7926 1300 7932 1352
rect 7984 1300 7990 1352
rect 4706 1272 4712 1284
rect 2700 1244 3188 1272
rect 3252 1244 3832 1272
rect 3988 1244 4712 1272
rect 1578 1164 1584 1216
rect 1636 1164 1642 1216
rect 2317 1207 2375 1213
rect 2317 1173 2329 1207
rect 2363 1204 2375 1207
rect 3252 1204 3280 1244
rect 3804 1216 3832 1244
rect 4706 1232 4712 1244
rect 4764 1232 4770 1284
rect 8036 1272 8064 1380
rect 8220 1352 8248 1380
rect 12084 1380 12480 1408
rect 8110 1300 8116 1352
rect 8168 1300 8174 1352
rect 8202 1300 8208 1352
rect 8260 1300 8266 1352
rect 8294 1300 8300 1352
rect 8352 1300 8358 1352
rect 8570 1300 8576 1352
rect 8628 1300 8634 1352
rect 9030 1300 9036 1352
rect 9088 1300 9094 1352
rect 9398 1300 9404 1352
rect 9456 1300 9462 1352
rect 9766 1300 9772 1352
rect 9824 1300 9830 1352
rect 10134 1300 10140 1352
rect 10192 1300 10198 1352
rect 10502 1300 10508 1352
rect 10560 1300 10566 1352
rect 10870 1300 10876 1352
rect 10928 1300 10934 1352
rect 11146 1300 11152 1352
rect 11204 1300 11210 1352
rect 11606 1300 11612 1352
rect 11664 1300 11670 1352
rect 11974 1300 11980 1352
rect 12032 1300 12038 1352
rect 4816 1244 6132 1272
rect 2363 1176 3280 1204
rect 2363 1173 2375 1176
rect 2317 1167 2375 1173
rect 3602 1164 3608 1216
rect 3660 1164 3666 1216
rect 3786 1164 3792 1216
rect 3844 1164 3850 1216
rect 4062 1164 4068 1216
rect 4120 1164 4126 1216
rect 4430 1164 4436 1216
rect 4488 1164 4494 1216
rect 4816 1213 4844 1244
rect 6104 1216 6132 1244
rect 6196 1244 8064 1272
rect 4801 1207 4859 1213
rect 4801 1173 4813 1207
rect 4847 1173 4859 1207
rect 4801 1167 4859 1173
rect 5166 1164 5172 1216
rect 5224 1164 5230 1216
rect 5537 1207 5595 1213
rect 5537 1173 5549 1207
rect 5583 1204 5595 1207
rect 5810 1204 5816 1216
rect 5583 1176 5816 1204
rect 5583 1173 5595 1176
rect 5537 1167 5595 1173
rect 5810 1164 5816 1176
rect 5868 1164 5874 1216
rect 5902 1164 5908 1216
rect 5960 1164 5966 1216
rect 6086 1164 6092 1216
rect 6144 1164 6150 1216
rect 6196 1213 6224 1244
rect 6181 1207 6239 1213
rect 6181 1173 6193 1207
rect 6227 1173 6239 1207
rect 6181 1167 6239 1173
rect 6638 1164 6644 1216
rect 6696 1164 6702 1216
rect 7006 1164 7012 1216
rect 7064 1164 7070 1216
rect 7377 1207 7435 1213
rect 7377 1173 7389 1207
rect 7423 1204 7435 1207
rect 7650 1204 7656 1216
rect 7423 1176 7656 1204
rect 7423 1173 7435 1176
rect 7377 1167 7435 1173
rect 7650 1164 7656 1176
rect 7708 1164 7714 1216
rect 7742 1164 7748 1216
rect 7800 1164 7806 1216
rect 8128 1213 8156 1300
rect 10410 1272 10416 1284
rect 8496 1244 10416 1272
rect 8496 1213 8524 1244
rect 10410 1232 10416 1244
rect 10468 1232 10474 1284
rect 12084 1272 12112 1380
rect 12158 1300 12164 1352
rect 12216 1340 12222 1352
rect 12345 1343 12403 1349
rect 12345 1340 12357 1343
rect 12216 1312 12357 1340
rect 12216 1300 12222 1312
rect 12345 1309 12357 1312
rect 12391 1309 12403 1343
rect 12452 1340 12480 1380
rect 13648 1380 13860 1408
rect 12526 1340 12532 1352
rect 12452 1312 12532 1340
rect 12345 1303 12403 1309
rect 12526 1300 12532 1312
rect 12584 1300 12590 1352
rect 12618 1300 12624 1352
rect 12676 1300 12682 1352
rect 12894 1300 12900 1352
rect 12952 1300 12958 1352
rect 13170 1300 13176 1352
rect 13228 1300 13234 1352
rect 13446 1300 13452 1352
rect 13504 1300 13510 1352
rect 13648 1340 13676 1380
rect 13556 1312 13676 1340
rect 13556 1272 13584 1312
rect 13722 1300 13728 1352
rect 13780 1300 13786 1352
rect 13832 1340 13860 1380
rect 15672 1380 15884 1408
rect 13998 1340 14004 1352
rect 13832 1312 14004 1340
rect 13998 1300 14004 1312
rect 14056 1300 14062 1352
rect 14093 1343 14151 1349
rect 14093 1309 14105 1343
rect 14139 1309 14151 1343
rect 14093 1303 14151 1309
rect 14369 1343 14427 1349
rect 14369 1309 14381 1343
rect 14415 1340 14427 1343
rect 14550 1340 14556 1352
rect 14415 1312 14556 1340
rect 14415 1309 14427 1312
rect 14369 1303 14427 1309
rect 14108 1272 14136 1303
rect 14550 1300 14556 1312
rect 14608 1300 14614 1352
rect 14645 1343 14703 1349
rect 14645 1309 14657 1343
rect 14691 1309 14703 1343
rect 14645 1303 14703 1309
rect 14921 1343 14979 1349
rect 14921 1309 14933 1343
rect 14967 1340 14979 1343
rect 15102 1340 15108 1352
rect 14967 1312 15108 1340
rect 14967 1309 14979 1312
rect 14921 1303 14979 1309
rect 14458 1272 14464 1284
rect 11808 1244 12112 1272
rect 12406 1244 13584 1272
rect 13648 1244 14044 1272
rect 14108 1244 14464 1272
rect 8113 1207 8171 1213
rect 8113 1173 8125 1207
rect 8159 1173 8171 1207
rect 8113 1167 8171 1173
rect 8481 1207 8539 1213
rect 8481 1173 8493 1207
rect 8527 1173 8539 1207
rect 8481 1167 8539 1173
rect 8754 1164 8760 1216
rect 8812 1164 8818 1216
rect 9214 1164 9220 1216
rect 9272 1164 9278 1216
rect 9582 1164 9588 1216
rect 9640 1164 9646 1216
rect 9950 1164 9956 1216
rect 10008 1164 10014 1216
rect 10318 1164 10324 1216
rect 10376 1164 10382 1216
rect 10686 1164 10692 1216
rect 10744 1164 10750 1216
rect 11054 1164 11060 1216
rect 11112 1164 11118 1216
rect 11330 1164 11336 1216
rect 11388 1164 11394 1216
rect 11808 1213 11836 1244
rect 11793 1207 11851 1213
rect 11793 1173 11805 1207
rect 11839 1173 11851 1207
rect 11793 1167 11851 1173
rect 12161 1207 12219 1213
rect 12161 1173 12173 1207
rect 12207 1204 12219 1207
rect 12406 1204 12434 1244
rect 12207 1176 12434 1204
rect 12207 1173 12219 1176
rect 12161 1167 12219 1173
rect 12526 1164 12532 1216
rect 12584 1164 12590 1216
rect 12802 1164 12808 1216
rect 12860 1164 12866 1216
rect 13078 1164 13084 1216
rect 13136 1164 13142 1216
rect 13262 1164 13268 1216
rect 13320 1204 13326 1216
rect 13648 1213 13676 1244
rect 13357 1207 13415 1213
rect 13357 1204 13369 1207
rect 13320 1176 13369 1204
rect 13320 1164 13326 1176
rect 13357 1173 13369 1176
rect 13403 1173 13415 1207
rect 13357 1167 13415 1173
rect 13633 1207 13691 1213
rect 13633 1173 13645 1207
rect 13679 1173 13691 1207
rect 13633 1167 13691 1173
rect 13906 1164 13912 1216
rect 13964 1164 13970 1216
rect 14016 1204 14044 1244
rect 14458 1232 14464 1244
rect 14516 1232 14522 1284
rect 14660 1272 14688 1303
rect 15102 1300 15108 1312
rect 15160 1300 15166 1352
rect 15197 1343 15255 1349
rect 15197 1309 15209 1343
rect 15243 1340 15255 1343
rect 15378 1340 15384 1352
rect 15243 1312 15384 1340
rect 15243 1309 15255 1312
rect 15197 1303 15255 1309
rect 15378 1300 15384 1312
rect 15436 1300 15442 1352
rect 15473 1343 15531 1349
rect 15473 1309 15485 1343
rect 15519 1340 15531 1343
rect 15672 1340 15700 1380
rect 15856 1352 15884 1380
rect 17126 1368 17132 1420
rect 17184 1408 17190 1420
rect 17184 1380 17632 1408
rect 17184 1368 17190 1380
rect 15519 1312 15700 1340
rect 15749 1343 15807 1349
rect 15519 1309 15531 1312
rect 15473 1303 15531 1309
rect 15749 1309 15761 1343
rect 15795 1309 15807 1343
rect 15749 1303 15807 1309
rect 15010 1272 15016 1284
rect 14660 1244 15016 1272
rect 15010 1232 15016 1244
rect 15068 1232 15074 1284
rect 15764 1272 15792 1303
rect 15838 1300 15844 1352
rect 15896 1300 15902 1352
rect 15930 1300 15936 1352
rect 15988 1300 15994 1352
rect 16022 1300 16028 1352
rect 16080 1300 16086 1352
rect 16301 1343 16359 1349
rect 16301 1309 16313 1343
rect 16347 1340 16359 1343
rect 16482 1340 16488 1352
rect 16347 1312 16488 1340
rect 16347 1309 16359 1312
rect 16301 1303 16359 1309
rect 16482 1300 16488 1312
rect 16540 1300 16546 1352
rect 16758 1300 16764 1352
rect 16816 1300 16822 1352
rect 17037 1343 17095 1349
rect 17037 1309 17049 1343
rect 17083 1309 17095 1343
rect 17037 1303 17095 1309
rect 15120 1244 15792 1272
rect 14090 1204 14096 1216
rect 14016 1176 14096 1204
rect 14090 1164 14096 1176
rect 14148 1164 14154 1216
rect 14829 1207 14887 1213
rect 14829 1173 14841 1207
rect 14875 1204 14887 1207
rect 15120 1204 15148 1244
rect 15948 1213 15976 1300
rect 17052 1272 17080 1303
rect 17310 1300 17316 1352
rect 17368 1300 17374 1352
rect 17494 1300 17500 1352
rect 17552 1300 17558 1352
rect 17604 1340 17632 1380
rect 18892 1380 19196 1408
rect 18892 1352 18920 1380
rect 17773 1343 17831 1349
rect 17773 1340 17785 1343
rect 17604 1312 17785 1340
rect 17773 1309 17785 1312
rect 17819 1309 17831 1343
rect 17773 1303 17831 1309
rect 18230 1300 18236 1352
rect 18288 1300 18294 1352
rect 18506 1300 18512 1352
rect 18564 1300 18570 1352
rect 18782 1300 18788 1352
rect 18840 1300 18846 1352
rect 18874 1300 18880 1352
rect 18932 1300 18938 1352
rect 18966 1300 18972 1352
rect 19024 1300 19030 1352
rect 19058 1300 19064 1352
rect 19116 1300 19122 1352
rect 19168 1340 19196 1380
rect 19812 1380 20668 1408
rect 19812 1352 19840 1380
rect 19245 1343 19303 1349
rect 19245 1340 19257 1343
rect 19168 1312 19257 1340
rect 19245 1309 19257 1312
rect 19291 1309 19303 1343
rect 19521 1343 19579 1349
rect 19521 1340 19533 1343
rect 19245 1303 19303 1309
rect 19352 1312 19533 1340
rect 16224 1244 17080 1272
rect 16224 1213 16252 1244
rect 14875 1176 15148 1204
rect 15933 1207 15991 1213
rect 14875 1173 14887 1176
rect 14829 1167 14887 1173
rect 15933 1173 15945 1207
rect 15979 1173 15991 1207
rect 15933 1167 15991 1173
rect 16209 1207 16267 1213
rect 16209 1173 16221 1207
rect 16255 1173 16267 1207
rect 16209 1167 16267 1173
rect 17221 1207 17279 1213
rect 17221 1173 17233 1207
rect 17267 1204 17279 1207
rect 17328 1204 17356 1300
rect 18984 1272 19012 1300
rect 19352 1272 19380 1312
rect 19521 1309 19533 1312
rect 19567 1309 19579 1343
rect 19521 1303 19579 1309
rect 19794 1300 19800 1352
rect 19852 1300 19858 1352
rect 19889 1343 19947 1349
rect 19889 1309 19901 1343
rect 19935 1309 19947 1343
rect 19889 1303 19947 1309
rect 19904 1272 19932 1303
rect 19978 1300 19984 1352
rect 20036 1340 20042 1352
rect 20257 1343 20315 1349
rect 20257 1340 20269 1343
rect 20036 1312 20269 1340
rect 20036 1300 20042 1312
rect 20257 1309 20269 1312
rect 20303 1309 20315 1343
rect 20640 1340 20668 1380
rect 21361 1343 21419 1349
rect 21361 1340 21373 1343
rect 20640 1312 21373 1340
rect 20257 1303 20315 1309
rect 21361 1309 21373 1312
rect 21407 1309 21419 1343
rect 21361 1303 21419 1309
rect 21450 1300 21456 1352
rect 21508 1340 21514 1352
rect 21821 1343 21879 1349
rect 21821 1340 21833 1343
rect 21508 1312 21833 1340
rect 21508 1300 21514 1312
rect 21821 1309 21833 1312
rect 21867 1309 21879 1343
rect 22020 1340 22048 1448
rect 22278 1436 22284 1488
rect 22336 1476 22342 1488
rect 22336 1448 23980 1476
rect 22336 1436 22342 1448
rect 22462 1368 22468 1420
rect 22520 1368 22526 1420
rect 22572 1380 22876 1408
rect 22572 1340 22600 1380
rect 22848 1349 22876 1380
rect 23566 1368 23572 1420
rect 23624 1368 23630 1420
rect 23952 1408 23980 1448
rect 24486 1436 24492 1488
rect 24544 1436 24550 1488
rect 24688 1476 24716 1516
rect 24762 1504 24768 1556
rect 24820 1544 24826 1556
rect 25041 1547 25099 1553
rect 25041 1544 25053 1547
rect 24820 1516 25053 1544
rect 24820 1504 24826 1516
rect 25041 1513 25053 1516
rect 25087 1513 25099 1547
rect 25041 1507 25099 1513
rect 25406 1504 25412 1556
rect 25464 1544 25470 1556
rect 27246 1544 27252 1556
rect 25464 1516 27252 1544
rect 25464 1504 25470 1516
rect 27246 1504 27252 1516
rect 27304 1504 27310 1556
rect 27338 1504 27344 1556
rect 27396 1544 27402 1556
rect 27893 1547 27951 1553
rect 27893 1544 27905 1547
rect 27396 1516 27905 1544
rect 27396 1504 27402 1516
rect 27893 1513 27905 1516
rect 27939 1513 27951 1547
rect 27893 1507 27951 1513
rect 28810 1504 28816 1556
rect 28868 1544 28874 1556
rect 29733 1547 29791 1553
rect 29733 1544 29745 1547
rect 28868 1516 29745 1544
rect 28868 1504 28874 1516
rect 29733 1513 29745 1516
rect 29779 1513 29791 1547
rect 29733 1507 29791 1513
rect 30006 1504 30012 1556
rect 30064 1544 30070 1556
rect 31021 1547 31079 1553
rect 31021 1544 31033 1547
rect 30064 1516 31033 1544
rect 30064 1504 30070 1516
rect 31021 1513 31033 1516
rect 31067 1513 31079 1547
rect 31021 1507 31079 1513
rect 31846 1504 31852 1556
rect 31904 1544 31910 1556
rect 32309 1547 32367 1553
rect 32309 1544 32321 1547
rect 31904 1516 32321 1544
rect 31904 1504 31910 1516
rect 32309 1513 32321 1516
rect 32355 1513 32367 1547
rect 32309 1507 32367 1513
rect 32766 1504 32772 1556
rect 32824 1544 32830 1556
rect 33413 1547 33471 1553
rect 33413 1544 33425 1547
rect 32824 1516 33425 1544
rect 32824 1504 32830 1516
rect 33413 1513 33425 1516
rect 33459 1513 33471 1547
rect 33413 1507 33471 1513
rect 33965 1547 34023 1553
rect 33965 1513 33977 1547
rect 34011 1513 34023 1547
rect 33965 1507 34023 1513
rect 24688 1448 31892 1476
rect 24504 1408 24532 1436
rect 23952 1380 24072 1408
rect 24504 1380 24808 1408
rect 22020 1312 22600 1340
rect 22833 1343 22891 1349
rect 21821 1303 21879 1309
rect 22833 1309 22845 1343
rect 22879 1309 22891 1343
rect 23937 1343 23995 1349
rect 23937 1340 23949 1343
rect 22833 1303 22891 1309
rect 22940 1312 23949 1340
rect 18984 1244 19380 1272
rect 19444 1244 19932 1272
rect 19444 1213 19472 1244
rect 20162 1232 20168 1284
rect 20220 1272 20226 1284
rect 20717 1275 20775 1281
rect 20717 1272 20729 1275
rect 20220 1244 20729 1272
rect 20220 1232 20226 1244
rect 20717 1241 20729 1244
rect 20763 1241 20775 1275
rect 20717 1235 20775 1241
rect 20898 1232 20904 1284
rect 20956 1272 20962 1284
rect 22189 1275 22247 1281
rect 22189 1272 22201 1275
rect 20956 1244 22201 1272
rect 20956 1232 20962 1244
rect 22189 1241 22201 1244
rect 22235 1241 22247 1275
rect 22940 1272 22968 1312
rect 23937 1309 23949 1312
rect 23983 1309 23995 1343
rect 24044 1340 24072 1380
rect 24489 1343 24547 1349
rect 24489 1340 24501 1343
rect 24044 1312 24501 1340
rect 23937 1303 23995 1309
rect 24489 1309 24501 1312
rect 24535 1309 24547 1343
rect 24780 1340 24808 1380
rect 24854 1368 24860 1420
rect 24912 1408 24918 1420
rect 24912 1380 25820 1408
rect 24912 1368 24918 1380
rect 25792 1349 25820 1380
rect 26418 1368 26424 1420
rect 26476 1368 26482 1420
rect 26878 1368 26884 1420
rect 26936 1408 26942 1420
rect 28166 1408 28172 1420
rect 26936 1380 28172 1408
rect 26936 1368 26942 1380
rect 28166 1368 28172 1380
rect 28224 1368 28230 1420
rect 28442 1368 28448 1420
rect 28500 1408 28506 1420
rect 28905 1411 28963 1417
rect 28905 1408 28917 1411
rect 28500 1380 28917 1408
rect 28500 1368 28506 1380
rect 28905 1377 28917 1380
rect 28951 1377 28963 1411
rect 28905 1371 28963 1377
rect 29546 1368 29552 1420
rect 29604 1408 29610 1420
rect 29604 1380 30328 1408
rect 29604 1368 29610 1380
rect 25409 1343 25467 1349
rect 25409 1340 25421 1343
rect 24780 1312 25421 1340
rect 24489 1303 24547 1309
rect 25409 1309 25421 1312
rect 25455 1309 25467 1343
rect 25409 1303 25467 1309
rect 25777 1343 25835 1349
rect 25777 1309 25789 1343
rect 25823 1309 25835 1343
rect 25777 1303 25835 1309
rect 26510 1300 26516 1352
rect 26568 1340 26574 1352
rect 26697 1343 26755 1349
rect 26697 1340 26709 1343
rect 26568 1312 26709 1340
rect 26568 1300 26574 1312
rect 26697 1309 26709 1312
rect 26743 1309 26755 1343
rect 26697 1303 26755 1309
rect 26786 1300 26792 1352
rect 26844 1340 26850 1352
rect 26973 1343 27031 1349
rect 26973 1340 26985 1343
rect 26844 1312 26985 1340
rect 26844 1300 26850 1312
rect 26973 1309 26985 1312
rect 27019 1309 27031 1343
rect 26973 1303 27031 1309
rect 27154 1300 27160 1352
rect 27212 1340 27218 1352
rect 27341 1343 27399 1349
rect 27341 1340 27353 1343
rect 27212 1312 27353 1340
rect 27212 1300 27218 1312
rect 27341 1309 27353 1312
rect 27387 1309 27399 1343
rect 27341 1303 27399 1309
rect 27706 1300 27712 1352
rect 27764 1340 27770 1352
rect 27801 1343 27859 1349
rect 27801 1340 27813 1343
rect 27764 1312 27813 1340
rect 27764 1300 27770 1312
rect 27801 1309 27813 1312
rect 27847 1309 27859 1343
rect 27801 1303 27859 1309
rect 27982 1300 27988 1352
rect 28040 1340 28046 1352
rect 28261 1343 28319 1349
rect 28261 1340 28273 1343
rect 28040 1312 28273 1340
rect 28040 1300 28046 1312
rect 28261 1309 28273 1312
rect 28307 1309 28319 1343
rect 28261 1303 28319 1309
rect 29178 1300 29184 1352
rect 29236 1300 29242 1352
rect 29270 1300 29276 1352
rect 29328 1340 29334 1352
rect 29641 1343 29699 1349
rect 29641 1340 29653 1343
rect 29328 1312 29653 1340
rect 29328 1300 29334 1312
rect 29641 1309 29653 1312
rect 29687 1309 29699 1343
rect 30300 1340 30328 1380
rect 30374 1368 30380 1420
rect 30432 1408 30438 1420
rect 31757 1411 31815 1417
rect 31757 1408 31769 1411
rect 30432 1380 31769 1408
rect 30432 1368 30438 1380
rect 31757 1377 31769 1380
rect 31803 1377 31815 1411
rect 31864 1408 31892 1448
rect 32950 1436 32956 1488
rect 33008 1476 33014 1488
rect 33980 1476 34008 1507
rect 34054 1504 34060 1556
rect 34112 1504 34118 1556
rect 34238 1504 34244 1556
rect 34296 1544 34302 1556
rect 34885 1547 34943 1553
rect 34885 1544 34897 1547
rect 34296 1516 34897 1544
rect 34296 1504 34302 1516
rect 34885 1513 34897 1516
rect 34931 1513 34943 1547
rect 34885 1507 34943 1513
rect 35437 1547 35495 1553
rect 35437 1513 35449 1547
rect 35483 1513 35495 1547
rect 35437 1507 35495 1513
rect 33008 1448 34008 1476
rect 33008 1436 33014 1448
rect 34072 1408 34100 1504
rect 34698 1436 34704 1488
rect 34756 1476 34762 1488
rect 35452 1476 35480 1507
rect 35802 1504 35808 1556
rect 35860 1544 35866 1556
rect 35989 1547 36047 1553
rect 35989 1544 36001 1547
rect 35860 1516 36001 1544
rect 35860 1504 35866 1516
rect 35989 1513 36001 1516
rect 36035 1513 36047 1547
rect 35989 1507 36047 1513
rect 36541 1547 36599 1553
rect 36541 1513 36553 1547
rect 36587 1513 36599 1547
rect 36541 1507 36599 1513
rect 34756 1448 35480 1476
rect 34756 1436 34762 1448
rect 35710 1436 35716 1488
rect 35768 1476 35774 1488
rect 36556 1476 36584 1507
rect 36998 1504 37004 1556
rect 37056 1544 37062 1556
rect 38013 1547 38071 1553
rect 38013 1544 38025 1547
rect 37056 1516 38025 1544
rect 37056 1504 37062 1516
rect 38013 1513 38025 1516
rect 38059 1513 38071 1547
rect 38013 1507 38071 1513
rect 38286 1504 38292 1556
rect 38344 1544 38350 1556
rect 39117 1547 39175 1553
rect 39117 1544 39129 1547
rect 38344 1516 39129 1544
rect 38344 1504 38350 1516
rect 39117 1513 39129 1516
rect 39163 1513 39175 1547
rect 39117 1507 39175 1513
rect 39206 1504 39212 1556
rect 39264 1544 39270 1556
rect 40405 1547 40463 1553
rect 40405 1544 40417 1547
rect 39264 1516 40417 1544
rect 39264 1504 39270 1516
rect 40405 1513 40417 1516
rect 40451 1513 40463 1547
rect 40405 1507 40463 1513
rect 42426 1504 42432 1556
rect 42484 1504 42490 1556
rect 42518 1504 42524 1556
rect 42576 1544 42582 1556
rect 44637 1547 44695 1553
rect 44637 1544 44649 1547
rect 42576 1516 44649 1544
rect 42576 1504 42582 1516
rect 44637 1513 44649 1516
rect 44683 1513 44695 1547
rect 44637 1507 44695 1513
rect 35768 1448 36584 1476
rect 35768 1436 35774 1448
rect 37366 1436 37372 1488
rect 37424 1476 37430 1488
rect 38657 1479 38715 1485
rect 38657 1476 38669 1479
rect 37424 1448 38669 1476
rect 37424 1436 37430 1448
rect 38657 1445 38669 1448
rect 38703 1445 38715 1479
rect 38657 1439 38715 1445
rect 38838 1436 38844 1488
rect 38896 1476 38902 1488
rect 40129 1479 40187 1485
rect 40129 1476 40141 1479
rect 38896 1448 40141 1476
rect 38896 1436 38902 1448
rect 40129 1445 40141 1448
rect 40175 1445 40187 1479
rect 40129 1439 40187 1445
rect 41340 1448 43116 1476
rect 31864 1380 34100 1408
rect 31757 1371 31815 1377
rect 35802 1368 35808 1420
rect 35860 1408 35866 1420
rect 37645 1411 37703 1417
rect 37645 1408 37657 1411
rect 35860 1380 37657 1408
rect 35860 1368 35866 1380
rect 37645 1377 37657 1380
rect 37691 1377 37703 1411
rect 37645 1371 37703 1377
rect 37918 1368 37924 1420
rect 37976 1408 37982 1420
rect 41340 1408 41368 1448
rect 37976 1380 41368 1408
rect 41892 1380 42104 1408
rect 37976 1368 37982 1380
rect 30300 1312 30420 1340
rect 29641 1303 29699 1309
rect 22189 1235 22247 1241
rect 22296 1244 22968 1272
rect 17267 1176 17356 1204
rect 19429 1207 19487 1213
rect 17267 1173 17279 1176
rect 17221 1167 17279 1173
rect 19429 1173 19441 1207
rect 19475 1173 19487 1207
rect 19429 1167 19487 1173
rect 19702 1164 19708 1216
rect 19760 1164 19766 1216
rect 20070 1164 20076 1216
rect 20128 1164 20134 1216
rect 20438 1164 20444 1216
rect 20496 1164 20502 1216
rect 20806 1164 20812 1216
rect 20864 1164 20870 1216
rect 21542 1164 21548 1216
rect 21600 1164 21606 1216
rect 22005 1207 22063 1213
rect 22005 1173 22017 1207
rect 22051 1204 22063 1207
rect 22296 1204 22324 1244
rect 23106 1232 23112 1284
rect 23164 1272 23170 1284
rect 23293 1275 23351 1281
rect 23293 1272 23305 1275
rect 23164 1244 23305 1272
rect 23164 1232 23170 1244
rect 23293 1241 23305 1244
rect 23339 1241 23351 1275
rect 23293 1235 23351 1241
rect 24578 1232 24584 1284
rect 24636 1272 24642 1284
rect 24636 1244 24808 1272
rect 24636 1232 24642 1244
rect 22051 1176 22324 1204
rect 22051 1173 22063 1176
rect 22005 1167 22063 1173
rect 23014 1164 23020 1216
rect 23072 1164 23078 1216
rect 24118 1164 24124 1216
rect 24176 1164 24182 1216
rect 24670 1164 24676 1216
rect 24728 1164 24734 1216
rect 24780 1204 24808 1244
rect 24946 1232 24952 1284
rect 25004 1232 25010 1284
rect 25056 1244 28580 1272
rect 25056 1204 25084 1244
rect 24780 1176 25084 1204
rect 25130 1164 25136 1216
rect 25188 1204 25194 1216
rect 25593 1207 25651 1213
rect 25593 1204 25605 1207
rect 25188 1176 25605 1204
rect 25188 1164 25194 1176
rect 25593 1173 25605 1176
rect 25639 1173 25651 1207
rect 25593 1167 25651 1173
rect 25682 1164 25688 1216
rect 25740 1204 25746 1216
rect 25961 1207 26019 1213
rect 25961 1204 25973 1207
rect 25740 1176 25973 1204
rect 25740 1164 25746 1176
rect 25961 1173 25973 1176
rect 26007 1173 26019 1207
rect 25961 1167 26019 1173
rect 26602 1164 26608 1216
rect 26660 1204 26666 1216
rect 27157 1207 27215 1213
rect 27157 1204 27169 1207
rect 26660 1176 27169 1204
rect 26660 1164 26666 1176
rect 27157 1173 27169 1176
rect 27203 1173 27215 1207
rect 27157 1167 27215 1173
rect 27246 1164 27252 1216
rect 27304 1204 27310 1216
rect 27525 1207 27583 1213
rect 27525 1204 27537 1207
rect 27304 1176 27537 1204
rect 27304 1164 27310 1176
rect 27525 1173 27537 1176
rect 27571 1173 27583 1207
rect 27525 1167 27583 1173
rect 27706 1164 27712 1216
rect 27764 1204 27770 1216
rect 28445 1207 28503 1213
rect 28445 1204 28457 1207
rect 27764 1176 28457 1204
rect 27764 1164 27770 1176
rect 28445 1173 28457 1176
rect 28491 1173 28503 1207
rect 28552 1204 28580 1244
rect 29546 1232 29552 1284
rect 29604 1272 29610 1284
rect 30285 1275 30343 1281
rect 30285 1272 30297 1275
rect 29604 1244 30297 1272
rect 29604 1232 29610 1244
rect 30285 1241 30297 1244
rect 30331 1241 30343 1275
rect 30392 1272 30420 1312
rect 30466 1300 30472 1352
rect 30524 1340 30530 1352
rect 30653 1343 30711 1349
rect 30653 1340 30665 1343
rect 30524 1312 30665 1340
rect 30524 1300 30530 1312
rect 30653 1309 30665 1312
rect 30699 1309 30711 1343
rect 30653 1303 30711 1309
rect 30742 1300 30748 1352
rect 30800 1340 30806 1352
rect 30929 1343 30987 1349
rect 30929 1340 30941 1343
rect 30800 1312 30941 1340
rect 30800 1300 30806 1312
rect 30929 1309 30941 1312
rect 30975 1309 30987 1343
rect 30929 1303 30987 1309
rect 31018 1300 31024 1352
rect 31076 1340 31082 1352
rect 31481 1343 31539 1349
rect 31481 1340 31493 1343
rect 31076 1312 31493 1340
rect 31076 1300 31082 1312
rect 31481 1309 31493 1312
rect 31527 1309 31539 1343
rect 31481 1303 31539 1309
rect 31938 1300 31944 1352
rect 31996 1340 32002 1352
rect 32217 1343 32275 1349
rect 32217 1340 32229 1343
rect 31996 1312 32229 1340
rect 31996 1300 32002 1312
rect 32217 1309 32229 1312
rect 32263 1309 32275 1343
rect 32217 1303 32275 1309
rect 32677 1343 32735 1349
rect 32677 1309 32689 1343
rect 32723 1309 32735 1343
rect 32677 1303 32735 1309
rect 32692 1272 32720 1303
rect 35158 1300 35164 1352
rect 35216 1340 35222 1352
rect 35897 1343 35955 1349
rect 35897 1340 35909 1343
rect 35216 1312 35909 1340
rect 35216 1300 35222 1312
rect 35897 1309 35909 1312
rect 35943 1309 35955 1343
rect 35897 1303 35955 1309
rect 37090 1300 37096 1352
rect 37148 1340 37154 1352
rect 37148 1312 38608 1340
rect 37148 1300 37154 1312
rect 30392 1244 32720 1272
rect 30285 1235 30343 1241
rect 33318 1232 33324 1284
rect 33376 1232 33382 1284
rect 33410 1232 33416 1284
rect 33468 1272 33474 1284
rect 33873 1275 33931 1281
rect 33873 1272 33885 1275
rect 33468 1244 33885 1272
rect 33468 1232 33474 1244
rect 33873 1241 33885 1244
rect 33919 1241 33931 1275
rect 33873 1235 33931 1241
rect 34790 1232 34796 1284
rect 34848 1232 34854 1284
rect 34882 1232 34888 1284
rect 34940 1272 34946 1284
rect 35345 1275 35403 1281
rect 35345 1272 35357 1275
rect 34940 1244 35357 1272
rect 34940 1232 34946 1244
rect 35345 1241 35357 1244
rect 35391 1241 35403 1275
rect 35345 1235 35403 1241
rect 35434 1232 35440 1284
rect 35492 1272 35498 1284
rect 36449 1275 36507 1281
rect 36449 1272 36461 1275
rect 35492 1244 36461 1272
rect 35492 1232 35498 1244
rect 36449 1241 36461 1244
rect 36495 1241 36507 1275
rect 36449 1235 36507 1241
rect 37369 1275 37427 1281
rect 37369 1241 37381 1275
rect 37415 1272 37427 1275
rect 37458 1272 37464 1284
rect 37415 1244 37464 1272
rect 37415 1241 37427 1244
rect 37369 1235 37427 1241
rect 37458 1232 37464 1244
rect 37516 1232 37522 1284
rect 37826 1232 37832 1284
rect 37884 1272 37890 1284
rect 37921 1275 37979 1281
rect 37921 1272 37933 1275
rect 37884 1244 37933 1272
rect 37884 1232 37890 1244
rect 37921 1241 37933 1244
rect 37967 1241 37979 1275
rect 37921 1235 37979 1241
rect 38102 1232 38108 1284
rect 38160 1272 38166 1284
rect 38473 1275 38531 1281
rect 38473 1272 38485 1275
rect 38160 1244 38485 1272
rect 38160 1232 38166 1244
rect 38473 1241 38485 1244
rect 38519 1241 38531 1275
rect 38580 1272 38608 1312
rect 38746 1300 38752 1352
rect 38804 1340 38810 1352
rect 39669 1343 39727 1349
rect 39669 1340 39681 1343
rect 38804 1312 39681 1340
rect 38804 1300 38810 1312
rect 39669 1309 39681 1312
rect 39715 1309 39727 1343
rect 40589 1343 40647 1349
rect 40589 1340 40601 1343
rect 39669 1303 39727 1309
rect 39868 1312 40601 1340
rect 39025 1275 39083 1281
rect 39025 1272 39037 1275
rect 38580 1244 39037 1272
rect 38473 1235 38531 1241
rect 39025 1241 39037 1244
rect 39071 1241 39083 1275
rect 39025 1235 39083 1241
rect 39206 1232 39212 1284
rect 39264 1272 39270 1284
rect 39868 1272 39896 1312
rect 40589 1309 40601 1312
rect 40635 1309 40647 1343
rect 40589 1303 40647 1309
rect 40865 1343 40923 1349
rect 40865 1309 40877 1343
rect 40911 1309 40923 1343
rect 40865 1303 40923 1309
rect 39264 1244 39896 1272
rect 39945 1275 40003 1281
rect 39264 1232 39270 1244
rect 39945 1241 39957 1275
rect 39991 1241 40003 1275
rect 40880 1272 40908 1303
rect 41138 1300 41144 1352
rect 41196 1300 41202 1352
rect 41230 1300 41236 1352
rect 41288 1340 41294 1352
rect 41892 1340 41920 1380
rect 41288 1312 41920 1340
rect 41288 1300 41294 1312
rect 41966 1300 41972 1352
rect 42024 1300 42030 1352
rect 42076 1340 42104 1380
rect 42702 1368 42708 1420
rect 42760 1408 42766 1420
rect 43088 1408 43116 1448
rect 43530 1436 43536 1488
rect 43588 1436 43594 1488
rect 43806 1436 43812 1488
rect 43864 1436 43870 1488
rect 44174 1436 44180 1488
rect 44232 1476 44238 1488
rect 44361 1479 44419 1485
rect 44361 1476 44373 1479
rect 44232 1448 44373 1476
rect 44232 1436 44238 1448
rect 44361 1445 44373 1448
rect 44407 1445 44419 1479
rect 44361 1439 44419 1445
rect 45005 1479 45063 1485
rect 45005 1445 45017 1479
rect 45051 1445 45063 1479
rect 45005 1439 45063 1445
rect 45020 1408 45048 1439
rect 42760 1380 43024 1408
rect 43088 1380 45048 1408
rect 42760 1368 42766 1380
rect 42245 1343 42303 1349
rect 42245 1340 42257 1343
rect 42076 1312 42257 1340
rect 42245 1309 42257 1312
rect 42291 1309 42303 1343
rect 42613 1343 42671 1349
rect 42613 1340 42625 1343
rect 42245 1303 42303 1309
rect 42352 1312 42625 1340
rect 41322 1272 41328 1284
rect 40880 1244 41328 1272
rect 39945 1235 40003 1241
rect 29638 1204 29644 1216
rect 28552 1176 29644 1204
rect 28445 1167 28503 1173
rect 29638 1164 29644 1176
rect 29696 1164 29702 1216
rect 31754 1164 31760 1216
rect 31812 1204 31818 1216
rect 32861 1207 32919 1213
rect 32861 1204 32873 1207
rect 31812 1176 32873 1204
rect 31812 1164 31818 1176
rect 32861 1173 32873 1176
rect 32907 1173 32919 1207
rect 32861 1167 32919 1173
rect 32950 1164 32956 1216
rect 33008 1204 33014 1216
rect 39298 1204 39304 1216
rect 33008 1176 39304 1204
rect 33008 1164 33014 1176
rect 39298 1164 39304 1176
rect 39356 1164 39362 1216
rect 39390 1164 39396 1216
rect 39448 1204 39454 1216
rect 39485 1207 39543 1213
rect 39485 1204 39497 1207
rect 39448 1176 39497 1204
rect 39448 1164 39454 1176
rect 39485 1173 39497 1176
rect 39531 1173 39543 1207
rect 39485 1167 39543 1173
rect 39666 1164 39672 1216
rect 39724 1204 39730 1216
rect 39960 1204 39988 1235
rect 41322 1232 41328 1244
rect 41380 1232 41386 1284
rect 41690 1232 41696 1284
rect 41748 1272 41754 1284
rect 42352 1272 42380 1312
rect 42613 1309 42625 1312
rect 42659 1309 42671 1343
rect 42889 1343 42947 1349
rect 42889 1340 42901 1343
rect 42613 1303 42671 1309
rect 42720 1312 42901 1340
rect 42720 1272 42748 1312
rect 42889 1309 42901 1312
rect 42935 1309 42947 1343
rect 42996 1340 43024 1380
rect 43165 1343 43223 1349
rect 43165 1340 43177 1343
rect 42996 1312 43177 1340
rect 42889 1303 42947 1309
rect 43165 1309 43177 1312
rect 43211 1309 43223 1343
rect 43441 1343 43499 1349
rect 43441 1340 43453 1343
rect 43165 1303 43223 1309
rect 43272 1312 43453 1340
rect 41748 1244 42380 1272
rect 42444 1244 42748 1272
rect 41748 1232 41754 1244
rect 39724 1176 39988 1204
rect 39724 1164 39730 1176
rect 40034 1164 40040 1216
rect 40092 1204 40098 1216
rect 41785 1207 41843 1213
rect 41785 1204 41797 1207
rect 40092 1176 41797 1204
rect 40092 1164 40098 1176
rect 41785 1173 41797 1176
rect 41831 1173 41843 1207
rect 41785 1167 41843 1173
rect 42058 1164 42064 1216
rect 42116 1164 42122 1216
rect 42334 1164 42340 1216
rect 42392 1204 42398 1216
rect 42444 1204 42472 1244
rect 42794 1232 42800 1284
rect 42852 1272 42858 1284
rect 43272 1272 43300 1312
rect 43441 1309 43453 1312
rect 43487 1309 43499 1343
rect 43717 1343 43775 1349
rect 43717 1340 43729 1343
rect 43441 1303 43499 1309
rect 43548 1312 43729 1340
rect 42852 1244 43300 1272
rect 42852 1232 42858 1244
rect 43346 1232 43352 1284
rect 43404 1272 43410 1284
rect 43548 1272 43576 1312
rect 43717 1309 43729 1312
rect 43763 1309 43775 1343
rect 43717 1303 43775 1309
rect 43993 1343 44051 1349
rect 43993 1309 44005 1343
rect 44039 1309 44051 1343
rect 43993 1303 44051 1309
rect 43404 1244 43576 1272
rect 43404 1232 43410 1244
rect 43622 1232 43628 1284
rect 43680 1272 43686 1284
rect 44008 1272 44036 1303
rect 44266 1300 44272 1352
rect 44324 1300 44330 1352
rect 44542 1300 44548 1352
rect 44600 1300 44606 1352
rect 44818 1300 44824 1352
rect 44876 1300 44882 1352
rect 45189 1343 45247 1349
rect 45189 1309 45201 1343
rect 45235 1309 45247 1343
rect 45189 1303 45247 1309
rect 43680 1244 44036 1272
rect 43680 1232 43686 1244
rect 44726 1232 44732 1284
rect 44784 1272 44790 1284
rect 45204 1272 45232 1303
rect 44784 1244 45232 1272
rect 44784 1232 44790 1244
rect 42392 1176 42472 1204
rect 42392 1164 42398 1176
rect 42518 1164 42524 1216
rect 42576 1204 42582 1216
rect 42705 1207 42763 1213
rect 42705 1204 42717 1207
rect 42576 1176 42717 1204
rect 42576 1164 42582 1176
rect 42705 1173 42717 1176
rect 42751 1173 42763 1207
rect 42705 1167 42763 1173
rect 42978 1164 42984 1216
rect 43036 1164 43042 1216
rect 43070 1164 43076 1216
rect 43128 1204 43134 1216
rect 43257 1207 43315 1213
rect 43257 1204 43269 1207
rect 43128 1176 43269 1204
rect 43128 1164 43134 1176
rect 43257 1173 43269 1176
rect 43303 1173 43315 1207
rect 43257 1167 43315 1173
rect 44082 1164 44088 1216
rect 44140 1164 44146 1216
rect 1104 1114 45696 1136
rect 1104 1062 12058 1114
rect 12110 1062 12122 1114
rect 12174 1062 12186 1114
rect 12238 1062 12250 1114
rect 12302 1062 12314 1114
rect 12366 1062 23166 1114
rect 23218 1062 23230 1114
rect 23282 1062 23294 1114
rect 23346 1062 23358 1114
rect 23410 1062 23422 1114
rect 23474 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 34530 1114
rect 34582 1062 45382 1114
rect 45434 1062 45446 1114
rect 45498 1062 45510 1114
rect 45562 1062 45574 1114
rect 45626 1062 45638 1114
rect 45690 1062 45696 1114
rect 1104 1040 45696 1062
rect 3602 960 3608 1012
rect 3660 1000 3666 1012
rect 5534 1000 5540 1012
rect 3660 972 5540 1000
rect 3660 960 3666 972
rect 5534 960 5540 972
rect 5592 960 5598 1012
rect 6638 960 6644 1012
rect 6696 1000 6702 1012
rect 10962 1000 10968 1012
rect 6696 972 10968 1000
rect 6696 960 6702 972
rect 10962 960 10968 972
rect 11020 960 11026 1012
rect 11330 960 11336 1012
rect 11388 1000 11394 1012
rect 24578 1000 24584 1012
rect 11388 972 24584 1000
rect 11388 960 11394 972
rect 24578 960 24584 972
rect 24636 960 24642 1012
rect 25406 1000 25412 1012
rect 24872 972 25412 1000
rect 4430 892 4436 944
rect 4488 892 4494 944
rect 5166 892 5172 944
rect 5224 932 5230 944
rect 5224 904 12434 932
rect 5224 892 5230 904
rect 4448 796 4476 892
rect 5902 824 5908 876
rect 5960 864 5966 876
rect 9858 864 9864 876
rect 5960 836 9864 864
rect 5960 824 5966 836
rect 9858 824 9864 836
rect 9916 824 9922 876
rect 9950 824 9956 876
rect 10008 824 10014 876
rect 10410 824 10416 876
rect 10468 824 10474 876
rect 4448 768 6040 796
rect 5810 688 5816 740
rect 5868 688 5874 740
rect 5828 524 5856 688
rect 6012 592 6040 768
rect 6086 756 6092 808
rect 6144 796 6150 808
rect 8938 796 8944 808
rect 6144 768 8944 796
rect 6144 756 6150 768
rect 8938 756 8944 768
rect 8996 756 9002 808
rect 9968 660 9996 824
rect 10428 728 10456 824
rect 12406 796 12434 904
rect 13078 892 13084 944
rect 13136 892 13142 944
rect 17678 892 17684 944
rect 17736 932 17742 944
rect 24872 932 24900 972
rect 25406 960 25412 972
rect 25464 960 25470 1012
rect 27522 960 27528 1012
rect 27580 960 27586 1012
rect 30374 960 30380 1012
rect 30432 1000 30438 1012
rect 30650 1000 30656 1012
rect 30432 972 30656 1000
rect 30432 960 30438 972
rect 30650 960 30656 972
rect 30708 960 30714 1012
rect 31386 960 31392 1012
rect 31444 1000 31450 1012
rect 35434 1000 35440 1012
rect 31444 972 35440 1000
rect 31444 960 31450 972
rect 35434 960 35440 972
rect 35492 960 35498 1012
rect 40034 1000 40040 1012
rect 35866 972 40040 1000
rect 27540 932 27568 960
rect 17736 904 24900 932
rect 24964 904 27568 932
rect 17736 892 17742 904
rect 13096 864 13124 892
rect 13096 836 17540 864
rect 12986 796 12992 808
rect 12406 768 12992 796
rect 12986 756 12992 768
rect 13044 756 13050 808
rect 13078 756 13084 808
rect 13136 796 13142 808
rect 13354 796 13360 808
rect 13136 768 13360 796
rect 13136 756 13142 768
rect 13354 756 13360 768
rect 13412 756 13418 808
rect 16758 756 16764 808
rect 16816 796 16822 808
rect 17402 796 17408 808
rect 16816 768 17408 796
rect 16816 756 16822 768
rect 17402 756 17408 768
rect 17460 756 17466 808
rect 17512 796 17540 836
rect 17862 824 17868 876
rect 17920 864 17926 876
rect 24964 864 24992 904
rect 30098 892 30104 944
rect 30156 932 30162 944
rect 35866 932 35894 972
rect 40034 960 40040 972
rect 40092 960 40098 1012
rect 40586 960 40592 1012
rect 40644 1000 40650 1012
rect 41966 1000 41972 1012
rect 40644 972 41972 1000
rect 40644 960 40650 972
rect 41966 960 41972 972
rect 42024 960 42030 1012
rect 42518 960 42524 1012
rect 42576 960 42582 1012
rect 43070 960 43076 1012
rect 43128 960 43134 1012
rect 30156 904 35894 932
rect 30156 892 30162 904
rect 39298 892 39304 944
rect 39356 932 39362 944
rect 42536 932 42564 960
rect 39356 904 42564 932
rect 39356 892 39362 904
rect 17920 836 24992 864
rect 17920 824 17926 836
rect 27062 824 27068 876
rect 27120 864 27126 876
rect 43088 864 43116 960
rect 27120 836 43116 864
rect 27120 824 27126 836
rect 25774 796 25780 808
rect 17512 768 25780 796
rect 25774 756 25780 768
rect 25832 756 25838 808
rect 39390 796 39396 808
rect 26896 768 39396 796
rect 10428 700 17264 728
rect 17236 660 17264 700
rect 17310 688 17316 740
rect 17368 728 17374 740
rect 26896 728 26924 768
rect 39390 756 39396 768
rect 39448 756 39454 808
rect 42058 756 42064 808
rect 42116 756 42122 808
rect 42978 756 42984 808
rect 43036 756 43042 808
rect 17368 700 26924 728
rect 17368 688 17374 700
rect 28626 688 28632 740
rect 28684 728 28690 740
rect 32950 728 32956 740
rect 28684 700 32956 728
rect 28684 688 28690 700
rect 32950 688 32956 700
rect 33008 688 33014 740
rect 27798 660 27804 672
rect 9968 632 17172 660
rect 17236 632 27804 660
rect 6012 564 7696 592
rect 5828 496 7328 524
rect 7006 416 7012 468
rect 7064 416 7070 468
rect 1578 212 1584 264
rect 1636 212 1642 264
rect 1596 116 1624 212
rect 7024 184 7052 416
rect 7300 252 7328 496
rect 7668 456 7696 564
rect 11054 552 11060 604
rect 11112 592 11118 604
rect 11112 564 15240 592
rect 11112 552 11118 564
rect 7742 484 7748 536
rect 7800 524 7806 536
rect 11238 524 11244 536
rect 7800 496 11244 524
rect 7800 484 7806 496
rect 11238 484 11244 496
rect 11296 484 11302 536
rect 15212 524 15240 564
rect 15746 552 15752 604
rect 15804 592 15810 604
rect 17034 592 17040 604
rect 15804 564 17040 592
rect 15804 552 15810 564
rect 17034 552 17040 564
rect 17092 552 17098 604
rect 17144 592 17172 632
rect 27798 620 27804 632
rect 27856 620 27862 672
rect 27890 620 27896 672
rect 27948 660 27954 672
rect 42076 660 42104 756
rect 27948 632 42104 660
rect 27948 620 27954 632
rect 23566 592 23572 604
rect 17144 564 23572 592
rect 23566 552 23572 564
rect 23624 552 23630 604
rect 28994 552 29000 604
rect 29052 592 29058 604
rect 33410 592 33416 604
rect 29052 564 33416 592
rect 29052 552 29058 564
rect 33410 552 33416 564
rect 33468 552 33474 604
rect 28350 524 28356 536
rect 15212 496 28356 524
rect 28350 484 28356 496
rect 28408 484 28414 536
rect 12066 456 12072 468
rect 7668 428 12072 456
rect 12066 416 12072 428
rect 12124 416 12130 468
rect 13998 416 14004 468
rect 14056 456 14062 468
rect 17678 456 17684 468
rect 14056 428 17684 456
rect 14056 416 14062 428
rect 17678 416 17684 428
rect 17736 416 17742 468
rect 20254 416 20260 468
rect 20312 416 20318 468
rect 25222 416 25228 468
rect 25280 456 25286 468
rect 42996 456 43024 756
rect 25280 428 28396 456
rect 25280 416 25286 428
rect 7650 348 7656 400
rect 7708 388 7714 400
rect 13630 388 13636 400
rect 7708 360 13636 388
rect 7708 348 7714 360
rect 13630 348 13636 360
rect 13688 348 13694 400
rect 13906 348 13912 400
rect 13964 388 13970 400
rect 20272 388 20300 416
rect 13964 360 20300 388
rect 22066 360 26924 388
rect 13964 348 13970 360
rect 12526 280 12532 332
rect 12584 320 12590 332
rect 22066 320 22094 360
rect 26896 332 26924 360
rect 26694 320 26700 332
rect 12584 292 22094 320
rect 24504 292 26700 320
rect 12584 280 12590 292
rect 12710 252 12716 264
rect 7300 224 12716 252
rect 12710 212 12716 224
rect 12768 212 12774 264
rect 13262 212 13268 264
rect 13320 252 13326 264
rect 24504 252 24532 292
rect 26694 280 26700 292
rect 26752 280 26758 332
rect 26878 280 26884 332
rect 26936 280 26942 332
rect 28368 320 28396 428
rect 32876 428 43024 456
rect 28534 348 28540 400
rect 28592 388 28598 400
rect 28994 388 29000 400
rect 28592 360 29000 388
rect 28592 348 28598 360
rect 28994 348 29000 360
rect 29052 348 29058 400
rect 32876 320 32904 428
rect 34882 348 34888 400
rect 34940 348 34946 400
rect 36262 348 36268 400
rect 36320 388 36326 400
rect 44082 388 44088 400
rect 36320 360 44088 388
rect 36320 348 36326 360
rect 44082 348 44088 360
rect 44140 348 44146 400
rect 28368 292 32904 320
rect 33318 280 33324 332
rect 33376 280 33382 332
rect 13320 224 24532 252
rect 13320 212 13326 224
rect 26050 212 26056 264
rect 26108 252 26114 264
rect 33336 252 33364 280
rect 26108 224 33364 252
rect 26108 212 26114 224
rect 18322 184 18328 196
rect 7024 156 18328 184
rect 18322 144 18328 156
rect 18380 144 18386 196
rect 25038 144 25044 196
rect 25096 184 25102 196
rect 34900 184 34928 348
rect 25096 156 34928 184
rect 25096 144 25102 156
rect 11698 116 11704 128
rect 1596 88 11704 116
rect 11698 76 11704 88
rect 11756 76 11762 128
rect 11790 76 11796 128
rect 11848 76 11854 128
rect 12066 76 12072 128
rect 12124 116 12130 128
rect 12124 88 12434 116
rect 12124 76 12130 88
rect 4062 8 4068 60
rect 4120 48 4126 60
rect 11808 48 11836 76
rect 4120 20 11836 48
rect 12406 48 12434 88
rect 23566 76 23572 128
rect 23624 116 23630 128
rect 30374 116 30380 128
rect 23624 88 30380 116
rect 23624 76 23630 88
rect 30374 76 30380 88
rect 30432 76 30438 128
rect 13078 48 13084 60
rect 12406 20 13084 48
rect 4120 8 4126 20
rect 13078 8 13084 20
rect 13136 8 13142 60
<< via1 >>
rect 17316 8916 17368 8968
rect 22376 8916 22428 8968
rect 8208 8848 8260 8900
rect 22928 8848 22980 8900
rect 4068 8780 4120 8832
rect 23664 8780 23716 8832
rect 12058 8678 12110 8730
rect 12122 8678 12174 8730
rect 12186 8678 12238 8730
rect 12250 8678 12302 8730
rect 12314 8678 12366 8730
rect 23166 8678 23218 8730
rect 23230 8678 23282 8730
rect 23294 8678 23346 8730
rect 23358 8678 23410 8730
rect 23422 8678 23474 8730
rect 34274 8678 34326 8730
rect 34338 8678 34390 8730
rect 34402 8678 34454 8730
rect 34466 8678 34518 8730
rect 34530 8678 34582 8730
rect 45382 8678 45434 8730
rect 45446 8678 45498 8730
rect 45510 8678 45562 8730
rect 45574 8678 45626 8730
rect 45638 8678 45690 8730
rect 3424 8576 3476 8628
rect 5632 8619 5684 8628
rect 5632 8585 5641 8619
rect 5641 8585 5675 8619
rect 5675 8585 5684 8619
rect 5632 8576 5684 8585
rect 7840 8576 7892 8628
rect 10048 8576 10100 8628
rect 14464 8576 14516 8628
rect 1400 8551 1452 8560
rect 1400 8517 1409 8551
rect 1409 8517 1443 8551
rect 1443 8517 1452 8551
rect 1400 8508 1452 8517
rect 4068 8483 4120 8492
rect 4068 8449 4077 8483
rect 4077 8449 4111 8483
rect 4111 8449 4120 8483
rect 4068 8440 4120 8449
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 12164 8551 12216 8560
rect 12164 8517 12173 8551
rect 12173 8517 12207 8551
rect 12207 8517 12216 8551
rect 12164 8508 12216 8517
rect 17316 8576 17368 8628
rect 18880 8576 18932 8628
rect 21088 8576 21140 8628
rect 25504 8576 25556 8628
rect 27712 8619 27764 8628
rect 27712 8585 27721 8619
rect 27721 8585 27755 8619
rect 27755 8585 27764 8619
rect 27712 8576 27764 8585
rect 29920 8576 29972 8628
rect 32128 8576 32180 8628
rect 34152 8576 34204 8628
rect 36544 8576 36596 8628
rect 38752 8619 38804 8628
rect 38752 8585 38761 8619
rect 38761 8585 38795 8619
rect 38795 8585 38804 8619
rect 38752 8576 38804 8585
rect 40960 8576 41012 8628
rect 43168 8576 43220 8628
rect 45284 8576 45336 8628
rect 16672 8551 16724 8560
rect 16672 8517 16681 8551
rect 16681 8517 16715 8551
rect 16715 8517 16724 8551
rect 16672 8508 16724 8517
rect 13820 8440 13872 8492
rect 20628 8508 20680 8560
rect 23020 8508 23072 8560
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 19248 8440 19300 8492
rect 19340 8483 19392 8492
rect 19340 8449 19349 8483
rect 19349 8449 19383 8483
rect 19383 8449 19392 8483
rect 19340 8440 19392 8449
rect 21456 8483 21508 8492
rect 21456 8449 21465 8483
rect 21465 8449 21499 8483
rect 21499 8449 21508 8483
rect 21456 8440 21508 8449
rect 23572 8483 23624 8492
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 25872 8483 25924 8492
rect 25872 8449 25881 8483
rect 25881 8449 25915 8483
rect 25915 8449 25924 8483
rect 25872 8440 25924 8449
rect 27988 8483 28040 8492
rect 27988 8449 27997 8483
rect 27997 8449 28031 8483
rect 28031 8449 28040 8483
rect 27988 8440 28040 8449
rect 30380 8440 30432 8492
rect 32496 8483 32548 8492
rect 32496 8449 32505 8483
rect 32505 8449 32539 8483
rect 32539 8449 32548 8483
rect 32496 8440 32548 8449
rect 34796 8483 34848 8492
rect 34796 8449 34805 8483
rect 34805 8449 34839 8483
rect 34839 8449 34848 8483
rect 34796 8440 34848 8449
rect 36912 8483 36964 8492
rect 36912 8449 36921 8483
rect 36921 8449 36955 8483
rect 36955 8449 36964 8483
rect 36912 8440 36964 8449
rect 39028 8483 39080 8492
rect 39028 8449 39037 8483
rect 39037 8449 39071 8483
rect 39071 8449 39080 8483
rect 39028 8440 39080 8449
rect 41328 8483 41380 8492
rect 41328 8449 41337 8483
rect 41337 8449 41371 8483
rect 41371 8449 41380 8483
rect 41328 8440 41380 8449
rect 43536 8483 43588 8492
rect 43536 8449 43545 8483
rect 43545 8449 43579 8483
rect 43579 8449 43588 8483
rect 43536 8440 43588 8449
rect 44548 8483 44600 8492
rect 44548 8449 44557 8483
rect 44557 8449 44591 8483
rect 44591 8449 44600 8483
rect 44548 8440 44600 8449
rect 23020 8372 23072 8424
rect 19248 8304 19300 8356
rect 24400 8304 24452 8356
rect 6504 8134 6556 8186
rect 6568 8134 6620 8186
rect 6632 8134 6684 8186
rect 6696 8134 6748 8186
rect 6760 8134 6812 8186
rect 17612 8134 17664 8186
rect 17676 8134 17728 8186
rect 17740 8134 17792 8186
rect 17804 8134 17856 8186
rect 17868 8134 17920 8186
rect 28720 8134 28772 8186
rect 28784 8134 28836 8186
rect 28848 8134 28900 8186
rect 28912 8134 28964 8186
rect 28976 8134 29028 8186
rect 39828 8134 39880 8186
rect 39892 8134 39944 8186
rect 39956 8134 40008 8186
rect 40020 8134 40072 8186
rect 40084 8134 40136 8186
rect 12058 7590 12110 7642
rect 12122 7590 12174 7642
rect 12186 7590 12238 7642
rect 12250 7590 12302 7642
rect 12314 7590 12366 7642
rect 23166 7590 23218 7642
rect 23230 7590 23282 7642
rect 23294 7590 23346 7642
rect 23358 7590 23410 7642
rect 23422 7590 23474 7642
rect 34274 7590 34326 7642
rect 34338 7590 34390 7642
rect 34402 7590 34454 7642
rect 34466 7590 34518 7642
rect 34530 7590 34582 7642
rect 45382 7590 45434 7642
rect 45446 7590 45498 7642
rect 45510 7590 45562 7642
rect 45574 7590 45626 7642
rect 45638 7590 45690 7642
rect 6504 7046 6556 7098
rect 6568 7046 6620 7098
rect 6632 7046 6684 7098
rect 6696 7046 6748 7098
rect 6760 7046 6812 7098
rect 17612 7046 17664 7098
rect 17676 7046 17728 7098
rect 17740 7046 17792 7098
rect 17804 7046 17856 7098
rect 17868 7046 17920 7098
rect 28720 7046 28772 7098
rect 28784 7046 28836 7098
rect 28848 7046 28900 7098
rect 28912 7046 28964 7098
rect 28976 7046 29028 7098
rect 39828 7046 39880 7098
rect 39892 7046 39944 7098
rect 39956 7046 40008 7098
rect 40020 7046 40072 7098
rect 40084 7046 40136 7098
rect 12058 6502 12110 6554
rect 12122 6502 12174 6554
rect 12186 6502 12238 6554
rect 12250 6502 12302 6554
rect 12314 6502 12366 6554
rect 23166 6502 23218 6554
rect 23230 6502 23282 6554
rect 23294 6502 23346 6554
rect 23358 6502 23410 6554
rect 23422 6502 23474 6554
rect 34274 6502 34326 6554
rect 34338 6502 34390 6554
rect 34402 6502 34454 6554
rect 34466 6502 34518 6554
rect 34530 6502 34582 6554
rect 45382 6502 45434 6554
rect 45446 6502 45498 6554
rect 45510 6502 45562 6554
rect 45574 6502 45626 6554
rect 45638 6502 45690 6554
rect 6504 5958 6556 6010
rect 6568 5958 6620 6010
rect 6632 5958 6684 6010
rect 6696 5958 6748 6010
rect 6760 5958 6812 6010
rect 17612 5958 17664 6010
rect 17676 5958 17728 6010
rect 17740 5958 17792 6010
rect 17804 5958 17856 6010
rect 17868 5958 17920 6010
rect 28720 5958 28772 6010
rect 28784 5958 28836 6010
rect 28848 5958 28900 6010
rect 28912 5958 28964 6010
rect 28976 5958 29028 6010
rect 39828 5958 39880 6010
rect 39892 5958 39944 6010
rect 39956 5958 40008 6010
rect 40020 5958 40072 6010
rect 40084 5958 40136 6010
rect 12058 5414 12110 5466
rect 12122 5414 12174 5466
rect 12186 5414 12238 5466
rect 12250 5414 12302 5466
rect 12314 5414 12366 5466
rect 23166 5414 23218 5466
rect 23230 5414 23282 5466
rect 23294 5414 23346 5466
rect 23358 5414 23410 5466
rect 23422 5414 23474 5466
rect 34274 5414 34326 5466
rect 34338 5414 34390 5466
rect 34402 5414 34454 5466
rect 34466 5414 34518 5466
rect 34530 5414 34582 5466
rect 45382 5414 45434 5466
rect 45446 5414 45498 5466
rect 45510 5414 45562 5466
rect 45574 5414 45626 5466
rect 45638 5414 45690 5466
rect 6504 4870 6556 4922
rect 6568 4870 6620 4922
rect 6632 4870 6684 4922
rect 6696 4870 6748 4922
rect 6760 4870 6812 4922
rect 17612 4870 17664 4922
rect 17676 4870 17728 4922
rect 17740 4870 17792 4922
rect 17804 4870 17856 4922
rect 17868 4870 17920 4922
rect 28720 4870 28772 4922
rect 28784 4870 28836 4922
rect 28848 4870 28900 4922
rect 28912 4870 28964 4922
rect 28976 4870 29028 4922
rect 39828 4870 39880 4922
rect 39892 4870 39944 4922
rect 39956 4870 40008 4922
rect 40020 4870 40072 4922
rect 40084 4870 40136 4922
rect 5540 4496 5592 4548
rect 24308 4496 24360 4548
rect 2320 4428 2372 4480
rect 26608 4428 26660 4480
rect 12058 4326 12110 4378
rect 12122 4326 12174 4378
rect 12186 4326 12238 4378
rect 12250 4326 12302 4378
rect 12314 4326 12366 4378
rect 23166 4326 23218 4378
rect 23230 4326 23282 4378
rect 23294 4326 23346 4378
rect 23358 4326 23410 4378
rect 23422 4326 23474 4378
rect 34274 4326 34326 4378
rect 34338 4326 34390 4378
rect 34402 4326 34454 4378
rect 34466 4326 34518 4378
rect 34530 4326 34582 4378
rect 45382 4326 45434 4378
rect 45446 4326 45498 4378
rect 45510 4326 45562 4378
rect 45574 4326 45626 4378
rect 45638 4326 45690 4378
rect 18512 4224 18564 4276
rect 42432 4224 42484 4276
rect 16948 4156 17000 4208
rect 41144 4156 41196 4208
rect 6504 3782 6556 3834
rect 6568 3782 6620 3834
rect 6632 3782 6684 3834
rect 6696 3782 6748 3834
rect 6760 3782 6812 3834
rect 17612 3782 17664 3834
rect 17676 3782 17728 3834
rect 17740 3782 17792 3834
rect 17804 3782 17856 3834
rect 17868 3782 17920 3834
rect 28720 3782 28772 3834
rect 28784 3782 28836 3834
rect 28848 3782 28900 3834
rect 28912 3782 28964 3834
rect 28976 3782 29028 3834
rect 39828 3782 39880 3834
rect 39892 3782 39944 3834
rect 39956 3782 40008 3834
rect 40020 3782 40072 3834
rect 40084 3782 40136 3834
rect 16212 3612 16264 3664
rect 35256 3612 35308 3664
rect 8116 3408 8168 3460
rect 22744 3476 22796 3528
rect 23020 3476 23072 3528
rect 25504 3476 25556 3528
rect 20444 3408 20496 3460
rect 28632 3408 28684 3460
rect 17500 3340 17552 3392
rect 25044 3340 25096 3392
rect 12058 3238 12110 3290
rect 12122 3238 12174 3290
rect 12186 3238 12238 3290
rect 12250 3238 12302 3290
rect 12314 3238 12366 3290
rect 23166 3238 23218 3290
rect 23230 3238 23282 3290
rect 23294 3238 23346 3290
rect 23358 3238 23410 3290
rect 23422 3238 23474 3290
rect 34274 3238 34326 3290
rect 34338 3238 34390 3290
rect 34402 3238 34454 3290
rect 34466 3238 34518 3290
rect 34530 3238 34582 3290
rect 45382 3238 45434 3290
rect 45446 3238 45498 3290
rect 45510 3238 45562 3290
rect 45574 3238 45626 3290
rect 45638 3238 45690 3290
rect 13636 3136 13688 3188
rect 19248 3136 19300 3188
rect 39672 3136 39724 3188
rect 12532 3068 12584 3120
rect 29092 3068 29144 3120
rect 8208 3000 8260 3052
rect 12992 2932 13044 2984
rect 14096 2864 14148 2916
rect 30104 3000 30156 3052
rect 16856 2796 16908 2848
rect 19432 2796 19484 2848
rect 22284 2796 22336 2848
rect 23480 2864 23532 2916
rect 23204 2839 23256 2848
rect 23204 2805 23213 2839
rect 23213 2805 23247 2839
rect 23247 2805 23256 2839
rect 23204 2796 23256 2805
rect 30288 2796 30340 2848
rect 32864 2796 32916 2848
rect 6504 2694 6556 2746
rect 6568 2694 6620 2746
rect 6632 2694 6684 2746
rect 6696 2694 6748 2746
rect 6760 2694 6812 2746
rect 17612 2694 17664 2746
rect 17676 2694 17728 2746
rect 17740 2694 17792 2746
rect 17804 2694 17856 2746
rect 17868 2694 17920 2746
rect 28720 2694 28772 2746
rect 28784 2694 28836 2746
rect 28848 2694 28900 2746
rect 28912 2694 28964 2746
rect 28976 2694 29028 2746
rect 39828 2694 39880 2746
rect 39892 2694 39944 2746
rect 39956 2694 40008 2746
rect 40020 2694 40072 2746
rect 40084 2694 40136 2746
rect 17040 2635 17092 2644
rect 17040 2601 17049 2635
rect 17049 2601 17083 2635
rect 17083 2601 17092 2635
rect 17040 2592 17092 2601
rect 19524 2592 19576 2644
rect 20628 2635 20680 2644
rect 20628 2601 20637 2635
rect 20637 2601 20671 2635
rect 20671 2601 20680 2635
rect 20628 2592 20680 2601
rect 21456 2592 21508 2644
rect 10968 2456 11020 2508
rect 18144 2524 18196 2576
rect 22008 2592 22060 2644
rect 22376 2635 22428 2644
rect 22376 2601 22385 2635
rect 22385 2601 22419 2635
rect 22419 2601 22428 2635
rect 22376 2592 22428 2601
rect 22744 2592 22796 2644
rect 23020 2592 23072 2644
rect 19800 2456 19852 2508
rect 22192 2456 22244 2508
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 18788 2431 18840 2440
rect 18788 2397 18797 2431
rect 18797 2397 18831 2431
rect 18831 2397 18840 2431
rect 18788 2388 18840 2397
rect 19156 2388 19208 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 19708 2388 19760 2440
rect 19892 2431 19944 2440
rect 19892 2397 19901 2431
rect 19901 2397 19935 2431
rect 19935 2397 19944 2431
rect 19892 2388 19944 2397
rect 11244 2320 11296 2372
rect 18052 2320 18104 2372
rect 18328 2320 18380 2372
rect 15292 2252 15344 2304
rect 18880 2252 18932 2304
rect 18972 2295 19024 2304
rect 18972 2261 18981 2295
rect 18981 2261 19015 2295
rect 19015 2261 19024 2295
rect 18972 2252 19024 2261
rect 19984 2252 20036 2304
rect 20168 2252 20220 2304
rect 20996 2252 21048 2304
rect 21364 2388 21416 2440
rect 21824 2431 21876 2440
rect 21824 2397 21833 2431
rect 21833 2397 21867 2431
rect 21867 2397 21876 2431
rect 21824 2388 21876 2397
rect 22100 2431 22152 2440
rect 22100 2397 22109 2431
rect 22109 2397 22143 2431
rect 22143 2397 22152 2431
rect 22100 2388 22152 2397
rect 22744 2456 22796 2508
rect 23112 2524 23164 2576
rect 23572 2524 23624 2576
rect 24400 2635 24452 2644
rect 24400 2601 24409 2635
rect 24409 2601 24443 2635
rect 24443 2601 24452 2635
rect 24400 2592 24452 2601
rect 25872 2592 25924 2644
rect 28080 2592 28132 2644
rect 29184 2635 29236 2644
rect 29184 2601 29193 2635
rect 29193 2601 29227 2635
rect 29227 2601 29236 2635
rect 29184 2592 29236 2601
rect 30380 2635 30432 2644
rect 30380 2601 30389 2635
rect 30389 2601 30423 2635
rect 30423 2601 30432 2635
rect 30380 2592 30432 2601
rect 30472 2592 30524 2644
rect 27896 2524 27948 2576
rect 30288 2524 30340 2576
rect 32496 2592 32548 2644
rect 34796 2635 34848 2644
rect 34796 2601 34805 2635
rect 34805 2601 34839 2635
rect 34839 2601 34848 2635
rect 34796 2592 34848 2601
rect 35072 2524 35124 2576
rect 36912 2592 36964 2644
rect 39028 2592 39080 2644
rect 41328 2635 41380 2644
rect 41328 2601 41337 2635
rect 41337 2601 41371 2635
rect 41371 2601 41380 2635
rect 41328 2592 41380 2601
rect 43536 2592 43588 2644
rect 44548 2635 44600 2644
rect 44548 2601 44557 2635
rect 44557 2601 44591 2635
rect 44591 2601 44600 2635
rect 44548 2592 44600 2601
rect 22192 2252 22244 2304
rect 22284 2295 22336 2304
rect 22284 2261 22293 2295
rect 22293 2261 22327 2295
rect 22327 2261 22336 2295
rect 22284 2252 22336 2261
rect 22652 2431 22704 2440
rect 22652 2397 22661 2431
rect 22661 2397 22695 2431
rect 22695 2397 22704 2431
rect 22652 2388 22704 2397
rect 23112 2431 23164 2440
rect 25780 2456 25832 2508
rect 30472 2456 30524 2508
rect 23112 2397 23129 2431
rect 23129 2397 23163 2431
rect 23163 2397 23164 2431
rect 23112 2388 23164 2397
rect 23204 2252 23256 2304
rect 23848 2388 23900 2440
rect 24124 2431 24176 2440
rect 24124 2397 24133 2431
rect 24133 2397 24167 2431
rect 24167 2397 24176 2431
rect 24124 2388 24176 2397
rect 24584 2431 24636 2440
rect 24584 2397 24593 2431
rect 24593 2397 24627 2431
rect 24627 2397 24636 2431
rect 24584 2388 24636 2397
rect 26148 2431 26200 2440
rect 26148 2397 26157 2431
rect 26157 2397 26191 2431
rect 26191 2397 26200 2431
rect 26148 2388 26200 2397
rect 27804 2431 27856 2440
rect 27804 2397 27813 2431
rect 27813 2397 27847 2431
rect 27847 2397 27856 2431
rect 27804 2388 27856 2397
rect 29184 2388 29236 2440
rect 32128 2456 32180 2508
rect 36636 2456 36688 2508
rect 40408 2524 40460 2576
rect 40684 2456 40736 2508
rect 23756 2363 23808 2372
rect 23756 2329 23765 2363
rect 23765 2329 23799 2363
rect 23799 2329 23808 2363
rect 23756 2320 23808 2329
rect 24216 2320 24268 2372
rect 29276 2320 29328 2372
rect 30656 2431 30708 2440
rect 30656 2397 30665 2431
rect 30665 2397 30699 2431
rect 30699 2397 30708 2431
rect 30656 2388 30708 2397
rect 30932 2431 30984 2440
rect 30932 2397 30941 2431
rect 30941 2397 30975 2431
rect 30975 2397 30984 2431
rect 30932 2388 30984 2397
rect 31208 2431 31260 2440
rect 31208 2397 31217 2431
rect 31217 2397 31251 2431
rect 31251 2397 31260 2431
rect 31208 2388 31260 2397
rect 32312 2388 32364 2440
rect 32772 2431 32824 2440
rect 32772 2397 32781 2431
rect 32781 2397 32815 2431
rect 32815 2397 32824 2431
rect 32772 2388 32824 2397
rect 34980 2431 35032 2440
rect 34980 2397 34989 2431
rect 34989 2397 35023 2431
rect 35023 2397 35032 2431
rect 34980 2388 35032 2397
rect 37188 2431 37240 2440
rect 37188 2397 37197 2431
rect 37197 2397 37231 2431
rect 37231 2397 37240 2431
rect 37188 2388 37240 2397
rect 39304 2431 39356 2440
rect 39304 2397 39313 2431
rect 39313 2397 39347 2431
rect 39347 2397 39356 2431
rect 39304 2388 39356 2397
rect 41512 2431 41564 2440
rect 41512 2397 41521 2431
rect 41521 2397 41555 2431
rect 41555 2397 41564 2431
rect 41512 2388 41564 2397
rect 43996 2431 44048 2440
rect 43996 2397 44005 2431
rect 44005 2397 44039 2431
rect 44039 2397 44048 2431
rect 43996 2388 44048 2397
rect 44364 2431 44416 2440
rect 44364 2397 44373 2431
rect 44373 2397 44407 2431
rect 44407 2397 44416 2431
rect 44364 2388 44416 2397
rect 45100 2388 45152 2440
rect 46112 2388 46164 2440
rect 43536 2320 43588 2372
rect 24032 2252 24084 2304
rect 30564 2252 30616 2304
rect 30840 2295 30892 2304
rect 30840 2261 30849 2295
rect 30849 2261 30883 2295
rect 30883 2261 30892 2295
rect 30840 2252 30892 2261
rect 31116 2295 31168 2304
rect 31116 2261 31125 2295
rect 31125 2261 31159 2295
rect 31159 2261 31168 2295
rect 31116 2252 31168 2261
rect 31944 2252 31996 2304
rect 32036 2252 32088 2304
rect 35072 2252 35124 2304
rect 35348 2252 35400 2304
rect 44180 2252 44232 2304
rect 44640 2295 44692 2304
rect 44640 2261 44649 2295
rect 44649 2261 44683 2295
rect 44683 2261 44692 2295
rect 44640 2252 44692 2261
rect 45008 2295 45060 2304
rect 45008 2261 45017 2295
rect 45017 2261 45051 2295
rect 45051 2261 45060 2295
rect 45008 2252 45060 2261
rect 12058 2150 12110 2202
rect 12122 2150 12174 2202
rect 12186 2150 12238 2202
rect 12250 2150 12302 2202
rect 12314 2150 12366 2202
rect 23166 2150 23218 2202
rect 23230 2150 23282 2202
rect 23294 2150 23346 2202
rect 23358 2150 23410 2202
rect 23422 2150 23474 2202
rect 34274 2150 34326 2202
rect 34338 2150 34390 2202
rect 34402 2150 34454 2202
rect 34466 2150 34518 2202
rect 34530 2150 34582 2202
rect 45382 2150 45434 2202
rect 45446 2150 45498 2202
rect 45510 2150 45562 2202
rect 45574 2150 45626 2202
rect 45638 2150 45690 2202
rect 480 1912 532 1964
rect 848 1844 900 1896
rect 2320 1955 2372 1964
rect 2320 1921 2329 1955
rect 2329 1921 2363 1955
rect 2363 1921 2372 1955
rect 2320 1912 2372 1921
rect 3148 1955 3200 1964
rect 3148 1921 3157 1955
rect 3157 1921 3191 1955
rect 3191 1921 3200 1955
rect 3148 1912 3200 1921
rect 2044 1887 2096 1896
rect 2044 1853 2053 1887
rect 2053 1853 2087 1887
rect 2087 1853 2096 1887
rect 2044 1844 2096 1853
rect 13820 2048 13872 2100
rect 7564 1980 7616 2032
rect 16212 2091 16264 2100
rect 16212 2057 16221 2091
rect 16221 2057 16255 2091
rect 16255 2057 16264 2091
rect 16212 2048 16264 2057
rect 16488 2091 16540 2100
rect 16488 2057 16497 2091
rect 16497 2057 16531 2091
rect 16531 2057 16540 2091
rect 16488 2048 16540 2057
rect 17132 2048 17184 2100
rect 17500 2048 17552 2100
rect 18144 2091 18196 2100
rect 18144 2057 18153 2091
rect 18153 2057 18187 2091
rect 18187 2057 18196 2091
rect 18144 2048 18196 2057
rect 19156 2048 19208 2100
rect 19248 2091 19300 2100
rect 19248 2057 19257 2091
rect 19257 2057 19291 2091
rect 19291 2057 19300 2091
rect 19248 2048 19300 2057
rect 19800 2048 19852 2100
rect 20812 2048 20864 2100
rect 20904 2091 20956 2100
rect 20904 2057 20913 2091
rect 20913 2057 20947 2091
rect 20947 2057 20956 2091
rect 20904 2048 20956 2057
rect 20996 2048 21048 2100
rect 17868 1980 17920 2032
rect 18052 1980 18104 2032
rect 23112 2048 23164 2100
rect 15016 1955 15068 1964
rect 15016 1921 15025 1955
rect 15025 1921 15059 1955
rect 15059 1921 15068 1955
rect 15016 1912 15068 1921
rect 15660 1912 15712 1964
rect 14832 1844 14884 1896
rect 15108 1844 15160 1896
rect 16028 1955 16080 1964
rect 16028 1921 16037 1955
rect 16037 1921 16071 1955
rect 16071 1921 16080 1955
rect 16028 1912 16080 1921
rect 16304 1955 16356 1964
rect 16304 1921 16313 1955
rect 16313 1921 16347 1955
rect 16347 1921 16356 1955
rect 16304 1912 16356 1921
rect 16488 1912 16540 1964
rect 17132 1955 17184 1964
rect 17132 1921 17141 1955
rect 17141 1921 17175 1955
rect 17175 1921 17184 1955
rect 17132 1912 17184 1921
rect 17408 1955 17460 1964
rect 17408 1921 17417 1955
rect 17417 1921 17451 1955
rect 17451 1921 17460 1955
rect 17408 1912 17460 1921
rect 17500 1912 17552 1964
rect 18144 1912 18196 1964
rect 18420 1912 18472 1964
rect 18512 1955 18564 1964
rect 18512 1921 18521 1955
rect 18521 1921 18555 1955
rect 18555 1921 18564 1955
rect 18512 1912 18564 1921
rect 18696 1912 18748 1964
rect 18788 1955 18840 1964
rect 18788 1921 18797 1955
rect 18797 1921 18831 1955
rect 18831 1921 18840 1955
rect 18788 1912 18840 1921
rect 18880 1912 18932 1964
rect 22192 1980 22244 2032
rect 23756 2048 23808 2100
rect 24124 2048 24176 2100
rect 26148 2048 26200 2100
rect 24584 1980 24636 2032
rect 24860 1980 24912 2032
rect 19524 1912 19576 1964
rect 19708 1912 19760 1964
rect 20260 1912 20312 1964
rect 20444 1955 20496 1964
rect 20444 1921 20453 1955
rect 20453 1921 20487 1955
rect 20487 1921 20496 1955
rect 20444 1912 20496 1921
rect 20720 1955 20772 1964
rect 20720 1921 20729 1955
rect 20729 1921 20763 1955
rect 20763 1921 20772 1955
rect 20720 1912 20772 1921
rect 21548 1912 21600 1964
rect 22468 1955 22520 1964
rect 22468 1921 22477 1955
rect 22477 1921 22511 1955
rect 22511 1921 22520 1955
rect 22468 1912 22520 1921
rect 22560 1912 22612 1964
rect 23572 1955 23624 1964
rect 23572 1921 23581 1955
rect 23581 1921 23615 1955
rect 23615 1921 23624 1955
rect 23572 1912 23624 1921
rect 16856 1776 16908 1828
rect 1584 1751 1636 1760
rect 1584 1717 1593 1751
rect 1593 1717 1627 1751
rect 1627 1717 1636 1751
rect 1584 1708 1636 1717
rect 15200 1751 15252 1760
rect 15200 1717 15209 1751
rect 15209 1717 15243 1751
rect 15243 1717 15252 1751
rect 15200 1708 15252 1717
rect 24032 1844 24084 1896
rect 24308 1955 24360 1964
rect 24308 1921 24317 1955
rect 24317 1921 24351 1955
rect 24351 1921 24360 1955
rect 24308 1912 24360 1921
rect 24676 1955 24728 1964
rect 24676 1921 24685 1955
rect 24685 1921 24719 1955
rect 24719 1921 24728 1955
rect 24676 1912 24728 1921
rect 25136 1955 25188 1964
rect 25136 1921 25145 1955
rect 25145 1921 25179 1955
rect 25179 1921 25188 1955
rect 25136 1912 25188 1921
rect 25504 1955 25556 1964
rect 25504 1921 25513 1955
rect 25513 1921 25547 1955
rect 25547 1921 25556 1955
rect 25504 1912 25556 1921
rect 26332 1955 26384 1964
rect 26332 1921 26341 1955
rect 26341 1921 26375 1955
rect 26375 1921 26384 1955
rect 26332 1912 26384 1921
rect 26608 1955 26660 1964
rect 26608 1921 26617 1955
rect 26617 1921 26651 1955
rect 26651 1921 26660 1955
rect 26608 1912 26660 1921
rect 26700 1912 26752 1964
rect 27068 1912 27120 1964
rect 27620 1912 27672 1964
rect 28172 1912 28224 1964
rect 28448 2048 28500 2100
rect 18052 1708 18104 1760
rect 18696 1708 18748 1760
rect 20996 1776 21048 1828
rect 19708 1708 19760 1760
rect 19800 1751 19852 1760
rect 19800 1717 19809 1751
rect 19809 1717 19843 1751
rect 19843 1717 19852 1751
rect 19800 1708 19852 1717
rect 20352 1751 20404 1760
rect 20352 1717 20361 1751
rect 20361 1717 20395 1751
rect 20395 1717 20404 1751
rect 20352 1708 20404 1717
rect 21180 1751 21232 1760
rect 21180 1717 21189 1751
rect 21189 1717 21223 1751
rect 21223 1717 21232 1751
rect 21180 1708 21232 1717
rect 23020 1776 23072 1828
rect 24952 1776 25004 1828
rect 25780 1776 25832 1828
rect 29092 1955 29144 1964
rect 29092 1921 29101 1955
rect 29101 1921 29135 1955
rect 29135 1921 29144 1955
rect 29092 1912 29144 1921
rect 29368 1955 29420 1964
rect 29368 1921 29377 1955
rect 29377 1921 29411 1955
rect 29411 1921 29420 1955
rect 29368 1912 29420 1921
rect 29644 1955 29696 1964
rect 29644 1921 29653 1955
rect 29653 1921 29687 1955
rect 29687 1921 29696 1955
rect 29644 1912 29696 1921
rect 29828 1912 29880 1964
rect 30840 2048 30892 2100
rect 30564 1955 30616 1964
rect 30564 1921 30573 1955
rect 30573 1921 30607 1955
rect 30607 1921 30616 1955
rect 30564 1912 30616 1921
rect 30840 1955 30892 1964
rect 30840 1921 30849 1955
rect 30849 1921 30883 1955
rect 30883 1921 30892 1955
rect 30840 1912 30892 1921
rect 31116 2048 31168 2100
rect 31852 2091 31904 2100
rect 31852 2057 31861 2091
rect 31861 2057 31895 2091
rect 31895 2057 31904 2091
rect 31852 2048 31904 2057
rect 32128 2091 32180 2100
rect 32128 2057 32137 2091
rect 32137 2057 32171 2091
rect 32171 2057 32180 2091
rect 32128 2048 32180 2057
rect 32772 2048 32824 2100
rect 34980 2048 35032 2100
rect 35256 2048 35308 2100
rect 32312 1955 32364 1964
rect 32312 1921 32321 1955
rect 32321 1921 32355 1955
rect 32355 1921 32364 1955
rect 32312 1912 32364 1921
rect 32864 1955 32916 1964
rect 32864 1921 32873 1955
rect 32873 1921 32907 1955
rect 32907 1921 32916 1955
rect 32864 1912 32916 1921
rect 36268 1980 36320 2032
rect 36636 2048 36688 2100
rect 37188 2048 37240 2100
rect 39304 2048 39356 2100
rect 40132 2091 40184 2100
rect 40132 2057 40141 2091
rect 40141 2057 40175 2091
rect 40175 2057 40184 2091
rect 40132 2048 40184 2057
rect 40408 2091 40460 2100
rect 40408 2057 40417 2091
rect 40417 2057 40451 2091
rect 40451 2057 40460 2091
rect 40408 2048 40460 2057
rect 40684 2091 40736 2100
rect 40684 2057 40693 2091
rect 40693 2057 40727 2091
rect 40727 2057 40736 2091
rect 40684 2048 40736 2057
rect 41512 2048 41564 2100
rect 43996 2048 44048 2100
rect 44640 2048 44692 2100
rect 45008 2048 45060 2100
rect 33508 1912 33560 1964
rect 34060 1912 34112 1964
rect 35348 1955 35400 1964
rect 35348 1921 35357 1955
rect 35357 1921 35391 1955
rect 35391 1921 35400 1955
rect 35348 1912 35400 1921
rect 35440 1955 35492 1964
rect 35440 1921 35449 1955
rect 35449 1921 35483 1955
rect 35483 1921 35492 1955
rect 35440 1912 35492 1921
rect 37924 1912 37976 1964
rect 38016 1955 38068 1964
rect 38016 1921 38025 1955
rect 38025 1921 38059 1955
rect 38059 1921 38068 1955
rect 38016 1912 38068 1921
rect 38384 1955 38436 1964
rect 38384 1921 38393 1955
rect 38393 1921 38427 1955
rect 38427 1921 38436 1955
rect 38384 1912 38436 1921
rect 39212 1844 39264 1896
rect 22100 1751 22152 1760
rect 22100 1717 22109 1751
rect 22109 1717 22143 1751
rect 22143 1717 22152 1751
rect 22100 1708 22152 1717
rect 22652 1751 22704 1760
rect 22652 1717 22661 1751
rect 22661 1717 22695 1751
rect 22695 1717 22704 1751
rect 22652 1708 22704 1717
rect 23756 1751 23808 1760
rect 23756 1717 23765 1751
rect 23765 1717 23799 1751
rect 23799 1717 23808 1751
rect 23756 1708 23808 1717
rect 24492 1751 24544 1760
rect 24492 1717 24501 1751
rect 24501 1717 24535 1751
rect 24535 1717 24544 1751
rect 24492 1708 24544 1717
rect 24860 1751 24912 1760
rect 24860 1717 24869 1751
rect 24869 1717 24903 1751
rect 24903 1717 24912 1751
rect 24860 1708 24912 1717
rect 26056 1708 26108 1760
rect 26148 1751 26200 1760
rect 26148 1717 26157 1751
rect 26157 1717 26191 1751
rect 26191 1717 26200 1751
rect 26148 1708 26200 1717
rect 26516 1751 26568 1760
rect 26516 1717 26525 1751
rect 26525 1717 26559 1751
rect 26559 1717 26568 1751
rect 26516 1708 26568 1717
rect 26792 1751 26844 1760
rect 26792 1717 26801 1751
rect 26801 1717 26835 1751
rect 26835 1717 26844 1751
rect 26792 1708 26844 1717
rect 27160 1751 27212 1760
rect 27160 1717 27169 1751
rect 27169 1717 27203 1751
rect 27203 1717 27212 1751
rect 27160 1708 27212 1717
rect 27252 1708 27304 1760
rect 29092 1776 29144 1828
rect 27712 1751 27764 1760
rect 27712 1717 27721 1751
rect 27721 1717 27755 1751
rect 27755 1717 27764 1751
rect 27712 1708 27764 1717
rect 27988 1751 28040 1760
rect 27988 1717 27997 1751
rect 27997 1717 28031 1751
rect 28031 1717 28040 1751
rect 27988 1708 28040 1717
rect 28080 1708 28132 1760
rect 29184 1708 29236 1760
rect 29276 1751 29328 1760
rect 29276 1717 29285 1751
rect 29285 1717 29319 1751
rect 29319 1717 29328 1751
rect 29276 1708 29328 1717
rect 29552 1751 29604 1760
rect 29552 1717 29561 1751
rect 29561 1717 29595 1751
rect 29595 1717 29604 1751
rect 29552 1708 29604 1717
rect 29828 1751 29880 1760
rect 29828 1717 29837 1751
rect 29837 1717 29871 1751
rect 29871 1717 29880 1751
rect 29828 1708 29880 1717
rect 30840 1776 30892 1828
rect 31852 1776 31904 1828
rect 30472 1751 30524 1760
rect 30472 1717 30481 1751
rect 30481 1717 30515 1751
rect 30515 1717 30524 1751
rect 30472 1708 30524 1717
rect 30748 1751 30800 1760
rect 30748 1717 30757 1751
rect 30757 1717 30791 1751
rect 30791 1717 30800 1751
rect 30748 1708 30800 1717
rect 31024 1751 31076 1760
rect 31024 1717 31033 1751
rect 31033 1717 31067 1751
rect 31067 1717 31076 1751
rect 31024 1708 31076 1717
rect 31300 1751 31352 1760
rect 31300 1717 31309 1751
rect 31309 1717 31343 1751
rect 31343 1717 31352 1751
rect 31300 1708 31352 1717
rect 31484 1708 31536 1760
rect 32404 1708 32456 1760
rect 33232 1776 33284 1828
rect 33508 1708 33560 1760
rect 33876 1751 33928 1760
rect 33876 1717 33885 1751
rect 33885 1717 33919 1751
rect 33919 1717 33928 1751
rect 33876 1708 33928 1717
rect 37648 1776 37700 1828
rect 34980 1708 35032 1760
rect 36452 1751 36504 1760
rect 36452 1717 36461 1751
rect 36461 1717 36495 1751
rect 36495 1717 36504 1751
rect 36452 1708 36504 1717
rect 37556 1708 37608 1760
rect 39580 1844 39632 1896
rect 40592 1955 40644 1964
rect 40592 1921 40601 1955
rect 40601 1921 40635 1955
rect 40635 1921 40644 1955
rect 40592 1912 40644 1921
rect 40500 1776 40552 1828
rect 44364 1912 44416 1964
rect 42524 1844 42576 1896
rect 45744 1912 45796 1964
rect 43812 1708 43864 1760
rect 6504 1606 6556 1658
rect 6568 1606 6620 1658
rect 6632 1606 6684 1658
rect 6696 1606 6748 1658
rect 6760 1606 6812 1658
rect 17612 1606 17664 1658
rect 17676 1606 17728 1658
rect 17740 1606 17792 1658
rect 17804 1606 17856 1658
rect 17868 1606 17920 1658
rect 28720 1606 28772 1658
rect 28784 1606 28836 1658
rect 28848 1606 28900 1658
rect 28912 1606 28964 1658
rect 28976 1606 29028 1658
rect 39828 1606 39880 1658
rect 39892 1606 39944 1658
rect 39956 1606 40008 1658
rect 40020 1606 40072 1658
rect 40084 1606 40136 1658
rect 1584 1504 1636 1556
rect 7564 1504 7616 1556
rect 15016 1504 15068 1556
rect 15108 1547 15160 1556
rect 15108 1513 15117 1547
rect 15117 1513 15151 1547
rect 15151 1513 15160 1547
rect 15108 1504 15160 1513
rect 15292 1504 15344 1556
rect 16028 1504 16080 1556
rect 16304 1504 16356 1556
rect 16488 1547 16540 1556
rect 16488 1513 16497 1547
rect 16497 1513 16531 1547
rect 16531 1513 16540 1547
rect 16488 1504 16540 1513
rect 17132 1504 17184 1556
rect 17224 1504 17276 1556
rect 17408 1504 17460 1556
rect 17500 1504 17552 1556
rect 18144 1504 18196 1556
rect 18420 1504 18472 1556
rect 18696 1504 18748 1556
rect 18788 1504 18840 1556
rect 1860 1479 1912 1488
rect 1860 1445 1869 1479
rect 1869 1445 1903 1479
rect 1903 1445 1912 1479
rect 1860 1436 1912 1445
rect 20904 1436 20956 1488
rect 1216 1300 1268 1352
rect 1676 1343 1728 1352
rect 1676 1309 1685 1343
rect 1685 1309 1719 1343
rect 1719 1309 1728 1343
rect 1676 1300 1728 1309
rect 2412 1343 2464 1352
rect 2412 1309 2421 1343
rect 2421 1309 2455 1343
rect 2455 1309 2464 1343
rect 2412 1300 2464 1309
rect 2504 1232 2556 1284
rect 3424 1343 3476 1352
rect 3424 1309 3433 1343
rect 3433 1309 3467 1343
rect 3467 1309 3476 1343
rect 3424 1300 3476 1309
rect 3884 1343 3936 1352
rect 3884 1309 3893 1343
rect 3893 1309 3927 1343
rect 3927 1309 3936 1343
rect 3884 1300 3936 1309
rect 4252 1343 4304 1352
rect 4252 1309 4261 1343
rect 4261 1309 4295 1343
rect 4295 1309 4304 1343
rect 4252 1300 4304 1309
rect 4620 1343 4672 1352
rect 4620 1309 4629 1343
rect 4629 1309 4663 1343
rect 4663 1309 4672 1343
rect 4620 1300 4672 1309
rect 4988 1343 5040 1352
rect 4988 1309 4997 1343
rect 4997 1309 5031 1343
rect 5031 1309 5040 1343
rect 4988 1300 5040 1309
rect 5356 1343 5408 1352
rect 5356 1309 5365 1343
rect 5365 1309 5399 1343
rect 5399 1309 5408 1343
rect 5356 1300 5408 1309
rect 5724 1343 5776 1352
rect 5724 1309 5733 1343
rect 5733 1309 5767 1343
rect 5767 1309 5776 1343
rect 5724 1300 5776 1309
rect 6000 1343 6052 1352
rect 6000 1309 6009 1343
rect 6009 1309 6043 1343
rect 6043 1309 6052 1343
rect 6000 1300 6052 1309
rect 6460 1343 6512 1352
rect 6460 1309 6469 1343
rect 6469 1309 6503 1343
rect 6503 1309 6512 1343
rect 6460 1300 6512 1309
rect 6828 1343 6880 1352
rect 6828 1309 6837 1343
rect 6837 1309 6871 1343
rect 6871 1309 6880 1343
rect 6828 1300 6880 1309
rect 7196 1343 7248 1352
rect 7196 1309 7205 1343
rect 7205 1309 7239 1343
rect 7239 1309 7248 1343
rect 7196 1300 7248 1309
rect 7564 1343 7616 1352
rect 7564 1309 7573 1343
rect 7573 1309 7607 1343
rect 7607 1309 7616 1343
rect 7564 1300 7616 1309
rect 7932 1343 7984 1352
rect 7932 1309 7941 1343
rect 7941 1309 7975 1343
rect 7975 1309 7984 1343
rect 7932 1300 7984 1309
rect 1584 1207 1636 1216
rect 1584 1173 1593 1207
rect 1593 1173 1627 1207
rect 1627 1173 1636 1207
rect 1584 1164 1636 1173
rect 4712 1232 4764 1284
rect 8116 1300 8168 1352
rect 8208 1300 8260 1352
rect 8300 1343 8352 1352
rect 8300 1309 8309 1343
rect 8309 1309 8343 1343
rect 8343 1309 8352 1343
rect 8300 1300 8352 1309
rect 8576 1343 8628 1352
rect 8576 1309 8585 1343
rect 8585 1309 8619 1343
rect 8619 1309 8628 1343
rect 8576 1300 8628 1309
rect 9036 1343 9088 1352
rect 9036 1309 9045 1343
rect 9045 1309 9079 1343
rect 9079 1309 9088 1343
rect 9036 1300 9088 1309
rect 9404 1343 9456 1352
rect 9404 1309 9413 1343
rect 9413 1309 9447 1343
rect 9447 1309 9456 1343
rect 9404 1300 9456 1309
rect 9772 1343 9824 1352
rect 9772 1309 9781 1343
rect 9781 1309 9815 1343
rect 9815 1309 9824 1343
rect 9772 1300 9824 1309
rect 10140 1343 10192 1352
rect 10140 1309 10149 1343
rect 10149 1309 10183 1343
rect 10183 1309 10192 1343
rect 10140 1300 10192 1309
rect 10508 1343 10560 1352
rect 10508 1309 10517 1343
rect 10517 1309 10551 1343
rect 10551 1309 10560 1343
rect 10508 1300 10560 1309
rect 10876 1343 10928 1352
rect 10876 1309 10885 1343
rect 10885 1309 10919 1343
rect 10919 1309 10928 1343
rect 10876 1300 10928 1309
rect 11152 1343 11204 1352
rect 11152 1309 11161 1343
rect 11161 1309 11195 1343
rect 11195 1309 11204 1343
rect 11152 1300 11204 1309
rect 11612 1343 11664 1352
rect 11612 1309 11621 1343
rect 11621 1309 11655 1343
rect 11655 1309 11664 1343
rect 11612 1300 11664 1309
rect 11980 1343 12032 1352
rect 11980 1309 11989 1343
rect 11989 1309 12023 1343
rect 12023 1309 12032 1343
rect 11980 1300 12032 1309
rect 3608 1207 3660 1216
rect 3608 1173 3617 1207
rect 3617 1173 3651 1207
rect 3651 1173 3660 1207
rect 3608 1164 3660 1173
rect 3792 1164 3844 1216
rect 4068 1207 4120 1216
rect 4068 1173 4077 1207
rect 4077 1173 4111 1207
rect 4111 1173 4120 1207
rect 4068 1164 4120 1173
rect 4436 1207 4488 1216
rect 4436 1173 4445 1207
rect 4445 1173 4479 1207
rect 4479 1173 4488 1207
rect 4436 1164 4488 1173
rect 5172 1207 5224 1216
rect 5172 1173 5181 1207
rect 5181 1173 5215 1207
rect 5215 1173 5224 1207
rect 5172 1164 5224 1173
rect 5816 1164 5868 1216
rect 5908 1207 5960 1216
rect 5908 1173 5917 1207
rect 5917 1173 5951 1207
rect 5951 1173 5960 1207
rect 5908 1164 5960 1173
rect 6092 1164 6144 1216
rect 6644 1207 6696 1216
rect 6644 1173 6653 1207
rect 6653 1173 6687 1207
rect 6687 1173 6696 1207
rect 6644 1164 6696 1173
rect 7012 1207 7064 1216
rect 7012 1173 7021 1207
rect 7021 1173 7055 1207
rect 7055 1173 7064 1207
rect 7012 1164 7064 1173
rect 7656 1164 7708 1216
rect 7748 1207 7800 1216
rect 7748 1173 7757 1207
rect 7757 1173 7791 1207
rect 7791 1173 7800 1207
rect 7748 1164 7800 1173
rect 10416 1232 10468 1284
rect 12164 1300 12216 1352
rect 12532 1300 12584 1352
rect 12624 1343 12676 1352
rect 12624 1309 12633 1343
rect 12633 1309 12667 1343
rect 12667 1309 12676 1343
rect 12624 1300 12676 1309
rect 12900 1343 12952 1352
rect 12900 1309 12909 1343
rect 12909 1309 12943 1343
rect 12943 1309 12952 1343
rect 12900 1300 12952 1309
rect 13176 1343 13228 1352
rect 13176 1309 13185 1343
rect 13185 1309 13219 1343
rect 13219 1309 13228 1343
rect 13176 1300 13228 1309
rect 13452 1343 13504 1352
rect 13452 1309 13461 1343
rect 13461 1309 13495 1343
rect 13495 1309 13504 1343
rect 13452 1300 13504 1309
rect 13728 1343 13780 1352
rect 13728 1309 13737 1343
rect 13737 1309 13771 1343
rect 13771 1309 13780 1343
rect 13728 1300 13780 1309
rect 14004 1300 14056 1352
rect 14556 1300 14608 1352
rect 8760 1207 8812 1216
rect 8760 1173 8769 1207
rect 8769 1173 8803 1207
rect 8803 1173 8812 1207
rect 8760 1164 8812 1173
rect 9220 1207 9272 1216
rect 9220 1173 9229 1207
rect 9229 1173 9263 1207
rect 9263 1173 9272 1207
rect 9220 1164 9272 1173
rect 9588 1207 9640 1216
rect 9588 1173 9597 1207
rect 9597 1173 9631 1207
rect 9631 1173 9640 1207
rect 9588 1164 9640 1173
rect 9956 1207 10008 1216
rect 9956 1173 9965 1207
rect 9965 1173 9999 1207
rect 9999 1173 10008 1207
rect 9956 1164 10008 1173
rect 10324 1207 10376 1216
rect 10324 1173 10333 1207
rect 10333 1173 10367 1207
rect 10367 1173 10376 1207
rect 10324 1164 10376 1173
rect 10692 1207 10744 1216
rect 10692 1173 10701 1207
rect 10701 1173 10735 1207
rect 10735 1173 10744 1207
rect 10692 1164 10744 1173
rect 11060 1207 11112 1216
rect 11060 1173 11069 1207
rect 11069 1173 11103 1207
rect 11103 1173 11112 1207
rect 11060 1164 11112 1173
rect 11336 1207 11388 1216
rect 11336 1173 11345 1207
rect 11345 1173 11379 1207
rect 11379 1173 11388 1207
rect 11336 1164 11388 1173
rect 12532 1207 12584 1216
rect 12532 1173 12541 1207
rect 12541 1173 12575 1207
rect 12575 1173 12584 1207
rect 12532 1164 12584 1173
rect 12808 1207 12860 1216
rect 12808 1173 12817 1207
rect 12817 1173 12851 1207
rect 12851 1173 12860 1207
rect 12808 1164 12860 1173
rect 13084 1207 13136 1216
rect 13084 1173 13093 1207
rect 13093 1173 13127 1207
rect 13127 1173 13136 1207
rect 13084 1164 13136 1173
rect 13268 1164 13320 1216
rect 13912 1207 13964 1216
rect 13912 1173 13921 1207
rect 13921 1173 13955 1207
rect 13955 1173 13964 1207
rect 13912 1164 13964 1173
rect 14464 1232 14516 1284
rect 15108 1300 15160 1352
rect 15384 1300 15436 1352
rect 17132 1368 17184 1420
rect 15016 1232 15068 1284
rect 15844 1300 15896 1352
rect 15936 1300 15988 1352
rect 16028 1343 16080 1352
rect 16028 1309 16037 1343
rect 16037 1309 16071 1343
rect 16071 1309 16080 1343
rect 16028 1300 16080 1309
rect 16488 1300 16540 1352
rect 16764 1343 16816 1352
rect 16764 1309 16773 1343
rect 16773 1309 16807 1343
rect 16807 1309 16816 1343
rect 16764 1300 16816 1309
rect 14096 1164 14148 1216
rect 17316 1300 17368 1352
rect 17500 1343 17552 1352
rect 17500 1309 17509 1343
rect 17509 1309 17543 1343
rect 17543 1309 17552 1343
rect 17500 1300 17552 1309
rect 18236 1343 18288 1352
rect 18236 1309 18245 1343
rect 18245 1309 18279 1343
rect 18279 1309 18288 1343
rect 18236 1300 18288 1309
rect 18512 1343 18564 1352
rect 18512 1309 18521 1343
rect 18521 1309 18555 1343
rect 18555 1309 18564 1343
rect 18512 1300 18564 1309
rect 18788 1343 18840 1352
rect 18788 1309 18797 1343
rect 18797 1309 18831 1343
rect 18831 1309 18840 1343
rect 18788 1300 18840 1309
rect 18880 1300 18932 1352
rect 18972 1300 19024 1352
rect 19064 1343 19116 1352
rect 19064 1309 19073 1343
rect 19073 1309 19107 1343
rect 19107 1309 19116 1343
rect 19064 1300 19116 1309
rect 19800 1300 19852 1352
rect 19984 1300 20036 1352
rect 21456 1300 21508 1352
rect 22284 1436 22336 1488
rect 22468 1411 22520 1420
rect 22468 1377 22477 1411
rect 22477 1377 22511 1411
rect 22511 1377 22520 1411
rect 22468 1368 22520 1377
rect 23572 1411 23624 1420
rect 23572 1377 23581 1411
rect 23581 1377 23615 1411
rect 23615 1377 23624 1411
rect 23572 1368 23624 1377
rect 24492 1436 24544 1488
rect 24768 1504 24820 1556
rect 25412 1504 25464 1556
rect 27252 1504 27304 1556
rect 27344 1504 27396 1556
rect 28816 1504 28868 1556
rect 30012 1504 30064 1556
rect 31852 1504 31904 1556
rect 32772 1504 32824 1556
rect 20168 1232 20220 1284
rect 20904 1232 20956 1284
rect 24860 1368 24912 1420
rect 26424 1411 26476 1420
rect 26424 1377 26433 1411
rect 26433 1377 26467 1411
rect 26467 1377 26476 1411
rect 26424 1368 26476 1377
rect 26884 1368 26936 1420
rect 28172 1368 28224 1420
rect 28448 1368 28500 1420
rect 29552 1368 29604 1420
rect 26516 1300 26568 1352
rect 26792 1300 26844 1352
rect 27160 1300 27212 1352
rect 27712 1300 27764 1352
rect 27988 1300 28040 1352
rect 29184 1343 29236 1352
rect 29184 1309 29193 1343
rect 29193 1309 29227 1343
rect 29227 1309 29236 1343
rect 29184 1300 29236 1309
rect 29276 1300 29328 1352
rect 30380 1368 30432 1420
rect 32956 1436 33008 1488
rect 34060 1504 34112 1556
rect 34244 1504 34296 1556
rect 34704 1436 34756 1488
rect 35808 1504 35860 1556
rect 35716 1436 35768 1488
rect 37004 1504 37056 1556
rect 38292 1504 38344 1556
rect 39212 1504 39264 1556
rect 42432 1547 42484 1556
rect 42432 1513 42441 1547
rect 42441 1513 42475 1547
rect 42475 1513 42484 1547
rect 42432 1504 42484 1513
rect 42524 1504 42576 1556
rect 37372 1436 37424 1488
rect 38844 1436 38896 1488
rect 35808 1368 35860 1420
rect 37924 1368 37976 1420
rect 19708 1207 19760 1216
rect 19708 1173 19717 1207
rect 19717 1173 19751 1207
rect 19751 1173 19760 1207
rect 19708 1164 19760 1173
rect 20076 1207 20128 1216
rect 20076 1173 20085 1207
rect 20085 1173 20119 1207
rect 20119 1173 20128 1207
rect 20076 1164 20128 1173
rect 20444 1207 20496 1216
rect 20444 1173 20453 1207
rect 20453 1173 20487 1207
rect 20487 1173 20496 1207
rect 20444 1164 20496 1173
rect 20812 1207 20864 1216
rect 20812 1173 20821 1207
rect 20821 1173 20855 1207
rect 20855 1173 20864 1207
rect 20812 1164 20864 1173
rect 21548 1207 21600 1216
rect 21548 1173 21557 1207
rect 21557 1173 21591 1207
rect 21591 1173 21600 1207
rect 21548 1164 21600 1173
rect 23112 1232 23164 1284
rect 24584 1232 24636 1284
rect 23020 1207 23072 1216
rect 23020 1173 23029 1207
rect 23029 1173 23063 1207
rect 23063 1173 23072 1207
rect 23020 1164 23072 1173
rect 24124 1207 24176 1216
rect 24124 1173 24133 1207
rect 24133 1173 24167 1207
rect 24167 1173 24176 1207
rect 24124 1164 24176 1173
rect 24676 1207 24728 1216
rect 24676 1173 24685 1207
rect 24685 1173 24719 1207
rect 24719 1173 24728 1207
rect 24676 1164 24728 1173
rect 24952 1275 25004 1284
rect 24952 1241 24961 1275
rect 24961 1241 24995 1275
rect 24995 1241 25004 1275
rect 24952 1232 25004 1241
rect 25136 1164 25188 1216
rect 25688 1164 25740 1216
rect 26608 1164 26660 1216
rect 27252 1164 27304 1216
rect 27712 1164 27764 1216
rect 29552 1232 29604 1284
rect 30472 1300 30524 1352
rect 30748 1300 30800 1352
rect 31024 1300 31076 1352
rect 31944 1300 31996 1352
rect 35164 1300 35216 1352
rect 37096 1300 37148 1352
rect 33324 1275 33376 1284
rect 33324 1241 33333 1275
rect 33333 1241 33367 1275
rect 33367 1241 33376 1275
rect 33324 1232 33376 1241
rect 33416 1232 33468 1284
rect 34796 1275 34848 1284
rect 34796 1241 34805 1275
rect 34805 1241 34839 1275
rect 34839 1241 34848 1275
rect 34796 1232 34848 1241
rect 34888 1232 34940 1284
rect 35440 1232 35492 1284
rect 37464 1232 37516 1284
rect 37832 1232 37884 1284
rect 38108 1232 38160 1284
rect 38752 1300 38804 1352
rect 39212 1232 39264 1284
rect 41144 1343 41196 1352
rect 41144 1309 41153 1343
rect 41153 1309 41187 1343
rect 41187 1309 41196 1343
rect 41144 1300 41196 1309
rect 41236 1300 41288 1352
rect 41972 1343 42024 1352
rect 41972 1309 41981 1343
rect 41981 1309 42015 1343
rect 42015 1309 42024 1343
rect 41972 1300 42024 1309
rect 42708 1368 42760 1420
rect 43536 1479 43588 1488
rect 43536 1445 43545 1479
rect 43545 1445 43579 1479
rect 43579 1445 43588 1479
rect 43536 1436 43588 1445
rect 43812 1479 43864 1488
rect 43812 1445 43821 1479
rect 43821 1445 43855 1479
rect 43855 1445 43864 1479
rect 43812 1436 43864 1445
rect 44180 1436 44232 1488
rect 29644 1164 29696 1216
rect 31760 1164 31812 1216
rect 32956 1164 33008 1216
rect 39304 1164 39356 1216
rect 39396 1164 39448 1216
rect 39672 1164 39724 1216
rect 41328 1232 41380 1284
rect 41696 1232 41748 1284
rect 40040 1164 40092 1216
rect 42064 1207 42116 1216
rect 42064 1173 42073 1207
rect 42073 1173 42107 1207
rect 42107 1173 42116 1207
rect 42064 1164 42116 1173
rect 42340 1164 42392 1216
rect 42800 1232 42852 1284
rect 43352 1232 43404 1284
rect 43628 1232 43680 1284
rect 44272 1343 44324 1352
rect 44272 1309 44281 1343
rect 44281 1309 44315 1343
rect 44315 1309 44324 1343
rect 44272 1300 44324 1309
rect 44548 1343 44600 1352
rect 44548 1309 44557 1343
rect 44557 1309 44591 1343
rect 44591 1309 44600 1343
rect 44548 1300 44600 1309
rect 44824 1343 44876 1352
rect 44824 1309 44833 1343
rect 44833 1309 44867 1343
rect 44867 1309 44876 1343
rect 44824 1300 44876 1309
rect 44732 1232 44784 1284
rect 42524 1164 42576 1216
rect 42984 1207 43036 1216
rect 42984 1173 42993 1207
rect 42993 1173 43027 1207
rect 43027 1173 43036 1207
rect 42984 1164 43036 1173
rect 43076 1164 43128 1216
rect 44088 1207 44140 1216
rect 44088 1173 44097 1207
rect 44097 1173 44131 1207
rect 44131 1173 44140 1207
rect 44088 1164 44140 1173
rect 12058 1062 12110 1114
rect 12122 1062 12174 1114
rect 12186 1062 12238 1114
rect 12250 1062 12302 1114
rect 12314 1062 12366 1114
rect 23166 1062 23218 1114
rect 23230 1062 23282 1114
rect 23294 1062 23346 1114
rect 23358 1062 23410 1114
rect 23422 1062 23474 1114
rect 34274 1062 34326 1114
rect 34338 1062 34390 1114
rect 34402 1062 34454 1114
rect 34466 1062 34518 1114
rect 34530 1062 34582 1114
rect 45382 1062 45434 1114
rect 45446 1062 45498 1114
rect 45510 1062 45562 1114
rect 45574 1062 45626 1114
rect 45638 1062 45690 1114
rect 3608 960 3660 1012
rect 5540 960 5592 1012
rect 6644 960 6696 1012
rect 10968 960 11020 1012
rect 11336 960 11388 1012
rect 24584 960 24636 1012
rect 4436 892 4488 944
rect 5172 892 5224 944
rect 5908 824 5960 876
rect 9864 824 9916 876
rect 9956 824 10008 876
rect 10416 824 10468 876
rect 5816 688 5868 740
rect 6092 756 6144 808
rect 8944 756 8996 808
rect 13084 892 13136 944
rect 17684 892 17736 944
rect 25412 960 25464 1012
rect 27528 960 27580 1012
rect 30380 960 30432 1012
rect 30656 960 30708 1012
rect 31392 960 31444 1012
rect 35440 960 35492 1012
rect 12992 756 13044 808
rect 13084 756 13136 808
rect 13360 756 13412 808
rect 16764 756 16816 808
rect 17408 756 17460 808
rect 17868 824 17920 876
rect 30104 892 30156 944
rect 40040 960 40092 1012
rect 40592 960 40644 1012
rect 41972 960 42024 1012
rect 42524 960 42576 1012
rect 43076 960 43128 1012
rect 39304 892 39356 944
rect 27068 824 27120 876
rect 25780 756 25832 808
rect 17316 688 17368 740
rect 39396 756 39448 808
rect 42064 756 42116 808
rect 42984 756 43036 808
rect 28632 688 28684 740
rect 32956 688 33008 740
rect 7012 416 7064 468
rect 1584 212 1636 264
rect 11060 552 11112 604
rect 7748 484 7800 536
rect 11244 484 11296 536
rect 15752 552 15804 604
rect 17040 552 17092 604
rect 27804 620 27856 672
rect 27896 620 27948 672
rect 23572 552 23624 604
rect 29000 552 29052 604
rect 33416 552 33468 604
rect 28356 484 28408 536
rect 12072 416 12124 468
rect 14004 416 14056 468
rect 17684 416 17736 468
rect 20260 416 20312 468
rect 25228 416 25280 468
rect 7656 348 7708 400
rect 13636 348 13688 400
rect 13912 348 13964 400
rect 12532 280 12584 332
rect 12716 212 12768 264
rect 13268 212 13320 264
rect 26700 280 26752 332
rect 26884 280 26936 332
rect 28540 348 28592 400
rect 29000 348 29052 400
rect 34888 348 34940 400
rect 36268 348 36320 400
rect 44088 348 44140 400
rect 33324 280 33376 332
rect 26056 212 26108 264
rect 18328 144 18380 196
rect 25044 144 25096 196
rect 11704 76 11756 128
rect 11796 76 11848 128
rect 12072 76 12124 128
rect 4068 8 4120 60
rect 23572 76 23624 128
rect 30380 76 30432 128
rect 13084 8 13136 60
<< metal2 >>
rect 1214 9840 1270 10300
rect 3422 9840 3478 10300
rect 5630 9840 5686 10300
rect 7838 9840 7894 10300
rect 10046 9840 10102 10300
rect 11992 9846 12204 9874
rect 1228 9058 1256 9840
rect 1228 9030 1440 9058
rect 1412 8566 1440 9030
rect 3436 8634 3464 9840
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 4080 8498 4108 8774
rect 5644 8634 5672 9840
rect 7852 8634 7880 9840
rect 8208 8900 8260 8906
rect 8208 8842 8260 8848
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8220 8498 8248 8842
rect 10060 8634 10088 9840
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 11992 8548 12020 9846
rect 12176 9738 12204 9846
rect 12254 9840 12310 10300
rect 14462 9840 14518 10300
rect 16670 9840 16726 10300
rect 18878 9840 18934 10300
rect 21086 9840 21142 10300
rect 23032 9846 23244 9874
rect 12268 9738 12296 9840
rect 12176 9710 12296 9738
rect 12058 8732 12366 8741
rect 12058 8730 12064 8732
rect 12120 8730 12144 8732
rect 12200 8730 12224 8732
rect 12280 8730 12304 8732
rect 12360 8730 12366 8732
rect 12120 8678 12122 8730
rect 12302 8678 12304 8730
rect 12058 8676 12064 8678
rect 12120 8676 12144 8678
rect 12200 8676 12224 8678
rect 12280 8676 12304 8678
rect 12360 8676 12366 8678
rect 12058 8667 12366 8676
rect 14476 8634 14504 9840
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 16684 8566 16712 9840
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17328 8634 17356 8910
rect 18892 8634 18920 9840
rect 21100 8634 21128 9840
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 12164 8560 12216 8566
rect 11992 8520 12164 8548
rect 12164 8502 12216 8508
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 20628 8560 20680 8566
rect 20628 8502 20680 8508
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 6504 8188 6812 8197
rect 6504 8186 6510 8188
rect 6566 8186 6590 8188
rect 6646 8186 6670 8188
rect 6726 8186 6750 8188
rect 6806 8186 6812 8188
rect 6566 8134 6568 8186
rect 6748 8134 6750 8186
rect 6504 8132 6510 8134
rect 6566 8132 6590 8134
rect 6646 8132 6670 8134
rect 6726 8132 6750 8134
rect 6806 8132 6812 8134
rect 6504 8123 6812 8132
rect 12058 7644 12366 7653
rect 12058 7642 12064 7644
rect 12120 7642 12144 7644
rect 12200 7642 12224 7644
rect 12280 7642 12304 7644
rect 12360 7642 12366 7644
rect 12120 7590 12122 7642
rect 12302 7590 12304 7642
rect 12058 7588 12064 7590
rect 12120 7588 12144 7590
rect 12200 7588 12224 7590
rect 12280 7588 12304 7590
rect 12360 7588 12366 7590
rect 12058 7579 12366 7588
rect 6504 7100 6812 7109
rect 6504 7098 6510 7100
rect 6566 7098 6590 7100
rect 6646 7098 6670 7100
rect 6726 7098 6750 7100
rect 6806 7098 6812 7100
rect 6566 7046 6568 7098
rect 6748 7046 6750 7098
rect 6504 7044 6510 7046
rect 6566 7044 6590 7046
rect 6646 7044 6670 7046
rect 6726 7044 6750 7046
rect 6806 7044 6812 7046
rect 6504 7035 6812 7044
rect 12058 6556 12366 6565
rect 12058 6554 12064 6556
rect 12120 6554 12144 6556
rect 12200 6554 12224 6556
rect 12280 6554 12304 6556
rect 12360 6554 12366 6556
rect 12120 6502 12122 6554
rect 12302 6502 12304 6554
rect 12058 6500 12064 6502
rect 12120 6500 12144 6502
rect 12200 6500 12224 6502
rect 12280 6500 12304 6502
rect 12360 6500 12366 6502
rect 12058 6491 12366 6500
rect 6504 6012 6812 6021
rect 6504 6010 6510 6012
rect 6566 6010 6590 6012
rect 6646 6010 6670 6012
rect 6726 6010 6750 6012
rect 6806 6010 6812 6012
rect 6566 5958 6568 6010
rect 6748 5958 6750 6010
rect 6504 5956 6510 5958
rect 6566 5956 6590 5958
rect 6646 5956 6670 5958
rect 6726 5956 6750 5958
rect 6806 5956 6812 5958
rect 6504 5947 6812 5956
rect 12058 5468 12366 5477
rect 12058 5466 12064 5468
rect 12120 5466 12144 5468
rect 12200 5466 12224 5468
rect 12280 5466 12304 5468
rect 12360 5466 12366 5468
rect 12120 5414 12122 5466
rect 12302 5414 12304 5466
rect 12058 5412 12064 5414
rect 12120 5412 12144 5414
rect 12200 5412 12224 5414
rect 12280 5412 12304 5414
rect 12360 5412 12366 5414
rect 12058 5403 12366 5412
rect 6504 4924 6812 4933
rect 6504 4922 6510 4924
rect 6566 4922 6590 4924
rect 6646 4922 6670 4924
rect 6726 4922 6750 4924
rect 6806 4922 6812 4924
rect 6566 4870 6568 4922
rect 6748 4870 6750 4922
rect 6504 4868 6510 4870
rect 6566 4868 6590 4870
rect 6646 4868 6670 4870
rect 6726 4868 6750 4870
rect 6806 4868 6812 4870
rect 6504 4859 6812 4868
rect 4710 4584 4766 4593
rect 4710 4519 4766 4528
rect 5540 4548 5592 4554
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 1858 2544 1914 2553
rect 1858 2479 1914 2488
rect 480 1964 532 1970
rect 480 1906 532 1912
rect 492 160 520 1906
rect 848 1896 900 1902
rect 848 1838 900 1844
rect 860 160 888 1838
rect 1584 1760 1636 1766
rect 1584 1702 1636 1708
rect 1596 1562 1624 1702
rect 1584 1556 1636 1562
rect 1584 1498 1636 1504
rect 1872 1494 1900 2479
rect 2332 1970 2360 4422
rect 3790 4176 3846 4185
rect 3790 4111 3846 4120
rect 2320 1964 2372 1970
rect 2320 1906 2372 1912
rect 3148 1964 3200 1970
rect 3148 1906 3200 1912
rect 2044 1896 2096 1902
rect 2044 1838 2096 1844
rect 1860 1488 1912 1494
rect 1860 1430 1912 1436
rect 1216 1352 1268 1358
rect 1216 1294 1268 1300
rect 1676 1352 1728 1358
rect 1676 1294 1728 1300
rect 1228 160 1256 1294
rect 1584 1216 1636 1222
rect 1584 1158 1636 1164
rect 1596 270 1624 1158
rect 1584 264 1636 270
rect 1584 206 1636 212
rect 478 -300 534 160
rect 846 -300 902 160
rect 1214 -300 1270 160
rect 1582 82 1638 160
rect 1688 82 1716 1294
rect 1582 54 1716 82
rect 1950 82 2006 160
rect 2056 82 2084 1838
rect 2412 1352 2464 1358
rect 2412 1294 2464 1300
rect 1950 54 2084 82
rect 2318 82 2374 160
rect 2424 82 2452 1294
rect 2504 1284 2556 1290
rect 2504 1226 2556 1232
rect 2318 54 2452 82
rect 2516 82 2544 1226
rect 2686 82 2742 160
rect 2516 54 2742 82
rect 1582 -300 1638 54
rect 1950 -300 2006 54
rect 2318 -300 2374 54
rect 2686 -300 2742 54
rect 3054 82 3110 160
rect 3160 82 3188 1906
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 3436 160 3464 1294
rect 3804 1222 3832 4111
rect 3884 1352 3936 1358
rect 3884 1294 3936 1300
rect 4252 1352 4304 1358
rect 4252 1294 4304 1300
rect 4620 1352 4672 1358
rect 4620 1294 4672 1300
rect 3608 1216 3660 1222
rect 3608 1158 3660 1164
rect 3792 1216 3844 1222
rect 3792 1158 3844 1164
rect 3620 1018 3648 1158
rect 3608 1012 3660 1018
rect 3608 954 3660 960
rect 3054 54 3188 82
rect 3054 -300 3110 54
rect 3422 -300 3478 160
rect 3790 82 3846 160
rect 3896 82 3924 1294
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 3790 54 3924 82
rect 4080 66 4108 1158
rect 4158 82 4214 160
rect 4264 82 4292 1294
rect 4436 1216 4488 1222
rect 4436 1158 4488 1164
rect 4448 950 4476 1158
rect 4436 944 4488 950
rect 4436 886 4488 892
rect 4068 60 4120 66
rect 3790 -300 3846 54
rect 4068 2 4120 8
rect 4158 54 4292 82
rect 4526 82 4582 160
rect 4632 82 4660 1294
rect 4724 1290 4752 4519
rect 5540 4490 5592 4496
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 4712 1284 4764 1290
rect 4712 1226 4764 1232
rect 4526 54 4660 82
rect 4894 82 4950 160
rect 5000 82 5028 1294
rect 5172 1216 5224 1222
rect 5172 1158 5224 1164
rect 5184 950 5212 1158
rect 5172 944 5224 950
rect 5172 886 5224 892
rect 4894 54 5028 82
rect 5262 82 5318 160
rect 5368 82 5396 1294
rect 5552 1018 5580 4490
rect 12058 4380 12366 4389
rect 12058 4378 12064 4380
rect 12120 4378 12144 4380
rect 12200 4378 12224 4380
rect 12280 4378 12304 4380
rect 12360 4378 12366 4380
rect 12120 4326 12122 4378
rect 12302 4326 12304 4378
rect 12058 4324 12064 4326
rect 12120 4324 12144 4326
rect 12200 4324 12224 4326
rect 12280 4324 12304 4326
rect 12360 4324 12366 4326
rect 12058 4315 12366 4324
rect 11886 4040 11942 4049
rect 11886 3975 11942 3984
rect 6504 3836 6812 3845
rect 6504 3834 6510 3836
rect 6566 3834 6590 3836
rect 6646 3834 6670 3836
rect 6726 3834 6750 3836
rect 6806 3834 6812 3836
rect 6566 3782 6568 3834
rect 6748 3782 6750 3834
rect 6504 3780 6510 3782
rect 6566 3780 6590 3782
rect 6646 3780 6670 3782
rect 6726 3780 6750 3782
rect 6806 3780 6812 3782
rect 6504 3771 6812 3780
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 6504 2748 6812 2757
rect 6504 2746 6510 2748
rect 6566 2746 6590 2748
rect 6646 2746 6670 2748
rect 6726 2746 6750 2748
rect 6806 2746 6812 2748
rect 6566 2694 6568 2746
rect 6748 2694 6750 2746
rect 6504 2692 6510 2694
rect 6566 2692 6590 2694
rect 6646 2692 6670 2694
rect 6726 2692 6750 2694
rect 6806 2692 6812 2694
rect 6504 2683 6812 2692
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 6504 1660 6812 1669
rect 6504 1658 6510 1660
rect 6566 1658 6590 1660
rect 6646 1658 6670 1660
rect 6726 1658 6750 1660
rect 6806 1658 6812 1660
rect 6566 1606 6568 1658
rect 6748 1606 6750 1658
rect 6504 1604 6510 1606
rect 6566 1604 6590 1606
rect 6646 1604 6670 1606
rect 6726 1604 6750 1606
rect 6806 1604 6812 1606
rect 6504 1595 6812 1604
rect 7576 1562 7604 1974
rect 7564 1556 7616 1562
rect 7564 1498 7616 1504
rect 8128 1358 8156 3402
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 8220 1358 8248 2994
rect 11900 2774 11928 3975
rect 12058 3292 12366 3301
rect 12058 3290 12064 3292
rect 12120 3290 12144 3292
rect 12200 3290 12224 3292
rect 12280 3290 12304 3292
rect 12360 3290 12366 3292
rect 12120 3238 12122 3290
rect 12302 3238 12304 3290
rect 12058 3236 12064 3238
rect 12120 3236 12144 3238
rect 12200 3236 12224 3238
rect 12280 3236 12304 3238
rect 12360 3236 12366 3238
rect 12058 3227 12366 3236
rect 13358 3224 13414 3233
rect 13358 3159 13414 3168
rect 13636 3188 13688 3194
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 11808 2746 11928 2774
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 9954 2408 10010 2417
rect 9954 2343 10010 2352
rect 8942 2000 8998 2009
rect 8942 1935 8998 1944
rect 5724 1352 5776 1358
rect 5724 1294 5776 1300
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 6460 1352 6512 1358
rect 6460 1294 6512 1300
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 7564 1352 7616 1358
rect 7564 1294 7616 1300
rect 7932 1352 7984 1358
rect 7932 1294 7984 1300
rect 8116 1352 8168 1358
rect 8116 1294 8168 1300
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 8300 1352 8352 1358
rect 8300 1294 8352 1300
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 5540 1012 5592 1018
rect 5540 954 5592 960
rect 5262 54 5396 82
rect 5630 82 5686 160
rect 5736 82 5764 1294
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 5908 1216 5960 1222
rect 5908 1158 5960 1164
rect 5828 746 5856 1158
rect 5920 882 5948 1158
rect 5908 876 5960 882
rect 5908 818 5960 824
rect 5816 740 5868 746
rect 5816 682 5868 688
rect 6012 160 6040 1294
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6104 814 6132 1158
rect 6092 808 6144 814
rect 6092 750 6144 756
rect 5630 54 5764 82
rect 4158 -300 4214 54
rect 4526 -300 4582 54
rect 4894 -300 4950 54
rect 5262 -300 5318 54
rect 5630 -300 5686 54
rect 5998 -300 6054 160
rect 6366 82 6422 160
rect 6472 82 6500 1294
rect 6644 1216 6696 1222
rect 6644 1158 6696 1164
rect 6656 1018 6684 1158
rect 6644 1012 6696 1018
rect 6644 954 6696 960
rect 6366 54 6500 82
rect 6734 82 6790 160
rect 6840 82 6868 1294
rect 7012 1216 7064 1222
rect 7012 1158 7064 1164
rect 7024 474 7052 1158
rect 7012 468 7064 474
rect 7012 410 7064 416
rect 6734 54 6868 82
rect 7102 82 7158 160
rect 7208 82 7236 1294
rect 7102 54 7236 82
rect 7470 82 7526 160
rect 7576 82 7604 1294
rect 7656 1216 7708 1222
rect 7656 1158 7708 1164
rect 7748 1216 7800 1222
rect 7748 1158 7800 1164
rect 7668 406 7696 1158
rect 7760 542 7788 1158
rect 7748 536 7800 542
rect 7748 478 7800 484
rect 7656 400 7708 406
rect 7656 342 7708 348
rect 7470 54 7604 82
rect 7838 82 7894 160
rect 7944 82 7972 1294
rect 7838 54 7972 82
rect 8206 82 8262 160
rect 8312 82 8340 1294
rect 8588 160 8616 1294
rect 8760 1216 8812 1222
rect 8760 1158 8812 1164
rect 8772 921 8800 1158
rect 8758 912 8814 921
rect 8758 847 8814 856
rect 8956 814 8984 1935
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 9404 1352 9456 1358
rect 9404 1294 9456 1300
rect 9772 1352 9824 1358
rect 9968 1340 9996 2343
rect 9772 1294 9824 1300
rect 9876 1312 9996 1340
rect 10140 1352 10192 1358
rect 8944 808 8996 814
rect 8944 750 8996 756
rect 8206 54 8340 82
rect 6366 -300 6422 54
rect 6734 -300 6790 54
rect 7102 -300 7158 54
rect 7470 -300 7526 54
rect 7838 -300 7894 54
rect 8206 -300 8262 54
rect 8574 -300 8630 160
rect 8942 82 8998 160
rect 9048 82 9076 1294
rect 9220 1216 9272 1222
rect 9220 1158 9272 1164
rect 9232 649 9260 1158
rect 9218 640 9274 649
rect 9218 575 9274 584
rect 8942 54 9076 82
rect 9310 82 9366 160
rect 9416 82 9444 1294
rect 9588 1216 9640 1222
rect 9588 1158 9640 1164
rect 9600 513 9628 1158
rect 9586 504 9642 513
rect 9586 439 9642 448
rect 9310 54 9444 82
rect 9678 82 9734 160
rect 9784 82 9812 1294
rect 9876 882 9904 1312
rect 10140 1294 10192 1300
rect 10508 1352 10560 1358
rect 10508 1294 10560 1300
rect 10876 1352 10928 1358
rect 10876 1294 10928 1300
rect 9956 1216 10008 1222
rect 9956 1158 10008 1164
rect 9968 882 9996 1158
rect 9864 876 9916 882
rect 9864 818 9916 824
rect 9956 876 10008 882
rect 9956 818 10008 824
rect 9678 54 9812 82
rect 10046 82 10102 160
rect 10152 82 10180 1294
rect 10416 1284 10468 1290
rect 10416 1226 10468 1232
rect 10324 1216 10376 1222
rect 10324 1158 10376 1164
rect 10336 377 10364 1158
rect 10428 882 10456 1226
rect 10416 876 10468 882
rect 10416 818 10468 824
rect 10322 368 10378 377
rect 10322 303 10378 312
rect 10046 54 10180 82
rect 10414 82 10470 160
rect 10520 82 10548 1294
rect 10692 1216 10744 1222
rect 10692 1158 10744 1164
rect 10704 785 10732 1158
rect 10690 776 10746 785
rect 10690 711 10746 720
rect 10414 54 10548 82
rect 10782 82 10838 160
rect 10888 82 10916 1294
rect 10980 1018 11008 2450
rect 11244 2372 11296 2378
rect 11244 2314 11296 2320
rect 11152 1352 11204 1358
rect 11152 1294 11204 1300
rect 11060 1216 11112 1222
rect 11060 1158 11112 1164
rect 10968 1012 11020 1018
rect 10968 954 11020 960
rect 11072 610 11100 1158
rect 11060 604 11112 610
rect 11060 546 11112 552
rect 11164 160 11192 1294
rect 11256 542 11284 2314
rect 11612 1352 11664 1358
rect 11612 1294 11664 1300
rect 11702 1320 11758 1329
rect 11336 1216 11388 1222
rect 11336 1158 11388 1164
rect 11348 1018 11376 1158
rect 11336 1012 11388 1018
rect 11336 954 11388 960
rect 11244 536 11296 542
rect 11244 478 11296 484
rect 10782 54 10916 82
rect 8942 -300 8998 54
rect 9310 -300 9366 54
rect 9678 -300 9734 54
rect 10046 -300 10102 54
rect 10414 -300 10470 54
rect 10782 -300 10838 54
rect 11150 -300 11206 160
rect 11518 82 11574 160
rect 11624 82 11652 1294
rect 11702 1255 11758 1264
rect 11716 134 11744 1255
rect 11808 134 11836 2746
rect 12058 2204 12366 2213
rect 12058 2202 12064 2204
rect 12120 2202 12144 2204
rect 12200 2202 12224 2204
rect 12280 2202 12304 2204
rect 12360 2202 12366 2204
rect 12120 2150 12122 2202
rect 12302 2150 12304 2202
rect 12058 2148 12064 2150
rect 12120 2148 12144 2150
rect 12200 2148 12224 2150
rect 12280 2148 12304 2150
rect 12360 2148 12366 2150
rect 12058 2139 12366 2148
rect 12544 1358 12572 3062
rect 12992 2984 13044 2990
rect 12992 2926 13044 2932
rect 11980 1352 12032 1358
rect 11980 1294 12032 1300
rect 12164 1352 12216 1358
rect 12532 1352 12584 1358
rect 12216 1312 12296 1340
rect 12164 1294 12216 1300
rect 11518 54 11652 82
rect 11704 128 11756 134
rect 11704 70 11756 76
rect 11796 128 11848 134
rect 11796 70 11848 76
rect 11886 82 11942 160
rect 11992 82 12020 1294
rect 12268 1204 12296 1312
rect 12532 1294 12584 1300
rect 12624 1352 12676 1358
rect 12624 1294 12676 1300
rect 12900 1352 12952 1358
rect 12900 1294 12952 1300
rect 12532 1216 12584 1222
rect 12268 1176 12434 1204
rect 12058 1116 12366 1125
rect 12058 1114 12064 1116
rect 12120 1114 12144 1116
rect 12200 1114 12224 1116
rect 12280 1114 12304 1116
rect 12360 1114 12366 1116
rect 12120 1062 12122 1114
rect 12302 1062 12304 1114
rect 12058 1060 12064 1062
rect 12120 1060 12144 1062
rect 12200 1060 12224 1062
rect 12280 1060 12304 1062
rect 12360 1060 12366 1062
rect 12058 1051 12366 1060
rect 12406 932 12434 1176
rect 12532 1158 12584 1164
rect 12360 904 12434 932
rect 12072 468 12124 474
rect 12072 410 12124 416
rect 12084 134 12112 410
rect 11886 54 12020 82
rect 12072 128 12124 134
rect 12072 70 12124 76
rect 12254 82 12310 160
rect 12360 82 12388 904
rect 12544 338 12572 1158
rect 12532 332 12584 338
rect 12532 274 12584 280
rect 12636 160 12664 1294
rect 12808 1216 12860 1222
rect 12806 1184 12808 1193
rect 12860 1184 12862 1193
rect 12806 1119 12862 1128
rect 12714 1048 12770 1057
rect 12714 983 12770 992
rect 12728 270 12756 983
rect 12716 264 12768 270
rect 12716 206 12768 212
rect 12254 54 12388 82
rect 11518 -300 11574 54
rect 11886 -300 11942 54
rect 12254 -300 12310 54
rect 12622 -300 12678 160
rect 12912 82 12940 1294
rect 13004 814 13032 2926
rect 13176 1352 13228 1358
rect 13176 1294 13228 1300
rect 13084 1216 13136 1222
rect 13084 1158 13136 1164
rect 13096 950 13124 1158
rect 13084 944 13136 950
rect 13084 886 13136 892
rect 12992 808 13044 814
rect 12992 750 13044 756
rect 13084 808 13136 814
rect 13084 750 13136 756
rect 12990 82 13046 160
rect 12912 54 13046 82
rect 13096 66 13124 750
rect 13188 82 13216 1294
rect 13268 1216 13320 1222
rect 13268 1158 13320 1164
rect 13280 270 13308 1158
rect 13372 814 13400 3159
rect 13636 3130 13688 3136
rect 13452 1352 13504 1358
rect 13452 1294 13504 1300
rect 13360 808 13412 814
rect 13360 750 13412 756
rect 13268 264 13320 270
rect 13268 206 13320 212
rect 13358 82 13414 160
rect 12990 -300 13046 54
rect 13084 60 13136 66
rect 13188 54 13414 82
rect 13464 82 13492 1294
rect 13648 406 13676 3130
rect 13832 2106 13860 8434
rect 16948 4208 17000 4214
rect 16948 4150 17000 4156
rect 16212 3664 16264 3670
rect 15934 3632 15990 3641
rect 16212 3606 16264 3612
rect 15934 3567 15990 3576
rect 14096 2916 14148 2922
rect 14096 2858 14148 2864
rect 13820 2100 13872 2106
rect 13820 2042 13872 2048
rect 13728 1352 13780 1358
rect 14004 1352 14056 1358
rect 13780 1312 13860 1340
rect 13728 1294 13780 1300
rect 13636 400 13688 406
rect 13636 342 13688 348
rect 13648 190 13768 218
rect 13648 82 13676 190
rect 13740 160 13768 190
rect 13464 54 13676 82
rect 13084 2 13136 8
rect 13358 -300 13414 54
rect 13726 -300 13782 160
rect 13832 82 13860 1312
rect 14004 1294 14056 1300
rect 13912 1216 13964 1222
rect 13912 1158 13964 1164
rect 13924 406 13952 1158
rect 14016 474 14044 1294
rect 14108 1222 14136 2858
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15016 1964 15068 1970
rect 15016 1906 15068 1912
rect 14832 1896 14884 1902
rect 14832 1838 14884 1844
rect 14844 1465 14872 1838
rect 15028 1562 15056 1906
rect 15108 1896 15160 1902
rect 15108 1838 15160 1844
rect 15198 1864 15254 1873
rect 15120 1562 15148 1838
rect 15198 1799 15254 1808
rect 15212 1766 15240 1799
rect 15200 1760 15252 1766
rect 15200 1702 15252 1708
rect 15304 1562 15332 2246
rect 15660 1964 15712 1970
rect 15712 1924 15792 1952
rect 15660 1906 15712 1912
rect 15016 1556 15068 1562
rect 15016 1498 15068 1504
rect 15108 1556 15160 1562
rect 15108 1498 15160 1504
rect 15292 1556 15344 1562
rect 15292 1498 15344 1504
rect 14830 1456 14886 1465
rect 14830 1391 14886 1400
rect 14556 1352 14608 1358
rect 14556 1294 14608 1300
rect 15108 1352 15160 1358
rect 15384 1352 15436 1358
rect 15160 1312 15332 1340
rect 15108 1294 15160 1300
rect 14464 1284 14516 1290
rect 14464 1226 14516 1232
rect 14096 1216 14148 1222
rect 14096 1158 14148 1164
rect 14004 468 14056 474
rect 14004 410 14056 416
rect 13912 400 13964 406
rect 13912 342 13964 348
rect 14016 190 14136 218
rect 14016 82 14044 190
rect 14108 160 14136 190
rect 14476 160 14504 1226
rect 13832 54 14044 82
rect 14094 -300 14150 160
rect 14462 -300 14518 160
rect 14568 82 14596 1294
rect 15016 1284 15068 1290
rect 15016 1226 15068 1232
rect 15028 762 15056 1226
rect 15028 734 15240 762
rect 15212 160 15240 734
rect 14830 82 14886 160
rect 14568 54 14886 82
rect 14830 -300 14886 54
rect 15198 -300 15254 160
rect 15304 82 15332 1312
rect 15436 1312 15700 1340
rect 15384 1294 15436 1300
rect 15566 82 15622 160
rect 15304 54 15622 82
rect 15672 82 15700 1312
rect 15764 610 15792 1924
rect 15948 1358 15976 3567
rect 16224 2106 16252 3606
rect 16856 2848 16908 2854
rect 16856 2790 16908 2796
rect 16486 2272 16542 2281
rect 16486 2207 16542 2216
rect 16500 2106 16528 2207
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16488 2100 16540 2106
rect 16488 2042 16540 2048
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16488 1964 16540 1970
rect 16488 1906 16540 1912
rect 16040 1562 16068 1906
rect 16316 1562 16344 1906
rect 16500 1562 16528 1906
rect 16868 1834 16896 2790
rect 16856 1828 16908 1834
rect 16856 1770 16908 1776
rect 16028 1556 16080 1562
rect 16028 1498 16080 1504
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 16488 1556 16540 1562
rect 16488 1498 16540 1504
rect 16960 1442 16988 4150
rect 17052 2650 17080 8434
rect 19260 8362 19288 8434
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 17612 8188 17920 8197
rect 17612 8186 17618 8188
rect 17674 8186 17698 8188
rect 17754 8186 17778 8188
rect 17834 8186 17858 8188
rect 17914 8186 17920 8188
rect 17674 8134 17676 8186
rect 17856 8134 17858 8186
rect 17612 8132 17618 8134
rect 17674 8132 17698 8134
rect 17754 8132 17778 8134
rect 17834 8132 17858 8134
rect 17914 8132 17920 8134
rect 17612 8123 17920 8132
rect 17612 7100 17920 7109
rect 17612 7098 17618 7100
rect 17674 7098 17698 7100
rect 17754 7098 17778 7100
rect 17834 7098 17858 7100
rect 17914 7098 17920 7100
rect 17674 7046 17676 7098
rect 17856 7046 17858 7098
rect 17612 7044 17618 7046
rect 17674 7044 17698 7046
rect 17754 7044 17778 7046
rect 17834 7044 17858 7046
rect 17914 7044 17920 7046
rect 17612 7035 17920 7044
rect 17612 6012 17920 6021
rect 17612 6010 17618 6012
rect 17674 6010 17698 6012
rect 17754 6010 17778 6012
rect 17834 6010 17858 6012
rect 17914 6010 17920 6012
rect 17674 5958 17676 6010
rect 17856 5958 17858 6010
rect 17612 5956 17618 5958
rect 17674 5956 17698 5958
rect 17754 5956 17778 5958
rect 17834 5956 17858 5958
rect 17914 5956 17920 5958
rect 17612 5947 17920 5956
rect 19352 5658 19380 8434
rect 19352 5630 19564 5658
rect 17612 4924 17920 4933
rect 17612 4922 17618 4924
rect 17674 4922 17698 4924
rect 17754 4922 17778 4924
rect 17834 4922 17858 4924
rect 17914 4922 17920 4924
rect 17674 4870 17676 4922
rect 17856 4870 17858 4922
rect 17612 4868 17618 4870
rect 17674 4868 17698 4870
rect 17754 4868 17778 4870
rect 17834 4868 17858 4870
rect 17914 4868 17920 4870
rect 17612 4859 17920 4868
rect 18512 4276 18564 4282
rect 18512 4218 18564 4224
rect 17612 3836 17920 3845
rect 17612 3834 17618 3836
rect 17674 3834 17698 3836
rect 17754 3834 17778 3836
rect 17834 3834 17858 3836
rect 17914 3834 17920 3836
rect 17674 3782 17676 3834
rect 17856 3782 17858 3834
rect 17612 3780 17618 3782
rect 17674 3780 17698 3782
rect 17754 3780 17778 3782
rect 17834 3780 17858 3782
rect 17914 3780 17920 3782
rect 17612 3771 17920 3780
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17130 3088 17186 3097
rect 17130 3023 17186 3032
rect 17040 2644 17092 2650
rect 17040 2586 17092 2592
rect 17144 2106 17172 3023
rect 17314 2952 17370 2961
rect 17314 2887 17370 2896
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17132 2100 17184 2106
rect 17132 2042 17184 2048
rect 17132 1964 17184 1970
rect 17132 1906 17184 1912
rect 17144 1562 17172 1906
rect 17236 1562 17264 2382
rect 17132 1556 17184 1562
rect 17132 1498 17184 1504
rect 17224 1556 17276 1562
rect 17224 1498 17276 1504
rect 16960 1426 17172 1442
rect 16960 1420 17184 1426
rect 16960 1414 17132 1420
rect 17132 1362 17184 1368
rect 17328 1358 17356 2887
rect 17512 2106 17540 3334
rect 17612 2748 17920 2757
rect 17612 2746 17618 2748
rect 17674 2746 17698 2748
rect 17754 2746 17778 2748
rect 17834 2746 17858 2748
rect 17914 2746 17920 2748
rect 17674 2694 17676 2746
rect 17856 2694 17858 2746
rect 17612 2692 17618 2694
rect 17674 2692 17698 2694
rect 17754 2692 17778 2694
rect 17834 2692 17858 2694
rect 17914 2692 17920 2694
rect 17612 2683 17920 2692
rect 18050 2680 18106 2689
rect 17880 2624 18050 2632
rect 17880 2615 18106 2624
rect 17880 2604 18092 2615
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 17880 2038 17908 2604
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 18052 2372 18104 2378
rect 18052 2314 18104 2320
rect 18064 2038 18092 2314
rect 18156 2106 18184 2518
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 18144 2100 18196 2106
rect 18144 2042 18196 2048
rect 17868 2032 17920 2038
rect 17868 1974 17920 1980
rect 18052 2032 18104 2038
rect 18052 1974 18104 1980
rect 17408 1964 17460 1970
rect 17408 1906 17460 1912
rect 17500 1964 17552 1970
rect 17500 1906 17552 1912
rect 18144 1964 18196 1970
rect 18144 1906 18196 1912
rect 17420 1562 17448 1906
rect 17512 1562 17540 1906
rect 18052 1760 18104 1766
rect 18052 1702 18104 1708
rect 17612 1660 17920 1669
rect 17612 1658 17618 1660
rect 17674 1658 17698 1660
rect 17754 1658 17778 1660
rect 17834 1658 17858 1660
rect 17914 1658 17920 1660
rect 17674 1606 17676 1658
rect 17856 1606 17858 1658
rect 17612 1604 17618 1606
rect 17674 1604 17698 1606
rect 17754 1604 17778 1606
rect 17834 1604 17858 1606
rect 17914 1604 17920 1606
rect 17612 1595 17920 1604
rect 17408 1556 17460 1562
rect 17408 1498 17460 1504
rect 17500 1556 17552 1562
rect 17500 1498 17552 1504
rect 15844 1352 15896 1358
rect 15844 1294 15896 1300
rect 15936 1352 15988 1358
rect 15936 1294 15988 1300
rect 16028 1352 16080 1358
rect 16488 1352 16540 1358
rect 16080 1312 16436 1340
rect 16028 1294 16080 1300
rect 15752 604 15804 610
rect 15752 546 15804 552
rect 15856 218 15884 1294
rect 15856 190 16068 218
rect 15934 82 15990 160
rect 15672 54 15990 82
rect 16040 82 16068 190
rect 16224 190 16344 218
rect 16224 82 16252 190
rect 16316 160 16344 190
rect 16040 54 16252 82
rect 15566 -300 15622 54
rect 15934 -300 15990 54
rect 16302 -300 16358 160
rect 16408 82 16436 1312
rect 16764 1352 16816 1358
rect 16540 1312 16620 1340
rect 16488 1294 16540 1300
rect 16592 218 16620 1312
rect 16764 1294 16816 1300
rect 17316 1352 17368 1358
rect 17316 1294 17368 1300
rect 17500 1352 17552 1358
rect 17500 1294 17552 1300
rect 16776 814 16804 1294
rect 16764 808 16816 814
rect 16764 750 16816 756
rect 17408 808 17460 814
rect 17408 750 17460 756
rect 17316 740 17368 746
rect 17316 682 17368 688
rect 17328 626 17356 682
rect 17052 610 17356 626
rect 17040 604 17356 610
rect 17092 598 17356 604
rect 17040 546 17092 552
rect 16592 190 16804 218
rect 16670 82 16726 160
rect 16408 54 16726 82
rect 16776 82 16804 190
rect 16960 190 17080 218
rect 16960 82 16988 190
rect 17052 160 17080 190
rect 17420 160 17448 750
rect 16776 54 16988 82
rect 16670 -300 16726 54
rect 17038 -300 17094 160
rect 17406 -300 17462 160
rect 17512 82 17540 1294
rect 18064 1193 18092 1702
rect 18156 1562 18184 1906
rect 18144 1556 18196 1562
rect 18144 1498 18196 1504
rect 18236 1352 18288 1358
rect 18236 1294 18288 1300
rect 17866 1184 17922 1193
rect 17866 1119 17922 1128
rect 18050 1184 18106 1193
rect 18050 1119 18106 1128
rect 17684 944 17736 950
rect 17684 886 17736 892
rect 17696 474 17724 886
rect 17880 882 17908 1119
rect 17868 876 17920 882
rect 17868 818 17920 824
rect 17684 468 17736 474
rect 17684 410 17736 416
rect 17696 190 17816 218
rect 17696 82 17724 190
rect 17788 160 17816 190
rect 17512 54 17724 82
rect 17774 -300 17830 160
rect 18142 82 18198 160
rect 18248 82 18276 1294
rect 18340 202 18368 2314
rect 18524 1970 18552 4218
rect 18694 3496 18750 3505
rect 18694 3431 18750 3440
rect 18708 1970 18736 3431
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 18786 2544 18842 2553
rect 18786 2479 18842 2488
rect 18800 2446 18828 2479
rect 18788 2440 18840 2446
rect 18788 2382 18840 2388
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18892 1970 18920 2246
rect 18420 1964 18472 1970
rect 18420 1906 18472 1912
rect 18512 1964 18564 1970
rect 18512 1906 18564 1912
rect 18696 1964 18748 1970
rect 18696 1906 18748 1912
rect 18788 1964 18840 1970
rect 18788 1906 18840 1912
rect 18880 1964 18932 1970
rect 18880 1906 18932 1912
rect 18432 1562 18460 1906
rect 18696 1760 18748 1766
rect 18696 1702 18748 1708
rect 18708 1562 18736 1702
rect 18800 1562 18828 1906
rect 18420 1556 18472 1562
rect 18420 1498 18472 1504
rect 18696 1556 18748 1562
rect 18696 1498 18748 1504
rect 18788 1556 18840 1562
rect 18788 1498 18840 1504
rect 18984 1358 19012 2246
rect 19168 2106 19196 2382
rect 19260 2360 19288 3130
rect 19432 2848 19484 2854
rect 19432 2790 19484 2796
rect 19444 2530 19472 2790
rect 19536 2650 19564 5630
rect 20534 3904 20590 3913
rect 20534 3839 20590 3848
rect 20444 3460 20496 3466
rect 20444 3402 20496 3408
rect 19890 2680 19946 2689
rect 19524 2644 19576 2650
rect 19890 2615 19946 2624
rect 19524 2586 19576 2592
rect 19444 2502 19656 2530
rect 19628 2446 19656 2502
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 19260 2332 19564 2360
rect 19156 2100 19208 2106
rect 19156 2042 19208 2048
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 19260 2009 19288 2042
rect 19246 2000 19302 2009
rect 19536 1970 19564 2332
rect 19720 1970 19748 2382
rect 19812 2106 19840 2450
rect 19904 2446 19932 2615
rect 19892 2440 19944 2446
rect 19892 2382 19944 2388
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 19800 2100 19852 2106
rect 19800 2042 19852 2048
rect 19246 1935 19302 1944
rect 19524 1964 19576 1970
rect 19524 1906 19576 1912
rect 19708 1964 19760 1970
rect 19708 1906 19760 1912
rect 19708 1760 19760 1766
rect 19706 1728 19708 1737
rect 19800 1760 19852 1766
rect 19760 1728 19762 1737
rect 19800 1702 19852 1708
rect 19706 1663 19762 1672
rect 19812 1358 19840 1702
rect 19996 1358 20024 2246
rect 18512 1352 18564 1358
rect 18512 1294 18564 1300
rect 18788 1352 18840 1358
rect 18880 1352 18932 1358
rect 18788 1294 18840 1300
rect 18878 1320 18880 1329
rect 18972 1352 19024 1358
rect 18932 1320 18934 1329
rect 18328 196 18380 202
rect 18524 160 18552 1294
rect 18328 138 18380 144
rect 18142 54 18276 82
rect 18142 -300 18198 54
rect 18510 -300 18566 160
rect 18800 82 18828 1294
rect 18972 1294 19024 1300
rect 19064 1352 19116 1358
rect 19800 1352 19852 1358
rect 19116 1312 19288 1340
rect 19064 1294 19116 1300
rect 18878 1255 18934 1264
rect 19260 160 19288 1312
rect 19800 1294 19852 1300
rect 19984 1352 20036 1358
rect 19984 1294 20036 1300
rect 20180 1290 20208 2246
rect 20456 1970 20484 3402
rect 20548 2394 20576 3839
rect 20640 2650 20668 8502
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21468 2650 21496 8434
rect 22098 3224 22154 3233
rect 22098 3159 22154 3168
rect 22006 2680 22062 2689
rect 20628 2644 20680 2650
rect 20628 2586 20680 2592
rect 21456 2644 21508 2650
rect 22006 2615 22008 2624
rect 21456 2586 21508 2592
rect 22060 2615 22062 2624
rect 22008 2586 22060 2592
rect 21546 2544 21602 2553
rect 21546 2479 21602 2488
rect 21364 2440 21416 2446
rect 20718 2408 20774 2417
rect 20548 2366 20668 2394
rect 20640 2281 20668 2366
rect 20718 2343 20774 2352
rect 21100 2400 21364 2428
rect 20626 2272 20682 2281
rect 20626 2207 20682 2216
rect 20732 1970 20760 2343
rect 20996 2304 21048 2310
rect 20996 2246 21048 2252
rect 21008 2106 21036 2246
rect 20812 2100 20864 2106
rect 20812 2042 20864 2048
rect 20904 2100 20956 2106
rect 20904 2042 20956 2048
rect 20996 2100 21048 2106
rect 20996 2042 21048 2048
rect 20260 1964 20312 1970
rect 20260 1906 20312 1912
rect 20444 1964 20496 1970
rect 20444 1906 20496 1912
rect 20720 1964 20772 1970
rect 20720 1906 20772 1912
rect 20168 1284 20220 1290
rect 20168 1226 20220 1232
rect 19708 1216 19760 1222
rect 19628 1176 19708 1204
rect 19628 160 19656 1176
rect 19708 1158 19760 1164
rect 20076 1216 20128 1222
rect 20076 1158 20128 1164
rect 18878 82 18934 160
rect 18800 54 18934 82
rect 18878 -300 18934 54
rect 19246 -300 19302 160
rect 19614 -300 19670 160
rect 19982 82 20038 160
rect 20088 82 20116 1158
rect 20272 474 20300 1906
rect 20352 1760 20404 1766
rect 20352 1702 20404 1708
rect 20364 1465 20392 1702
rect 20350 1456 20406 1465
rect 20350 1391 20406 1400
rect 20824 1306 20852 2042
rect 20916 1494 20944 2042
rect 21100 1850 21128 2400
rect 21364 2382 21416 2388
rect 21454 2136 21510 2145
rect 21454 2071 21510 2080
rect 21008 1834 21128 1850
rect 20996 1828 21128 1834
rect 21048 1822 21128 1828
rect 20996 1770 21048 1776
rect 21180 1760 21232 1766
rect 21180 1702 21232 1708
rect 20904 1488 20956 1494
rect 20904 1430 20956 1436
rect 20824 1290 20944 1306
rect 20824 1284 20956 1290
rect 20824 1278 20904 1284
rect 20904 1226 20956 1232
rect 20444 1216 20496 1222
rect 20364 1176 20444 1204
rect 20260 468 20312 474
rect 20260 410 20312 416
rect 20364 160 20392 1176
rect 20812 1216 20864 1222
rect 20444 1158 20496 1164
rect 20732 1176 20812 1204
rect 20732 160 20760 1176
rect 20812 1158 20864 1164
rect 19982 54 20116 82
rect 19982 -300 20038 54
rect 20350 -300 20406 160
rect 20718 -300 20774 160
rect 21086 82 21142 160
rect 21192 82 21220 1702
rect 21468 1358 21496 2071
rect 21560 1970 21588 2479
rect 22112 2446 22140 3159
rect 22284 2848 22336 2854
rect 22284 2790 22336 2796
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 22100 2440 22152 2446
rect 22204 2417 22232 2450
rect 22100 2382 22152 2388
rect 22190 2408 22246 2417
rect 21548 1964 21600 1970
rect 21548 1906 21600 1912
rect 21836 1850 21864 2382
rect 22296 2394 22324 2790
rect 22388 2650 22416 8910
rect 22928 8900 22980 8906
rect 22928 8842 22980 8848
rect 22558 4040 22614 4049
rect 22558 3975 22614 3984
rect 22376 2644 22428 2650
rect 22376 2586 22428 2592
rect 22296 2366 22508 2394
rect 22190 2343 22246 2352
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22284 2304 22336 2310
rect 22284 2246 22336 2252
rect 22204 2038 22232 2246
rect 22192 2032 22244 2038
rect 22192 1974 22244 1980
rect 21744 1822 21864 1850
rect 21456 1352 21508 1358
rect 21456 1294 21508 1300
rect 21548 1216 21600 1222
rect 21468 1176 21548 1204
rect 21468 160 21496 1176
rect 21548 1158 21600 1164
rect 21744 1057 21772 1822
rect 22100 1760 22152 1766
rect 21836 1720 22100 1748
rect 21730 1048 21786 1057
rect 21730 983 21786 992
rect 21836 160 21864 1720
rect 22100 1702 22152 1708
rect 22296 1494 22324 2246
rect 22480 1970 22508 2366
rect 22572 1970 22600 3975
rect 22744 3528 22796 3534
rect 22744 3470 22796 3476
rect 22650 2816 22706 2825
rect 22650 2751 22706 2760
rect 22664 2446 22692 2751
rect 22756 2650 22784 3470
rect 22744 2644 22796 2650
rect 22940 2632 22968 8842
rect 23032 8566 23060 9846
rect 23216 9738 23244 9846
rect 23294 9840 23350 10300
rect 25502 9840 25558 10300
rect 27710 9840 27766 10300
rect 29918 9840 29974 10300
rect 32126 9840 32182 10300
rect 34334 9840 34390 10300
rect 36542 9840 36598 10300
rect 38750 9840 38806 10300
rect 40958 9840 41014 10300
rect 43166 9840 43222 10300
rect 45374 9840 45430 10300
rect 23308 9738 23336 9840
rect 23216 9710 23336 9738
rect 23664 8832 23716 8838
rect 23664 8774 23716 8780
rect 23166 8732 23474 8741
rect 23166 8730 23172 8732
rect 23228 8730 23252 8732
rect 23308 8730 23332 8732
rect 23388 8730 23412 8732
rect 23468 8730 23474 8732
rect 23228 8678 23230 8730
rect 23410 8678 23412 8730
rect 23166 8676 23172 8678
rect 23228 8676 23252 8678
rect 23308 8676 23332 8678
rect 23388 8676 23412 8678
rect 23468 8676 23474 8678
rect 23166 8667 23474 8676
rect 23020 8560 23072 8566
rect 23020 8502 23072 8508
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 23032 3534 23060 8366
rect 23166 7644 23474 7653
rect 23166 7642 23172 7644
rect 23228 7642 23252 7644
rect 23308 7642 23332 7644
rect 23388 7642 23412 7644
rect 23468 7642 23474 7644
rect 23228 7590 23230 7642
rect 23410 7590 23412 7642
rect 23166 7588 23172 7590
rect 23228 7588 23252 7590
rect 23308 7588 23332 7590
rect 23388 7588 23412 7590
rect 23468 7588 23474 7590
rect 23166 7579 23474 7588
rect 23166 6556 23474 6565
rect 23166 6554 23172 6556
rect 23228 6554 23252 6556
rect 23308 6554 23332 6556
rect 23388 6554 23412 6556
rect 23468 6554 23474 6556
rect 23228 6502 23230 6554
rect 23410 6502 23412 6554
rect 23166 6500 23172 6502
rect 23228 6500 23252 6502
rect 23308 6500 23332 6502
rect 23388 6500 23412 6502
rect 23468 6500 23474 6502
rect 23166 6491 23474 6500
rect 23166 5468 23474 5477
rect 23166 5466 23172 5468
rect 23228 5466 23252 5468
rect 23308 5466 23332 5468
rect 23388 5466 23412 5468
rect 23468 5466 23474 5468
rect 23228 5414 23230 5466
rect 23410 5414 23412 5466
rect 23166 5412 23172 5414
rect 23228 5412 23252 5414
rect 23308 5412 23332 5414
rect 23388 5412 23412 5414
rect 23468 5412 23474 5414
rect 23166 5403 23474 5412
rect 23166 4380 23474 4389
rect 23166 4378 23172 4380
rect 23228 4378 23252 4380
rect 23308 4378 23332 4380
rect 23388 4378 23412 4380
rect 23468 4378 23474 4380
rect 23228 4326 23230 4378
rect 23410 4326 23412 4378
rect 23166 4324 23172 4326
rect 23228 4324 23252 4326
rect 23308 4324 23332 4326
rect 23388 4324 23412 4326
rect 23468 4324 23474 4326
rect 23166 4315 23474 4324
rect 23020 3528 23072 3534
rect 23020 3470 23072 3476
rect 23166 3292 23474 3301
rect 23166 3290 23172 3292
rect 23228 3290 23252 3292
rect 23308 3290 23332 3292
rect 23388 3290 23412 3292
rect 23468 3290 23474 3292
rect 23228 3238 23230 3290
rect 23410 3238 23412 3290
rect 23166 3236 23172 3238
rect 23228 3236 23252 3238
rect 23308 3236 23332 3238
rect 23388 3236 23412 3238
rect 23468 3236 23474 3238
rect 23166 3227 23474 3236
rect 23480 2916 23532 2922
rect 23480 2858 23532 2864
rect 23204 2848 23256 2854
rect 23204 2790 23256 2796
rect 23020 2644 23072 2650
rect 22940 2604 23020 2632
rect 22744 2586 22796 2592
rect 23020 2586 23072 2592
rect 23112 2576 23164 2582
rect 22756 2524 23112 2530
rect 22756 2518 23164 2524
rect 22756 2514 23152 2518
rect 22744 2508 23152 2514
rect 22796 2502 23152 2508
rect 22744 2450 22796 2456
rect 22652 2440 22704 2446
rect 23112 2440 23164 2446
rect 22652 2382 22704 2388
rect 23032 2400 23112 2428
rect 22468 1964 22520 1970
rect 22468 1906 22520 1912
rect 22560 1964 22612 1970
rect 22560 1906 22612 1912
rect 23032 1834 23060 2400
rect 23112 2382 23164 2388
rect 23216 2310 23244 2790
rect 23492 2394 23520 2858
rect 23584 2582 23612 8434
rect 23676 2774 23704 8774
rect 25516 8634 25544 9840
rect 27724 8634 27752 9840
rect 29932 8634 29960 9840
rect 32140 8634 32168 9840
rect 34348 9058 34376 9840
rect 34164 9030 34376 9058
rect 34164 8634 34192 9030
rect 34274 8732 34582 8741
rect 34274 8730 34280 8732
rect 34336 8730 34360 8732
rect 34416 8730 34440 8732
rect 34496 8730 34520 8732
rect 34576 8730 34582 8732
rect 34336 8678 34338 8730
rect 34518 8678 34520 8730
rect 34274 8676 34280 8678
rect 34336 8676 34360 8678
rect 34416 8676 34440 8678
rect 34496 8676 34520 8678
rect 34576 8676 34582 8678
rect 34274 8667 34582 8676
rect 36556 8634 36584 9840
rect 38764 8634 38792 9840
rect 40972 8634 41000 9840
rect 43180 8634 43208 9840
rect 45388 8922 45416 9840
rect 45296 8894 45416 8922
rect 45296 8634 45324 8894
rect 45382 8732 45690 8741
rect 45382 8730 45388 8732
rect 45444 8730 45468 8732
rect 45524 8730 45548 8732
rect 45604 8730 45628 8732
rect 45684 8730 45690 8732
rect 45444 8678 45446 8730
rect 45626 8678 45628 8730
rect 45382 8676 45388 8678
rect 45444 8676 45468 8678
rect 45524 8676 45548 8678
rect 45604 8676 45628 8678
rect 45684 8676 45690 8678
rect 45382 8667 45690 8676
rect 25504 8628 25556 8634
rect 25504 8570 25556 8576
rect 27712 8628 27764 8634
rect 27712 8570 27764 8576
rect 29920 8628 29972 8634
rect 29920 8570 29972 8576
rect 32128 8628 32180 8634
rect 32128 8570 32180 8576
rect 34152 8628 34204 8634
rect 34152 8570 34204 8576
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 38752 8628 38804 8634
rect 38752 8570 38804 8576
rect 40960 8628 41012 8634
rect 40960 8570 41012 8576
rect 43168 8628 43220 8634
rect 43168 8570 43220 8576
rect 45284 8628 45336 8634
rect 45284 8570 45336 8576
rect 25872 8492 25924 8498
rect 25872 8434 25924 8440
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 30380 8492 30432 8498
rect 30380 8434 30432 8440
rect 32496 8492 32548 8498
rect 32496 8434 32548 8440
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 36912 8492 36964 8498
rect 36912 8434 36964 8440
rect 39028 8492 39080 8498
rect 39028 8434 39080 8440
rect 41328 8492 41380 8498
rect 41328 8434 41380 8440
rect 43536 8492 43588 8498
rect 43536 8434 43588 8440
rect 44548 8492 44600 8498
rect 44548 8434 44600 8440
rect 24400 8356 24452 8362
rect 24400 8298 24452 8304
rect 24308 4548 24360 4554
rect 24308 4490 24360 4496
rect 23676 2746 23888 2774
rect 23572 2576 23624 2582
rect 23572 2518 23624 2524
rect 23860 2446 23888 2746
rect 24214 2680 24270 2689
rect 24214 2615 24270 2624
rect 23848 2440 23900 2446
rect 23492 2366 23612 2394
rect 23848 2382 23900 2388
rect 24124 2440 24176 2446
rect 24124 2382 24176 2388
rect 23204 2304 23256 2310
rect 23204 2246 23256 2252
rect 23166 2204 23474 2213
rect 23166 2202 23172 2204
rect 23228 2202 23252 2204
rect 23308 2202 23332 2204
rect 23388 2202 23412 2204
rect 23468 2202 23474 2204
rect 23228 2150 23230 2202
rect 23410 2150 23412 2202
rect 23166 2148 23172 2150
rect 23228 2148 23252 2150
rect 23308 2148 23332 2150
rect 23388 2148 23412 2150
rect 23468 2148 23474 2150
rect 23166 2139 23474 2148
rect 23112 2100 23164 2106
rect 23112 2042 23164 2048
rect 23020 1828 23072 1834
rect 23020 1770 23072 1776
rect 22652 1760 22704 1766
rect 22572 1720 22652 1748
rect 22284 1488 22336 1494
rect 22284 1430 22336 1436
rect 22468 1420 22520 1426
rect 22468 1362 22520 1368
rect 21086 54 21220 82
rect 21086 -300 21142 54
rect 21454 -300 21510 160
rect 21822 -300 21878 160
rect 22190 82 22246 160
rect 22480 82 22508 1362
rect 22572 160 22600 1720
rect 22652 1702 22704 1708
rect 23124 1290 23152 2042
rect 23584 1970 23612 2366
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 23768 2106 23796 2314
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 23756 2100 23808 2106
rect 23756 2042 23808 2048
rect 23572 1964 23624 1970
rect 23572 1906 23624 1912
rect 24044 1902 24072 2246
rect 24136 2106 24164 2382
rect 24228 2378 24256 2615
rect 24216 2372 24268 2378
rect 24216 2314 24268 2320
rect 24124 2100 24176 2106
rect 24124 2042 24176 2048
rect 24320 1970 24348 4490
rect 24412 2650 24440 8298
rect 24858 4176 24914 4185
rect 24858 4111 24914 4120
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 24584 2440 24636 2446
rect 24584 2382 24636 2388
rect 24596 2038 24624 2382
rect 24872 2038 24900 4111
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25044 3392 25096 3398
rect 25044 3334 25096 3340
rect 24584 2032 24636 2038
rect 24584 1974 24636 1980
rect 24860 2032 24912 2038
rect 24860 1974 24912 1980
rect 24308 1964 24360 1970
rect 24308 1906 24360 1912
rect 24676 1964 24728 1970
rect 24676 1906 24728 1912
rect 24032 1896 24084 1902
rect 24032 1838 24084 1844
rect 23756 1760 23808 1766
rect 23756 1702 23808 1708
rect 24492 1760 24544 1766
rect 24492 1702 24544 1708
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 23112 1284 23164 1290
rect 23112 1226 23164 1232
rect 23020 1216 23072 1222
rect 23020 1158 23072 1164
rect 22190 54 22508 82
rect 22190 -300 22246 54
rect 22558 -300 22614 160
rect 22926 82 22982 160
rect 23032 82 23060 1158
rect 23166 1116 23474 1125
rect 23166 1114 23172 1116
rect 23228 1114 23252 1116
rect 23308 1114 23332 1116
rect 23388 1114 23412 1116
rect 23468 1114 23474 1116
rect 23228 1062 23230 1114
rect 23410 1062 23412 1114
rect 23166 1060 23172 1062
rect 23228 1060 23252 1062
rect 23308 1060 23332 1062
rect 23388 1060 23412 1062
rect 23468 1060 23474 1062
rect 23166 1051 23474 1060
rect 23584 898 23612 1362
rect 23308 870 23612 898
rect 23308 160 23336 870
rect 23572 604 23624 610
rect 23572 546 23624 552
rect 22926 54 23060 82
rect 22926 -300 22982 54
rect 23294 -300 23350 160
rect 23584 134 23612 546
rect 23572 128 23624 134
rect 23572 70 23624 76
rect 23662 82 23718 160
rect 23768 82 23796 1702
rect 24504 1494 24532 1702
rect 24688 1601 24716 1906
rect 24952 1828 25004 1834
rect 24952 1770 25004 1776
rect 24860 1760 24912 1766
rect 24860 1702 24912 1708
rect 24674 1592 24730 1601
rect 24674 1527 24730 1536
rect 24768 1556 24820 1562
rect 24768 1498 24820 1504
rect 24492 1488 24544 1494
rect 24492 1430 24544 1436
rect 24584 1284 24636 1290
rect 24584 1226 24636 1232
rect 24124 1216 24176 1222
rect 24124 1158 24176 1164
rect 23662 54 23796 82
rect 24030 82 24086 160
rect 24136 82 24164 1158
rect 24596 1018 24624 1226
rect 24676 1216 24728 1222
rect 24676 1158 24728 1164
rect 24584 1012 24636 1018
rect 24584 954 24636 960
rect 24030 54 24164 82
rect 24398 82 24454 160
rect 24688 82 24716 1158
rect 24780 160 24808 1498
rect 24872 1426 24900 1702
rect 24860 1420 24912 1426
rect 24860 1362 24912 1368
rect 24964 1290 24992 1770
rect 24952 1284 25004 1290
rect 24952 1226 25004 1232
rect 25056 202 25084 3334
rect 25516 1970 25544 3470
rect 25778 2816 25834 2825
rect 25778 2751 25834 2760
rect 25792 2514 25820 2751
rect 25884 2650 25912 8434
rect 26330 4584 26386 4593
rect 26330 4519 26386 4528
rect 25872 2644 25924 2650
rect 25872 2586 25924 2592
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26160 2106 26188 2382
rect 26148 2100 26200 2106
rect 26148 2042 26200 2048
rect 26344 1970 26372 4519
rect 26608 4480 26660 4486
rect 26608 4422 26660 4428
rect 26620 1970 26648 4422
rect 28000 2632 28028 8434
rect 28720 8188 29028 8197
rect 28720 8186 28726 8188
rect 28782 8186 28806 8188
rect 28862 8186 28886 8188
rect 28942 8186 28966 8188
rect 29022 8186 29028 8188
rect 28782 8134 28784 8186
rect 28964 8134 28966 8186
rect 28720 8132 28726 8134
rect 28782 8132 28806 8134
rect 28862 8132 28886 8134
rect 28942 8132 28966 8134
rect 29022 8132 29028 8134
rect 28720 8123 29028 8132
rect 28720 7100 29028 7109
rect 28720 7098 28726 7100
rect 28782 7098 28806 7100
rect 28862 7098 28886 7100
rect 28942 7098 28966 7100
rect 29022 7098 29028 7100
rect 28782 7046 28784 7098
rect 28964 7046 28966 7098
rect 28720 7044 28726 7046
rect 28782 7044 28806 7046
rect 28862 7044 28886 7046
rect 28942 7044 28966 7046
rect 29022 7044 29028 7046
rect 28720 7035 29028 7044
rect 28720 6012 29028 6021
rect 28720 6010 28726 6012
rect 28782 6010 28806 6012
rect 28862 6010 28886 6012
rect 28942 6010 28966 6012
rect 29022 6010 29028 6012
rect 28782 5958 28784 6010
rect 28964 5958 28966 6010
rect 28720 5956 28726 5958
rect 28782 5956 28806 5958
rect 28862 5956 28886 5958
rect 28942 5956 28966 5958
rect 29022 5956 29028 5958
rect 28720 5947 29028 5956
rect 28720 4924 29028 4933
rect 28720 4922 28726 4924
rect 28782 4922 28806 4924
rect 28862 4922 28886 4924
rect 28942 4922 28966 4924
rect 29022 4922 29028 4924
rect 28782 4870 28784 4922
rect 28964 4870 28966 4922
rect 28720 4868 28726 4870
rect 28782 4868 28806 4870
rect 28862 4868 28886 4870
rect 28942 4868 28966 4870
rect 29022 4868 29028 4870
rect 28720 4859 29028 4868
rect 28720 3836 29028 3845
rect 28720 3834 28726 3836
rect 28782 3834 28806 3836
rect 28862 3834 28886 3836
rect 28942 3834 28966 3836
rect 29022 3834 29028 3836
rect 28782 3782 28784 3834
rect 28964 3782 28966 3834
rect 28720 3780 28726 3782
rect 28782 3780 28806 3782
rect 28862 3780 28886 3782
rect 28942 3780 28966 3782
rect 29022 3780 29028 3782
rect 28720 3771 29028 3780
rect 28632 3460 28684 3466
rect 28632 3402 28684 3408
rect 28080 2644 28132 2650
rect 28000 2604 28080 2632
rect 28080 2586 28132 2592
rect 27896 2576 27948 2582
rect 27896 2518 27948 2524
rect 27804 2440 27856 2446
rect 27804 2382 27856 2388
rect 25136 1964 25188 1970
rect 25136 1906 25188 1912
rect 25504 1964 25556 1970
rect 25504 1906 25556 1912
rect 26332 1964 26384 1970
rect 26332 1906 26384 1912
rect 26608 1964 26660 1970
rect 26608 1906 26660 1912
rect 26700 1964 26752 1970
rect 26700 1906 26752 1912
rect 27068 1964 27120 1970
rect 27068 1906 27120 1912
rect 27620 1964 27672 1970
rect 27620 1906 27672 1912
rect 25148 1306 25176 1906
rect 25780 1828 25832 1834
rect 25780 1770 25832 1776
rect 25412 1556 25464 1562
rect 25412 1498 25464 1504
rect 25148 1278 25268 1306
rect 25136 1216 25188 1222
rect 25136 1158 25188 1164
rect 25044 196 25096 202
rect 24398 54 24716 82
rect 23662 -300 23718 54
rect 24030 -300 24086 54
rect 24398 -300 24454 54
rect 24766 -300 24822 160
rect 25148 160 25176 1158
rect 25240 474 25268 1278
rect 25424 1018 25452 1498
rect 25688 1216 25740 1222
rect 25516 1176 25688 1204
rect 25412 1012 25464 1018
rect 25412 954 25464 960
rect 25228 468 25280 474
rect 25228 410 25280 416
rect 25516 160 25544 1176
rect 25688 1158 25740 1164
rect 25792 814 25820 1770
rect 26056 1760 26108 1766
rect 26056 1702 26108 1708
rect 26148 1760 26200 1766
rect 26148 1702 26200 1708
rect 26516 1760 26568 1766
rect 26516 1702 26568 1708
rect 25780 808 25832 814
rect 25780 750 25832 756
rect 26068 270 26096 1702
rect 26056 264 26108 270
rect 26056 206 26108 212
rect 25044 138 25096 144
rect 25134 -300 25190 160
rect 25502 -300 25558 160
rect 25870 82 25926 160
rect 26160 82 26188 1702
rect 26424 1420 26476 1426
rect 26424 1362 26476 1368
rect 26330 1048 26386 1057
rect 26330 983 26386 992
rect 26344 649 26372 983
rect 26330 640 26386 649
rect 26330 575 26386 584
rect 25870 54 26188 82
rect 26238 82 26294 160
rect 26436 82 26464 1362
rect 26528 1358 26556 1702
rect 26516 1352 26568 1358
rect 26516 1294 26568 1300
rect 26608 1216 26660 1222
rect 26608 1158 26660 1164
rect 26620 160 26648 1158
rect 26712 338 26740 1906
rect 26792 1760 26844 1766
rect 26792 1702 26844 1708
rect 26804 1358 26832 1702
rect 26884 1420 26936 1426
rect 26884 1362 26936 1368
rect 26792 1352 26844 1358
rect 26792 1294 26844 1300
rect 26896 338 26924 1362
rect 27080 882 27108 1906
rect 27632 1850 27660 1906
rect 27540 1822 27660 1850
rect 27160 1760 27212 1766
rect 27160 1702 27212 1708
rect 27252 1760 27304 1766
rect 27252 1702 27304 1708
rect 27172 1358 27200 1702
rect 27264 1562 27292 1702
rect 27252 1556 27304 1562
rect 27252 1498 27304 1504
rect 27344 1556 27396 1562
rect 27344 1498 27396 1504
rect 27160 1352 27212 1358
rect 27160 1294 27212 1300
rect 27252 1216 27304 1222
rect 27252 1158 27304 1164
rect 27068 876 27120 882
rect 27068 818 27120 824
rect 26700 332 26752 338
rect 26700 274 26752 280
rect 26884 332 26936 338
rect 26884 274 26936 280
rect 26988 190 27108 218
rect 26988 160 27016 190
rect 26238 54 26464 82
rect 25870 -300 25926 54
rect 26238 -300 26294 54
rect 26606 -300 26662 160
rect 26974 -300 27030 160
rect 27080 82 27108 190
rect 27264 82 27292 1158
rect 27356 160 27384 1498
rect 27540 1018 27568 1822
rect 27712 1760 27764 1766
rect 27712 1702 27764 1708
rect 27724 1358 27752 1702
rect 27712 1352 27764 1358
rect 27712 1294 27764 1300
rect 27712 1216 27764 1222
rect 27712 1158 27764 1164
rect 27528 1012 27580 1018
rect 27528 954 27580 960
rect 27724 160 27752 1158
rect 27816 678 27844 2382
rect 27908 678 27936 2518
rect 28448 2100 28500 2106
rect 28368 2060 28448 2088
rect 28172 1964 28224 1970
rect 28172 1906 28224 1912
rect 27988 1760 28040 1766
rect 27988 1702 28040 1708
rect 28080 1760 28132 1766
rect 28080 1702 28132 1708
rect 28000 1358 28028 1702
rect 27988 1352 28040 1358
rect 27988 1294 28040 1300
rect 27804 672 27856 678
rect 27804 614 27856 620
rect 27896 672 27948 678
rect 27896 614 27948 620
rect 28092 160 28120 1702
rect 28184 1426 28212 1906
rect 28172 1420 28224 1426
rect 28172 1362 28224 1368
rect 28368 542 28396 2060
rect 28448 2042 28500 2048
rect 28538 1728 28594 1737
rect 28538 1663 28594 1672
rect 28448 1420 28500 1426
rect 28448 1362 28500 1368
rect 28356 536 28408 542
rect 28356 478 28408 484
rect 28460 160 28488 1362
rect 28552 406 28580 1663
rect 28644 746 28672 3402
rect 29092 3120 29144 3126
rect 29092 3062 29144 3068
rect 28720 2748 29028 2757
rect 28720 2746 28726 2748
rect 28782 2746 28806 2748
rect 28862 2746 28886 2748
rect 28942 2746 28966 2748
rect 29022 2746 29028 2748
rect 28782 2694 28784 2746
rect 28964 2694 28966 2746
rect 28720 2692 28726 2694
rect 28782 2692 28806 2694
rect 28862 2692 28886 2694
rect 28942 2692 28966 2694
rect 29022 2692 29028 2694
rect 28720 2683 29028 2692
rect 29104 1970 29132 3062
rect 30104 3052 30156 3058
rect 30104 2994 30156 3000
rect 29184 2644 29236 2650
rect 29184 2586 29236 2592
rect 29196 2446 29224 2586
rect 29184 2440 29236 2446
rect 29184 2382 29236 2388
rect 29276 2372 29328 2378
rect 29276 2314 29328 2320
rect 29288 2145 29316 2314
rect 29274 2136 29330 2145
rect 29274 2071 29330 2080
rect 29092 1964 29144 1970
rect 29092 1906 29144 1912
rect 29368 1964 29420 1970
rect 29368 1906 29420 1912
rect 29644 1964 29696 1970
rect 29644 1906 29696 1912
rect 29828 1964 29880 1970
rect 29828 1906 29880 1912
rect 29092 1828 29144 1834
rect 29092 1770 29144 1776
rect 28720 1660 29028 1669
rect 28720 1658 28726 1660
rect 28782 1658 28806 1660
rect 28862 1658 28886 1660
rect 28942 1658 28966 1660
rect 29022 1658 29028 1660
rect 28782 1606 28784 1658
rect 28964 1606 28966 1658
rect 28720 1604 28726 1606
rect 28782 1604 28806 1606
rect 28862 1604 28886 1606
rect 28942 1604 28966 1606
rect 29022 1604 29028 1606
rect 28720 1595 29028 1604
rect 28816 1556 28868 1562
rect 28816 1498 28868 1504
rect 28632 740 28684 746
rect 28632 682 28684 688
rect 28540 400 28592 406
rect 28540 342 28592 348
rect 28828 160 28856 1498
rect 29000 604 29052 610
rect 29000 546 29052 552
rect 29012 406 29040 546
rect 29000 400 29052 406
rect 29000 342 29052 348
rect 27080 54 27292 82
rect 27342 -300 27398 160
rect 27710 -300 27766 160
rect 28078 -300 28134 160
rect 28446 -300 28502 160
rect 28814 -300 28870 160
rect 29104 82 29132 1770
rect 29184 1760 29236 1766
rect 29184 1702 29236 1708
rect 29276 1760 29328 1766
rect 29276 1702 29328 1708
rect 29196 1358 29224 1702
rect 29288 1358 29316 1702
rect 29184 1352 29236 1358
rect 29184 1294 29236 1300
rect 29276 1352 29328 1358
rect 29276 1294 29328 1300
rect 29380 1193 29408 1906
rect 29552 1760 29604 1766
rect 29552 1702 29604 1708
rect 29564 1426 29592 1702
rect 29552 1420 29604 1426
rect 29552 1362 29604 1368
rect 29552 1284 29604 1290
rect 29552 1226 29604 1232
rect 29366 1184 29422 1193
rect 29366 1119 29422 1128
rect 29564 160 29592 1226
rect 29656 1222 29684 1906
rect 29840 1766 29868 1906
rect 29828 1760 29880 1766
rect 29828 1702 29880 1708
rect 30012 1556 30064 1562
rect 29932 1516 30012 1544
rect 29644 1216 29696 1222
rect 29644 1158 29696 1164
rect 29932 160 29960 1516
rect 30012 1498 30064 1504
rect 30116 950 30144 2994
rect 30288 2848 30340 2854
rect 30288 2790 30340 2796
rect 30300 2582 30328 2790
rect 30392 2650 30420 8434
rect 31390 2952 31446 2961
rect 31390 2887 31446 2896
rect 30380 2644 30432 2650
rect 30380 2586 30432 2592
rect 30472 2644 30524 2650
rect 30472 2586 30524 2592
rect 30288 2576 30340 2582
rect 30288 2518 30340 2524
rect 30484 2514 30512 2586
rect 30472 2508 30524 2514
rect 30472 2450 30524 2456
rect 30656 2440 30708 2446
rect 30656 2382 30708 2388
rect 30932 2440 30984 2446
rect 31208 2440 31260 2446
rect 30984 2400 31064 2428
rect 30932 2382 30984 2388
rect 30564 2304 30616 2310
rect 30562 2272 30564 2281
rect 30616 2272 30618 2281
rect 30562 2207 30618 2216
rect 30564 1964 30616 1970
rect 30564 1906 30616 1912
rect 30472 1760 30524 1766
rect 30472 1702 30524 1708
rect 30380 1420 30432 1426
rect 30380 1362 30432 1368
rect 30392 1306 30420 1362
rect 30484 1358 30512 1702
rect 30300 1278 30420 1306
rect 30472 1352 30524 1358
rect 30472 1294 30524 1300
rect 30104 944 30156 950
rect 30104 886 30156 892
rect 30300 160 30328 1278
rect 30380 1012 30432 1018
rect 30380 954 30432 960
rect 29182 82 29238 160
rect 29104 54 29238 82
rect 29182 -300 29238 54
rect 29550 -300 29606 160
rect 29918 -300 29974 160
rect 30286 -300 30342 160
rect 30392 134 30420 954
rect 30576 785 30604 1906
rect 30668 1018 30696 2382
rect 30840 2304 30892 2310
rect 30840 2246 30892 2252
rect 30852 2106 30880 2246
rect 30840 2100 30892 2106
rect 30840 2042 30892 2048
rect 30852 1970 30972 1986
rect 30840 1964 30972 1970
rect 30892 1958 30972 1964
rect 30840 1906 30892 1912
rect 30840 1828 30892 1834
rect 30840 1770 30892 1776
rect 30748 1760 30800 1766
rect 30748 1702 30800 1708
rect 30760 1358 30788 1702
rect 30748 1352 30800 1358
rect 30748 1294 30800 1300
rect 30656 1012 30708 1018
rect 30656 954 30708 960
rect 30852 898 30880 1770
rect 30668 870 30880 898
rect 30562 776 30618 785
rect 30562 711 30618 720
rect 30668 160 30696 870
rect 30944 377 30972 1958
rect 31036 1850 31064 2400
rect 31208 2382 31260 2388
rect 31116 2304 31168 2310
rect 31116 2246 31168 2252
rect 31128 2106 31156 2246
rect 31116 2100 31168 2106
rect 31116 2042 31168 2048
rect 31036 1822 31156 1850
rect 31024 1760 31076 1766
rect 31024 1702 31076 1708
rect 31036 1358 31064 1702
rect 31024 1352 31076 1358
rect 31024 1294 31076 1300
rect 31128 649 31156 1822
rect 31220 1193 31248 2382
rect 31300 1760 31352 1766
rect 31300 1702 31352 1708
rect 31206 1184 31262 1193
rect 31206 1119 31262 1128
rect 31114 640 31170 649
rect 31114 575 31170 584
rect 30930 368 30986 377
rect 30930 303 30986 312
rect 30380 128 30432 134
rect 30380 70 30432 76
rect 30654 -300 30710 160
rect 31022 82 31078 160
rect 31312 82 31340 1702
rect 31404 1018 31432 2887
rect 32508 2650 32536 8434
rect 34274 7644 34582 7653
rect 34274 7642 34280 7644
rect 34336 7642 34360 7644
rect 34416 7642 34440 7644
rect 34496 7642 34520 7644
rect 34576 7642 34582 7644
rect 34336 7590 34338 7642
rect 34518 7590 34520 7642
rect 34274 7588 34280 7590
rect 34336 7588 34360 7590
rect 34416 7588 34440 7590
rect 34496 7588 34520 7590
rect 34576 7588 34582 7590
rect 34274 7579 34582 7588
rect 34274 6556 34582 6565
rect 34274 6554 34280 6556
rect 34336 6554 34360 6556
rect 34416 6554 34440 6556
rect 34496 6554 34520 6556
rect 34576 6554 34582 6556
rect 34336 6502 34338 6554
rect 34518 6502 34520 6554
rect 34274 6500 34280 6502
rect 34336 6500 34360 6502
rect 34416 6500 34440 6502
rect 34496 6500 34520 6502
rect 34576 6500 34582 6502
rect 34274 6491 34582 6500
rect 34274 5468 34582 5477
rect 34274 5466 34280 5468
rect 34336 5466 34360 5468
rect 34416 5466 34440 5468
rect 34496 5466 34520 5468
rect 34576 5466 34582 5468
rect 34336 5414 34338 5466
rect 34518 5414 34520 5466
rect 34274 5412 34280 5414
rect 34336 5412 34360 5414
rect 34416 5412 34440 5414
rect 34496 5412 34520 5414
rect 34576 5412 34582 5414
rect 34274 5403 34582 5412
rect 34274 4380 34582 4389
rect 34274 4378 34280 4380
rect 34336 4378 34360 4380
rect 34416 4378 34440 4380
rect 34496 4378 34520 4380
rect 34576 4378 34582 4380
rect 34336 4326 34338 4378
rect 34518 4326 34520 4378
rect 34274 4324 34280 4326
rect 34336 4324 34360 4326
rect 34416 4324 34440 4326
rect 34496 4324 34520 4326
rect 34576 4324 34582 4326
rect 34274 4315 34582 4324
rect 34274 3292 34582 3301
rect 34274 3290 34280 3292
rect 34336 3290 34360 3292
rect 34416 3290 34440 3292
rect 34496 3290 34520 3292
rect 34576 3290 34582 3292
rect 34336 3238 34338 3290
rect 34518 3238 34520 3290
rect 34274 3236 34280 3238
rect 34336 3236 34360 3238
rect 34416 3236 34440 3238
rect 34496 3236 34520 3238
rect 34576 3236 34582 3238
rect 34274 3227 34582 3236
rect 32864 2848 32916 2854
rect 32864 2790 32916 2796
rect 32496 2644 32548 2650
rect 32496 2586 32548 2592
rect 32128 2508 32180 2514
rect 32128 2450 32180 2456
rect 31944 2304 31996 2310
rect 32036 2304 32088 2310
rect 31944 2246 31996 2252
rect 32034 2272 32036 2281
rect 32088 2272 32090 2281
rect 31482 2136 31538 2145
rect 31482 2071 31538 2080
rect 31852 2100 31904 2106
rect 31496 1766 31524 2071
rect 31852 2042 31904 2048
rect 31864 1834 31892 2042
rect 31852 1828 31904 1834
rect 31852 1770 31904 1776
rect 31484 1760 31536 1766
rect 31484 1702 31536 1708
rect 31852 1556 31904 1562
rect 31852 1498 31904 1504
rect 31864 1442 31892 1498
rect 31680 1414 31892 1442
rect 31392 1012 31444 1018
rect 31392 954 31444 960
rect 31022 54 31340 82
rect 31390 82 31446 160
rect 31680 82 31708 1414
rect 31956 1358 31984 2246
rect 32034 2207 32090 2216
rect 32140 2106 32168 2450
rect 32312 2440 32364 2446
rect 32312 2382 32364 2388
rect 32772 2440 32824 2446
rect 32772 2382 32824 2388
rect 32128 2100 32180 2106
rect 32128 2042 32180 2048
rect 32324 1970 32352 2382
rect 32784 2106 32812 2382
rect 32772 2100 32824 2106
rect 32772 2042 32824 2048
rect 32876 1970 32904 2790
rect 34808 2650 34836 8434
rect 35256 3664 35308 3670
rect 35256 3606 35308 3612
rect 35162 3088 35218 3097
rect 35162 3023 35218 3032
rect 34796 2644 34848 2650
rect 34796 2586 34848 2592
rect 35072 2576 35124 2582
rect 35072 2518 35124 2524
rect 34980 2440 35032 2446
rect 34980 2382 35032 2388
rect 34274 2204 34582 2213
rect 34274 2202 34280 2204
rect 34336 2202 34360 2204
rect 34416 2202 34440 2204
rect 34496 2202 34520 2204
rect 34576 2202 34582 2204
rect 34336 2150 34338 2202
rect 34518 2150 34520 2202
rect 34274 2148 34280 2150
rect 34336 2148 34360 2150
rect 34416 2148 34440 2150
rect 34496 2148 34520 2150
rect 34576 2148 34582 2150
rect 34274 2139 34582 2148
rect 34992 2106 35020 2382
rect 35084 2310 35112 2518
rect 35072 2304 35124 2310
rect 35072 2246 35124 2252
rect 34980 2100 35032 2106
rect 34980 2042 35032 2048
rect 32312 1964 32364 1970
rect 32312 1906 32364 1912
rect 32864 1964 32916 1970
rect 32864 1906 32916 1912
rect 33508 1964 33560 1970
rect 33508 1906 33560 1912
rect 34060 1964 34112 1970
rect 34060 1906 34112 1912
rect 33232 1828 33284 1834
rect 33232 1770 33284 1776
rect 32404 1760 32456 1766
rect 32404 1702 32456 1708
rect 31944 1352 31996 1358
rect 31944 1294 31996 1300
rect 31760 1216 31812 1222
rect 31760 1158 31812 1164
rect 31772 160 31800 1158
rect 31390 54 31708 82
rect 31022 -300 31078 54
rect 31390 -300 31446 54
rect 31758 -300 31814 160
rect 32126 82 32182 160
rect 32416 82 32444 1702
rect 32772 1556 32824 1562
rect 32772 1498 32824 1504
rect 32126 54 32444 82
rect 32494 82 32550 160
rect 32784 82 32812 1498
rect 32956 1488 33008 1494
rect 32876 1448 32956 1476
rect 32876 160 32904 1448
rect 32956 1430 33008 1436
rect 32956 1216 33008 1222
rect 32956 1158 33008 1164
rect 32968 746 32996 1158
rect 32956 740 33008 746
rect 32956 682 33008 688
rect 33244 160 33272 1770
rect 33520 1766 33548 1906
rect 33508 1760 33560 1766
rect 33508 1702 33560 1708
rect 33876 1760 33928 1766
rect 33876 1702 33928 1708
rect 33324 1284 33376 1290
rect 33324 1226 33376 1232
rect 33416 1284 33468 1290
rect 33416 1226 33468 1232
rect 33336 338 33364 1226
rect 33428 610 33456 1226
rect 33416 604 33468 610
rect 33416 546 33468 552
rect 33324 332 33376 338
rect 33324 274 33376 280
rect 32494 54 32812 82
rect 32126 -300 32182 54
rect 32494 -300 32550 54
rect 32862 -300 32918 160
rect 33230 -300 33286 160
rect 33598 82 33654 160
rect 33888 82 33916 1702
rect 34072 1562 34100 1906
rect 34980 1760 35032 1766
rect 34980 1702 35032 1708
rect 34164 1562 34284 1578
rect 34060 1556 34112 1562
rect 34060 1498 34112 1504
rect 34164 1556 34296 1562
rect 34164 1550 34244 1556
rect 33598 54 33916 82
rect 33966 82 34022 160
rect 34164 82 34192 1550
rect 34244 1498 34296 1504
rect 34704 1488 34756 1494
rect 34624 1448 34704 1476
rect 34274 1116 34582 1125
rect 34274 1114 34280 1116
rect 34336 1114 34360 1116
rect 34416 1114 34440 1116
rect 34496 1114 34520 1116
rect 34576 1114 34582 1116
rect 34336 1062 34338 1114
rect 34518 1062 34520 1114
rect 34274 1060 34280 1062
rect 34336 1060 34360 1062
rect 34416 1060 34440 1062
rect 34496 1060 34520 1062
rect 34576 1060 34582 1062
rect 34274 1051 34582 1060
rect 34624 932 34652 1448
rect 34704 1430 34756 1436
rect 34794 1320 34850 1329
rect 34794 1255 34796 1264
rect 34848 1255 34850 1264
rect 34888 1284 34940 1290
rect 34796 1226 34848 1232
rect 34888 1226 34940 1232
rect 34440 904 34652 932
rect 33966 54 34192 82
rect 34334 82 34390 160
rect 34440 82 34468 904
rect 34900 406 34928 1226
rect 34888 400 34940 406
rect 34888 342 34940 348
rect 34334 54 34468 82
rect 34702 82 34758 160
rect 34992 82 35020 1702
rect 35176 1358 35204 3023
rect 35268 2106 35296 3606
rect 36924 2650 36952 8434
rect 37278 4040 37334 4049
rect 37334 3998 37504 4026
rect 37278 3975 37334 3984
rect 36912 2644 36964 2650
rect 36912 2586 36964 2592
rect 36636 2508 36688 2514
rect 36636 2450 36688 2456
rect 35438 2408 35494 2417
rect 35438 2343 35494 2352
rect 35348 2304 35400 2310
rect 35348 2246 35400 2252
rect 35256 2100 35308 2106
rect 35256 2042 35308 2048
rect 35360 1970 35388 2246
rect 35452 1970 35480 2343
rect 36648 2106 36676 2450
rect 37188 2440 37240 2446
rect 37188 2382 37240 2388
rect 37200 2106 37228 2382
rect 36636 2100 36688 2106
rect 36636 2042 36688 2048
rect 37188 2100 37240 2106
rect 37188 2042 37240 2048
rect 36268 2032 36320 2038
rect 36268 1974 36320 1980
rect 35348 1964 35400 1970
rect 35348 1906 35400 1912
rect 35440 1964 35492 1970
rect 35440 1906 35492 1912
rect 35360 1562 35848 1578
rect 35360 1556 35860 1562
rect 35360 1550 35808 1556
rect 35164 1352 35216 1358
rect 35164 1294 35216 1300
rect 34702 54 35020 82
rect 35070 82 35126 160
rect 35360 82 35388 1550
rect 35808 1498 35860 1504
rect 35716 1488 35768 1494
rect 35716 1430 35768 1436
rect 35440 1284 35492 1290
rect 35440 1226 35492 1232
rect 35452 1018 35480 1226
rect 35440 1012 35492 1018
rect 35440 954 35492 960
rect 35452 190 35572 218
rect 35452 160 35480 190
rect 35070 54 35388 82
rect 33598 -300 33654 54
rect 33966 -300 34022 54
rect 34334 -300 34390 54
rect 34702 -300 34758 54
rect 35070 -300 35126 54
rect 35438 -300 35494 160
rect 35544 82 35572 190
rect 35728 82 35756 1430
rect 35808 1420 35860 1426
rect 35808 1362 35860 1368
rect 35820 160 35848 1362
rect 36280 406 36308 1974
rect 36452 1760 36504 1766
rect 36452 1702 36504 1708
rect 36268 400 36320 406
rect 36268 342 36320 348
rect 35544 54 35756 82
rect 35806 -300 35862 160
rect 36174 82 36230 160
rect 36464 82 36492 1702
rect 37004 1556 37056 1562
rect 37004 1498 37056 1504
rect 37016 1442 37044 1498
rect 37372 1488 37424 1494
rect 36832 1414 37044 1442
rect 37094 1456 37150 1465
rect 36174 54 36492 82
rect 36542 82 36598 160
rect 36832 82 36860 1414
rect 37094 1391 37150 1400
rect 37200 1448 37372 1476
rect 37108 1358 37136 1391
rect 37096 1352 37148 1358
rect 37096 1294 37148 1300
rect 36542 54 36860 82
rect 36910 82 36966 160
rect 37200 82 37228 1448
rect 37372 1430 37424 1436
rect 37476 1290 37504 3998
rect 38106 3632 38162 3641
rect 38106 3567 38162 3576
rect 37830 3496 37886 3505
rect 37830 3431 37886 3440
rect 37648 1828 37700 1834
rect 37648 1770 37700 1776
rect 37556 1760 37608 1766
rect 37556 1702 37608 1708
rect 37464 1284 37516 1290
rect 37464 1226 37516 1232
rect 36910 54 37228 82
rect 37278 82 37334 160
rect 37568 82 37596 1702
rect 37660 160 37688 1770
rect 37844 1290 37872 3431
rect 37924 1964 37976 1970
rect 37924 1906 37976 1912
rect 38016 1964 38068 1970
rect 38016 1906 38068 1912
rect 37936 1426 37964 1906
rect 38028 1873 38056 1906
rect 38014 1864 38070 1873
rect 38014 1799 38070 1808
rect 37924 1420 37976 1426
rect 37924 1362 37976 1368
rect 38120 1290 38148 3567
rect 39040 2650 39068 8434
rect 39828 8188 40136 8197
rect 39828 8186 39834 8188
rect 39890 8186 39914 8188
rect 39970 8186 39994 8188
rect 40050 8186 40074 8188
rect 40130 8186 40136 8188
rect 39890 8134 39892 8186
rect 40072 8134 40074 8186
rect 39828 8132 39834 8134
rect 39890 8132 39914 8134
rect 39970 8132 39994 8134
rect 40050 8132 40074 8134
rect 40130 8132 40136 8134
rect 39828 8123 40136 8132
rect 39828 7100 40136 7109
rect 39828 7098 39834 7100
rect 39890 7098 39914 7100
rect 39970 7098 39994 7100
rect 40050 7098 40074 7100
rect 40130 7098 40136 7100
rect 39890 7046 39892 7098
rect 40072 7046 40074 7098
rect 39828 7044 39834 7046
rect 39890 7044 39914 7046
rect 39970 7044 39994 7046
rect 40050 7044 40074 7046
rect 40130 7044 40136 7046
rect 39828 7035 40136 7044
rect 39828 6012 40136 6021
rect 39828 6010 39834 6012
rect 39890 6010 39914 6012
rect 39970 6010 39994 6012
rect 40050 6010 40074 6012
rect 40130 6010 40136 6012
rect 39890 5958 39892 6010
rect 40072 5958 40074 6010
rect 39828 5956 39834 5958
rect 39890 5956 39914 5958
rect 39970 5956 39994 5958
rect 40050 5956 40074 5958
rect 40130 5956 40136 5958
rect 39828 5947 40136 5956
rect 39828 4924 40136 4933
rect 39828 4922 39834 4924
rect 39890 4922 39914 4924
rect 39970 4922 39994 4924
rect 40050 4922 40074 4924
rect 40130 4922 40136 4924
rect 39890 4870 39892 4922
rect 40072 4870 40074 4922
rect 39828 4868 39834 4870
rect 39890 4868 39914 4870
rect 39970 4868 39994 4870
rect 40050 4868 40074 4870
rect 40130 4868 40136 4870
rect 39828 4859 40136 4868
rect 41144 4208 41196 4214
rect 41144 4150 41196 4156
rect 39828 3836 40136 3845
rect 39828 3834 39834 3836
rect 39890 3834 39914 3836
rect 39970 3834 39994 3836
rect 40050 3834 40074 3836
rect 40130 3834 40136 3836
rect 39890 3782 39892 3834
rect 40072 3782 40074 3834
rect 39828 3780 39834 3782
rect 39890 3780 39914 3782
rect 39970 3780 39994 3782
rect 40050 3780 40074 3782
rect 40130 3780 40136 3782
rect 39828 3771 40136 3780
rect 39672 3188 39724 3194
rect 39672 3130 39724 3136
rect 39028 2644 39080 2650
rect 39028 2586 39080 2592
rect 39304 2440 39356 2446
rect 39304 2382 39356 2388
rect 39316 2106 39344 2382
rect 39304 2100 39356 2106
rect 39304 2042 39356 2048
rect 38382 2000 38438 2009
rect 38382 1935 38384 1944
rect 38436 1935 38438 1944
rect 38384 1906 38436 1912
rect 39212 1896 39264 1902
rect 39212 1838 39264 1844
rect 39580 1896 39632 1902
rect 39580 1838 39632 1844
rect 39224 1562 39252 1838
rect 38292 1556 38344 1562
rect 38292 1498 38344 1504
rect 39212 1556 39264 1562
rect 39212 1498 39264 1504
rect 37832 1284 37884 1290
rect 37832 1226 37884 1232
rect 38108 1284 38160 1290
rect 38108 1226 38160 1232
rect 38028 190 38148 218
rect 38028 160 38056 190
rect 37278 54 37596 82
rect 36174 -300 36230 54
rect 36542 -300 36598 54
rect 36910 -300 36966 54
rect 37278 -300 37334 54
rect 37646 -300 37702 160
rect 38014 -300 38070 160
rect 38120 82 38148 190
rect 38304 82 38332 1498
rect 38844 1488 38896 1494
rect 38396 1448 38844 1476
rect 38396 160 38424 1448
rect 38844 1430 38896 1436
rect 38752 1352 38804 1358
rect 38752 1294 38804 1300
rect 38764 160 38792 1294
rect 39212 1284 39264 1290
rect 39132 1244 39212 1272
rect 39132 160 39160 1244
rect 39212 1226 39264 1232
rect 39304 1216 39356 1222
rect 39304 1158 39356 1164
rect 39396 1216 39448 1222
rect 39396 1158 39448 1164
rect 39316 950 39344 1158
rect 39304 944 39356 950
rect 39304 886 39356 892
rect 39408 814 39436 1158
rect 39592 1034 39620 1838
rect 39684 1222 39712 3130
rect 39828 2748 40136 2757
rect 39828 2746 39834 2748
rect 39890 2746 39914 2748
rect 39970 2746 39994 2748
rect 40050 2746 40074 2748
rect 40130 2746 40136 2748
rect 39890 2694 39892 2746
rect 40072 2694 40074 2746
rect 39828 2692 39834 2694
rect 39890 2692 39914 2694
rect 39970 2692 39994 2694
rect 40050 2692 40074 2694
rect 40130 2692 40136 2694
rect 39828 2683 40136 2692
rect 40408 2576 40460 2582
rect 40130 2544 40186 2553
rect 40408 2518 40460 2524
rect 40130 2479 40186 2488
rect 40144 2106 40172 2479
rect 40420 2106 40448 2518
rect 40684 2508 40736 2514
rect 40684 2450 40736 2456
rect 40696 2106 40724 2450
rect 40132 2100 40184 2106
rect 40132 2042 40184 2048
rect 40408 2100 40460 2106
rect 40408 2042 40460 2048
rect 40684 2100 40736 2106
rect 40684 2042 40736 2048
rect 40592 1964 40644 1970
rect 40328 1924 40592 1952
rect 39828 1660 40136 1669
rect 39828 1658 39834 1660
rect 39890 1658 39914 1660
rect 39970 1658 39994 1660
rect 40050 1658 40074 1660
rect 40130 1658 40136 1660
rect 39890 1606 39892 1658
rect 40072 1606 40074 1658
rect 39828 1604 39834 1606
rect 39890 1604 39914 1606
rect 39970 1604 39994 1606
rect 40050 1604 40074 1606
rect 40130 1604 40136 1606
rect 39828 1595 40136 1604
rect 40328 1442 40356 1924
rect 40592 1906 40644 1912
rect 40500 1828 40552 1834
rect 40500 1770 40552 1776
rect 39868 1414 40356 1442
rect 39672 1216 39724 1222
rect 39672 1158 39724 1164
rect 39500 1006 39620 1034
rect 39396 808 39448 814
rect 39396 750 39448 756
rect 39500 160 39528 1006
rect 39868 160 39896 1414
rect 40040 1216 40092 1222
rect 40040 1158 40092 1164
rect 40052 1018 40080 1158
rect 40040 1012 40092 1018
rect 40040 954 40092 960
rect 38120 54 38332 82
rect 38382 -300 38438 160
rect 38750 -300 38806 160
rect 39118 -300 39174 160
rect 39486 -300 39542 160
rect 39854 -300 39910 160
rect 40222 82 40278 160
rect 40512 82 40540 1770
rect 41156 1358 41184 4150
rect 41340 2650 41368 8434
rect 42432 4276 42484 4282
rect 42432 4218 42484 4224
rect 41328 2644 41380 2650
rect 41328 2586 41380 2592
rect 41512 2440 41564 2446
rect 41512 2382 41564 2388
rect 41524 2106 41552 2382
rect 41512 2100 41564 2106
rect 41512 2042 41564 2048
rect 42444 1562 42472 4218
rect 43548 2650 43576 8434
rect 44560 2650 44588 8434
rect 45382 7644 45690 7653
rect 45382 7642 45388 7644
rect 45444 7642 45468 7644
rect 45524 7642 45548 7644
rect 45604 7642 45628 7644
rect 45684 7642 45690 7644
rect 45444 7590 45446 7642
rect 45626 7590 45628 7642
rect 45382 7588 45388 7590
rect 45444 7588 45468 7590
rect 45524 7588 45548 7590
rect 45604 7588 45628 7590
rect 45684 7588 45690 7590
rect 45382 7579 45690 7588
rect 45382 6556 45690 6565
rect 45382 6554 45388 6556
rect 45444 6554 45468 6556
rect 45524 6554 45548 6556
rect 45604 6554 45628 6556
rect 45684 6554 45690 6556
rect 45444 6502 45446 6554
rect 45626 6502 45628 6554
rect 45382 6500 45388 6502
rect 45444 6500 45468 6502
rect 45524 6500 45548 6502
rect 45604 6500 45628 6502
rect 45684 6500 45690 6502
rect 45382 6491 45690 6500
rect 45382 5468 45690 5477
rect 45382 5466 45388 5468
rect 45444 5466 45468 5468
rect 45524 5466 45548 5468
rect 45604 5466 45628 5468
rect 45684 5466 45690 5468
rect 45444 5414 45446 5466
rect 45626 5414 45628 5466
rect 45382 5412 45388 5414
rect 45444 5412 45468 5414
rect 45524 5412 45548 5414
rect 45604 5412 45628 5414
rect 45684 5412 45690 5414
rect 45382 5403 45690 5412
rect 45382 4380 45690 4389
rect 45382 4378 45388 4380
rect 45444 4378 45468 4380
rect 45524 4378 45548 4380
rect 45604 4378 45628 4380
rect 45684 4378 45690 4380
rect 45444 4326 45446 4378
rect 45626 4326 45628 4378
rect 45382 4324 45388 4326
rect 45444 4324 45468 4326
rect 45524 4324 45548 4326
rect 45604 4324 45628 4326
rect 45684 4324 45690 4326
rect 45382 4315 45690 4324
rect 45382 3292 45690 3301
rect 45382 3290 45388 3292
rect 45444 3290 45468 3292
rect 45524 3290 45548 3292
rect 45604 3290 45628 3292
rect 45684 3290 45690 3292
rect 45444 3238 45446 3290
rect 45626 3238 45628 3290
rect 45382 3236 45388 3238
rect 45444 3236 45468 3238
rect 45524 3236 45548 3238
rect 45604 3236 45628 3238
rect 45684 3236 45690 3238
rect 45382 3227 45690 3236
rect 43536 2644 43588 2650
rect 43536 2586 43588 2592
rect 44548 2644 44600 2650
rect 44548 2586 44600 2592
rect 43996 2440 44048 2446
rect 43996 2382 44048 2388
rect 44364 2440 44416 2446
rect 44364 2382 44416 2388
rect 45100 2440 45152 2446
rect 45100 2382 45152 2388
rect 46112 2440 46164 2446
rect 46112 2382 46164 2388
rect 43536 2372 43588 2378
rect 43536 2314 43588 2320
rect 42524 1896 42576 1902
rect 42524 1838 42576 1844
rect 42536 1562 42564 1838
rect 42432 1556 42484 1562
rect 42432 1498 42484 1504
rect 42524 1556 42576 1562
rect 42524 1498 42576 1504
rect 43548 1494 43576 2314
rect 44008 2106 44036 2382
rect 44180 2304 44232 2310
rect 44180 2246 44232 2252
rect 43996 2100 44048 2106
rect 43996 2042 44048 2048
rect 43812 1760 43864 1766
rect 43812 1702 43864 1708
rect 43824 1494 43852 1702
rect 44192 1494 44220 2246
rect 44376 1970 44404 2382
rect 44640 2304 44692 2310
rect 44640 2246 44692 2252
rect 45008 2304 45060 2310
rect 45008 2246 45060 2252
rect 44652 2106 44680 2246
rect 45020 2106 45048 2246
rect 44640 2100 44692 2106
rect 44640 2042 44692 2048
rect 45008 2100 45060 2106
rect 45008 2042 45060 2048
rect 44364 1964 44416 1970
rect 44364 1906 44416 1912
rect 43536 1488 43588 1494
rect 43536 1430 43588 1436
rect 43812 1488 43864 1494
rect 43812 1430 43864 1436
rect 44180 1488 44232 1494
rect 44180 1430 44232 1436
rect 42708 1420 42760 1426
rect 42708 1362 42760 1368
rect 41144 1352 41196 1358
rect 41144 1294 41196 1300
rect 41236 1352 41288 1358
rect 41236 1294 41288 1300
rect 41972 1352 42024 1358
rect 41972 1294 42024 1300
rect 40592 1012 40644 1018
rect 40592 954 40644 960
rect 40604 160 40632 954
rect 40222 54 40540 82
rect 40222 -300 40278 54
rect 40590 -300 40646 160
rect 40958 82 41014 160
rect 41248 82 41276 1294
rect 41328 1284 41380 1290
rect 41328 1226 41380 1232
rect 41696 1284 41748 1290
rect 41696 1226 41748 1232
rect 41340 160 41368 1226
rect 41708 160 41736 1226
rect 41984 1018 42012 1294
rect 42064 1216 42116 1222
rect 42064 1158 42116 1164
rect 42340 1216 42392 1222
rect 42340 1158 42392 1164
rect 42524 1216 42576 1222
rect 42524 1158 42576 1164
rect 41972 1012 42024 1018
rect 41972 954 42024 960
rect 42076 814 42104 1158
rect 42064 808 42116 814
rect 42064 750 42116 756
rect 40958 54 41276 82
rect 40958 -300 41014 54
rect 41326 -300 41382 160
rect 41694 -300 41750 160
rect 42062 82 42118 160
rect 42352 82 42380 1158
rect 42536 1018 42564 1158
rect 42524 1012 42576 1018
rect 42524 954 42576 960
rect 42062 54 42380 82
rect 42430 82 42486 160
rect 42720 82 42748 1362
rect 44272 1352 44324 1358
rect 44272 1294 44324 1300
rect 44548 1352 44600 1358
rect 44548 1294 44600 1300
rect 44824 1352 44876 1358
rect 44824 1294 44876 1300
rect 42800 1284 42852 1290
rect 43352 1284 43404 1290
rect 42800 1226 42852 1232
rect 43180 1244 43352 1272
rect 42812 160 42840 1226
rect 42984 1216 43036 1222
rect 42984 1158 43036 1164
rect 43076 1216 43128 1222
rect 43076 1158 43128 1164
rect 42996 814 43024 1158
rect 43088 1018 43116 1158
rect 43076 1012 43128 1018
rect 43076 954 43128 960
rect 42984 808 43036 814
rect 42984 750 43036 756
rect 43180 160 43208 1244
rect 43628 1284 43680 1290
rect 43352 1226 43404 1232
rect 43548 1244 43628 1272
rect 43548 160 43576 1244
rect 43628 1226 43680 1232
rect 44088 1216 44140 1222
rect 44088 1158 44140 1164
rect 44100 406 44128 1158
rect 44284 490 44312 1294
rect 44192 462 44312 490
rect 44088 400 44140 406
rect 44088 342 44140 348
rect 42430 54 42748 82
rect 42062 -300 42118 54
rect 42430 -300 42486 54
rect 42798 -300 42854 160
rect 43166 -300 43222 160
rect 43534 -300 43590 160
rect 43902 82 43958 160
rect 44192 82 44220 462
rect 44284 190 44404 218
rect 44284 160 44312 190
rect 43902 54 44220 82
rect 43902 -300 43958 54
rect 44270 -300 44326 160
rect 44376 82 44404 190
rect 44560 82 44588 1294
rect 44732 1284 44784 1290
rect 44732 1226 44784 1232
rect 44376 54 44588 82
rect 44638 82 44694 160
rect 44744 82 44772 1226
rect 44638 54 44772 82
rect 44836 82 44864 1294
rect 45006 82 45062 160
rect 44836 54 45062 82
rect 45112 82 45140 2382
rect 45382 2204 45690 2213
rect 45382 2202 45388 2204
rect 45444 2202 45468 2204
rect 45524 2202 45548 2204
rect 45604 2202 45628 2204
rect 45684 2202 45690 2204
rect 45444 2150 45446 2202
rect 45626 2150 45628 2202
rect 45382 2148 45388 2150
rect 45444 2148 45468 2150
rect 45524 2148 45548 2150
rect 45604 2148 45628 2150
rect 45684 2148 45690 2150
rect 45382 2139 45690 2148
rect 45744 1964 45796 1970
rect 45744 1906 45796 1912
rect 45382 1116 45690 1125
rect 45382 1114 45388 1116
rect 45444 1114 45468 1116
rect 45524 1114 45548 1116
rect 45604 1114 45628 1116
rect 45684 1114 45690 1116
rect 45444 1062 45446 1114
rect 45626 1062 45628 1114
rect 45382 1060 45388 1062
rect 45444 1060 45468 1062
rect 45524 1060 45548 1062
rect 45604 1060 45628 1062
rect 45684 1060 45690 1062
rect 45382 1051 45690 1060
rect 45756 160 45784 1906
rect 46124 160 46152 2382
rect 45374 82 45430 160
rect 45112 54 45430 82
rect 44638 -300 44694 54
rect 45006 -300 45062 54
rect 45374 -300 45430 54
rect 45742 -300 45798 160
rect 46110 -300 46166 160
<< via2 >>
rect 12064 8730 12120 8732
rect 12144 8730 12200 8732
rect 12224 8730 12280 8732
rect 12304 8730 12360 8732
rect 12064 8678 12110 8730
rect 12110 8678 12120 8730
rect 12144 8678 12174 8730
rect 12174 8678 12186 8730
rect 12186 8678 12200 8730
rect 12224 8678 12238 8730
rect 12238 8678 12250 8730
rect 12250 8678 12280 8730
rect 12304 8678 12314 8730
rect 12314 8678 12360 8730
rect 12064 8676 12120 8678
rect 12144 8676 12200 8678
rect 12224 8676 12280 8678
rect 12304 8676 12360 8678
rect 6510 8186 6566 8188
rect 6590 8186 6646 8188
rect 6670 8186 6726 8188
rect 6750 8186 6806 8188
rect 6510 8134 6556 8186
rect 6556 8134 6566 8186
rect 6590 8134 6620 8186
rect 6620 8134 6632 8186
rect 6632 8134 6646 8186
rect 6670 8134 6684 8186
rect 6684 8134 6696 8186
rect 6696 8134 6726 8186
rect 6750 8134 6760 8186
rect 6760 8134 6806 8186
rect 6510 8132 6566 8134
rect 6590 8132 6646 8134
rect 6670 8132 6726 8134
rect 6750 8132 6806 8134
rect 12064 7642 12120 7644
rect 12144 7642 12200 7644
rect 12224 7642 12280 7644
rect 12304 7642 12360 7644
rect 12064 7590 12110 7642
rect 12110 7590 12120 7642
rect 12144 7590 12174 7642
rect 12174 7590 12186 7642
rect 12186 7590 12200 7642
rect 12224 7590 12238 7642
rect 12238 7590 12250 7642
rect 12250 7590 12280 7642
rect 12304 7590 12314 7642
rect 12314 7590 12360 7642
rect 12064 7588 12120 7590
rect 12144 7588 12200 7590
rect 12224 7588 12280 7590
rect 12304 7588 12360 7590
rect 6510 7098 6566 7100
rect 6590 7098 6646 7100
rect 6670 7098 6726 7100
rect 6750 7098 6806 7100
rect 6510 7046 6556 7098
rect 6556 7046 6566 7098
rect 6590 7046 6620 7098
rect 6620 7046 6632 7098
rect 6632 7046 6646 7098
rect 6670 7046 6684 7098
rect 6684 7046 6696 7098
rect 6696 7046 6726 7098
rect 6750 7046 6760 7098
rect 6760 7046 6806 7098
rect 6510 7044 6566 7046
rect 6590 7044 6646 7046
rect 6670 7044 6726 7046
rect 6750 7044 6806 7046
rect 12064 6554 12120 6556
rect 12144 6554 12200 6556
rect 12224 6554 12280 6556
rect 12304 6554 12360 6556
rect 12064 6502 12110 6554
rect 12110 6502 12120 6554
rect 12144 6502 12174 6554
rect 12174 6502 12186 6554
rect 12186 6502 12200 6554
rect 12224 6502 12238 6554
rect 12238 6502 12250 6554
rect 12250 6502 12280 6554
rect 12304 6502 12314 6554
rect 12314 6502 12360 6554
rect 12064 6500 12120 6502
rect 12144 6500 12200 6502
rect 12224 6500 12280 6502
rect 12304 6500 12360 6502
rect 6510 6010 6566 6012
rect 6590 6010 6646 6012
rect 6670 6010 6726 6012
rect 6750 6010 6806 6012
rect 6510 5958 6556 6010
rect 6556 5958 6566 6010
rect 6590 5958 6620 6010
rect 6620 5958 6632 6010
rect 6632 5958 6646 6010
rect 6670 5958 6684 6010
rect 6684 5958 6696 6010
rect 6696 5958 6726 6010
rect 6750 5958 6760 6010
rect 6760 5958 6806 6010
rect 6510 5956 6566 5958
rect 6590 5956 6646 5958
rect 6670 5956 6726 5958
rect 6750 5956 6806 5958
rect 12064 5466 12120 5468
rect 12144 5466 12200 5468
rect 12224 5466 12280 5468
rect 12304 5466 12360 5468
rect 12064 5414 12110 5466
rect 12110 5414 12120 5466
rect 12144 5414 12174 5466
rect 12174 5414 12186 5466
rect 12186 5414 12200 5466
rect 12224 5414 12238 5466
rect 12238 5414 12250 5466
rect 12250 5414 12280 5466
rect 12304 5414 12314 5466
rect 12314 5414 12360 5466
rect 12064 5412 12120 5414
rect 12144 5412 12200 5414
rect 12224 5412 12280 5414
rect 12304 5412 12360 5414
rect 6510 4922 6566 4924
rect 6590 4922 6646 4924
rect 6670 4922 6726 4924
rect 6750 4922 6806 4924
rect 6510 4870 6556 4922
rect 6556 4870 6566 4922
rect 6590 4870 6620 4922
rect 6620 4870 6632 4922
rect 6632 4870 6646 4922
rect 6670 4870 6684 4922
rect 6684 4870 6696 4922
rect 6696 4870 6726 4922
rect 6750 4870 6760 4922
rect 6760 4870 6806 4922
rect 6510 4868 6566 4870
rect 6590 4868 6646 4870
rect 6670 4868 6726 4870
rect 6750 4868 6806 4870
rect 4710 4528 4766 4584
rect 1858 2488 1914 2544
rect 3790 4120 3846 4176
rect 12064 4378 12120 4380
rect 12144 4378 12200 4380
rect 12224 4378 12280 4380
rect 12304 4378 12360 4380
rect 12064 4326 12110 4378
rect 12110 4326 12120 4378
rect 12144 4326 12174 4378
rect 12174 4326 12186 4378
rect 12186 4326 12200 4378
rect 12224 4326 12238 4378
rect 12238 4326 12250 4378
rect 12250 4326 12280 4378
rect 12304 4326 12314 4378
rect 12314 4326 12360 4378
rect 12064 4324 12120 4326
rect 12144 4324 12200 4326
rect 12224 4324 12280 4326
rect 12304 4324 12360 4326
rect 11886 3984 11942 4040
rect 6510 3834 6566 3836
rect 6590 3834 6646 3836
rect 6670 3834 6726 3836
rect 6750 3834 6806 3836
rect 6510 3782 6556 3834
rect 6556 3782 6566 3834
rect 6590 3782 6620 3834
rect 6620 3782 6632 3834
rect 6632 3782 6646 3834
rect 6670 3782 6684 3834
rect 6684 3782 6696 3834
rect 6696 3782 6726 3834
rect 6750 3782 6760 3834
rect 6760 3782 6806 3834
rect 6510 3780 6566 3782
rect 6590 3780 6646 3782
rect 6670 3780 6726 3782
rect 6750 3780 6806 3782
rect 6510 2746 6566 2748
rect 6590 2746 6646 2748
rect 6670 2746 6726 2748
rect 6750 2746 6806 2748
rect 6510 2694 6556 2746
rect 6556 2694 6566 2746
rect 6590 2694 6620 2746
rect 6620 2694 6632 2746
rect 6632 2694 6646 2746
rect 6670 2694 6684 2746
rect 6684 2694 6696 2746
rect 6696 2694 6726 2746
rect 6750 2694 6760 2746
rect 6760 2694 6806 2746
rect 6510 2692 6566 2694
rect 6590 2692 6646 2694
rect 6670 2692 6726 2694
rect 6750 2692 6806 2694
rect 6510 1658 6566 1660
rect 6590 1658 6646 1660
rect 6670 1658 6726 1660
rect 6750 1658 6806 1660
rect 6510 1606 6556 1658
rect 6556 1606 6566 1658
rect 6590 1606 6620 1658
rect 6620 1606 6632 1658
rect 6632 1606 6646 1658
rect 6670 1606 6684 1658
rect 6684 1606 6696 1658
rect 6696 1606 6726 1658
rect 6750 1606 6760 1658
rect 6760 1606 6806 1658
rect 6510 1604 6566 1606
rect 6590 1604 6646 1606
rect 6670 1604 6726 1606
rect 6750 1604 6806 1606
rect 12064 3290 12120 3292
rect 12144 3290 12200 3292
rect 12224 3290 12280 3292
rect 12304 3290 12360 3292
rect 12064 3238 12110 3290
rect 12110 3238 12120 3290
rect 12144 3238 12174 3290
rect 12174 3238 12186 3290
rect 12186 3238 12200 3290
rect 12224 3238 12238 3290
rect 12238 3238 12250 3290
rect 12250 3238 12280 3290
rect 12304 3238 12314 3290
rect 12314 3238 12360 3290
rect 12064 3236 12120 3238
rect 12144 3236 12200 3238
rect 12224 3236 12280 3238
rect 12304 3236 12360 3238
rect 13358 3168 13414 3224
rect 9954 2352 10010 2408
rect 8942 1944 8998 2000
rect 8758 856 8814 912
rect 9218 584 9274 640
rect 9586 448 9642 504
rect 10322 312 10378 368
rect 10690 720 10746 776
rect 11702 1264 11758 1320
rect 12064 2202 12120 2204
rect 12144 2202 12200 2204
rect 12224 2202 12280 2204
rect 12304 2202 12360 2204
rect 12064 2150 12110 2202
rect 12110 2150 12120 2202
rect 12144 2150 12174 2202
rect 12174 2150 12186 2202
rect 12186 2150 12200 2202
rect 12224 2150 12238 2202
rect 12238 2150 12250 2202
rect 12250 2150 12280 2202
rect 12304 2150 12314 2202
rect 12314 2150 12360 2202
rect 12064 2148 12120 2150
rect 12144 2148 12200 2150
rect 12224 2148 12280 2150
rect 12304 2148 12360 2150
rect 12064 1114 12120 1116
rect 12144 1114 12200 1116
rect 12224 1114 12280 1116
rect 12304 1114 12360 1116
rect 12064 1062 12110 1114
rect 12110 1062 12120 1114
rect 12144 1062 12174 1114
rect 12174 1062 12186 1114
rect 12186 1062 12200 1114
rect 12224 1062 12238 1114
rect 12238 1062 12250 1114
rect 12250 1062 12280 1114
rect 12304 1062 12314 1114
rect 12314 1062 12360 1114
rect 12064 1060 12120 1062
rect 12144 1060 12200 1062
rect 12224 1060 12280 1062
rect 12304 1060 12360 1062
rect 12806 1164 12808 1184
rect 12808 1164 12860 1184
rect 12860 1164 12862 1184
rect 12806 1128 12862 1164
rect 12714 992 12770 1048
rect 15934 3576 15990 3632
rect 15198 1808 15254 1864
rect 14830 1400 14886 1456
rect 16486 2216 16542 2272
rect 17618 8186 17674 8188
rect 17698 8186 17754 8188
rect 17778 8186 17834 8188
rect 17858 8186 17914 8188
rect 17618 8134 17664 8186
rect 17664 8134 17674 8186
rect 17698 8134 17728 8186
rect 17728 8134 17740 8186
rect 17740 8134 17754 8186
rect 17778 8134 17792 8186
rect 17792 8134 17804 8186
rect 17804 8134 17834 8186
rect 17858 8134 17868 8186
rect 17868 8134 17914 8186
rect 17618 8132 17674 8134
rect 17698 8132 17754 8134
rect 17778 8132 17834 8134
rect 17858 8132 17914 8134
rect 17618 7098 17674 7100
rect 17698 7098 17754 7100
rect 17778 7098 17834 7100
rect 17858 7098 17914 7100
rect 17618 7046 17664 7098
rect 17664 7046 17674 7098
rect 17698 7046 17728 7098
rect 17728 7046 17740 7098
rect 17740 7046 17754 7098
rect 17778 7046 17792 7098
rect 17792 7046 17804 7098
rect 17804 7046 17834 7098
rect 17858 7046 17868 7098
rect 17868 7046 17914 7098
rect 17618 7044 17674 7046
rect 17698 7044 17754 7046
rect 17778 7044 17834 7046
rect 17858 7044 17914 7046
rect 17618 6010 17674 6012
rect 17698 6010 17754 6012
rect 17778 6010 17834 6012
rect 17858 6010 17914 6012
rect 17618 5958 17664 6010
rect 17664 5958 17674 6010
rect 17698 5958 17728 6010
rect 17728 5958 17740 6010
rect 17740 5958 17754 6010
rect 17778 5958 17792 6010
rect 17792 5958 17804 6010
rect 17804 5958 17834 6010
rect 17858 5958 17868 6010
rect 17868 5958 17914 6010
rect 17618 5956 17674 5958
rect 17698 5956 17754 5958
rect 17778 5956 17834 5958
rect 17858 5956 17914 5958
rect 17618 4922 17674 4924
rect 17698 4922 17754 4924
rect 17778 4922 17834 4924
rect 17858 4922 17914 4924
rect 17618 4870 17664 4922
rect 17664 4870 17674 4922
rect 17698 4870 17728 4922
rect 17728 4870 17740 4922
rect 17740 4870 17754 4922
rect 17778 4870 17792 4922
rect 17792 4870 17804 4922
rect 17804 4870 17834 4922
rect 17858 4870 17868 4922
rect 17868 4870 17914 4922
rect 17618 4868 17674 4870
rect 17698 4868 17754 4870
rect 17778 4868 17834 4870
rect 17858 4868 17914 4870
rect 17618 3834 17674 3836
rect 17698 3834 17754 3836
rect 17778 3834 17834 3836
rect 17858 3834 17914 3836
rect 17618 3782 17664 3834
rect 17664 3782 17674 3834
rect 17698 3782 17728 3834
rect 17728 3782 17740 3834
rect 17740 3782 17754 3834
rect 17778 3782 17792 3834
rect 17792 3782 17804 3834
rect 17804 3782 17834 3834
rect 17858 3782 17868 3834
rect 17868 3782 17914 3834
rect 17618 3780 17674 3782
rect 17698 3780 17754 3782
rect 17778 3780 17834 3782
rect 17858 3780 17914 3782
rect 17130 3032 17186 3088
rect 17314 2896 17370 2952
rect 17618 2746 17674 2748
rect 17698 2746 17754 2748
rect 17778 2746 17834 2748
rect 17858 2746 17914 2748
rect 17618 2694 17664 2746
rect 17664 2694 17674 2746
rect 17698 2694 17728 2746
rect 17728 2694 17740 2746
rect 17740 2694 17754 2746
rect 17778 2694 17792 2746
rect 17792 2694 17804 2746
rect 17804 2694 17834 2746
rect 17858 2694 17868 2746
rect 17868 2694 17914 2746
rect 17618 2692 17674 2694
rect 17698 2692 17754 2694
rect 17778 2692 17834 2694
rect 17858 2692 17914 2694
rect 18050 2624 18106 2680
rect 17618 1658 17674 1660
rect 17698 1658 17754 1660
rect 17778 1658 17834 1660
rect 17858 1658 17914 1660
rect 17618 1606 17664 1658
rect 17664 1606 17674 1658
rect 17698 1606 17728 1658
rect 17728 1606 17740 1658
rect 17740 1606 17754 1658
rect 17778 1606 17792 1658
rect 17792 1606 17804 1658
rect 17804 1606 17834 1658
rect 17858 1606 17868 1658
rect 17868 1606 17914 1658
rect 17618 1604 17674 1606
rect 17698 1604 17754 1606
rect 17778 1604 17834 1606
rect 17858 1604 17914 1606
rect 17866 1128 17922 1184
rect 18050 1128 18106 1184
rect 18694 3440 18750 3496
rect 18786 2488 18842 2544
rect 20534 3848 20590 3904
rect 19890 2624 19946 2680
rect 19246 1944 19302 2000
rect 19706 1708 19708 1728
rect 19708 1708 19760 1728
rect 19760 1708 19762 1728
rect 19706 1672 19762 1708
rect 18878 1300 18880 1320
rect 18880 1300 18932 1320
rect 18932 1300 18934 1320
rect 18878 1264 18934 1300
rect 22098 3168 22154 3224
rect 22006 2644 22062 2680
rect 22006 2624 22008 2644
rect 22008 2624 22060 2644
rect 22060 2624 22062 2644
rect 21546 2488 21602 2544
rect 20718 2352 20774 2408
rect 20626 2216 20682 2272
rect 20350 1400 20406 1456
rect 21454 2080 21510 2136
rect 22190 2352 22246 2408
rect 22558 3984 22614 4040
rect 21730 992 21786 1048
rect 22650 2760 22706 2816
rect 23172 8730 23228 8732
rect 23252 8730 23308 8732
rect 23332 8730 23388 8732
rect 23412 8730 23468 8732
rect 23172 8678 23218 8730
rect 23218 8678 23228 8730
rect 23252 8678 23282 8730
rect 23282 8678 23294 8730
rect 23294 8678 23308 8730
rect 23332 8678 23346 8730
rect 23346 8678 23358 8730
rect 23358 8678 23388 8730
rect 23412 8678 23422 8730
rect 23422 8678 23468 8730
rect 23172 8676 23228 8678
rect 23252 8676 23308 8678
rect 23332 8676 23388 8678
rect 23412 8676 23468 8678
rect 23172 7642 23228 7644
rect 23252 7642 23308 7644
rect 23332 7642 23388 7644
rect 23412 7642 23468 7644
rect 23172 7590 23218 7642
rect 23218 7590 23228 7642
rect 23252 7590 23282 7642
rect 23282 7590 23294 7642
rect 23294 7590 23308 7642
rect 23332 7590 23346 7642
rect 23346 7590 23358 7642
rect 23358 7590 23388 7642
rect 23412 7590 23422 7642
rect 23422 7590 23468 7642
rect 23172 7588 23228 7590
rect 23252 7588 23308 7590
rect 23332 7588 23388 7590
rect 23412 7588 23468 7590
rect 23172 6554 23228 6556
rect 23252 6554 23308 6556
rect 23332 6554 23388 6556
rect 23412 6554 23468 6556
rect 23172 6502 23218 6554
rect 23218 6502 23228 6554
rect 23252 6502 23282 6554
rect 23282 6502 23294 6554
rect 23294 6502 23308 6554
rect 23332 6502 23346 6554
rect 23346 6502 23358 6554
rect 23358 6502 23388 6554
rect 23412 6502 23422 6554
rect 23422 6502 23468 6554
rect 23172 6500 23228 6502
rect 23252 6500 23308 6502
rect 23332 6500 23388 6502
rect 23412 6500 23468 6502
rect 23172 5466 23228 5468
rect 23252 5466 23308 5468
rect 23332 5466 23388 5468
rect 23412 5466 23468 5468
rect 23172 5414 23218 5466
rect 23218 5414 23228 5466
rect 23252 5414 23282 5466
rect 23282 5414 23294 5466
rect 23294 5414 23308 5466
rect 23332 5414 23346 5466
rect 23346 5414 23358 5466
rect 23358 5414 23388 5466
rect 23412 5414 23422 5466
rect 23422 5414 23468 5466
rect 23172 5412 23228 5414
rect 23252 5412 23308 5414
rect 23332 5412 23388 5414
rect 23412 5412 23468 5414
rect 23172 4378 23228 4380
rect 23252 4378 23308 4380
rect 23332 4378 23388 4380
rect 23412 4378 23468 4380
rect 23172 4326 23218 4378
rect 23218 4326 23228 4378
rect 23252 4326 23282 4378
rect 23282 4326 23294 4378
rect 23294 4326 23308 4378
rect 23332 4326 23346 4378
rect 23346 4326 23358 4378
rect 23358 4326 23388 4378
rect 23412 4326 23422 4378
rect 23422 4326 23468 4378
rect 23172 4324 23228 4326
rect 23252 4324 23308 4326
rect 23332 4324 23388 4326
rect 23412 4324 23468 4326
rect 23172 3290 23228 3292
rect 23252 3290 23308 3292
rect 23332 3290 23388 3292
rect 23412 3290 23468 3292
rect 23172 3238 23218 3290
rect 23218 3238 23228 3290
rect 23252 3238 23282 3290
rect 23282 3238 23294 3290
rect 23294 3238 23308 3290
rect 23332 3238 23346 3290
rect 23346 3238 23358 3290
rect 23358 3238 23388 3290
rect 23412 3238 23422 3290
rect 23422 3238 23468 3290
rect 23172 3236 23228 3238
rect 23252 3236 23308 3238
rect 23332 3236 23388 3238
rect 23412 3236 23468 3238
rect 34280 8730 34336 8732
rect 34360 8730 34416 8732
rect 34440 8730 34496 8732
rect 34520 8730 34576 8732
rect 34280 8678 34326 8730
rect 34326 8678 34336 8730
rect 34360 8678 34390 8730
rect 34390 8678 34402 8730
rect 34402 8678 34416 8730
rect 34440 8678 34454 8730
rect 34454 8678 34466 8730
rect 34466 8678 34496 8730
rect 34520 8678 34530 8730
rect 34530 8678 34576 8730
rect 34280 8676 34336 8678
rect 34360 8676 34416 8678
rect 34440 8676 34496 8678
rect 34520 8676 34576 8678
rect 45388 8730 45444 8732
rect 45468 8730 45524 8732
rect 45548 8730 45604 8732
rect 45628 8730 45684 8732
rect 45388 8678 45434 8730
rect 45434 8678 45444 8730
rect 45468 8678 45498 8730
rect 45498 8678 45510 8730
rect 45510 8678 45524 8730
rect 45548 8678 45562 8730
rect 45562 8678 45574 8730
rect 45574 8678 45604 8730
rect 45628 8678 45638 8730
rect 45638 8678 45684 8730
rect 45388 8676 45444 8678
rect 45468 8676 45524 8678
rect 45548 8676 45604 8678
rect 45628 8676 45684 8678
rect 24214 2624 24270 2680
rect 23172 2202 23228 2204
rect 23252 2202 23308 2204
rect 23332 2202 23388 2204
rect 23412 2202 23468 2204
rect 23172 2150 23218 2202
rect 23218 2150 23228 2202
rect 23252 2150 23282 2202
rect 23282 2150 23294 2202
rect 23294 2150 23308 2202
rect 23332 2150 23346 2202
rect 23346 2150 23358 2202
rect 23358 2150 23388 2202
rect 23412 2150 23422 2202
rect 23422 2150 23468 2202
rect 23172 2148 23228 2150
rect 23252 2148 23308 2150
rect 23332 2148 23388 2150
rect 23412 2148 23468 2150
rect 24858 4120 24914 4176
rect 23172 1114 23228 1116
rect 23252 1114 23308 1116
rect 23332 1114 23388 1116
rect 23412 1114 23468 1116
rect 23172 1062 23218 1114
rect 23218 1062 23228 1114
rect 23252 1062 23282 1114
rect 23282 1062 23294 1114
rect 23294 1062 23308 1114
rect 23332 1062 23346 1114
rect 23346 1062 23358 1114
rect 23358 1062 23388 1114
rect 23412 1062 23422 1114
rect 23422 1062 23468 1114
rect 23172 1060 23228 1062
rect 23252 1060 23308 1062
rect 23332 1060 23388 1062
rect 23412 1060 23468 1062
rect 24674 1536 24730 1592
rect 25778 2760 25834 2816
rect 26330 4528 26386 4584
rect 28726 8186 28782 8188
rect 28806 8186 28862 8188
rect 28886 8186 28942 8188
rect 28966 8186 29022 8188
rect 28726 8134 28772 8186
rect 28772 8134 28782 8186
rect 28806 8134 28836 8186
rect 28836 8134 28848 8186
rect 28848 8134 28862 8186
rect 28886 8134 28900 8186
rect 28900 8134 28912 8186
rect 28912 8134 28942 8186
rect 28966 8134 28976 8186
rect 28976 8134 29022 8186
rect 28726 8132 28782 8134
rect 28806 8132 28862 8134
rect 28886 8132 28942 8134
rect 28966 8132 29022 8134
rect 28726 7098 28782 7100
rect 28806 7098 28862 7100
rect 28886 7098 28942 7100
rect 28966 7098 29022 7100
rect 28726 7046 28772 7098
rect 28772 7046 28782 7098
rect 28806 7046 28836 7098
rect 28836 7046 28848 7098
rect 28848 7046 28862 7098
rect 28886 7046 28900 7098
rect 28900 7046 28912 7098
rect 28912 7046 28942 7098
rect 28966 7046 28976 7098
rect 28976 7046 29022 7098
rect 28726 7044 28782 7046
rect 28806 7044 28862 7046
rect 28886 7044 28942 7046
rect 28966 7044 29022 7046
rect 28726 6010 28782 6012
rect 28806 6010 28862 6012
rect 28886 6010 28942 6012
rect 28966 6010 29022 6012
rect 28726 5958 28772 6010
rect 28772 5958 28782 6010
rect 28806 5958 28836 6010
rect 28836 5958 28848 6010
rect 28848 5958 28862 6010
rect 28886 5958 28900 6010
rect 28900 5958 28912 6010
rect 28912 5958 28942 6010
rect 28966 5958 28976 6010
rect 28976 5958 29022 6010
rect 28726 5956 28782 5958
rect 28806 5956 28862 5958
rect 28886 5956 28942 5958
rect 28966 5956 29022 5958
rect 28726 4922 28782 4924
rect 28806 4922 28862 4924
rect 28886 4922 28942 4924
rect 28966 4922 29022 4924
rect 28726 4870 28772 4922
rect 28772 4870 28782 4922
rect 28806 4870 28836 4922
rect 28836 4870 28848 4922
rect 28848 4870 28862 4922
rect 28886 4870 28900 4922
rect 28900 4870 28912 4922
rect 28912 4870 28942 4922
rect 28966 4870 28976 4922
rect 28976 4870 29022 4922
rect 28726 4868 28782 4870
rect 28806 4868 28862 4870
rect 28886 4868 28942 4870
rect 28966 4868 29022 4870
rect 28726 3834 28782 3836
rect 28806 3834 28862 3836
rect 28886 3834 28942 3836
rect 28966 3834 29022 3836
rect 28726 3782 28772 3834
rect 28772 3782 28782 3834
rect 28806 3782 28836 3834
rect 28836 3782 28848 3834
rect 28848 3782 28862 3834
rect 28886 3782 28900 3834
rect 28900 3782 28912 3834
rect 28912 3782 28942 3834
rect 28966 3782 28976 3834
rect 28976 3782 29022 3834
rect 28726 3780 28782 3782
rect 28806 3780 28862 3782
rect 28886 3780 28942 3782
rect 28966 3780 29022 3782
rect 26330 992 26386 1048
rect 26330 584 26386 640
rect 28538 1672 28594 1728
rect 28726 2746 28782 2748
rect 28806 2746 28862 2748
rect 28886 2746 28942 2748
rect 28966 2746 29022 2748
rect 28726 2694 28772 2746
rect 28772 2694 28782 2746
rect 28806 2694 28836 2746
rect 28836 2694 28848 2746
rect 28848 2694 28862 2746
rect 28886 2694 28900 2746
rect 28900 2694 28912 2746
rect 28912 2694 28942 2746
rect 28966 2694 28976 2746
rect 28976 2694 29022 2746
rect 28726 2692 28782 2694
rect 28806 2692 28862 2694
rect 28886 2692 28942 2694
rect 28966 2692 29022 2694
rect 29274 2080 29330 2136
rect 28726 1658 28782 1660
rect 28806 1658 28862 1660
rect 28886 1658 28942 1660
rect 28966 1658 29022 1660
rect 28726 1606 28772 1658
rect 28772 1606 28782 1658
rect 28806 1606 28836 1658
rect 28836 1606 28848 1658
rect 28848 1606 28862 1658
rect 28886 1606 28900 1658
rect 28900 1606 28912 1658
rect 28912 1606 28942 1658
rect 28966 1606 28976 1658
rect 28976 1606 29022 1658
rect 28726 1604 28782 1606
rect 28806 1604 28862 1606
rect 28886 1604 28942 1606
rect 28966 1604 29022 1606
rect 29366 1128 29422 1184
rect 31390 2896 31446 2952
rect 30562 2252 30564 2272
rect 30564 2252 30616 2272
rect 30616 2252 30618 2272
rect 30562 2216 30618 2252
rect 30562 720 30618 776
rect 31206 1128 31262 1184
rect 31114 584 31170 640
rect 30930 312 30986 368
rect 34280 7642 34336 7644
rect 34360 7642 34416 7644
rect 34440 7642 34496 7644
rect 34520 7642 34576 7644
rect 34280 7590 34326 7642
rect 34326 7590 34336 7642
rect 34360 7590 34390 7642
rect 34390 7590 34402 7642
rect 34402 7590 34416 7642
rect 34440 7590 34454 7642
rect 34454 7590 34466 7642
rect 34466 7590 34496 7642
rect 34520 7590 34530 7642
rect 34530 7590 34576 7642
rect 34280 7588 34336 7590
rect 34360 7588 34416 7590
rect 34440 7588 34496 7590
rect 34520 7588 34576 7590
rect 34280 6554 34336 6556
rect 34360 6554 34416 6556
rect 34440 6554 34496 6556
rect 34520 6554 34576 6556
rect 34280 6502 34326 6554
rect 34326 6502 34336 6554
rect 34360 6502 34390 6554
rect 34390 6502 34402 6554
rect 34402 6502 34416 6554
rect 34440 6502 34454 6554
rect 34454 6502 34466 6554
rect 34466 6502 34496 6554
rect 34520 6502 34530 6554
rect 34530 6502 34576 6554
rect 34280 6500 34336 6502
rect 34360 6500 34416 6502
rect 34440 6500 34496 6502
rect 34520 6500 34576 6502
rect 34280 5466 34336 5468
rect 34360 5466 34416 5468
rect 34440 5466 34496 5468
rect 34520 5466 34576 5468
rect 34280 5414 34326 5466
rect 34326 5414 34336 5466
rect 34360 5414 34390 5466
rect 34390 5414 34402 5466
rect 34402 5414 34416 5466
rect 34440 5414 34454 5466
rect 34454 5414 34466 5466
rect 34466 5414 34496 5466
rect 34520 5414 34530 5466
rect 34530 5414 34576 5466
rect 34280 5412 34336 5414
rect 34360 5412 34416 5414
rect 34440 5412 34496 5414
rect 34520 5412 34576 5414
rect 34280 4378 34336 4380
rect 34360 4378 34416 4380
rect 34440 4378 34496 4380
rect 34520 4378 34576 4380
rect 34280 4326 34326 4378
rect 34326 4326 34336 4378
rect 34360 4326 34390 4378
rect 34390 4326 34402 4378
rect 34402 4326 34416 4378
rect 34440 4326 34454 4378
rect 34454 4326 34466 4378
rect 34466 4326 34496 4378
rect 34520 4326 34530 4378
rect 34530 4326 34576 4378
rect 34280 4324 34336 4326
rect 34360 4324 34416 4326
rect 34440 4324 34496 4326
rect 34520 4324 34576 4326
rect 34280 3290 34336 3292
rect 34360 3290 34416 3292
rect 34440 3290 34496 3292
rect 34520 3290 34576 3292
rect 34280 3238 34326 3290
rect 34326 3238 34336 3290
rect 34360 3238 34390 3290
rect 34390 3238 34402 3290
rect 34402 3238 34416 3290
rect 34440 3238 34454 3290
rect 34454 3238 34466 3290
rect 34466 3238 34496 3290
rect 34520 3238 34530 3290
rect 34530 3238 34576 3290
rect 34280 3236 34336 3238
rect 34360 3236 34416 3238
rect 34440 3236 34496 3238
rect 34520 3236 34576 3238
rect 32034 2252 32036 2272
rect 32036 2252 32088 2272
rect 32088 2252 32090 2272
rect 31482 2080 31538 2136
rect 32034 2216 32090 2252
rect 35162 3032 35218 3088
rect 34280 2202 34336 2204
rect 34360 2202 34416 2204
rect 34440 2202 34496 2204
rect 34520 2202 34576 2204
rect 34280 2150 34326 2202
rect 34326 2150 34336 2202
rect 34360 2150 34390 2202
rect 34390 2150 34402 2202
rect 34402 2150 34416 2202
rect 34440 2150 34454 2202
rect 34454 2150 34466 2202
rect 34466 2150 34496 2202
rect 34520 2150 34530 2202
rect 34530 2150 34576 2202
rect 34280 2148 34336 2150
rect 34360 2148 34416 2150
rect 34440 2148 34496 2150
rect 34520 2148 34576 2150
rect 34280 1114 34336 1116
rect 34360 1114 34416 1116
rect 34440 1114 34496 1116
rect 34520 1114 34576 1116
rect 34280 1062 34326 1114
rect 34326 1062 34336 1114
rect 34360 1062 34390 1114
rect 34390 1062 34402 1114
rect 34402 1062 34416 1114
rect 34440 1062 34454 1114
rect 34454 1062 34466 1114
rect 34466 1062 34496 1114
rect 34520 1062 34530 1114
rect 34530 1062 34576 1114
rect 34280 1060 34336 1062
rect 34360 1060 34416 1062
rect 34440 1060 34496 1062
rect 34520 1060 34576 1062
rect 34794 1284 34850 1320
rect 34794 1264 34796 1284
rect 34796 1264 34848 1284
rect 34848 1264 34850 1284
rect 37278 3984 37334 4040
rect 35438 2352 35494 2408
rect 37094 1400 37150 1456
rect 38106 3576 38162 3632
rect 37830 3440 37886 3496
rect 38014 1808 38070 1864
rect 39834 8186 39890 8188
rect 39914 8186 39970 8188
rect 39994 8186 40050 8188
rect 40074 8186 40130 8188
rect 39834 8134 39880 8186
rect 39880 8134 39890 8186
rect 39914 8134 39944 8186
rect 39944 8134 39956 8186
rect 39956 8134 39970 8186
rect 39994 8134 40008 8186
rect 40008 8134 40020 8186
rect 40020 8134 40050 8186
rect 40074 8134 40084 8186
rect 40084 8134 40130 8186
rect 39834 8132 39890 8134
rect 39914 8132 39970 8134
rect 39994 8132 40050 8134
rect 40074 8132 40130 8134
rect 39834 7098 39890 7100
rect 39914 7098 39970 7100
rect 39994 7098 40050 7100
rect 40074 7098 40130 7100
rect 39834 7046 39880 7098
rect 39880 7046 39890 7098
rect 39914 7046 39944 7098
rect 39944 7046 39956 7098
rect 39956 7046 39970 7098
rect 39994 7046 40008 7098
rect 40008 7046 40020 7098
rect 40020 7046 40050 7098
rect 40074 7046 40084 7098
rect 40084 7046 40130 7098
rect 39834 7044 39890 7046
rect 39914 7044 39970 7046
rect 39994 7044 40050 7046
rect 40074 7044 40130 7046
rect 39834 6010 39890 6012
rect 39914 6010 39970 6012
rect 39994 6010 40050 6012
rect 40074 6010 40130 6012
rect 39834 5958 39880 6010
rect 39880 5958 39890 6010
rect 39914 5958 39944 6010
rect 39944 5958 39956 6010
rect 39956 5958 39970 6010
rect 39994 5958 40008 6010
rect 40008 5958 40020 6010
rect 40020 5958 40050 6010
rect 40074 5958 40084 6010
rect 40084 5958 40130 6010
rect 39834 5956 39890 5958
rect 39914 5956 39970 5958
rect 39994 5956 40050 5958
rect 40074 5956 40130 5958
rect 39834 4922 39890 4924
rect 39914 4922 39970 4924
rect 39994 4922 40050 4924
rect 40074 4922 40130 4924
rect 39834 4870 39880 4922
rect 39880 4870 39890 4922
rect 39914 4870 39944 4922
rect 39944 4870 39956 4922
rect 39956 4870 39970 4922
rect 39994 4870 40008 4922
rect 40008 4870 40020 4922
rect 40020 4870 40050 4922
rect 40074 4870 40084 4922
rect 40084 4870 40130 4922
rect 39834 4868 39890 4870
rect 39914 4868 39970 4870
rect 39994 4868 40050 4870
rect 40074 4868 40130 4870
rect 39834 3834 39890 3836
rect 39914 3834 39970 3836
rect 39994 3834 40050 3836
rect 40074 3834 40130 3836
rect 39834 3782 39880 3834
rect 39880 3782 39890 3834
rect 39914 3782 39944 3834
rect 39944 3782 39956 3834
rect 39956 3782 39970 3834
rect 39994 3782 40008 3834
rect 40008 3782 40020 3834
rect 40020 3782 40050 3834
rect 40074 3782 40084 3834
rect 40084 3782 40130 3834
rect 39834 3780 39890 3782
rect 39914 3780 39970 3782
rect 39994 3780 40050 3782
rect 40074 3780 40130 3782
rect 38382 1964 38438 2000
rect 38382 1944 38384 1964
rect 38384 1944 38436 1964
rect 38436 1944 38438 1964
rect 39834 2746 39890 2748
rect 39914 2746 39970 2748
rect 39994 2746 40050 2748
rect 40074 2746 40130 2748
rect 39834 2694 39880 2746
rect 39880 2694 39890 2746
rect 39914 2694 39944 2746
rect 39944 2694 39956 2746
rect 39956 2694 39970 2746
rect 39994 2694 40008 2746
rect 40008 2694 40020 2746
rect 40020 2694 40050 2746
rect 40074 2694 40084 2746
rect 40084 2694 40130 2746
rect 39834 2692 39890 2694
rect 39914 2692 39970 2694
rect 39994 2692 40050 2694
rect 40074 2692 40130 2694
rect 40130 2488 40186 2544
rect 39834 1658 39890 1660
rect 39914 1658 39970 1660
rect 39994 1658 40050 1660
rect 40074 1658 40130 1660
rect 39834 1606 39880 1658
rect 39880 1606 39890 1658
rect 39914 1606 39944 1658
rect 39944 1606 39956 1658
rect 39956 1606 39970 1658
rect 39994 1606 40008 1658
rect 40008 1606 40020 1658
rect 40020 1606 40050 1658
rect 40074 1606 40084 1658
rect 40084 1606 40130 1658
rect 39834 1604 39890 1606
rect 39914 1604 39970 1606
rect 39994 1604 40050 1606
rect 40074 1604 40130 1606
rect 45388 7642 45444 7644
rect 45468 7642 45524 7644
rect 45548 7642 45604 7644
rect 45628 7642 45684 7644
rect 45388 7590 45434 7642
rect 45434 7590 45444 7642
rect 45468 7590 45498 7642
rect 45498 7590 45510 7642
rect 45510 7590 45524 7642
rect 45548 7590 45562 7642
rect 45562 7590 45574 7642
rect 45574 7590 45604 7642
rect 45628 7590 45638 7642
rect 45638 7590 45684 7642
rect 45388 7588 45444 7590
rect 45468 7588 45524 7590
rect 45548 7588 45604 7590
rect 45628 7588 45684 7590
rect 45388 6554 45444 6556
rect 45468 6554 45524 6556
rect 45548 6554 45604 6556
rect 45628 6554 45684 6556
rect 45388 6502 45434 6554
rect 45434 6502 45444 6554
rect 45468 6502 45498 6554
rect 45498 6502 45510 6554
rect 45510 6502 45524 6554
rect 45548 6502 45562 6554
rect 45562 6502 45574 6554
rect 45574 6502 45604 6554
rect 45628 6502 45638 6554
rect 45638 6502 45684 6554
rect 45388 6500 45444 6502
rect 45468 6500 45524 6502
rect 45548 6500 45604 6502
rect 45628 6500 45684 6502
rect 45388 5466 45444 5468
rect 45468 5466 45524 5468
rect 45548 5466 45604 5468
rect 45628 5466 45684 5468
rect 45388 5414 45434 5466
rect 45434 5414 45444 5466
rect 45468 5414 45498 5466
rect 45498 5414 45510 5466
rect 45510 5414 45524 5466
rect 45548 5414 45562 5466
rect 45562 5414 45574 5466
rect 45574 5414 45604 5466
rect 45628 5414 45638 5466
rect 45638 5414 45684 5466
rect 45388 5412 45444 5414
rect 45468 5412 45524 5414
rect 45548 5412 45604 5414
rect 45628 5412 45684 5414
rect 45388 4378 45444 4380
rect 45468 4378 45524 4380
rect 45548 4378 45604 4380
rect 45628 4378 45684 4380
rect 45388 4326 45434 4378
rect 45434 4326 45444 4378
rect 45468 4326 45498 4378
rect 45498 4326 45510 4378
rect 45510 4326 45524 4378
rect 45548 4326 45562 4378
rect 45562 4326 45574 4378
rect 45574 4326 45604 4378
rect 45628 4326 45638 4378
rect 45638 4326 45684 4378
rect 45388 4324 45444 4326
rect 45468 4324 45524 4326
rect 45548 4324 45604 4326
rect 45628 4324 45684 4326
rect 45388 3290 45444 3292
rect 45468 3290 45524 3292
rect 45548 3290 45604 3292
rect 45628 3290 45684 3292
rect 45388 3238 45434 3290
rect 45434 3238 45444 3290
rect 45468 3238 45498 3290
rect 45498 3238 45510 3290
rect 45510 3238 45524 3290
rect 45548 3238 45562 3290
rect 45562 3238 45574 3290
rect 45574 3238 45604 3290
rect 45628 3238 45638 3290
rect 45638 3238 45684 3290
rect 45388 3236 45444 3238
rect 45468 3236 45524 3238
rect 45548 3236 45604 3238
rect 45628 3236 45684 3238
rect 45388 2202 45444 2204
rect 45468 2202 45524 2204
rect 45548 2202 45604 2204
rect 45628 2202 45684 2204
rect 45388 2150 45434 2202
rect 45434 2150 45444 2202
rect 45468 2150 45498 2202
rect 45498 2150 45510 2202
rect 45510 2150 45524 2202
rect 45548 2150 45562 2202
rect 45562 2150 45574 2202
rect 45574 2150 45604 2202
rect 45628 2150 45638 2202
rect 45638 2150 45684 2202
rect 45388 2148 45444 2150
rect 45468 2148 45524 2150
rect 45548 2148 45604 2150
rect 45628 2148 45684 2150
rect 45388 1114 45444 1116
rect 45468 1114 45524 1116
rect 45548 1114 45604 1116
rect 45628 1114 45684 1116
rect 45388 1062 45434 1114
rect 45434 1062 45444 1114
rect 45468 1062 45498 1114
rect 45498 1062 45510 1114
rect 45510 1062 45524 1114
rect 45548 1062 45562 1114
rect 45562 1062 45574 1114
rect 45574 1062 45604 1114
rect 45628 1062 45638 1114
rect 45638 1062 45684 1114
rect 45388 1060 45444 1062
rect 45468 1060 45524 1062
rect 45548 1060 45604 1062
rect 45628 1060 45684 1062
<< metal3 >>
rect 12054 8736 12370 8737
rect 12054 8672 12060 8736
rect 12124 8672 12140 8736
rect 12204 8672 12220 8736
rect 12284 8672 12300 8736
rect 12364 8672 12370 8736
rect 12054 8671 12370 8672
rect 23162 8736 23478 8737
rect 23162 8672 23168 8736
rect 23232 8672 23248 8736
rect 23312 8672 23328 8736
rect 23392 8672 23408 8736
rect 23472 8672 23478 8736
rect 23162 8671 23478 8672
rect 34270 8736 34586 8737
rect 34270 8672 34276 8736
rect 34340 8672 34356 8736
rect 34420 8672 34436 8736
rect 34500 8672 34516 8736
rect 34580 8672 34586 8736
rect 34270 8671 34586 8672
rect 45378 8736 45694 8737
rect 45378 8672 45384 8736
rect 45448 8672 45464 8736
rect 45528 8672 45544 8736
rect 45608 8672 45624 8736
rect 45688 8672 45694 8736
rect 45378 8671 45694 8672
rect 6500 8192 6816 8193
rect 6500 8128 6506 8192
rect 6570 8128 6586 8192
rect 6650 8128 6666 8192
rect 6730 8128 6746 8192
rect 6810 8128 6816 8192
rect 6500 8127 6816 8128
rect 17608 8192 17924 8193
rect 17608 8128 17614 8192
rect 17678 8128 17694 8192
rect 17758 8128 17774 8192
rect 17838 8128 17854 8192
rect 17918 8128 17924 8192
rect 17608 8127 17924 8128
rect 28716 8192 29032 8193
rect 28716 8128 28722 8192
rect 28786 8128 28802 8192
rect 28866 8128 28882 8192
rect 28946 8128 28962 8192
rect 29026 8128 29032 8192
rect 28716 8127 29032 8128
rect 39824 8192 40140 8193
rect 39824 8128 39830 8192
rect 39894 8128 39910 8192
rect 39974 8128 39990 8192
rect 40054 8128 40070 8192
rect 40134 8128 40140 8192
rect 39824 8127 40140 8128
rect 12054 7648 12370 7649
rect 12054 7584 12060 7648
rect 12124 7584 12140 7648
rect 12204 7584 12220 7648
rect 12284 7584 12300 7648
rect 12364 7584 12370 7648
rect 12054 7583 12370 7584
rect 23162 7648 23478 7649
rect 23162 7584 23168 7648
rect 23232 7584 23248 7648
rect 23312 7584 23328 7648
rect 23392 7584 23408 7648
rect 23472 7584 23478 7648
rect 23162 7583 23478 7584
rect 34270 7648 34586 7649
rect 34270 7584 34276 7648
rect 34340 7584 34356 7648
rect 34420 7584 34436 7648
rect 34500 7584 34516 7648
rect 34580 7584 34586 7648
rect 34270 7583 34586 7584
rect 45378 7648 45694 7649
rect 45378 7584 45384 7648
rect 45448 7584 45464 7648
rect 45528 7584 45544 7648
rect 45608 7584 45624 7648
rect 45688 7584 45694 7648
rect 45378 7583 45694 7584
rect 6500 7104 6816 7105
rect 6500 7040 6506 7104
rect 6570 7040 6586 7104
rect 6650 7040 6666 7104
rect 6730 7040 6746 7104
rect 6810 7040 6816 7104
rect 6500 7039 6816 7040
rect 17608 7104 17924 7105
rect 17608 7040 17614 7104
rect 17678 7040 17694 7104
rect 17758 7040 17774 7104
rect 17838 7040 17854 7104
rect 17918 7040 17924 7104
rect 17608 7039 17924 7040
rect 28716 7104 29032 7105
rect 28716 7040 28722 7104
rect 28786 7040 28802 7104
rect 28866 7040 28882 7104
rect 28946 7040 28962 7104
rect 29026 7040 29032 7104
rect 28716 7039 29032 7040
rect 39824 7104 40140 7105
rect 39824 7040 39830 7104
rect 39894 7040 39910 7104
rect 39974 7040 39990 7104
rect 40054 7040 40070 7104
rect 40134 7040 40140 7104
rect 39824 7039 40140 7040
rect 12054 6560 12370 6561
rect 12054 6496 12060 6560
rect 12124 6496 12140 6560
rect 12204 6496 12220 6560
rect 12284 6496 12300 6560
rect 12364 6496 12370 6560
rect 12054 6495 12370 6496
rect 23162 6560 23478 6561
rect 23162 6496 23168 6560
rect 23232 6496 23248 6560
rect 23312 6496 23328 6560
rect 23392 6496 23408 6560
rect 23472 6496 23478 6560
rect 23162 6495 23478 6496
rect 34270 6560 34586 6561
rect 34270 6496 34276 6560
rect 34340 6496 34356 6560
rect 34420 6496 34436 6560
rect 34500 6496 34516 6560
rect 34580 6496 34586 6560
rect 34270 6495 34586 6496
rect 45378 6560 45694 6561
rect 45378 6496 45384 6560
rect 45448 6496 45464 6560
rect 45528 6496 45544 6560
rect 45608 6496 45624 6560
rect 45688 6496 45694 6560
rect 45378 6495 45694 6496
rect 6500 6016 6816 6017
rect 6500 5952 6506 6016
rect 6570 5952 6586 6016
rect 6650 5952 6666 6016
rect 6730 5952 6746 6016
rect 6810 5952 6816 6016
rect 6500 5951 6816 5952
rect 17608 6016 17924 6017
rect 17608 5952 17614 6016
rect 17678 5952 17694 6016
rect 17758 5952 17774 6016
rect 17838 5952 17854 6016
rect 17918 5952 17924 6016
rect 17608 5951 17924 5952
rect 28716 6016 29032 6017
rect 28716 5952 28722 6016
rect 28786 5952 28802 6016
rect 28866 5952 28882 6016
rect 28946 5952 28962 6016
rect 29026 5952 29032 6016
rect 28716 5951 29032 5952
rect 39824 6016 40140 6017
rect 39824 5952 39830 6016
rect 39894 5952 39910 6016
rect 39974 5952 39990 6016
rect 40054 5952 40070 6016
rect 40134 5952 40140 6016
rect 39824 5951 40140 5952
rect 12054 5472 12370 5473
rect 12054 5408 12060 5472
rect 12124 5408 12140 5472
rect 12204 5408 12220 5472
rect 12284 5408 12300 5472
rect 12364 5408 12370 5472
rect 12054 5407 12370 5408
rect 23162 5472 23478 5473
rect 23162 5408 23168 5472
rect 23232 5408 23248 5472
rect 23312 5408 23328 5472
rect 23392 5408 23408 5472
rect 23472 5408 23478 5472
rect 23162 5407 23478 5408
rect 34270 5472 34586 5473
rect 34270 5408 34276 5472
rect 34340 5408 34356 5472
rect 34420 5408 34436 5472
rect 34500 5408 34516 5472
rect 34580 5408 34586 5472
rect 34270 5407 34586 5408
rect 45378 5472 45694 5473
rect 45378 5408 45384 5472
rect 45448 5408 45464 5472
rect 45528 5408 45544 5472
rect 45608 5408 45624 5472
rect 45688 5408 45694 5472
rect 45378 5407 45694 5408
rect 6500 4928 6816 4929
rect 6500 4864 6506 4928
rect 6570 4864 6586 4928
rect 6650 4864 6666 4928
rect 6730 4864 6746 4928
rect 6810 4864 6816 4928
rect 6500 4863 6816 4864
rect 17608 4928 17924 4929
rect 17608 4864 17614 4928
rect 17678 4864 17694 4928
rect 17758 4864 17774 4928
rect 17838 4864 17854 4928
rect 17918 4864 17924 4928
rect 17608 4863 17924 4864
rect 28716 4928 29032 4929
rect 28716 4864 28722 4928
rect 28786 4864 28802 4928
rect 28866 4864 28882 4928
rect 28946 4864 28962 4928
rect 29026 4864 29032 4928
rect 28716 4863 29032 4864
rect 39824 4928 40140 4929
rect 39824 4864 39830 4928
rect 39894 4864 39910 4928
rect 39974 4864 39990 4928
rect 40054 4864 40070 4928
rect 40134 4864 40140 4928
rect 39824 4863 40140 4864
rect 4705 4586 4771 4589
rect 26325 4586 26391 4589
rect 4705 4584 26391 4586
rect 4705 4528 4710 4584
rect 4766 4528 26330 4584
rect 26386 4528 26391 4584
rect 4705 4526 26391 4528
rect 4705 4523 4771 4526
rect 26325 4523 26391 4526
rect 12054 4384 12370 4385
rect 12054 4320 12060 4384
rect 12124 4320 12140 4384
rect 12204 4320 12220 4384
rect 12284 4320 12300 4384
rect 12364 4320 12370 4384
rect 12054 4319 12370 4320
rect 23162 4384 23478 4385
rect 23162 4320 23168 4384
rect 23232 4320 23248 4384
rect 23312 4320 23328 4384
rect 23392 4320 23408 4384
rect 23472 4320 23478 4384
rect 23162 4319 23478 4320
rect 34270 4384 34586 4385
rect 34270 4320 34276 4384
rect 34340 4320 34356 4384
rect 34420 4320 34436 4384
rect 34500 4320 34516 4384
rect 34580 4320 34586 4384
rect 34270 4319 34586 4320
rect 45378 4384 45694 4385
rect 45378 4320 45384 4384
rect 45448 4320 45464 4384
rect 45528 4320 45544 4384
rect 45608 4320 45624 4384
rect 45688 4320 45694 4384
rect 45378 4319 45694 4320
rect 3785 4178 3851 4181
rect 24853 4178 24919 4181
rect 3785 4176 24919 4178
rect 3785 4120 3790 4176
rect 3846 4120 24858 4176
rect 24914 4120 24919 4176
rect 3785 4118 24919 4120
rect 3785 4115 3851 4118
rect 24853 4115 24919 4118
rect 11881 4042 11947 4045
rect 22553 4042 22619 4045
rect 37273 4042 37339 4045
rect 11881 4040 22619 4042
rect 11881 3984 11886 4040
rect 11942 3984 22558 4040
rect 22614 3984 22619 4040
rect 11881 3982 22619 3984
rect 11881 3979 11947 3982
rect 22553 3979 22619 3982
rect 26190 4040 37339 4042
rect 26190 3984 37278 4040
rect 37334 3984 37339 4040
rect 26190 3982 37339 3984
rect 20529 3906 20595 3909
rect 26190 3906 26250 3982
rect 37273 3979 37339 3982
rect 20529 3904 26250 3906
rect 20529 3848 20534 3904
rect 20590 3848 26250 3904
rect 20529 3846 26250 3848
rect 20529 3843 20595 3846
rect 6500 3840 6816 3841
rect 6500 3776 6506 3840
rect 6570 3776 6586 3840
rect 6650 3776 6666 3840
rect 6730 3776 6746 3840
rect 6810 3776 6816 3840
rect 6500 3775 6816 3776
rect 17608 3840 17924 3841
rect 17608 3776 17614 3840
rect 17678 3776 17694 3840
rect 17758 3776 17774 3840
rect 17838 3776 17854 3840
rect 17918 3776 17924 3840
rect 17608 3775 17924 3776
rect 28716 3840 29032 3841
rect 28716 3776 28722 3840
rect 28786 3776 28802 3840
rect 28866 3776 28882 3840
rect 28946 3776 28962 3840
rect 29026 3776 29032 3840
rect 28716 3775 29032 3776
rect 39824 3840 40140 3841
rect 39824 3776 39830 3840
rect 39894 3776 39910 3840
rect 39974 3776 39990 3840
rect 40054 3776 40070 3840
rect 40134 3776 40140 3840
rect 39824 3775 40140 3776
rect 15929 3634 15995 3637
rect 38101 3634 38167 3637
rect 15929 3632 38167 3634
rect 15929 3576 15934 3632
rect 15990 3576 38106 3632
rect 38162 3576 38167 3632
rect 15929 3574 38167 3576
rect 15929 3571 15995 3574
rect 38101 3571 38167 3574
rect 18689 3498 18755 3501
rect 37825 3498 37891 3501
rect 18689 3496 37891 3498
rect 18689 3440 18694 3496
rect 18750 3440 37830 3496
rect 37886 3440 37891 3496
rect 18689 3438 37891 3440
rect 18689 3435 18755 3438
rect 37825 3435 37891 3438
rect 12054 3296 12370 3297
rect 12054 3232 12060 3296
rect 12124 3232 12140 3296
rect 12204 3232 12220 3296
rect 12284 3232 12300 3296
rect 12364 3232 12370 3296
rect 12054 3231 12370 3232
rect 23162 3296 23478 3297
rect 23162 3232 23168 3296
rect 23232 3232 23248 3296
rect 23312 3232 23328 3296
rect 23392 3232 23408 3296
rect 23472 3232 23478 3296
rect 23162 3231 23478 3232
rect 34270 3296 34586 3297
rect 34270 3232 34276 3296
rect 34340 3232 34356 3296
rect 34420 3232 34436 3296
rect 34500 3232 34516 3296
rect 34580 3232 34586 3296
rect 34270 3231 34586 3232
rect 45378 3296 45694 3297
rect 45378 3232 45384 3296
rect 45448 3232 45464 3296
rect 45528 3232 45544 3296
rect 45608 3232 45624 3296
rect 45688 3232 45694 3296
rect 45378 3231 45694 3232
rect 13353 3226 13419 3229
rect 22093 3226 22159 3229
rect 13353 3224 22159 3226
rect 13353 3168 13358 3224
rect 13414 3168 22098 3224
rect 22154 3168 22159 3224
rect 13353 3166 22159 3168
rect 13353 3163 13419 3166
rect 22093 3163 22159 3166
rect 17125 3090 17191 3093
rect 35157 3090 35223 3093
rect 17125 3088 35223 3090
rect 17125 3032 17130 3088
rect 17186 3032 35162 3088
rect 35218 3032 35223 3088
rect 17125 3030 35223 3032
rect 17125 3027 17191 3030
rect 35157 3027 35223 3030
rect 17309 2954 17375 2957
rect 31385 2954 31451 2957
rect 17309 2952 31451 2954
rect 17309 2896 17314 2952
rect 17370 2896 31390 2952
rect 31446 2896 31451 2952
rect 17309 2894 31451 2896
rect 17309 2891 17375 2894
rect 31385 2891 31451 2894
rect 22645 2818 22711 2821
rect 25773 2818 25839 2821
rect 22645 2816 25839 2818
rect 22645 2760 22650 2816
rect 22706 2760 25778 2816
rect 25834 2760 25839 2816
rect 22645 2758 25839 2760
rect 22645 2755 22711 2758
rect 25773 2755 25839 2758
rect 6500 2752 6816 2753
rect 6500 2688 6506 2752
rect 6570 2688 6586 2752
rect 6650 2688 6666 2752
rect 6730 2688 6746 2752
rect 6810 2688 6816 2752
rect 6500 2687 6816 2688
rect 17608 2752 17924 2753
rect 17608 2688 17614 2752
rect 17678 2688 17694 2752
rect 17758 2688 17774 2752
rect 17838 2688 17854 2752
rect 17918 2688 17924 2752
rect 17608 2687 17924 2688
rect 28716 2752 29032 2753
rect 28716 2688 28722 2752
rect 28786 2688 28802 2752
rect 28866 2688 28882 2752
rect 28946 2688 28962 2752
rect 29026 2688 29032 2752
rect 28716 2687 29032 2688
rect 39824 2752 40140 2753
rect 39824 2688 39830 2752
rect 39894 2688 39910 2752
rect 39974 2688 39990 2752
rect 40054 2688 40070 2752
rect 40134 2688 40140 2752
rect 39824 2687 40140 2688
rect 18045 2682 18111 2685
rect 19885 2682 19951 2685
rect 18045 2680 19951 2682
rect 18045 2624 18050 2680
rect 18106 2624 19890 2680
rect 19946 2624 19951 2680
rect 18045 2622 19951 2624
rect 18045 2619 18111 2622
rect 19885 2619 19951 2622
rect 22001 2682 22067 2685
rect 24209 2682 24275 2685
rect 22001 2680 24275 2682
rect 22001 2624 22006 2680
rect 22062 2624 24214 2680
rect 24270 2624 24275 2680
rect 22001 2622 24275 2624
rect 22001 2619 22067 2622
rect 24209 2619 24275 2622
rect 1853 2546 1919 2549
rect 18781 2546 18847 2549
rect 1853 2544 18847 2546
rect 1853 2488 1858 2544
rect 1914 2488 18786 2544
rect 18842 2488 18847 2544
rect 1853 2486 18847 2488
rect 1853 2483 1919 2486
rect 18781 2483 18847 2486
rect 21541 2546 21607 2549
rect 40125 2546 40191 2549
rect 21541 2544 40191 2546
rect 21541 2488 21546 2544
rect 21602 2488 40130 2544
rect 40186 2488 40191 2544
rect 21541 2486 40191 2488
rect 21541 2483 21607 2486
rect 40125 2483 40191 2486
rect 9949 2410 10015 2413
rect 20713 2410 20779 2413
rect 9949 2408 20779 2410
rect 9949 2352 9954 2408
rect 10010 2352 20718 2408
rect 20774 2352 20779 2408
rect 9949 2350 20779 2352
rect 9949 2347 10015 2350
rect 20713 2347 20779 2350
rect 22185 2410 22251 2413
rect 35433 2410 35499 2413
rect 22185 2408 35499 2410
rect 22185 2352 22190 2408
rect 22246 2352 35438 2408
rect 35494 2352 35499 2408
rect 22185 2350 35499 2352
rect 22185 2347 22251 2350
rect 35433 2347 35499 2350
rect 16481 2274 16547 2277
rect 20621 2274 20687 2277
rect 16481 2272 20687 2274
rect 16481 2216 16486 2272
rect 16542 2216 20626 2272
rect 20682 2216 20687 2272
rect 16481 2214 20687 2216
rect 16481 2211 16547 2214
rect 20621 2211 20687 2214
rect 30557 2274 30623 2277
rect 32029 2274 32095 2277
rect 30557 2272 32095 2274
rect 30557 2216 30562 2272
rect 30618 2216 32034 2272
rect 32090 2216 32095 2272
rect 30557 2214 32095 2216
rect 30557 2211 30623 2214
rect 32029 2211 32095 2214
rect 12054 2208 12370 2209
rect 12054 2144 12060 2208
rect 12124 2144 12140 2208
rect 12204 2144 12220 2208
rect 12284 2144 12300 2208
rect 12364 2144 12370 2208
rect 12054 2143 12370 2144
rect 23162 2208 23478 2209
rect 23162 2144 23168 2208
rect 23232 2144 23248 2208
rect 23312 2144 23328 2208
rect 23392 2144 23408 2208
rect 23472 2144 23478 2208
rect 23162 2143 23478 2144
rect 34270 2208 34586 2209
rect 34270 2144 34276 2208
rect 34340 2144 34356 2208
rect 34420 2144 34436 2208
rect 34500 2144 34516 2208
rect 34580 2144 34586 2208
rect 34270 2143 34586 2144
rect 45378 2208 45694 2209
rect 45378 2144 45384 2208
rect 45448 2144 45464 2208
rect 45528 2144 45544 2208
rect 45608 2144 45624 2208
rect 45688 2144 45694 2208
rect 45378 2143 45694 2144
rect 21449 2138 21515 2141
rect 17128 2136 21515 2138
rect 17128 2080 21454 2136
rect 21510 2080 21515 2136
rect 17128 2078 21515 2080
rect 8937 2002 9003 2005
rect 17128 2002 17188 2078
rect 21449 2075 21515 2078
rect 29269 2138 29335 2141
rect 31477 2138 31543 2141
rect 29269 2136 31543 2138
rect 29269 2080 29274 2136
rect 29330 2080 31482 2136
rect 31538 2080 31543 2136
rect 29269 2078 31543 2080
rect 29269 2075 29335 2078
rect 31477 2075 31543 2078
rect 8937 2000 17188 2002
rect 8937 1944 8942 2000
rect 8998 1944 17188 2000
rect 8937 1942 17188 1944
rect 19241 2002 19307 2005
rect 38377 2002 38443 2005
rect 19241 2000 38443 2002
rect 19241 1944 19246 2000
rect 19302 1944 38382 2000
rect 38438 1944 38443 2000
rect 19241 1942 38443 1944
rect 8937 1939 9003 1942
rect 19241 1939 19307 1942
rect 38377 1939 38443 1942
rect 15193 1866 15259 1869
rect 38009 1866 38075 1869
rect 15193 1864 38075 1866
rect 15193 1808 15198 1864
rect 15254 1808 38014 1864
rect 38070 1808 38075 1864
rect 15193 1806 38075 1808
rect 15193 1803 15259 1806
rect 38009 1803 38075 1806
rect 19701 1730 19767 1733
rect 28533 1730 28599 1733
rect 19701 1728 28599 1730
rect 19701 1672 19706 1728
rect 19762 1672 28538 1728
rect 28594 1672 28599 1728
rect 19701 1670 28599 1672
rect 19701 1667 19767 1670
rect 28533 1667 28599 1670
rect 6500 1664 6816 1665
rect 6500 1600 6506 1664
rect 6570 1600 6586 1664
rect 6650 1600 6666 1664
rect 6730 1600 6746 1664
rect 6810 1600 6816 1664
rect 6500 1599 6816 1600
rect 17608 1664 17924 1665
rect 17608 1600 17614 1664
rect 17678 1600 17694 1664
rect 17758 1600 17774 1664
rect 17838 1600 17854 1664
rect 17918 1600 17924 1664
rect 17608 1599 17924 1600
rect 28716 1664 29032 1665
rect 28716 1600 28722 1664
rect 28786 1600 28802 1664
rect 28866 1600 28882 1664
rect 28946 1600 28962 1664
rect 29026 1600 29032 1664
rect 28716 1599 29032 1600
rect 39824 1664 40140 1665
rect 39824 1600 39830 1664
rect 39894 1600 39910 1664
rect 39974 1600 39990 1664
rect 40054 1600 40070 1664
rect 40134 1600 40140 1664
rect 39824 1599 40140 1600
rect 24669 1594 24735 1597
rect 18094 1592 24735 1594
rect 18094 1536 24674 1592
rect 24730 1536 24735 1592
rect 18094 1534 24735 1536
rect 14825 1458 14891 1461
rect 18094 1458 18154 1534
rect 24669 1531 24735 1534
rect 14825 1456 18154 1458
rect 14825 1400 14830 1456
rect 14886 1400 18154 1456
rect 14825 1398 18154 1400
rect 20345 1458 20411 1461
rect 37089 1458 37155 1461
rect 20345 1456 37155 1458
rect 20345 1400 20350 1456
rect 20406 1400 37094 1456
rect 37150 1400 37155 1456
rect 20345 1398 37155 1400
rect 14825 1395 14891 1398
rect 20345 1395 20411 1398
rect 37089 1395 37155 1398
rect 11697 1322 11763 1325
rect 18873 1322 18939 1325
rect 34789 1322 34855 1325
rect 11697 1320 18939 1322
rect 11697 1264 11702 1320
rect 11758 1264 18878 1320
rect 18934 1264 18939 1320
rect 11697 1262 18939 1264
rect 11697 1259 11763 1262
rect 18873 1259 18939 1262
rect 22050 1320 34855 1322
rect 22050 1264 34794 1320
rect 34850 1264 34855 1320
rect 22050 1262 34855 1264
rect 12801 1186 12867 1189
rect 17861 1186 17927 1189
rect 12801 1184 17927 1186
rect 12801 1128 12806 1184
rect 12862 1128 17866 1184
rect 17922 1128 17927 1184
rect 12801 1126 17927 1128
rect 12801 1123 12867 1126
rect 17861 1123 17927 1126
rect 18045 1186 18111 1189
rect 22050 1186 22110 1262
rect 34789 1259 34855 1262
rect 29361 1186 29427 1189
rect 31201 1186 31267 1189
rect 18045 1184 22110 1186
rect 18045 1128 18050 1184
rect 18106 1128 22110 1184
rect 18045 1126 22110 1128
rect 25638 1184 29427 1186
rect 25638 1128 29366 1184
rect 29422 1128 29427 1184
rect 25638 1126 29427 1128
rect 18045 1123 18111 1126
rect 12054 1120 12370 1121
rect 12054 1056 12060 1120
rect 12124 1056 12140 1120
rect 12204 1056 12220 1120
rect 12284 1056 12300 1120
rect 12364 1056 12370 1120
rect 12054 1055 12370 1056
rect 23162 1120 23478 1121
rect 23162 1056 23168 1120
rect 23232 1056 23248 1120
rect 23312 1056 23328 1120
rect 23392 1056 23408 1120
rect 23472 1056 23478 1120
rect 23162 1055 23478 1056
rect 12709 1050 12775 1053
rect 21725 1050 21791 1053
rect 12709 1048 21791 1050
rect 12709 992 12714 1048
rect 12770 992 21730 1048
rect 21786 992 21791 1048
rect 12709 990 21791 992
rect 12709 987 12775 990
rect 21725 987 21791 990
rect 8753 914 8819 917
rect 25638 914 25698 1126
rect 29361 1123 29427 1126
rect 29502 1184 31267 1186
rect 29502 1128 31206 1184
rect 31262 1128 31267 1184
rect 29502 1126 31267 1128
rect 26325 1050 26391 1053
rect 29502 1050 29562 1126
rect 31201 1123 31267 1126
rect 34270 1120 34586 1121
rect 34270 1056 34276 1120
rect 34340 1056 34356 1120
rect 34420 1056 34436 1120
rect 34500 1056 34516 1120
rect 34580 1056 34586 1120
rect 34270 1055 34586 1056
rect 45378 1120 45694 1121
rect 45378 1056 45384 1120
rect 45448 1056 45464 1120
rect 45528 1056 45544 1120
rect 45608 1056 45624 1120
rect 45688 1056 45694 1120
rect 45378 1055 45694 1056
rect 26325 1048 29562 1050
rect 26325 992 26330 1048
rect 26386 992 29562 1048
rect 26325 990 29562 992
rect 26325 987 26391 990
rect 8753 912 25698 914
rect 8753 856 8758 912
rect 8814 856 25698 912
rect 8753 854 25698 856
rect 8753 851 8819 854
rect 10685 778 10751 781
rect 30557 778 30623 781
rect 10685 776 30623 778
rect 10685 720 10690 776
rect 10746 720 30562 776
rect 30618 720 30623 776
rect 10685 718 30623 720
rect 10685 715 10751 718
rect 30557 715 30623 718
rect 9213 642 9279 645
rect 26325 642 26391 645
rect 31109 642 31175 645
rect 9213 640 26391 642
rect 9213 584 9218 640
rect 9274 584 26330 640
rect 26386 584 26391 640
rect 9213 582 26391 584
rect 9213 579 9279 582
rect 26325 579 26391 582
rect 26558 640 31175 642
rect 26558 584 31114 640
rect 31170 584 31175 640
rect 26558 582 31175 584
rect 9581 506 9647 509
rect 26558 506 26618 582
rect 31109 579 31175 582
rect 9581 504 26618 506
rect 9581 448 9586 504
rect 9642 448 26618 504
rect 9581 446 26618 448
rect 9581 443 9647 446
rect 10317 370 10383 373
rect 30925 370 30991 373
rect 10317 368 30991 370
rect 10317 312 10322 368
rect 10378 312 30930 368
rect 30986 312 30991 368
rect 10317 310 30991 312
rect 10317 307 10383 310
rect 30925 307 30991 310
<< via3 >>
rect 12060 8732 12124 8736
rect 12060 8676 12064 8732
rect 12064 8676 12120 8732
rect 12120 8676 12124 8732
rect 12060 8672 12124 8676
rect 12140 8732 12204 8736
rect 12140 8676 12144 8732
rect 12144 8676 12200 8732
rect 12200 8676 12204 8732
rect 12140 8672 12204 8676
rect 12220 8732 12284 8736
rect 12220 8676 12224 8732
rect 12224 8676 12280 8732
rect 12280 8676 12284 8732
rect 12220 8672 12284 8676
rect 12300 8732 12364 8736
rect 12300 8676 12304 8732
rect 12304 8676 12360 8732
rect 12360 8676 12364 8732
rect 12300 8672 12364 8676
rect 23168 8732 23232 8736
rect 23168 8676 23172 8732
rect 23172 8676 23228 8732
rect 23228 8676 23232 8732
rect 23168 8672 23232 8676
rect 23248 8732 23312 8736
rect 23248 8676 23252 8732
rect 23252 8676 23308 8732
rect 23308 8676 23312 8732
rect 23248 8672 23312 8676
rect 23328 8732 23392 8736
rect 23328 8676 23332 8732
rect 23332 8676 23388 8732
rect 23388 8676 23392 8732
rect 23328 8672 23392 8676
rect 23408 8732 23472 8736
rect 23408 8676 23412 8732
rect 23412 8676 23468 8732
rect 23468 8676 23472 8732
rect 23408 8672 23472 8676
rect 34276 8732 34340 8736
rect 34276 8676 34280 8732
rect 34280 8676 34336 8732
rect 34336 8676 34340 8732
rect 34276 8672 34340 8676
rect 34356 8732 34420 8736
rect 34356 8676 34360 8732
rect 34360 8676 34416 8732
rect 34416 8676 34420 8732
rect 34356 8672 34420 8676
rect 34436 8732 34500 8736
rect 34436 8676 34440 8732
rect 34440 8676 34496 8732
rect 34496 8676 34500 8732
rect 34436 8672 34500 8676
rect 34516 8732 34580 8736
rect 34516 8676 34520 8732
rect 34520 8676 34576 8732
rect 34576 8676 34580 8732
rect 34516 8672 34580 8676
rect 45384 8732 45448 8736
rect 45384 8676 45388 8732
rect 45388 8676 45444 8732
rect 45444 8676 45448 8732
rect 45384 8672 45448 8676
rect 45464 8732 45528 8736
rect 45464 8676 45468 8732
rect 45468 8676 45524 8732
rect 45524 8676 45528 8732
rect 45464 8672 45528 8676
rect 45544 8732 45608 8736
rect 45544 8676 45548 8732
rect 45548 8676 45604 8732
rect 45604 8676 45608 8732
rect 45544 8672 45608 8676
rect 45624 8732 45688 8736
rect 45624 8676 45628 8732
rect 45628 8676 45684 8732
rect 45684 8676 45688 8732
rect 45624 8672 45688 8676
rect 6506 8188 6570 8192
rect 6506 8132 6510 8188
rect 6510 8132 6566 8188
rect 6566 8132 6570 8188
rect 6506 8128 6570 8132
rect 6586 8188 6650 8192
rect 6586 8132 6590 8188
rect 6590 8132 6646 8188
rect 6646 8132 6650 8188
rect 6586 8128 6650 8132
rect 6666 8188 6730 8192
rect 6666 8132 6670 8188
rect 6670 8132 6726 8188
rect 6726 8132 6730 8188
rect 6666 8128 6730 8132
rect 6746 8188 6810 8192
rect 6746 8132 6750 8188
rect 6750 8132 6806 8188
rect 6806 8132 6810 8188
rect 6746 8128 6810 8132
rect 17614 8188 17678 8192
rect 17614 8132 17618 8188
rect 17618 8132 17674 8188
rect 17674 8132 17678 8188
rect 17614 8128 17678 8132
rect 17694 8188 17758 8192
rect 17694 8132 17698 8188
rect 17698 8132 17754 8188
rect 17754 8132 17758 8188
rect 17694 8128 17758 8132
rect 17774 8188 17838 8192
rect 17774 8132 17778 8188
rect 17778 8132 17834 8188
rect 17834 8132 17838 8188
rect 17774 8128 17838 8132
rect 17854 8188 17918 8192
rect 17854 8132 17858 8188
rect 17858 8132 17914 8188
rect 17914 8132 17918 8188
rect 17854 8128 17918 8132
rect 28722 8188 28786 8192
rect 28722 8132 28726 8188
rect 28726 8132 28782 8188
rect 28782 8132 28786 8188
rect 28722 8128 28786 8132
rect 28802 8188 28866 8192
rect 28802 8132 28806 8188
rect 28806 8132 28862 8188
rect 28862 8132 28866 8188
rect 28802 8128 28866 8132
rect 28882 8188 28946 8192
rect 28882 8132 28886 8188
rect 28886 8132 28942 8188
rect 28942 8132 28946 8188
rect 28882 8128 28946 8132
rect 28962 8188 29026 8192
rect 28962 8132 28966 8188
rect 28966 8132 29022 8188
rect 29022 8132 29026 8188
rect 28962 8128 29026 8132
rect 39830 8188 39894 8192
rect 39830 8132 39834 8188
rect 39834 8132 39890 8188
rect 39890 8132 39894 8188
rect 39830 8128 39894 8132
rect 39910 8188 39974 8192
rect 39910 8132 39914 8188
rect 39914 8132 39970 8188
rect 39970 8132 39974 8188
rect 39910 8128 39974 8132
rect 39990 8188 40054 8192
rect 39990 8132 39994 8188
rect 39994 8132 40050 8188
rect 40050 8132 40054 8188
rect 39990 8128 40054 8132
rect 40070 8188 40134 8192
rect 40070 8132 40074 8188
rect 40074 8132 40130 8188
rect 40130 8132 40134 8188
rect 40070 8128 40134 8132
rect 12060 7644 12124 7648
rect 12060 7588 12064 7644
rect 12064 7588 12120 7644
rect 12120 7588 12124 7644
rect 12060 7584 12124 7588
rect 12140 7644 12204 7648
rect 12140 7588 12144 7644
rect 12144 7588 12200 7644
rect 12200 7588 12204 7644
rect 12140 7584 12204 7588
rect 12220 7644 12284 7648
rect 12220 7588 12224 7644
rect 12224 7588 12280 7644
rect 12280 7588 12284 7644
rect 12220 7584 12284 7588
rect 12300 7644 12364 7648
rect 12300 7588 12304 7644
rect 12304 7588 12360 7644
rect 12360 7588 12364 7644
rect 12300 7584 12364 7588
rect 23168 7644 23232 7648
rect 23168 7588 23172 7644
rect 23172 7588 23228 7644
rect 23228 7588 23232 7644
rect 23168 7584 23232 7588
rect 23248 7644 23312 7648
rect 23248 7588 23252 7644
rect 23252 7588 23308 7644
rect 23308 7588 23312 7644
rect 23248 7584 23312 7588
rect 23328 7644 23392 7648
rect 23328 7588 23332 7644
rect 23332 7588 23388 7644
rect 23388 7588 23392 7644
rect 23328 7584 23392 7588
rect 23408 7644 23472 7648
rect 23408 7588 23412 7644
rect 23412 7588 23468 7644
rect 23468 7588 23472 7644
rect 23408 7584 23472 7588
rect 34276 7644 34340 7648
rect 34276 7588 34280 7644
rect 34280 7588 34336 7644
rect 34336 7588 34340 7644
rect 34276 7584 34340 7588
rect 34356 7644 34420 7648
rect 34356 7588 34360 7644
rect 34360 7588 34416 7644
rect 34416 7588 34420 7644
rect 34356 7584 34420 7588
rect 34436 7644 34500 7648
rect 34436 7588 34440 7644
rect 34440 7588 34496 7644
rect 34496 7588 34500 7644
rect 34436 7584 34500 7588
rect 34516 7644 34580 7648
rect 34516 7588 34520 7644
rect 34520 7588 34576 7644
rect 34576 7588 34580 7644
rect 34516 7584 34580 7588
rect 45384 7644 45448 7648
rect 45384 7588 45388 7644
rect 45388 7588 45444 7644
rect 45444 7588 45448 7644
rect 45384 7584 45448 7588
rect 45464 7644 45528 7648
rect 45464 7588 45468 7644
rect 45468 7588 45524 7644
rect 45524 7588 45528 7644
rect 45464 7584 45528 7588
rect 45544 7644 45608 7648
rect 45544 7588 45548 7644
rect 45548 7588 45604 7644
rect 45604 7588 45608 7644
rect 45544 7584 45608 7588
rect 45624 7644 45688 7648
rect 45624 7588 45628 7644
rect 45628 7588 45684 7644
rect 45684 7588 45688 7644
rect 45624 7584 45688 7588
rect 6506 7100 6570 7104
rect 6506 7044 6510 7100
rect 6510 7044 6566 7100
rect 6566 7044 6570 7100
rect 6506 7040 6570 7044
rect 6586 7100 6650 7104
rect 6586 7044 6590 7100
rect 6590 7044 6646 7100
rect 6646 7044 6650 7100
rect 6586 7040 6650 7044
rect 6666 7100 6730 7104
rect 6666 7044 6670 7100
rect 6670 7044 6726 7100
rect 6726 7044 6730 7100
rect 6666 7040 6730 7044
rect 6746 7100 6810 7104
rect 6746 7044 6750 7100
rect 6750 7044 6806 7100
rect 6806 7044 6810 7100
rect 6746 7040 6810 7044
rect 17614 7100 17678 7104
rect 17614 7044 17618 7100
rect 17618 7044 17674 7100
rect 17674 7044 17678 7100
rect 17614 7040 17678 7044
rect 17694 7100 17758 7104
rect 17694 7044 17698 7100
rect 17698 7044 17754 7100
rect 17754 7044 17758 7100
rect 17694 7040 17758 7044
rect 17774 7100 17838 7104
rect 17774 7044 17778 7100
rect 17778 7044 17834 7100
rect 17834 7044 17838 7100
rect 17774 7040 17838 7044
rect 17854 7100 17918 7104
rect 17854 7044 17858 7100
rect 17858 7044 17914 7100
rect 17914 7044 17918 7100
rect 17854 7040 17918 7044
rect 28722 7100 28786 7104
rect 28722 7044 28726 7100
rect 28726 7044 28782 7100
rect 28782 7044 28786 7100
rect 28722 7040 28786 7044
rect 28802 7100 28866 7104
rect 28802 7044 28806 7100
rect 28806 7044 28862 7100
rect 28862 7044 28866 7100
rect 28802 7040 28866 7044
rect 28882 7100 28946 7104
rect 28882 7044 28886 7100
rect 28886 7044 28942 7100
rect 28942 7044 28946 7100
rect 28882 7040 28946 7044
rect 28962 7100 29026 7104
rect 28962 7044 28966 7100
rect 28966 7044 29022 7100
rect 29022 7044 29026 7100
rect 28962 7040 29026 7044
rect 39830 7100 39894 7104
rect 39830 7044 39834 7100
rect 39834 7044 39890 7100
rect 39890 7044 39894 7100
rect 39830 7040 39894 7044
rect 39910 7100 39974 7104
rect 39910 7044 39914 7100
rect 39914 7044 39970 7100
rect 39970 7044 39974 7100
rect 39910 7040 39974 7044
rect 39990 7100 40054 7104
rect 39990 7044 39994 7100
rect 39994 7044 40050 7100
rect 40050 7044 40054 7100
rect 39990 7040 40054 7044
rect 40070 7100 40134 7104
rect 40070 7044 40074 7100
rect 40074 7044 40130 7100
rect 40130 7044 40134 7100
rect 40070 7040 40134 7044
rect 12060 6556 12124 6560
rect 12060 6500 12064 6556
rect 12064 6500 12120 6556
rect 12120 6500 12124 6556
rect 12060 6496 12124 6500
rect 12140 6556 12204 6560
rect 12140 6500 12144 6556
rect 12144 6500 12200 6556
rect 12200 6500 12204 6556
rect 12140 6496 12204 6500
rect 12220 6556 12284 6560
rect 12220 6500 12224 6556
rect 12224 6500 12280 6556
rect 12280 6500 12284 6556
rect 12220 6496 12284 6500
rect 12300 6556 12364 6560
rect 12300 6500 12304 6556
rect 12304 6500 12360 6556
rect 12360 6500 12364 6556
rect 12300 6496 12364 6500
rect 23168 6556 23232 6560
rect 23168 6500 23172 6556
rect 23172 6500 23228 6556
rect 23228 6500 23232 6556
rect 23168 6496 23232 6500
rect 23248 6556 23312 6560
rect 23248 6500 23252 6556
rect 23252 6500 23308 6556
rect 23308 6500 23312 6556
rect 23248 6496 23312 6500
rect 23328 6556 23392 6560
rect 23328 6500 23332 6556
rect 23332 6500 23388 6556
rect 23388 6500 23392 6556
rect 23328 6496 23392 6500
rect 23408 6556 23472 6560
rect 23408 6500 23412 6556
rect 23412 6500 23468 6556
rect 23468 6500 23472 6556
rect 23408 6496 23472 6500
rect 34276 6556 34340 6560
rect 34276 6500 34280 6556
rect 34280 6500 34336 6556
rect 34336 6500 34340 6556
rect 34276 6496 34340 6500
rect 34356 6556 34420 6560
rect 34356 6500 34360 6556
rect 34360 6500 34416 6556
rect 34416 6500 34420 6556
rect 34356 6496 34420 6500
rect 34436 6556 34500 6560
rect 34436 6500 34440 6556
rect 34440 6500 34496 6556
rect 34496 6500 34500 6556
rect 34436 6496 34500 6500
rect 34516 6556 34580 6560
rect 34516 6500 34520 6556
rect 34520 6500 34576 6556
rect 34576 6500 34580 6556
rect 34516 6496 34580 6500
rect 45384 6556 45448 6560
rect 45384 6500 45388 6556
rect 45388 6500 45444 6556
rect 45444 6500 45448 6556
rect 45384 6496 45448 6500
rect 45464 6556 45528 6560
rect 45464 6500 45468 6556
rect 45468 6500 45524 6556
rect 45524 6500 45528 6556
rect 45464 6496 45528 6500
rect 45544 6556 45608 6560
rect 45544 6500 45548 6556
rect 45548 6500 45604 6556
rect 45604 6500 45608 6556
rect 45544 6496 45608 6500
rect 45624 6556 45688 6560
rect 45624 6500 45628 6556
rect 45628 6500 45684 6556
rect 45684 6500 45688 6556
rect 45624 6496 45688 6500
rect 6506 6012 6570 6016
rect 6506 5956 6510 6012
rect 6510 5956 6566 6012
rect 6566 5956 6570 6012
rect 6506 5952 6570 5956
rect 6586 6012 6650 6016
rect 6586 5956 6590 6012
rect 6590 5956 6646 6012
rect 6646 5956 6650 6012
rect 6586 5952 6650 5956
rect 6666 6012 6730 6016
rect 6666 5956 6670 6012
rect 6670 5956 6726 6012
rect 6726 5956 6730 6012
rect 6666 5952 6730 5956
rect 6746 6012 6810 6016
rect 6746 5956 6750 6012
rect 6750 5956 6806 6012
rect 6806 5956 6810 6012
rect 6746 5952 6810 5956
rect 17614 6012 17678 6016
rect 17614 5956 17618 6012
rect 17618 5956 17674 6012
rect 17674 5956 17678 6012
rect 17614 5952 17678 5956
rect 17694 6012 17758 6016
rect 17694 5956 17698 6012
rect 17698 5956 17754 6012
rect 17754 5956 17758 6012
rect 17694 5952 17758 5956
rect 17774 6012 17838 6016
rect 17774 5956 17778 6012
rect 17778 5956 17834 6012
rect 17834 5956 17838 6012
rect 17774 5952 17838 5956
rect 17854 6012 17918 6016
rect 17854 5956 17858 6012
rect 17858 5956 17914 6012
rect 17914 5956 17918 6012
rect 17854 5952 17918 5956
rect 28722 6012 28786 6016
rect 28722 5956 28726 6012
rect 28726 5956 28782 6012
rect 28782 5956 28786 6012
rect 28722 5952 28786 5956
rect 28802 6012 28866 6016
rect 28802 5956 28806 6012
rect 28806 5956 28862 6012
rect 28862 5956 28866 6012
rect 28802 5952 28866 5956
rect 28882 6012 28946 6016
rect 28882 5956 28886 6012
rect 28886 5956 28942 6012
rect 28942 5956 28946 6012
rect 28882 5952 28946 5956
rect 28962 6012 29026 6016
rect 28962 5956 28966 6012
rect 28966 5956 29022 6012
rect 29022 5956 29026 6012
rect 28962 5952 29026 5956
rect 39830 6012 39894 6016
rect 39830 5956 39834 6012
rect 39834 5956 39890 6012
rect 39890 5956 39894 6012
rect 39830 5952 39894 5956
rect 39910 6012 39974 6016
rect 39910 5956 39914 6012
rect 39914 5956 39970 6012
rect 39970 5956 39974 6012
rect 39910 5952 39974 5956
rect 39990 6012 40054 6016
rect 39990 5956 39994 6012
rect 39994 5956 40050 6012
rect 40050 5956 40054 6012
rect 39990 5952 40054 5956
rect 40070 6012 40134 6016
rect 40070 5956 40074 6012
rect 40074 5956 40130 6012
rect 40130 5956 40134 6012
rect 40070 5952 40134 5956
rect 12060 5468 12124 5472
rect 12060 5412 12064 5468
rect 12064 5412 12120 5468
rect 12120 5412 12124 5468
rect 12060 5408 12124 5412
rect 12140 5468 12204 5472
rect 12140 5412 12144 5468
rect 12144 5412 12200 5468
rect 12200 5412 12204 5468
rect 12140 5408 12204 5412
rect 12220 5468 12284 5472
rect 12220 5412 12224 5468
rect 12224 5412 12280 5468
rect 12280 5412 12284 5468
rect 12220 5408 12284 5412
rect 12300 5468 12364 5472
rect 12300 5412 12304 5468
rect 12304 5412 12360 5468
rect 12360 5412 12364 5468
rect 12300 5408 12364 5412
rect 23168 5468 23232 5472
rect 23168 5412 23172 5468
rect 23172 5412 23228 5468
rect 23228 5412 23232 5468
rect 23168 5408 23232 5412
rect 23248 5468 23312 5472
rect 23248 5412 23252 5468
rect 23252 5412 23308 5468
rect 23308 5412 23312 5468
rect 23248 5408 23312 5412
rect 23328 5468 23392 5472
rect 23328 5412 23332 5468
rect 23332 5412 23388 5468
rect 23388 5412 23392 5468
rect 23328 5408 23392 5412
rect 23408 5468 23472 5472
rect 23408 5412 23412 5468
rect 23412 5412 23468 5468
rect 23468 5412 23472 5468
rect 23408 5408 23472 5412
rect 34276 5468 34340 5472
rect 34276 5412 34280 5468
rect 34280 5412 34336 5468
rect 34336 5412 34340 5468
rect 34276 5408 34340 5412
rect 34356 5468 34420 5472
rect 34356 5412 34360 5468
rect 34360 5412 34416 5468
rect 34416 5412 34420 5468
rect 34356 5408 34420 5412
rect 34436 5468 34500 5472
rect 34436 5412 34440 5468
rect 34440 5412 34496 5468
rect 34496 5412 34500 5468
rect 34436 5408 34500 5412
rect 34516 5468 34580 5472
rect 34516 5412 34520 5468
rect 34520 5412 34576 5468
rect 34576 5412 34580 5468
rect 34516 5408 34580 5412
rect 45384 5468 45448 5472
rect 45384 5412 45388 5468
rect 45388 5412 45444 5468
rect 45444 5412 45448 5468
rect 45384 5408 45448 5412
rect 45464 5468 45528 5472
rect 45464 5412 45468 5468
rect 45468 5412 45524 5468
rect 45524 5412 45528 5468
rect 45464 5408 45528 5412
rect 45544 5468 45608 5472
rect 45544 5412 45548 5468
rect 45548 5412 45604 5468
rect 45604 5412 45608 5468
rect 45544 5408 45608 5412
rect 45624 5468 45688 5472
rect 45624 5412 45628 5468
rect 45628 5412 45684 5468
rect 45684 5412 45688 5468
rect 45624 5408 45688 5412
rect 6506 4924 6570 4928
rect 6506 4868 6510 4924
rect 6510 4868 6566 4924
rect 6566 4868 6570 4924
rect 6506 4864 6570 4868
rect 6586 4924 6650 4928
rect 6586 4868 6590 4924
rect 6590 4868 6646 4924
rect 6646 4868 6650 4924
rect 6586 4864 6650 4868
rect 6666 4924 6730 4928
rect 6666 4868 6670 4924
rect 6670 4868 6726 4924
rect 6726 4868 6730 4924
rect 6666 4864 6730 4868
rect 6746 4924 6810 4928
rect 6746 4868 6750 4924
rect 6750 4868 6806 4924
rect 6806 4868 6810 4924
rect 6746 4864 6810 4868
rect 17614 4924 17678 4928
rect 17614 4868 17618 4924
rect 17618 4868 17674 4924
rect 17674 4868 17678 4924
rect 17614 4864 17678 4868
rect 17694 4924 17758 4928
rect 17694 4868 17698 4924
rect 17698 4868 17754 4924
rect 17754 4868 17758 4924
rect 17694 4864 17758 4868
rect 17774 4924 17838 4928
rect 17774 4868 17778 4924
rect 17778 4868 17834 4924
rect 17834 4868 17838 4924
rect 17774 4864 17838 4868
rect 17854 4924 17918 4928
rect 17854 4868 17858 4924
rect 17858 4868 17914 4924
rect 17914 4868 17918 4924
rect 17854 4864 17918 4868
rect 28722 4924 28786 4928
rect 28722 4868 28726 4924
rect 28726 4868 28782 4924
rect 28782 4868 28786 4924
rect 28722 4864 28786 4868
rect 28802 4924 28866 4928
rect 28802 4868 28806 4924
rect 28806 4868 28862 4924
rect 28862 4868 28866 4924
rect 28802 4864 28866 4868
rect 28882 4924 28946 4928
rect 28882 4868 28886 4924
rect 28886 4868 28942 4924
rect 28942 4868 28946 4924
rect 28882 4864 28946 4868
rect 28962 4924 29026 4928
rect 28962 4868 28966 4924
rect 28966 4868 29022 4924
rect 29022 4868 29026 4924
rect 28962 4864 29026 4868
rect 39830 4924 39894 4928
rect 39830 4868 39834 4924
rect 39834 4868 39890 4924
rect 39890 4868 39894 4924
rect 39830 4864 39894 4868
rect 39910 4924 39974 4928
rect 39910 4868 39914 4924
rect 39914 4868 39970 4924
rect 39970 4868 39974 4924
rect 39910 4864 39974 4868
rect 39990 4924 40054 4928
rect 39990 4868 39994 4924
rect 39994 4868 40050 4924
rect 40050 4868 40054 4924
rect 39990 4864 40054 4868
rect 40070 4924 40134 4928
rect 40070 4868 40074 4924
rect 40074 4868 40130 4924
rect 40130 4868 40134 4924
rect 40070 4864 40134 4868
rect 12060 4380 12124 4384
rect 12060 4324 12064 4380
rect 12064 4324 12120 4380
rect 12120 4324 12124 4380
rect 12060 4320 12124 4324
rect 12140 4380 12204 4384
rect 12140 4324 12144 4380
rect 12144 4324 12200 4380
rect 12200 4324 12204 4380
rect 12140 4320 12204 4324
rect 12220 4380 12284 4384
rect 12220 4324 12224 4380
rect 12224 4324 12280 4380
rect 12280 4324 12284 4380
rect 12220 4320 12284 4324
rect 12300 4380 12364 4384
rect 12300 4324 12304 4380
rect 12304 4324 12360 4380
rect 12360 4324 12364 4380
rect 12300 4320 12364 4324
rect 23168 4380 23232 4384
rect 23168 4324 23172 4380
rect 23172 4324 23228 4380
rect 23228 4324 23232 4380
rect 23168 4320 23232 4324
rect 23248 4380 23312 4384
rect 23248 4324 23252 4380
rect 23252 4324 23308 4380
rect 23308 4324 23312 4380
rect 23248 4320 23312 4324
rect 23328 4380 23392 4384
rect 23328 4324 23332 4380
rect 23332 4324 23388 4380
rect 23388 4324 23392 4380
rect 23328 4320 23392 4324
rect 23408 4380 23472 4384
rect 23408 4324 23412 4380
rect 23412 4324 23468 4380
rect 23468 4324 23472 4380
rect 23408 4320 23472 4324
rect 34276 4380 34340 4384
rect 34276 4324 34280 4380
rect 34280 4324 34336 4380
rect 34336 4324 34340 4380
rect 34276 4320 34340 4324
rect 34356 4380 34420 4384
rect 34356 4324 34360 4380
rect 34360 4324 34416 4380
rect 34416 4324 34420 4380
rect 34356 4320 34420 4324
rect 34436 4380 34500 4384
rect 34436 4324 34440 4380
rect 34440 4324 34496 4380
rect 34496 4324 34500 4380
rect 34436 4320 34500 4324
rect 34516 4380 34580 4384
rect 34516 4324 34520 4380
rect 34520 4324 34576 4380
rect 34576 4324 34580 4380
rect 34516 4320 34580 4324
rect 45384 4380 45448 4384
rect 45384 4324 45388 4380
rect 45388 4324 45444 4380
rect 45444 4324 45448 4380
rect 45384 4320 45448 4324
rect 45464 4380 45528 4384
rect 45464 4324 45468 4380
rect 45468 4324 45524 4380
rect 45524 4324 45528 4380
rect 45464 4320 45528 4324
rect 45544 4380 45608 4384
rect 45544 4324 45548 4380
rect 45548 4324 45604 4380
rect 45604 4324 45608 4380
rect 45544 4320 45608 4324
rect 45624 4380 45688 4384
rect 45624 4324 45628 4380
rect 45628 4324 45684 4380
rect 45684 4324 45688 4380
rect 45624 4320 45688 4324
rect 6506 3836 6570 3840
rect 6506 3780 6510 3836
rect 6510 3780 6566 3836
rect 6566 3780 6570 3836
rect 6506 3776 6570 3780
rect 6586 3836 6650 3840
rect 6586 3780 6590 3836
rect 6590 3780 6646 3836
rect 6646 3780 6650 3836
rect 6586 3776 6650 3780
rect 6666 3836 6730 3840
rect 6666 3780 6670 3836
rect 6670 3780 6726 3836
rect 6726 3780 6730 3836
rect 6666 3776 6730 3780
rect 6746 3836 6810 3840
rect 6746 3780 6750 3836
rect 6750 3780 6806 3836
rect 6806 3780 6810 3836
rect 6746 3776 6810 3780
rect 17614 3836 17678 3840
rect 17614 3780 17618 3836
rect 17618 3780 17674 3836
rect 17674 3780 17678 3836
rect 17614 3776 17678 3780
rect 17694 3836 17758 3840
rect 17694 3780 17698 3836
rect 17698 3780 17754 3836
rect 17754 3780 17758 3836
rect 17694 3776 17758 3780
rect 17774 3836 17838 3840
rect 17774 3780 17778 3836
rect 17778 3780 17834 3836
rect 17834 3780 17838 3836
rect 17774 3776 17838 3780
rect 17854 3836 17918 3840
rect 17854 3780 17858 3836
rect 17858 3780 17914 3836
rect 17914 3780 17918 3836
rect 17854 3776 17918 3780
rect 28722 3836 28786 3840
rect 28722 3780 28726 3836
rect 28726 3780 28782 3836
rect 28782 3780 28786 3836
rect 28722 3776 28786 3780
rect 28802 3836 28866 3840
rect 28802 3780 28806 3836
rect 28806 3780 28862 3836
rect 28862 3780 28866 3836
rect 28802 3776 28866 3780
rect 28882 3836 28946 3840
rect 28882 3780 28886 3836
rect 28886 3780 28942 3836
rect 28942 3780 28946 3836
rect 28882 3776 28946 3780
rect 28962 3836 29026 3840
rect 28962 3780 28966 3836
rect 28966 3780 29022 3836
rect 29022 3780 29026 3836
rect 28962 3776 29026 3780
rect 39830 3836 39894 3840
rect 39830 3780 39834 3836
rect 39834 3780 39890 3836
rect 39890 3780 39894 3836
rect 39830 3776 39894 3780
rect 39910 3836 39974 3840
rect 39910 3780 39914 3836
rect 39914 3780 39970 3836
rect 39970 3780 39974 3836
rect 39910 3776 39974 3780
rect 39990 3836 40054 3840
rect 39990 3780 39994 3836
rect 39994 3780 40050 3836
rect 40050 3780 40054 3836
rect 39990 3776 40054 3780
rect 40070 3836 40134 3840
rect 40070 3780 40074 3836
rect 40074 3780 40130 3836
rect 40130 3780 40134 3836
rect 40070 3776 40134 3780
rect 12060 3292 12124 3296
rect 12060 3236 12064 3292
rect 12064 3236 12120 3292
rect 12120 3236 12124 3292
rect 12060 3232 12124 3236
rect 12140 3292 12204 3296
rect 12140 3236 12144 3292
rect 12144 3236 12200 3292
rect 12200 3236 12204 3292
rect 12140 3232 12204 3236
rect 12220 3292 12284 3296
rect 12220 3236 12224 3292
rect 12224 3236 12280 3292
rect 12280 3236 12284 3292
rect 12220 3232 12284 3236
rect 12300 3292 12364 3296
rect 12300 3236 12304 3292
rect 12304 3236 12360 3292
rect 12360 3236 12364 3292
rect 12300 3232 12364 3236
rect 23168 3292 23232 3296
rect 23168 3236 23172 3292
rect 23172 3236 23228 3292
rect 23228 3236 23232 3292
rect 23168 3232 23232 3236
rect 23248 3292 23312 3296
rect 23248 3236 23252 3292
rect 23252 3236 23308 3292
rect 23308 3236 23312 3292
rect 23248 3232 23312 3236
rect 23328 3292 23392 3296
rect 23328 3236 23332 3292
rect 23332 3236 23388 3292
rect 23388 3236 23392 3292
rect 23328 3232 23392 3236
rect 23408 3292 23472 3296
rect 23408 3236 23412 3292
rect 23412 3236 23468 3292
rect 23468 3236 23472 3292
rect 23408 3232 23472 3236
rect 34276 3292 34340 3296
rect 34276 3236 34280 3292
rect 34280 3236 34336 3292
rect 34336 3236 34340 3292
rect 34276 3232 34340 3236
rect 34356 3292 34420 3296
rect 34356 3236 34360 3292
rect 34360 3236 34416 3292
rect 34416 3236 34420 3292
rect 34356 3232 34420 3236
rect 34436 3292 34500 3296
rect 34436 3236 34440 3292
rect 34440 3236 34496 3292
rect 34496 3236 34500 3292
rect 34436 3232 34500 3236
rect 34516 3292 34580 3296
rect 34516 3236 34520 3292
rect 34520 3236 34576 3292
rect 34576 3236 34580 3292
rect 34516 3232 34580 3236
rect 45384 3292 45448 3296
rect 45384 3236 45388 3292
rect 45388 3236 45444 3292
rect 45444 3236 45448 3292
rect 45384 3232 45448 3236
rect 45464 3292 45528 3296
rect 45464 3236 45468 3292
rect 45468 3236 45524 3292
rect 45524 3236 45528 3292
rect 45464 3232 45528 3236
rect 45544 3292 45608 3296
rect 45544 3236 45548 3292
rect 45548 3236 45604 3292
rect 45604 3236 45608 3292
rect 45544 3232 45608 3236
rect 45624 3292 45688 3296
rect 45624 3236 45628 3292
rect 45628 3236 45684 3292
rect 45684 3236 45688 3292
rect 45624 3232 45688 3236
rect 6506 2748 6570 2752
rect 6506 2692 6510 2748
rect 6510 2692 6566 2748
rect 6566 2692 6570 2748
rect 6506 2688 6570 2692
rect 6586 2748 6650 2752
rect 6586 2692 6590 2748
rect 6590 2692 6646 2748
rect 6646 2692 6650 2748
rect 6586 2688 6650 2692
rect 6666 2748 6730 2752
rect 6666 2692 6670 2748
rect 6670 2692 6726 2748
rect 6726 2692 6730 2748
rect 6666 2688 6730 2692
rect 6746 2748 6810 2752
rect 6746 2692 6750 2748
rect 6750 2692 6806 2748
rect 6806 2692 6810 2748
rect 6746 2688 6810 2692
rect 17614 2748 17678 2752
rect 17614 2692 17618 2748
rect 17618 2692 17674 2748
rect 17674 2692 17678 2748
rect 17614 2688 17678 2692
rect 17694 2748 17758 2752
rect 17694 2692 17698 2748
rect 17698 2692 17754 2748
rect 17754 2692 17758 2748
rect 17694 2688 17758 2692
rect 17774 2748 17838 2752
rect 17774 2692 17778 2748
rect 17778 2692 17834 2748
rect 17834 2692 17838 2748
rect 17774 2688 17838 2692
rect 17854 2748 17918 2752
rect 17854 2692 17858 2748
rect 17858 2692 17914 2748
rect 17914 2692 17918 2748
rect 17854 2688 17918 2692
rect 28722 2748 28786 2752
rect 28722 2692 28726 2748
rect 28726 2692 28782 2748
rect 28782 2692 28786 2748
rect 28722 2688 28786 2692
rect 28802 2748 28866 2752
rect 28802 2692 28806 2748
rect 28806 2692 28862 2748
rect 28862 2692 28866 2748
rect 28802 2688 28866 2692
rect 28882 2748 28946 2752
rect 28882 2692 28886 2748
rect 28886 2692 28942 2748
rect 28942 2692 28946 2748
rect 28882 2688 28946 2692
rect 28962 2748 29026 2752
rect 28962 2692 28966 2748
rect 28966 2692 29022 2748
rect 29022 2692 29026 2748
rect 28962 2688 29026 2692
rect 39830 2748 39894 2752
rect 39830 2692 39834 2748
rect 39834 2692 39890 2748
rect 39890 2692 39894 2748
rect 39830 2688 39894 2692
rect 39910 2748 39974 2752
rect 39910 2692 39914 2748
rect 39914 2692 39970 2748
rect 39970 2692 39974 2748
rect 39910 2688 39974 2692
rect 39990 2748 40054 2752
rect 39990 2692 39994 2748
rect 39994 2692 40050 2748
rect 40050 2692 40054 2748
rect 39990 2688 40054 2692
rect 40070 2748 40134 2752
rect 40070 2692 40074 2748
rect 40074 2692 40130 2748
rect 40130 2692 40134 2748
rect 40070 2688 40134 2692
rect 12060 2204 12124 2208
rect 12060 2148 12064 2204
rect 12064 2148 12120 2204
rect 12120 2148 12124 2204
rect 12060 2144 12124 2148
rect 12140 2204 12204 2208
rect 12140 2148 12144 2204
rect 12144 2148 12200 2204
rect 12200 2148 12204 2204
rect 12140 2144 12204 2148
rect 12220 2204 12284 2208
rect 12220 2148 12224 2204
rect 12224 2148 12280 2204
rect 12280 2148 12284 2204
rect 12220 2144 12284 2148
rect 12300 2204 12364 2208
rect 12300 2148 12304 2204
rect 12304 2148 12360 2204
rect 12360 2148 12364 2204
rect 12300 2144 12364 2148
rect 23168 2204 23232 2208
rect 23168 2148 23172 2204
rect 23172 2148 23228 2204
rect 23228 2148 23232 2204
rect 23168 2144 23232 2148
rect 23248 2204 23312 2208
rect 23248 2148 23252 2204
rect 23252 2148 23308 2204
rect 23308 2148 23312 2204
rect 23248 2144 23312 2148
rect 23328 2204 23392 2208
rect 23328 2148 23332 2204
rect 23332 2148 23388 2204
rect 23388 2148 23392 2204
rect 23328 2144 23392 2148
rect 23408 2204 23472 2208
rect 23408 2148 23412 2204
rect 23412 2148 23468 2204
rect 23468 2148 23472 2204
rect 23408 2144 23472 2148
rect 34276 2204 34340 2208
rect 34276 2148 34280 2204
rect 34280 2148 34336 2204
rect 34336 2148 34340 2204
rect 34276 2144 34340 2148
rect 34356 2204 34420 2208
rect 34356 2148 34360 2204
rect 34360 2148 34416 2204
rect 34416 2148 34420 2204
rect 34356 2144 34420 2148
rect 34436 2204 34500 2208
rect 34436 2148 34440 2204
rect 34440 2148 34496 2204
rect 34496 2148 34500 2204
rect 34436 2144 34500 2148
rect 34516 2204 34580 2208
rect 34516 2148 34520 2204
rect 34520 2148 34576 2204
rect 34576 2148 34580 2204
rect 34516 2144 34580 2148
rect 45384 2204 45448 2208
rect 45384 2148 45388 2204
rect 45388 2148 45444 2204
rect 45444 2148 45448 2204
rect 45384 2144 45448 2148
rect 45464 2204 45528 2208
rect 45464 2148 45468 2204
rect 45468 2148 45524 2204
rect 45524 2148 45528 2204
rect 45464 2144 45528 2148
rect 45544 2204 45608 2208
rect 45544 2148 45548 2204
rect 45548 2148 45604 2204
rect 45604 2148 45608 2204
rect 45544 2144 45608 2148
rect 45624 2204 45688 2208
rect 45624 2148 45628 2204
rect 45628 2148 45684 2204
rect 45684 2148 45688 2204
rect 45624 2144 45688 2148
rect 6506 1660 6570 1664
rect 6506 1604 6510 1660
rect 6510 1604 6566 1660
rect 6566 1604 6570 1660
rect 6506 1600 6570 1604
rect 6586 1660 6650 1664
rect 6586 1604 6590 1660
rect 6590 1604 6646 1660
rect 6646 1604 6650 1660
rect 6586 1600 6650 1604
rect 6666 1660 6730 1664
rect 6666 1604 6670 1660
rect 6670 1604 6726 1660
rect 6726 1604 6730 1660
rect 6666 1600 6730 1604
rect 6746 1660 6810 1664
rect 6746 1604 6750 1660
rect 6750 1604 6806 1660
rect 6806 1604 6810 1660
rect 6746 1600 6810 1604
rect 17614 1660 17678 1664
rect 17614 1604 17618 1660
rect 17618 1604 17674 1660
rect 17674 1604 17678 1660
rect 17614 1600 17678 1604
rect 17694 1660 17758 1664
rect 17694 1604 17698 1660
rect 17698 1604 17754 1660
rect 17754 1604 17758 1660
rect 17694 1600 17758 1604
rect 17774 1660 17838 1664
rect 17774 1604 17778 1660
rect 17778 1604 17834 1660
rect 17834 1604 17838 1660
rect 17774 1600 17838 1604
rect 17854 1660 17918 1664
rect 17854 1604 17858 1660
rect 17858 1604 17914 1660
rect 17914 1604 17918 1660
rect 17854 1600 17918 1604
rect 28722 1660 28786 1664
rect 28722 1604 28726 1660
rect 28726 1604 28782 1660
rect 28782 1604 28786 1660
rect 28722 1600 28786 1604
rect 28802 1660 28866 1664
rect 28802 1604 28806 1660
rect 28806 1604 28862 1660
rect 28862 1604 28866 1660
rect 28802 1600 28866 1604
rect 28882 1660 28946 1664
rect 28882 1604 28886 1660
rect 28886 1604 28942 1660
rect 28942 1604 28946 1660
rect 28882 1600 28946 1604
rect 28962 1660 29026 1664
rect 28962 1604 28966 1660
rect 28966 1604 29022 1660
rect 29022 1604 29026 1660
rect 28962 1600 29026 1604
rect 39830 1660 39894 1664
rect 39830 1604 39834 1660
rect 39834 1604 39890 1660
rect 39890 1604 39894 1660
rect 39830 1600 39894 1604
rect 39910 1660 39974 1664
rect 39910 1604 39914 1660
rect 39914 1604 39970 1660
rect 39970 1604 39974 1660
rect 39910 1600 39974 1604
rect 39990 1660 40054 1664
rect 39990 1604 39994 1660
rect 39994 1604 40050 1660
rect 40050 1604 40054 1660
rect 39990 1600 40054 1604
rect 40070 1660 40134 1664
rect 40070 1604 40074 1660
rect 40074 1604 40130 1660
rect 40130 1604 40134 1660
rect 40070 1600 40134 1604
rect 12060 1116 12124 1120
rect 12060 1060 12064 1116
rect 12064 1060 12120 1116
rect 12120 1060 12124 1116
rect 12060 1056 12124 1060
rect 12140 1116 12204 1120
rect 12140 1060 12144 1116
rect 12144 1060 12200 1116
rect 12200 1060 12204 1116
rect 12140 1056 12204 1060
rect 12220 1116 12284 1120
rect 12220 1060 12224 1116
rect 12224 1060 12280 1116
rect 12280 1060 12284 1116
rect 12220 1056 12284 1060
rect 12300 1116 12364 1120
rect 12300 1060 12304 1116
rect 12304 1060 12360 1116
rect 12360 1060 12364 1116
rect 12300 1056 12364 1060
rect 23168 1116 23232 1120
rect 23168 1060 23172 1116
rect 23172 1060 23228 1116
rect 23228 1060 23232 1116
rect 23168 1056 23232 1060
rect 23248 1116 23312 1120
rect 23248 1060 23252 1116
rect 23252 1060 23308 1116
rect 23308 1060 23312 1116
rect 23248 1056 23312 1060
rect 23328 1116 23392 1120
rect 23328 1060 23332 1116
rect 23332 1060 23388 1116
rect 23388 1060 23392 1116
rect 23328 1056 23392 1060
rect 23408 1116 23472 1120
rect 23408 1060 23412 1116
rect 23412 1060 23468 1116
rect 23468 1060 23472 1116
rect 23408 1056 23472 1060
rect 34276 1116 34340 1120
rect 34276 1060 34280 1116
rect 34280 1060 34336 1116
rect 34336 1060 34340 1116
rect 34276 1056 34340 1060
rect 34356 1116 34420 1120
rect 34356 1060 34360 1116
rect 34360 1060 34416 1116
rect 34416 1060 34420 1116
rect 34356 1056 34420 1060
rect 34436 1116 34500 1120
rect 34436 1060 34440 1116
rect 34440 1060 34496 1116
rect 34496 1060 34500 1116
rect 34436 1056 34500 1060
rect 34516 1116 34580 1120
rect 34516 1060 34520 1116
rect 34520 1060 34576 1116
rect 34576 1060 34580 1116
rect 34516 1056 34580 1060
rect 45384 1116 45448 1120
rect 45384 1060 45388 1116
rect 45388 1060 45444 1116
rect 45444 1060 45448 1116
rect 45384 1056 45448 1060
rect 45464 1116 45528 1120
rect 45464 1060 45468 1116
rect 45468 1060 45524 1116
rect 45524 1060 45528 1116
rect 45464 1056 45528 1060
rect 45544 1116 45608 1120
rect 45544 1060 45548 1116
rect 45548 1060 45604 1116
rect 45604 1060 45608 1116
rect 45544 1056 45608 1060
rect 45624 1116 45688 1120
rect 45624 1060 45628 1116
rect 45628 1060 45684 1116
rect 45684 1060 45688 1116
rect 45624 1056 45688 1060
<< metal4 >>
rect 6498 8192 6818 8752
rect 6498 8128 6506 8192
rect 6570 8128 6586 8192
rect 6650 8128 6666 8192
rect 6730 8128 6746 8192
rect 6810 8128 6818 8192
rect 6498 7104 6818 8128
rect 6498 7040 6506 7104
rect 6570 7040 6586 7104
rect 6650 7040 6666 7104
rect 6730 7040 6746 7104
rect 6810 7040 6818 7104
rect 6498 6016 6818 7040
rect 6498 5952 6506 6016
rect 6570 5952 6586 6016
rect 6650 5952 6666 6016
rect 6730 5952 6746 6016
rect 6810 5952 6818 6016
rect 6498 4928 6818 5952
rect 6498 4864 6506 4928
rect 6570 4864 6586 4928
rect 6650 4864 6666 4928
rect 6730 4864 6746 4928
rect 6810 4864 6818 4928
rect 6498 3840 6818 4864
rect 6498 3776 6506 3840
rect 6570 3776 6586 3840
rect 6650 3776 6666 3840
rect 6730 3776 6746 3840
rect 6810 3776 6818 3840
rect 6498 2752 6818 3776
rect 6498 2688 6506 2752
rect 6570 2688 6586 2752
rect 6650 2688 6666 2752
rect 6730 2688 6746 2752
rect 6810 2688 6818 2752
rect 6498 1664 6818 2688
rect 6498 1600 6506 1664
rect 6570 1600 6586 1664
rect 6650 1600 6666 1664
rect 6730 1600 6746 1664
rect 6810 1600 6818 1664
rect 6498 1040 6818 1600
rect 12052 8736 12372 8752
rect 12052 8672 12060 8736
rect 12124 8672 12140 8736
rect 12204 8672 12220 8736
rect 12284 8672 12300 8736
rect 12364 8672 12372 8736
rect 12052 7648 12372 8672
rect 12052 7584 12060 7648
rect 12124 7584 12140 7648
rect 12204 7584 12220 7648
rect 12284 7584 12300 7648
rect 12364 7584 12372 7648
rect 12052 6560 12372 7584
rect 12052 6496 12060 6560
rect 12124 6496 12140 6560
rect 12204 6496 12220 6560
rect 12284 6496 12300 6560
rect 12364 6496 12372 6560
rect 12052 5472 12372 6496
rect 12052 5408 12060 5472
rect 12124 5408 12140 5472
rect 12204 5408 12220 5472
rect 12284 5408 12300 5472
rect 12364 5408 12372 5472
rect 12052 4384 12372 5408
rect 12052 4320 12060 4384
rect 12124 4320 12140 4384
rect 12204 4320 12220 4384
rect 12284 4320 12300 4384
rect 12364 4320 12372 4384
rect 12052 3296 12372 4320
rect 12052 3232 12060 3296
rect 12124 3232 12140 3296
rect 12204 3232 12220 3296
rect 12284 3232 12300 3296
rect 12364 3232 12372 3296
rect 12052 2208 12372 3232
rect 12052 2144 12060 2208
rect 12124 2144 12140 2208
rect 12204 2144 12220 2208
rect 12284 2144 12300 2208
rect 12364 2144 12372 2208
rect 12052 1120 12372 2144
rect 12052 1056 12060 1120
rect 12124 1056 12140 1120
rect 12204 1056 12220 1120
rect 12284 1056 12300 1120
rect 12364 1056 12372 1120
rect 12052 1040 12372 1056
rect 17606 8192 17926 8752
rect 17606 8128 17614 8192
rect 17678 8128 17694 8192
rect 17758 8128 17774 8192
rect 17838 8128 17854 8192
rect 17918 8128 17926 8192
rect 17606 7104 17926 8128
rect 17606 7040 17614 7104
rect 17678 7040 17694 7104
rect 17758 7040 17774 7104
rect 17838 7040 17854 7104
rect 17918 7040 17926 7104
rect 17606 6016 17926 7040
rect 17606 5952 17614 6016
rect 17678 5952 17694 6016
rect 17758 5952 17774 6016
rect 17838 5952 17854 6016
rect 17918 5952 17926 6016
rect 17606 4928 17926 5952
rect 17606 4864 17614 4928
rect 17678 4864 17694 4928
rect 17758 4864 17774 4928
rect 17838 4864 17854 4928
rect 17918 4864 17926 4928
rect 17606 3840 17926 4864
rect 17606 3776 17614 3840
rect 17678 3776 17694 3840
rect 17758 3776 17774 3840
rect 17838 3776 17854 3840
rect 17918 3776 17926 3840
rect 17606 2752 17926 3776
rect 17606 2688 17614 2752
rect 17678 2688 17694 2752
rect 17758 2688 17774 2752
rect 17838 2688 17854 2752
rect 17918 2688 17926 2752
rect 17606 1664 17926 2688
rect 17606 1600 17614 1664
rect 17678 1600 17694 1664
rect 17758 1600 17774 1664
rect 17838 1600 17854 1664
rect 17918 1600 17926 1664
rect 17606 1040 17926 1600
rect 23160 8736 23480 8752
rect 23160 8672 23168 8736
rect 23232 8672 23248 8736
rect 23312 8672 23328 8736
rect 23392 8672 23408 8736
rect 23472 8672 23480 8736
rect 23160 7648 23480 8672
rect 23160 7584 23168 7648
rect 23232 7584 23248 7648
rect 23312 7584 23328 7648
rect 23392 7584 23408 7648
rect 23472 7584 23480 7648
rect 23160 6560 23480 7584
rect 23160 6496 23168 6560
rect 23232 6496 23248 6560
rect 23312 6496 23328 6560
rect 23392 6496 23408 6560
rect 23472 6496 23480 6560
rect 23160 5472 23480 6496
rect 23160 5408 23168 5472
rect 23232 5408 23248 5472
rect 23312 5408 23328 5472
rect 23392 5408 23408 5472
rect 23472 5408 23480 5472
rect 23160 4384 23480 5408
rect 23160 4320 23168 4384
rect 23232 4320 23248 4384
rect 23312 4320 23328 4384
rect 23392 4320 23408 4384
rect 23472 4320 23480 4384
rect 23160 3296 23480 4320
rect 23160 3232 23168 3296
rect 23232 3232 23248 3296
rect 23312 3232 23328 3296
rect 23392 3232 23408 3296
rect 23472 3232 23480 3296
rect 23160 2208 23480 3232
rect 23160 2144 23168 2208
rect 23232 2144 23248 2208
rect 23312 2144 23328 2208
rect 23392 2144 23408 2208
rect 23472 2144 23480 2208
rect 23160 1120 23480 2144
rect 23160 1056 23168 1120
rect 23232 1056 23248 1120
rect 23312 1056 23328 1120
rect 23392 1056 23408 1120
rect 23472 1056 23480 1120
rect 23160 1040 23480 1056
rect 28714 8192 29034 8752
rect 28714 8128 28722 8192
rect 28786 8128 28802 8192
rect 28866 8128 28882 8192
rect 28946 8128 28962 8192
rect 29026 8128 29034 8192
rect 28714 7104 29034 8128
rect 28714 7040 28722 7104
rect 28786 7040 28802 7104
rect 28866 7040 28882 7104
rect 28946 7040 28962 7104
rect 29026 7040 29034 7104
rect 28714 6016 29034 7040
rect 28714 5952 28722 6016
rect 28786 5952 28802 6016
rect 28866 5952 28882 6016
rect 28946 5952 28962 6016
rect 29026 5952 29034 6016
rect 28714 4928 29034 5952
rect 28714 4864 28722 4928
rect 28786 4864 28802 4928
rect 28866 4864 28882 4928
rect 28946 4864 28962 4928
rect 29026 4864 29034 4928
rect 28714 3840 29034 4864
rect 28714 3776 28722 3840
rect 28786 3776 28802 3840
rect 28866 3776 28882 3840
rect 28946 3776 28962 3840
rect 29026 3776 29034 3840
rect 28714 2752 29034 3776
rect 28714 2688 28722 2752
rect 28786 2688 28802 2752
rect 28866 2688 28882 2752
rect 28946 2688 28962 2752
rect 29026 2688 29034 2752
rect 28714 1664 29034 2688
rect 28714 1600 28722 1664
rect 28786 1600 28802 1664
rect 28866 1600 28882 1664
rect 28946 1600 28962 1664
rect 29026 1600 29034 1664
rect 28714 1040 29034 1600
rect 34268 8736 34588 8752
rect 34268 8672 34276 8736
rect 34340 8672 34356 8736
rect 34420 8672 34436 8736
rect 34500 8672 34516 8736
rect 34580 8672 34588 8736
rect 34268 7648 34588 8672
rect 34268 7584 34276 7648
rect 34340 7584 34356 7648
rect 34420 7584 34436 7648
rect 34500 7584 34516 7648
rect 34580 7584 34588 7648
rect 34268 6560 34588 7584
rect 34268 6496 34276 6560
rect 34340 6496 34356 6560
rect 34420 6496 34436 6560
rect 34500 6496 34516 6560
rect 34580 6496 34588 6560
rect 34268 5472 34588 6496
rect 34268 5408 34276 5472
rect 34340 5408 34356 5472
rect 34420 5408 34436 5472
rect 34500 5408 34516 5472
rect 34580 5408 34588 5472
rect 34268 4384 34588 5408
rect 34268 4320 34276 4384
rect 34340 4320 34356 4384
rect 34420 4320 34436 4384
rect 34500 4320 34516 4384
rect 34580 4320 34588 4384
rect 34268 3296 34588 4320
rect 34268 3232 34276 3296
rect 34340 3232 34356 3296
rect 34420 3232 34436 3296
rect 34500 3232 34516 3296
rect 34580 3232 34588 3296
rect 34268 2208 34588 3232
rect 34268 2144 34276 2208
rect 34340 2144 34356 2208
rect 34420 2144 34436 2208
rect 34500 2144 34516 2208
rect 34580 2144 34588 2208
rect 34268 1120 34588 2144
rect 34268 1056 34276 1120
rect 34340 1056 34356 1120
rect 34420 1056 34436 1120
rect 34500 1056 34516 1120
rect 34580 1056 34588 1120
rect 34268 1040 34588 1056
rect 39822 8192 40142 8752
rect 39822 8128 39830 8192
rect 39894 8128 39910 8192
rect 39974 8128 39990 8192
rect 40054 8128 40070 8192
rect 40134 8128 40142 8192
rect 39822 7104 40142 8128
rect 39822 7040 39830 7104
rect 39894 7040 39910 7104
rect 39974 7040 39990 7104
rect 40054 7040 40070 7104
rect 40134 7040 40142 7104
rect 39822 6016 40142 7040
rect 39822 5952 39830 6016
rect 39894 5952 39910 6016
rect 39974 5952 39990 6016
rect 40054 5952 40070 6016
rect 40134 5952 40142 6016
rect 39822 4928 40142 5952
rect 39822 4864 39830 4928
rect 39894 4864 39910 4928
rect 39974 4864 39990 4928
rect 40054 4864 40070 4928
rect 40134 4864 40142 4928
rect 39822 3840 40142 4864
rect 39822 3776 39830 3840
rect 39894 3776 39910 3840
rect 39974 3776 39990 3840
rect 40054 3776 40070 3840
rect 40134 3776 40142 3840
rect 39822 2752 40142 3776
rect 39822 2688 39830 2752
rect 39894 2688 39910 2752
rect 39974 2688 39990 2752
rect 40054 2688 40070 2752
rect 40134 2688 40142 2752
rect 39822 1664 40142 2688
rect 39822 1600 39830 1664
rect 39894 1600 39910 1664
rect 39974 1600 39990 1664
rect 40054 1600 40070 1664
rect 40134 1600 40142 1664
rect 39822 1040 40142 1600
rect 45376 8736 45696 8752
rect 45376 8672 45384 8736
rect 45448 8672 45464 8736
rect 45528 8672 45544 8736
rect 45608 8672 45624 8736
rect 45688 8672 45696 8736
rect 45376 7648 45696 8672
rect 45376 7584 45384 7648
rect 45448 7584 45464 7648
rect 45528 7584 45544 7648
rect 45608 7584 45624 7648
rect 45688 7584 45696 7648
rect 45376 6560 45696 7584
rect 45376 6496 45384 6560
rect 45448 6496 45464 6560
rect 45528 6496 45544 6560
rect 45608 6496 45624 6560
rect 45688 6496 45696 6560
rect 45376 5472 45696 6496
rect 45376 5408 45384 5472
rect 45448 5408 45464 5472
rect 45528 5408 45544 5472
rect 45608 5408 45624 5472
rect 45688 5408 45696 5472
rect 45376 4384 45696 5408
rect 45376 4320 45384 4384
rect 45448 4320 45464 4384
rect 45528 4320 45544 4384
rect 45608 4320 45624 4384
rect 45688 4320 45696 4384
rect 45376 3296 45696 4320
rect 45376 3232 45384 3296
rect 45448 3232 45464 3296
rect 45528 3232 45544 3296
rect 45608 3232 45624 3296
rect 45688 3232 45696 3296
rect 45376 2208 45696 3232
rect 45376 2144 45384 2208
rect 45448 2144 45464 2208
rect 45528 2144 45544 2208
rect 45608 2144 45624 2208
rect 45688 2144 45696 2208
rect 45376 1120 45696 2144
rect 45376 1056 45384 1120
rect 45448 1056 45464 1120
rect 45528 1056 45544 1120
rect 45608 1056 45624 1120
rect 45688 1056 45696 1120
rect 45376 1040 45696 1056
use sky130_fd_sc_hd__fill_2  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_33
timestamp 1688980957
transform 1 0 4140 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_45
timestamp 1688980957
transform 1 0 5244 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_49
timestamp 1688980957
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_61
timestamp 1688980957
transform 1 0 6716 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_73
timestamp 1688980957
transform 1 0 7820 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_77
timestamp 1688980957
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_89
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_93
timestamp 1688980957
transform 1 0 9660 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10764 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_117
timestamp 1688980957
transform 1 0 11868 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_182
timestamp 1688980957
transform 1 0 17848 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_218
timestamp 1688980957
transform 1 0 21160 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_234
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_246
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_272
timestamp 1688980957
transform 1 0 26128 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_315
timestamp 1688980957
transform 1 0 30084 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_347
timestamp 1688980957
transform 1 0 33028 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34316 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_430
timestamp 1688980957
transform 1 0 40664 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_9
timestamp 1688980957
transform 1 0 1932 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_20
timestamp 1688980957
transform 1 0 2944 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3404 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_37
timestamp 1688980957
transform 1 0 4508 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_158
timestamp 1688980957
transform 1 0 15640 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_220
timestamp 1688980957
transform 1 0 21344 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_236
timestamp 1688980957
transform 1 0 22816 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_248
timestamp 1688980957
transform 1 0 23920 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_255
timestamp 1688980957
transform 1 0 24564 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_268
timestamp 1688980957
transform 1 0 25760 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_296
timestamp 1688980957
transform 1 0 28336 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_340 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32384 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_344
timestamp 1688980957
transform 1 0 32752 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_352
timestamp 1688980957
transform 1 0 33488 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_364
timestamp 1688980957
transform 1 0 34592 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_377
timestamp 1688980957
transform 1 0 35788 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_381
timestamp 1688980957
transform 1 0 36156 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_388
timestamp 1688980957
transform 1 0 36800 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_397
timestamp 1688980957
transform 1 0 37628 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_409 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38732 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_422
timestamp 1688980957
transform 1 0 39928 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_433
timestamp 1688980957
transform 1 0 40940 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_441
timestamp 1688980957
transform 1 0 41676 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_445
timestamp 1688980957
transform 1 0 42044 0 -1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_469
timestamp 1688980957
transform 1 0 44252 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_476
timestamp 1688980957
transform 1 0 44896 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_176
timestamp 1688980957
transform 1 0 17296 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_188
timestamp 1688980957
transform 1 0 18400 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_207
timestamp 1688980957
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_215
timestamp 1688980957
transform 1 0 20884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_220
timestamp 1688980957
transform 1 0 21344 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_240
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_256
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_268
timestamp 1688980957
transform 1 0 25760 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_273
timestamp 1688980957
transform 1 0 26220 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_285
timestamp 1688980957
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_293
timestamp 1688980957
transform 1 0 28060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_297
timestamp 1688980957
transform 1 0 28428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_317
timestamp 1688980957
transform 1 0 30268 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_330
timestamp 1688980957
transform 1 0 31464 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_369
timestamp 1688980957
transform 1 0 35052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_381
timestamp 1688980957
transform 1 0 36156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_405
timestamp 1688980957
transform 1 0 38364 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_416
timestamp 1688980957
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_440
timestamp 1688980957
transform 1 0 41584 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_452
timestamp 1688980957
transform 1 0 42688 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_467
timestamp 1688980957
transform 1 0 44068 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_228
timestamp 1688980957
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_234
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_238
timestamp 1688980957
transform 1 0 23000 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_243
timestamp 1688980957
transform 1 0 23460 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_255
timestamp 1688980957
transform 1 0 24564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_267
timestamp 1688980957
transform 1 0 25668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_479
timestamp 1688980957
transform 1 0 45172 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_479
timestamp 1688980957
transform 1 0 45172 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_479
timestamp 1688980957
transform 1 0 45172 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_479
timestamp 1688980957
transform 1 0 45172 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_473
timestamp 1688980957
transform 1 0 44620 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_479
timestamp 1688980957
transform 1 0 45172 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 1688980957
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_21
timestamp 1688980957
transform 1 0 3036 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_33
timestamp 1688980957
transform 1 0 4140 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_45
timestamp 1688980957
transform 1 0 5244 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_73
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_78
timestamp 1688980957
transform 1 0 8280 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_97
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_119
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_126
timestamp 1688980957
transform 1 0 12696 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_138
timestamp 1688980957
transform 1 0 13800 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_150
timestamp 1688980957
transform 1 0 14904 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_162
timestamp 1688980957
transform 1 0 16008 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_175
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_187
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_195
timestamp 1688980957
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_203
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_215
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_246
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_265
timestamp 1688980957
transform 1 0 25484 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_270
timestamp 1688980957
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 1688980957
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_287
timestamp 1688980957
transform 1 0 27508 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_294
timestamp 1688980957
transform 1 0 28152 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_306
timestamp 1688980957
transform 1 0 29256 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_309
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_313
timestamp 1688980957
transform 1 0 29900 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_318
timestamp 1688980957
transform 1 0 30360 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_330
timestamp 1688980957
transform 1 0 31464 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_342
timestamp 1688980957
transform 1 0 32568 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_354
timestamp 1688980957
transform 1 0 33672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_362
timestamp 1688980957
transform 1 0 34408 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_371
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_383
timestamp 1688980957
transform 1 0 36340 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_390
timestamp 1688980957
transform 1 0 36984 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_414
timestamp 1688980957
transform 1 0 39192 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_421
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_433
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_438
timestamp 1688980957
transform 1 0 41400 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_446
timestamp 1688980957
transform 1 0 42136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_457
timestamp 1688980957
transform 1 0 43148 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_462
timestamp 1688980957
transform 1 0 43608 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_470
timestamp 1688980957
transform 1 0 44344 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_477
timestamp 1688980957
transform 1 0 44988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 40664 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1688980957
transform -1 0 43516 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1688980957
transform -1 0 43792 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform -1 0 44068 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform -1 0 44344 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform -1 0 44620 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 44620 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 44988 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform -1 0 40388 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 40664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform -1 0 40940 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform -1 0 42044 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform -1 0 42320 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40848 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform -1 0 42688 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 42964 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform -1 0 43240 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input21
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 1656 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 4968 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 5336 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 6440 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 1688980957
transform 1 0 6808 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 1688980957
transform 1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 7544 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1688980957
transform 1 0 2024 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1688980957
transform 1 0 2392 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 2116 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 3128 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 3864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 4232 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 4600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 11592 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 11960 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 9016 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 9384 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 9752 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 10488 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input55
timestamp 1688980957
transform 1 0 10856 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform -1 0 17020 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform 1 0 17296 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 18032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1688980957
transform 1 0 18584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1688980957
transform -1 0 13984 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1688980957
transform -1 0 14352 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1688980957
transform -1 0 14628 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1688980957
transform -1 0 14904 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1688980957
transform -1 0 15180 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1688980957
transform -1 0 15456 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1688980957
transform -1 0 15732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1688980957
transform -1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1688980957
transform -1 0 16560 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform -1 0 39744 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__00_
timestamp 1688980957
transform -1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__01_
timestamp 1688980957
transform -1 0 22356 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__02_
timestamp 1688980957
transform -1 0 23276 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__03_
timestamp 1688980957
transform -1 0 24564 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__04_
timestamp 1688980957
transform -1 0 24932 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__05_
timestamp 1688980957
transform -1 0 25484 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__06_
timestamp 1688980957
transform -1 0 26588 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__07_
timestamp 1688980957
transform -1 0 26864 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__08_
timestamp 1688980957
transform -1 0 19596 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__09_
timestamp 1688980957
transform -1 0 19872 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__10_
timestamp 1688980957
transform -1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__11_
timestamp 1688980957
transform -1 0 20148 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__12_
timestamp 1688980957
transform -1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__13_
timestamp 1688980957
transform -1 0 20976 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__14_
timestamp 1688980957
transform -1 0 22080 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__15_
timestamp 1688980957
transform -1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__16_
timestamp 1688980957
transform -1 0 27232 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__17_
timestamp 1688980957
transform -1 0 27784 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__18_
timestamp 1688980957
transform -1 0 30912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__19_
timestamp 1688980957
transform -1 0 31188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__20_
timestamp 1688980957
transform -1 0 31464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__21_
timestamp 1688980957
transform -1 0 29624 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__22_
timestamp 1688980957
transform -1 0 28060 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__23_
timestamp 1688980957
transform 1 0 25484 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__24_
timestamp 1688980957
transform -1 0 28060 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__25_
timestamp 1688980957
transform -1 0 28336 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__26_
timestamp 1688980957
transform -1 0 29072 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__27_
timestamp 1688980957
transform -1 0 29348 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__28_
timestamp 1688980957
transform -1 0 29900 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__29_
timestamp 1688980957
transform -1 0 30544 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__30_
timestamp 1688980957
transform -1 0 30820 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__31_
timestamp 1688980957
transform -1 0 31096 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__32_
timestamp 1688980957
transform 1 0 18768 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__33_
timestamp 1688980957
transform 1 0 18216 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__34_
timestamp 1688980957
transform 1 0 15732 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__35_
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__36_
timestamp 1688980957
transform 1 0 14996 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__37_
timestamp 1688980957
transform 1 0 19044 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__38_
timestamp 1688980957
transform 1 0 20148 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__39_
timestamp 1688980957
transform 1 0 22724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__40_
timestamp 1688980957
transform 1 0 17940 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__41_
timestamp 1688980957
transform 1 0 17664 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__42_
timestamp 1688980957
transform 1 0 17388 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__43_
timestamp 1688980957
transform 1 0 17112 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__44_
timestamp 1688980957
transform 1 0 16836 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__45_
timestamp 1688980957
transform 1 0 17020 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__46_
timestamp 1688980957
transform 1 0 16284 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_single2_switch_matrix__47_
timestamp 1688980957
transform 1 0 16008 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__48_
timestamp 1688980957
transform -1 0 19044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__49_
timestamp 1688980957
transform -1 0 19504 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__50_
timestamp 1688980957
transform -1 0 19872 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_single2_switch_matrix__51_
timestamp 1688980957
transform -1 0 20148 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4140 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1688980957
transform -1 0 25944 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output76 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28152 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1688980957
transform -1 0 30360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1688980957
transform -1 0 32568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform -1 0 36984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform -1 0 39192 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1688980957
transform -1 0 41400 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1688980957
transform -1 0 43608 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 44528 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform -1 0 6072 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1688980957
transform -1 0 8280 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1688980957
transform -1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform -1 0 12696 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1688980957
transform -1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform -1 0 17204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1688980957
transform -1 0 21528 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform -1 0 23736 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1688980957
transform 1 0 19872 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 20240 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 20608 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1688980957
transform 1 0 23920 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1688980957
transform 1 0 24472 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 24840 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 25392 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 25760 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1688980957
transform 1 0 25944 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform -1 0 26864 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1688980957
transform 1 0 20976 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1688980957
transform 1 0 21344 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 21896 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1688980957
transform 1 0 22448 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1688980957
transform 1 0 22816 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 23184 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 23552 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1688980957
transform 1 0 27324 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1688980957
transform 1 0 31648 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output116
timestamp 1688980957
transform 1 0 31096 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1688980957
transform 1 0 32660 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1688980957
transform 1 0 32844 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform 1 0 33212 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 27692 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1688980957
transform 1 0 28244 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1688980957
transform 1 0 28428 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform -1 0 29348 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1688980957
transform 1 0 29900 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform -1 0 30820 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output128
timestamp 1688980957
transform 1 0 30820 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 31372 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 33764 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform 1 0 37812 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 38364 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1688980957
transform 1 0 37996 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1688980957
transform 1 0 38364 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 38916 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1688980957
transform 1 0 34224 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output138
timestamp 1688980957
transform 1 0 33672 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 35236 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1688980957
transform 1 0 35420 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform 1 0 35788 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform 1 0 36340 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output145
timestamp 1688980957
transform 1 0 36248 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 45540 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 45540 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 45540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 45540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 45540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 45540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 45540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 45540 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 45540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 45540 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 45540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 45540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 45540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 45540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 24012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform -1 0 21712 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform -1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform -1 0 23552 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 23184 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 17572 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform -1 0 18768 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform -1 0 20700 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 24932 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 27232 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 33212 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 35144 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 37352 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 39652 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 41768 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 44344 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 44620 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_0__0_
timestamp 1688980957
transform -1 0 23920 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform -1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform -1 0 23552 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform -1 0 24656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform -1 0 22632 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform -1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 19320 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 21528 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 25944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 28152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 30360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 32568 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 34776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 36984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 39100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 41308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 43792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform -1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 44896 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 39118 -300 39174 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 42798 -300 42854 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 43166 -300 43222 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 43534 -300 43590 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 43902 -300 43958 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 44270 -300 44326 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 44638 -300 44694 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 45006 -300 45062 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 45374 -300 45430 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 45742 -300 45798 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 46110 -300 46166 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 39486 -300 39542 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 39854 -300 39910 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 40222 -300 40278 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 40590 -300 40646 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 40958 -300 41014 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 41326 -300 41382 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 41694 -300 41750 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 42062 -300 42118 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 42430 -300 42486 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 3422 9840 3478 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 25502 9840 25558 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 27710 9840 27766 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 29918 9840 29974 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 32126 9840 32182 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 34334 9840 34390 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 36542 9840 36598 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 38750 9840 38806 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 40958 9840 41014 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 43166 9840 43222 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 45374 9840 45430 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 5630 9840 5686 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 7838 9840 7894 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 10046 9840 10102 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 12254 9840 12310 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 14462 9840 14518 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 16670 9840 16726 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 18878 9840 18934 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 21086 9840 21142 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 23294 9840 23350 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 478 -300 534 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 846 -300 902 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 1214 -300 1270 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 1582 -300 1638 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 4894 -300 4950 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 5262 -300 5318 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 5630 -300 5686 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 5998 -300 6054 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 6366 -300 6422 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 6734 -300 6790 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 7102 -300 7158 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 7470 -300 7526 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 1950 -300 2006 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 2318 -300 2374 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 2686 -300 2742 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 3054 -300 3110 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 3422 -300 3478 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 3790 -300 3846 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 4158 -300 4214 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 4526 -300 4582 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 7838 -300 7894 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 11518 -300 11574 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 11886 -300 11942 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 12254 -300 12310 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 12622 -300 12678 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 12990 -300 13046 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 13358 -300 13414 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 8206 -300 8262 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 8574 -300 8630 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 8942 -300 8998 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 9310 -300 9366 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 9678 -300 9734 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 10046 -300 10102 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 10414 -300 10470 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 10782 -300 10838 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 11150 -300 11206 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 13726 -300 13782 160 0 FreeSans 224 90 0 0 NN4END[0]
port 76 nsew signal input
flabel metal2 s 17406 -300 17462 160 0 FreeSans 224 90 0 0 NN4END[10]
port 77 nsew signal input
flabel metal2 s 17774 -300 17830 160 0 FreeSans 224 90 0 0 NN4END[11]
port 78 nsew signal input
flabel metal2 s 18142 -300 18198 160 0 FreeSans 224 90 0 0 NN4END[12]
port 79 nsew signal input
flabel metal2 s 18510 -300 18566 160 0 FreeSans 224 90 0 0 NN4END[13]
port 80 nsew signal input
flabel metal2 s 18878 -300 18934 160 0 FreeSans 224 90 0 0 NN4END[14]
port 81 nsew signal input
flabel metal2 s 19246 -300 19302 160 0 FreeSans 224 90 0 0 NN4END[15]
port 82 nsew signal input
flabel metal2 s 14094 -300 14150 160 0 FreeSans 224 90 0 0 NN4END[1]
port 83 nsew signal input
flabel metal2 s 14462 -300 14518 160 0 FreeSans 224 90 0 0 NN4END[2]
port 84 nsew signal input
flabel metal2 s 14830 -300 14886 160 0 FreeSans 224 90 0 0 NN4END[3]
port 85 nsew signal input
flabel metal2 s 15198 -300 15254 160 0 FreeSans 224 90 0 0 NN4END[4]
port 86 nsew signal input
flabel metal2 s 15566 -300 15622 160 0 FreeSans 224 90 0 0 NN4END[5]
port 87 nsew signal input
flabel metal2 s 15934 -300 15990 160 0 FreeSans 224 90 0 0 NN4END[6]
port 88 nsew signal input
flabel metal2 s 16302 -300 16358 160 0 FreeSans 224 90 0 0 NN4END[7]
port 89 nsew signal input
flabel metal2 s 16670 -300 16726 160 0 FreeSans 224 90 0 0 NN4END[8]
port 90 nsew signal input
flabel metal2 s 17038 -300 17094 160 0 FreeSans 224 90 0 0 NN4END[9]
port 91 nsew signal input
flabel metal2 s 19614 -300 19670 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 92 nsew signal tristate
flabel metal2 s 19982 -300 20038 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 93 nsew signal tristate
flabel metal2 s 20350 -300 20406 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 94 nsew signal tristate
flabel metal2 s 20718 -300 20774 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 95 nsew signal tristate
flabel metal2 s 24030 -300 24086 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 96 nsew signal tristate
flabel metal2 s 24398 -300 24454 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 97 nsew signal tristate
flabel metal2 s 24766 -300 24822 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 98 nsew signal tristate
flabel metal2 s 25134 -300 25190 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 99 nsew signal tristate
flabel metal2 s 25502 -300 25558 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 100 nsew signal tristate
flabel metal2 s 25870 -300 25926 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 101 nsew signal tristate
flabel metal2 s 26238 -300 26294 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 102 nsew signal tristate
flabel metal2 s 26606 -300 26662 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 103 nsew signal tristate
flabel metal2 s 21086 -300 21142 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 104 nsew signal tristate
flabel metal2 s 21454 -300 21510 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 105 nsew signal tristate
flabel metal2 s 21822 -300 21878 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 106 nsew signal tristate
flabel metal2 s 22190 -300 22246 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 107 nsew signal tristate
flabel metal2 s 22558 -300 22614 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 108 nsew signal tristate
flabel metal2 s 22926 -300 22982 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 109 nsew signal tristate
flabel metal2 s 23294 -300 23350 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 110 nsew signal tristate
flabel metal2 s 23662 -300 23718 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 111 nsew signal tristate
flabel metal2 s 26974 -300 27030 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 112 nsew signal tristate
flabel metal2 s 30654 -300 30710 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 113 nsew signal tristate
flabel metal2 s 31022 -300 31078 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 114 nsew signal tristate
flabel metal2 s 31390 -300 31446 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 115 nsew signal tristate
flabel metal2 s 31758 -300 31814 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 116 nsew signal tristate
flabel metal2 s 32126 -300 32182 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 117 nsew signal tristate
flabel metal2 s 32494 -300 32550 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 118 nsew signal tristate
flabel metal2 s 27342 -300 27398 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 119 nsew signal tristate
flabel metal2 s 27710 -300 27766 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 120 nsew signal tristate
flabel metal2 s 28078 -300 28134 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 121 nsew signal tristate
flabel metal2 s 28446 -300 28502 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 122 nsew signal tristate
flabel metal2 s 28814 -300 28870 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 123 nsew signal tristate
flabel metal2 s 29182 -300 29238 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 124 nsew signal tristate
flabel metal2 s 29550 -300 29606 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 125 nsew signal tristate
flabel metal2 s 29918 -300 29974 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 126 nsew signal tristate
flabel metal2 s 30286 -300 30342 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 127 nsew signal tristate
flabel metal2 s 32862 -300 32918 160 0 FreeSans 224 90 0 0 SS4BEG[0]
port 128 nsew signal tristate
flabel metal2 s 36542 -300 36598 160 0 FreeSans 224 90 0 0 SS4BEG[10]
port 129 nsew signal tristate
flabel metal2 s 36910 -300 36966 160 0 FreeSans 224 90 0 0 SS4BEG[11]
port 130 nsew signal tristate
flabel metal2 s 37278 -300 37334 160 0 FreeSans 224 90 0 0 SS4BEG[12]
port 131 nsew signal tristate
flabel metal2 s 37646 -300 37702 160 0 FreeSans 224 90 0 0 SS4BEG[13]
port 132 nsew signal tristate
flabel metal2 s 38014 -300 38070 160 0 FreeSans 224 90 0 0 SS4BEG[14]
port 133 nsew signal tristate
flabel metal2 s 38382 -300 38438 160 0 FreeSans 224 90 0 0 SS4BEG[15]
port 134 nsew signal tristate
flabel metal2 s 33230 -300 33286 160 0 FreeSans 224 90 0 0 SS4BEG[1]
port 135 nsew signal tristate
flabel metal2 s 33598 -300 33654 160 0 FreeSans 224 90 0 0 SS4BEG[2]
port 136 nsew signal tristate
flabel metal2 s 33966 -300 34022 160 0 FreeSans 224 90 0 0 SS4BEG[3]
port 137 nsew signal tristate
flabel metal2 s 34334 -300 34390 160 0 FreeSans 224 90 0 0 SS4BEG[4]
port 138 nsew signal tristate
flabel metal2 s 34702 -300 34758 160 0 FreeSans 224 90 0 0 SS4BEG[5]
port 139 nsew signal tristate
flabel metal2 s 35070 -300 35126 160 0 FreeSans 224 90 0 0 SS4BEG[6]
port 140 nsew signal tristate
flabel metal2 s 35438 -300 35494 160 0 FreeSans 224 90 0 0 SS4BEG[7]
port 141 nsew signal tristate
flabel metal2 s 35806 -300 35862 160 0 FreeSans 224 90 0 0 SS4BEG[8]
port 142 nsew signal tristate
flabel metal2 s 36174 -300 36230 160 0 FreeSans 224 90 0 0 SS4BEG[9]
port 143 nsew signal tristate
flabel metal2 s 38750 -300 38806 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 1214 9840 1270 10300 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6498 1040 6818 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 17606 1040 17926 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 28714 1040 29034 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 39822 1040 40142 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 12052 1040 12372 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 23160 1040 23480 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 34268 1040 34588 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 45376 1040 45696 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 23322 8160 23322 8160 0 vccd1
rlabel via1 23400 8704 23400 8704 0 vssd1
rlabel metal2 39146 670 39146 670 0 FrameStrobe[0]
rlabel metal2 42826 670 42826 670 0 FrameStrobe[10]
rlabel metal2 43194 670 43194 670 0 FrameStrobe[11]
rlabel metal2 43562 670 43562 670 0 FrameStrobe[12]
rlabel metal2 44075 68 44075 68 0 FrameStrobe[13]
rlabel metal2 44298 143 44298 143 0 FrameStrobe[14]
rlabel metal2 44719 68 44719 68 0 FrameStrobe[15]
rlabel metal2 44935 68 44935 68 0 FrameStrobe[16]
rlabel metal2 45257 68 45257 68 0 FrameStrobe[17]
rlabel metal2 45770 1010 45770 1010 0 FrameStrobe[18]
rlabel metal2 46138 1248 46138 1248 0 FrameStrobe[19]
rlabel metal2 39514 551 39514 551 0 FrameStrobe[1]
rlabel metal2 39882 755 39882 755 0 FrameStrobe[2]
rlabel metal2 40395 68 40395 68 0 FrameStrobe[3]
rlabel metal2 40618 534 40618 534 0 FrameStrobe[4]
rlabel metal2 41131 68 41131 68 0 FrameStrobe[5]
rlabel metal2 41354 670 41354 670 0 FrameStrobe[6]
rlabel metal2 41722 670 41722 670 0 FrameStrobe[7]
rlabel metal2 42235 68 42235 68 0 FrameStrobe[8]
rlabel metal2 42603 68 42603 68 0 FrameStrobe[9]
rlabel metal1 3680 8602 3680 8602 0 FrameStrobe_O[0]
rlabel metal1 25622 8602 25622 8602 0 FrameStrobe_O[10]
rlabel metal2 27738 9224 27738 9224 0 FrameStrobe_O[11]
rlabel metal1 30038 8602 30038 8602 0 FrameStrobe_O[12]
rlabel metal1 32246 8602 32246 8602 0 FrameStrobe_O[13]
rlabel metal2 34362 9445 34362 9445 0 FrameStrobe_O[14]
rlabel metal1 36662 8602 36662 8602 0 FrameStrobe_O[15]
rlabel metal2 38778 9224 38778 9224 0 FrameStrobe_O[16]
rlabel metal1 41078 8602 41078 8602 0 FrameStrobe_O[17]
rlabel metal1 43286 8602 43286 8602 0 FrameStrobe_O[18]
rlabel metal1 45034 8602 45034 8602 0 FrameStrobe_O[19]
rlabel metal2 5658 9224 5658 9224 0 FrameStrobe_O[1]
rlabel metal1 7958 8602 7958 8602 0 FrameStrobe_O[2]
rlabel metal1 10166 8602 10166 8602 0 FrameStrobe_O[3]
rlabel metal2 12282 9785 12282 9785 0 FrameStrobe_O[4]
rlabel metal1 14582 8602 14582 8602 0 FrameStrobe_O[5]
rlabel metal2 16698 9190 16698 9190 0 FrameStrobe_O[6]
rlabel metal2 18906 9224 18906 9224 0 FrameStrobe_O[7]
rlabel metal1 21206 8602 21206 8602 0 FrameStrobe_O[8]
rlabel metal2 23322 9785 23322 9785 0 FrameStrobe_O[9]
rlabel metal1 23920 2074 23920 2074 0 FrameStrobe_O_i\[0\]
rlabel metal1 26726 2074 26726 2074 0 FrameStrobe_O_i\[10\]
rlabel metal1 28796 2414 28796 2414 0 FrameStrobe_O_i\[11\]
rlabel metal2 32154 2278 32154 2278 0 FrameStrobe_O_i\[12\]
rlabel metal1 33028 2074 33028 2074 0 FrameStrobe_O_i\[13\]
rlabel metal1 35098 2074 35098 2074 0 FrameStrobe_O_i\[14\]
rlabel metal1 37306 2074 37306 2074 0 FrameStrobe_O_i\[15\]
rlabel metal1 39514 2074 39514 2074 0 FrameStrobe_O_i\[16\]
rlabel metal1 41676 2074 41676 2074 0 FrameStrobe_O_i\[17\]
rlabel metal1 44206 2074 44206 2074 0 FrameStrobe_O_i\[18\]
rlabel metal1 44528 1802 44528 1802 0 FrameStrobe_O_i\[19\]
rlabel metal1 21666 1768 21666 1768 0 FrameStrobe_O_i\[1\]
rlabel metal1 23506 2448 23506 2448 0 FrameStrobe_O_i\[2\]
rlabel metal1 23506 2040 23506 2040 0 FrameStrobe_O_i\[3\]
rlabel metal1 22586 2346 22586 2346 0 FrameStrobe_O_i\[4\]
rlabel metal1 20976 2414 20976 2414 0 FrameStrobe_O_i\[5\]
rlabel metal1 17434 1462 17434 1462 0 FrameStrobe_O_i\[6\]
rlabel metal1 18952 2074 18952 2074 0 FrameStrobe_O_i\[7\]
rlabel metal1 20838 1802 20838 1802 0 FrameStrobe_O_i\[8\]
rlabel metal1 24564 2074 24564 2074 0 FrameStrobe_O_i\[9\]
rlabel metal2 506 1010 506 1010 0 N1END[0]
rlabel metal2 874 976 874 976 0 N1END[1]
rlabel metal2 1242 704 1242 704 0 N1END[2]
rlabel metal2 1663 68 1663 68 0 N1END[3]
rlabel metal2 4975 68 4975 68 0 N2END[0]
rlabel metal2 5343 68 5343 68 0 N2END[1]
rlabel metal2 5711 68 5711 68 0 N2END[2]
rlabel metal2 6026 704 6026 704 0 N2END[3]
rlabel metal2 6447 68 6447 68 0 N2END[4]
rlabel metal2 6815 68 6815 68 0 N2END[5]
rlabel metal2 7183 68 7183 68 0 N2END[6]
rlabel metal2 7551 68 7551 68 0 N2END[7]
rlabel metal2 2031 68 2031 68 0 N2MID[0]
rlabel metal2 2399 68 2399 68 0 N2MID[1]
rlabel metal2 2615 68 2615 68 0 N2MID[2]
rlabel metal2 3135 68 3135 68 0 N2MID[3]
rlabel metal2 3450 704 3450 704 0 N2MID[4]
rlabel metal2 3871 68 3871 68 0 N2MID[5]
rlabel metal2 4239 68 4239 68 0 N2MID[6]
rlabel metal2 4607 68 4607 68 0 N2MID[7]
rlabel metal2 7919 68 7919 68 0 N4END[0]
rlabel metal2 11599 68 11599 68 0 N4END[10]
rlabel metal2 11967 68 11967 68 0 N4END[11]
rlabel metal2 12335 68 12335 68 0 N4END[12]
rlabel metal2 12650 704 12650 704 0 N4END[13]
rlabel metal2 12965 68 12965 68 0 N4END[14]
rlabel metal2 13287 68 13287 68 0 N4END[15]
rlabel metal2 8287 68 8287 68 0 N4END[1]
rlabel metal2 8602 704 8602 704 0 N4END[2]
rlabel metal2 9023 68 9023 68 0 N4END[3]
rlabel metal2 9391 68 9391 68 0 N4END[4]
rlabel metal2 9759 68 9759 68 0 N4END[5]
rlabel metal2 10127 68 10127 68 0 N4END[6]
rlabel metal2 10495 68 10495 68 0 N4END[7]
rlabel metal2 10863 68 10863 68 0 N4END[8]
rlabel metal2 11178 704 11178 704 0 N4END[9]
rlabel metal2 13754 143 13754 143 0 NN4END[0]
rlabel metal2 17434 432 17434 432 0 NN4END[10]
rlabel metal2 17802 143 17802 143 0 NN4END[11]
rlabel metal2 18223 68 18223 68 0 NN4END[12]
rlabel metal2 18538 704 18538 704 0 NN4END[13]
rlabel metal2 18853 68 18853 68 0 NN4END[14]
rlabel metal2 19274 704 19274 704 0 NN4END[15]
rlabel metal2 14122 143 14122 143 0 NN4END[1]
rlabel metal2 14490 670 14490 670 0 NN4END[2]
rlabel metal2 14713 68 14713 68 0 NN4END[3]
rlabel metal2 15226 415 15226 415 0 NN4END[4]
rlabel metal2 15449 68 15449 68 0 NN4END[5]
rlabel metal2 15817 68 15817 68 0 NN4END[6]
rlabel metal2 16330 143 16330 143 0 NN4END[7]
rlabel metal2 16553 68 16553 68 0 NN4END[8]
rlabel metal2 17066 143 17066 143 0 NN4END[9]
rlabel metal2 19642 636 19642 636 0 S1BEG[0]
rlabel metal2 20063 68 20063 68 0 S1BEG[1]
rlabel metal2 20378 636 20378 636 0 S1BEG[2]
rlabel metal2 20746 636 20746 636 0 S1BEG[3]
rlabel metal2 24111 68 24111 68 0 S2BEG[0]
rlabel metal2 24571 68 24571 68 0 S2BEG[1]
rlabel metal2 24794 806 24794 806 0 S2BEG[2]
rlabel metal2 25162 636 25162 636 0 S2BEG[3]
rlabel metal2 25530 636 25530 636 0 S2BEG[4]
rlabel metal2 26043 68 26043 68 0 S2BEG[5]
rlabel metal2 26365 68 26365 68 0 S2BEG[6]
rlabel metal2 26634 636 26634 636 0 S2BEG[7]
rlabel metal2 21167 68 21167 68 0 S2BEGb[0]
rlabel metal2 21482 636 21482 636 0 S2BEGb[1]
rlabel metal2 21850 908 21850 908 0 S2BEGb[2]
rlabel metal2 22363 68 22363 68 0 S2BEGb[3]
rlabel metal2 22586 908 22586 908 0 S2BEGb[4]
rlabel metal2 23007 68 23007 68 0 S2BEGb[5]
rlabel metal2 23322 483 23322 483 0 S2BEGb[6]
rlabel metal2 23743 68 23743 68 0 S2BEGb[7]
rlabel metal2 27002 143 27002 143 0 S4BEG[0]
rlabel metal2 31878 1938 31878 1938 0 S4BEG[10]
rlabel metal2 31195 68 31195 68 0 S4BEG[11]
rlabel metal2 31878 1479 31878 1479 0 S4BEG[12]
rlabel metal2 31786 636 31786 636 0 S4BEG[13]
rlabel metal2 32299 68 32299 68 0 S4BEG[14]
rlabel metal2 32667 68 32667 68 0 S4BEG[15]
rlabel metal2 27370 806 27370 806 0 S4BEG[1]
rlabel metal2 27738 636 27738 636 0 S4BEG[2]
rlabel metal2 28106 908 28106 908 0 S4BEG[3]
rlabel metal2 28474 738 28474 738 0 S4BEG[4]
rlabel metal2 28842 806 28842 806 0 S4BEG[5]
rlabel metal2 29157 68 29157 68 0 S4BEG[6]
rlabel metal2 29578 670 29578 670 0 S4BEG[7]
rlabel metal2 29946 806 29946 806 0 S4BEG[8]
rlabel metal2 30314 687 30314 687 0 S4BEG[9]
rlabel metal2 32890 772 32890 772 0 SS4BEG[0]
rlabel metal2 36715 68 36715 68 0 SS4BEG[10]
rlabel metal2 37083 68 37083 68 0 SS4BEG[11]
rlabel metal2 37451 68 37451 68 0 SS4BEG[12]
rlabel metal2 37674 942 37674 942 0 SS4BEG[13]
rlabel metal2 38042 143 38042 143 0 SS4BEG[14]
rlabel metal2 38410 772 38410 772 0 SS4BEG[15]
rlabel metal2 33258 942 33258 942 0 SS4BEG[1]
rlabel metal2 33771 68 33771 68 0 SS4BEG[2]
rlabel metal2 34093 68 34093 68 0 SS4BEG[3]
rlabel metal2 34415 68 34415 68 0 SS4BEG[4]
rlabel metal2 34875 68 34875 68 0 SS4BEG[5]
rlabel metal2 35243 68 35243 68 0 SS4BEG[6]
rlabel metal1 36570 1496 36570 1496 0 SS4BEG[7]
rlabel metal2 35834 738 35834 738 0 SS4BEG[8]
rlabel metal2 36347 68 36347 68 0 SS4BEG[9]
rlabel metal2 38778 704 38778 704 0 UserCLK
rlabel metal2 1242 9445 1242 9445 0 UserCLKo
rlabel metal1 39836 1530 39836 1530 0 net1
rlabel metal1 44574 1904 44574 1904 0 net10
rlabel metal2 24978 1530 24978 1530 0 net100
rlabel metal1 25116 1326 25116 1326 0 net101
rlabel metal1 25806 1360 25806 1360 0 net102
rlabel metal1 25990 1904 25990 1904 0 net103
rlabel metal1 26634 1326 26634 1326 0 net104
rlabel metal1 26910 1326 26910 1326 0 net105
rlabel metal1 20976 1938 20976 1938 0 net106
rlabel metal1 21022 1326 21022 1326 0 net107
rlabel metal1 22034 2040 22034 2040 0 net108
rlabel via1 20930 1275 20930 1275 0 net109
rlabel metal1 44942 1938 44942 1938 0 net11
rlabel metal1 22172 2822 22172 2822 0 net110
rlabel metal1 22034 1394 22034 1394 0 net111
rlabel metal1 23230 1258 23230 1258 0 net112
rlabel metal1 23322 2890 23322 2890 0 net113
rlabel metal1 27278 1326 27278 1326 0 net114
rlabel metal1 31372 1938 31372 1938 0 net115
rlabel metal1 31188 2006 31188 2006 0 net116
rlabel metal1 32108 1326 32108 1326 0 net117
rlabel metal1 32706 1292 32706 1292 0 net118
rlabel metal2 30314 2686 30314 2686 0 net119
rlabel metal2 40158 2295 40158 2295 0 net12
rlabel metal1 33350 272 33350 272 0 net120
rlabel metal1 27784 1326 27784 1326 0 net121
rlabel metal1 28152 1326 28152 1326 0 net122
rlabel metal1 28428 1938 28428 1938 0 net123
rlabel metal2 29210 1530 29210 1530 0 net124
rlabel metal1 29486 1326 29486 1326 0 net125
rlabel metal1 29900 1938 29900 1938 0 net126
rlabel metal1 30590 1326 30590 1326 0 net127
rlabel metal1 30866 1326 30866 1326 0 net128
rlabel metal1 31280 1326 31280 1326 0 net129
rlabel metal2 40434 2312 40434 2312 0 net13
rlabel metal1 18998 1768 18998 1768 0 net130
rlabel metal1 37904 1258 37904 1258 0 net131
rlabel metal1 38318 1258 38318 1258 0 net132
rlabel metal2 38042 1887 38042 1887 0 net133
rlabel via2 38410 1955 38410 1955 0 net134
rlabel metal1 38824 1258 38824 1258 0 net135
rlabel metal1 39974 1224 39974 1224 0 net136
rlabel metal1 31878 1428 31878 1428 0 net137
rlabel metal1 33672 1938 33672 1938 0 net138
rlabel via2 34822 1275 34822 1275 0 net139
rlabel metal2 40710 2278 40710 2278 0 net14
rlabel metal1 34914 272 34914 272 0 net140
rlabel metal2 35466 2159 35466 2159 0 net141
rlabel metal2 35190 2193 35190 2193 0 net142
rlabel metal2 35466 1122 35466 1122 0 net143
rlabel metal1 37444 1258 37444 1258 0 net144
rlabel metal1 36386 2040 36386 2040 0 net145
rlabel metal1 10534 8500 10534 8500 0 net146
rlabel metal2 40066 1088 40066 1088 0 net15
rlabel metal1 42090 714 42090 714 0 net16
rlabel metal2 41170 2754 41170 2754 0 net17
rlabel metal2 42458 2890 42458 2890 0 net18
rlabel metal2 39330 1054 39330 1054 0 net19
rlabel metal1 43102 918 43102 918 0 net2
rlabel metal1 43010 612 43010 612 0 net20
rlabel metal2 1610 1632 1610 1632 0 net21
rlabel metal2 19550 2516 19550 2516 0 net22
rlabel via2 18906 1309 18906 1309 0 net23
rlabel metal2 18814 2465 18814 2465 0 net24
rlabel metal1 22402 2992 22402 2992 0 net25
rlabel metal2 12742 629 12742 629 0 net26
rlabel metal2 20746 2159 20746 2159 0 net27
rlabel metal1 15042 3026 15042 3026 0 net28
rlabel metal1 19734 2448 19734 2448 0 net29
rlabel metal2 43562 1904 43562 1904 0 net3
rlabel metal1 20378 2380 20378 2380 0 net30
rlabel metal2 19550 2142 19550 2142 0 net31
rlabel metal2 18078 2176 18078 2176 0 net32
rlabel metal2 2346 3196 2346 3196 0 net33
rlabel metal1 2714 1292 2714 1292 0 net34
rlabel metal3 14352 4148 14352 4148 0 net35
rlabel metal2 14858 1649 14858 1649 0 net36
rlabel metal1 14950 4522 14950 4522 0 net37
rlabel metal3 17250 4012 17250 4012 0 net38
rlabel metal2 13110 408 13110 408 0 net39
rlabel metal2 43838 1598 43838 1598 0 net4
rlabel metal3 17158 2040 17158 2040 0 net40
rlabel metal1 25530 3536 25530 3536 0 net41
rlabel metal1 12466 1360 12466 1360 0 net42
rlabel metal1 13570 1292 13570 1292 0 net43
rlabel metal2 12558 748 12558 748 0 net44
rlabel metal1 24978 884 24978 884 0 net45
rlabel metal2 25806 1292 25806 1292 0 net46
rlabel metal2 13294 714 13294 714 0 net47
rlabel metal1 17250 680 17250 680 0 net48
rlabel metal2 8786 1037 8786 1037 0 net49
rlabel metal2 44114 782 44114 782 0 net5
rlabel metal2 9246 901 9246 901 0 net50
rlabel metal2 9614 833 9614 833 0 net51
rlabel metal1 17158 612 17158 612 0 net52
rlabel metal2 10350 765 10350 765 0 net53
rlabel metal2 10718 969 10718 969 0 net54
rlabel metal2 28382 1292 28382 1292 0 net55
rlabel metal2 11362 1088 11362 1088 0 net56
rlabel metal1 22770 2958 22770 2958 0 net57
rlabel metal1 17066 1530 17066 1530 0 net58
rlabel metal1 17388 1530 17388 1530 0 net59
rlabel metal1 44298 1462 44298 1462 0 net6
rlabel metal1 17802 1530 17802 1530 0 net60
rlabel metal1 18262 1530 18262 1530 0 net61
rlabel metal1 18538 1530 18538 1530 0 net62
rlabel metal1 18860 1530 18860 1530 0 net63
rlabel metal2 13938 782 13938 782 0 net64
rlabel metal1 14812 1462 14812 1462 0 net65
rlabel metal1 14812 1530 14812 1530 0 net66
rlabel metal1 15778 1292 15778 1292 0 net67
rlabel metal2 15134 1700 15134 1700 0 net68
rlabel metal1 15732 1530 15732 1530 0 net69
rlabel metal1 45034 1428 45034 1428 0 net7
rlabel metal1 16008 1462 16008 1462 0 net70
rlabel metal1 17066 1292 17066 1292 0 net71
rlabel metal2 16514 1734 16514 1734 0 net72
rlabel metal2 39422 986 39422 986 0 net73
rlabel metal2 4094 8636 4094 8636 0 net74
rlabel metal1 25944 2618 25944 2618 0 net75
rlabel metal1 28152 2618 28152 2618 0 net76
rlabel metal1 30360 8466 30360 8466 0 net77
rlabel metal1 32568 2618 32568 2618 0 net78
rlabel metal2 34822 5542 34822 5542 0 net79
rlabel metal1 43608 1530 43608 1530 0 net8
rlabel metal1 36984 2618 36984 2618 0 net80
rlabel metal1 39100 2618 39100 2618 0 net81
rlabel metal2 41354 5542 41354 5542 0 net82
rlabel metal1 43700 2618 43700 2618 0 net83
rlabel metal2 44574 5542 44574 5542 0 net84
rlabel metal1 22908 3502 22908 3502 0 net85
rlabel metal2 8234 8670 8234 8670 0 net86
rlabel metal2 24426 5474 24426 5474 0 net87
rlabel metal1 14582 8534 14582 8534 0 net88
rlabel metal1 18814 8534 18814 8534 0 net89
rlabel metal1 41998 1972 41998 1972 0 net9
rlabel metal2 17066 5542 17066 5542 0 net90
rlabel metal1 19458 2618 19458 2618 0 net91
rlabel metal1 21528 2618 21528 2618 0 net92
rlabel metal1 23782 2550 23782 2550 0 net93
rlabel metal1 19458 1326 19458 1326 0 net94
rlabel metal1 19918 1292 19918 1292 0 net95
rlabel metal1 20148 1326 20148 1326 0 net96
rlabel metal1 20470 1258 20470 1258 0 net97
rlabel metal1 22310 1224 22310 1224 0 net98
rlabel metal1 24288 1326 24288 1326 0 net99
<< properties >>
string FIXED_BBOX 0 0 46700 10000
<< end >>
