magic
tech sky130A
magscale 1 2
timestamp 1733619042
<< viali >>
rect 2237 8585 2271 8619
rect 3433 8585 3467 8619
rect 4629 8585 4663 8619
rect 5917 8585 5951 8619
rect 7113 8585 7147 8619
rect 8309 8585 8343 8619
rect 9505 8585 9539 8619
rect 10701 8585 10735 8619
rect 11897 8585 11931 8619
rect 13093 8585 13127 8619
rect 14289 8585 14323 8619
rect 15485 8585 15519 8619
rect 17233 8585 17267 8619
rect 17785 8585 17819 8619
rect 19441 8585 19475 8619
rect 20177 8585 20211 8619
rect 21373 8585 21407 8619
rect 22569 8585 22603 8619
rect 23857 8585 23891 8619
rect 1409 8517 1443 8551
rect 16681 8517 16715 8551
rect 17049 8517 17083 8551
rect 1777 8449 1811 8483
rect 2421 8449 2455 8483
rect 3617 8449 3651 8483
rect 4813 8449 4847 8483
rect 5825 8449 5859 8483
rect 7021 8449 7055 8483
rect 8217 8449 8251 8483
rect 9321 8449 9355 8483
rect 10517 8449 10551 8483
rect 11713 8449 11747 8483
rect 12909 8449 12943 8483
rect 14105 8449 14139 8483
rect 15393 8449 15427 8483
rect 17417 8449 17451 8483
rect 17969 8449 18003 8483
rect 19349 8449 19383 8483
rect 20361 8449 20395 8483
rect 21557 8449 21591 8483
rect 22753 8449 22787 8483
rect 23489 8449 23523 8483
rect 23765 8449 23799 8483
rect 23213 8381 23247 8415
rect 16773 8041 16807 8075
rect 16589 7837 16623 7871
rect 9505 4097 9539 4131
rect 10701 4097 10735 4131
rect 11897 4097 11931 4131
rect 13093 4097 13127 4131
rect 19993 4097 20027 4131
rect 24041 4097 24075 4131
rect 19809 3961 19843 3995
rect 9321 3893 9355 3927
rect 10517 3893 10551 3927
rect 11713 3893 11747 3927
rect 12909 3893 12943 3927
rect 23857 3893 23891 3927
rect 9505 3689 9539 3723
rect 10609 3689 10643 3723
rect 11805 3689 11839 3723
rect 13001 3689 13035 3723
rect 14105 3689 14139 3723
rect 15301 3689 15335 3723
rect 19993 3689 20027 3723
rect 24041 3689 24075 3723
rect 23581 3621 23615 3655
rect 9689 3485 9723 3519
rect 10793 3485 10827 3519
rect 11989 3485 12023 3519
rect 13185 3485 13219 3519
rect 14289 3485 14323 3519
rect 14565 3485 14599 3519
rect 15485 3485 15519 3519
rect 20177 3485 20211 3519
rect 23489 3485 23523 3519
rect 23765 3485 23799 3519
rect 23857 3485 23891 3519
rect 14381 3349 14415 3383
rect 23305 3349 23339 3383
rect 8125 3145 8159 3179
rect 15393 3145 15427 3179
rect 22753 3145 22787 3179
rect 23213 3145 23247 3179
rect 8309 3009 8343 3043
rect 15577 3009 15611 3043
rect 22661 3009 22695 3043
rect 22937 3009 22971 3043
rect 23029 3009 23063 3043
rect 23305 3009 23339 3043
rect 23765 3009 23799 3043
rect 24041 3009 24075 3043
rect 22477 2873 22511 2907
rect 23489 2805 23523 2839
rect 23581 2805 23615 2839
rect 23857 2805 23891 2839
rect 1869 2601 1903 2635
rect 2145 2601 2179 2635
rect 8217 2601 8251 2635
rect 19257 2601 19291 2635
rect 23029 2601 23063 2635
rect 23673 2601 23707 2635
rect 1593 2533 1627 2567
rect 16957 2533 16991 2567
rect 17509 2533 17543 2567
rect 22201 2533 22235 2567
rect 22753 2533 22787 2567
rect 23949 2533 23983 2567
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 1961 2397 1995 2431
rect 8401 2397 8435 2431
rect 10701 2397 10735 2431
rect 11345 2397 11379 2431
rect 11713 2397 11747 2431
rect 12265 2397 12299 2431
rect 12541 2397 12575 2431
rect 14933 2397 14967 2431
rect 16129 2397 16163 2431
rect 16773 2397 16807 2431
rect 17049 2397 17083 2431
rect 17325 2397 17359 2431
rect 17785 2397 17819 2431
rect 18061 2397 18095 2431
rect 18429 2397 18463 2431
rect 19441 2397 19475 2431
rect 19993 2397 20027 2431
rect 22017 2397 22051 2431
rect 22477 2397 22511 2431
rect 22569 2397 22603 2431
rect 22845 2397 22879 2431
rect 23305 2397 23339 2431
rect 23397 2397 23431 2431
rect 23857 2397 23891 2431
rect 24133 2397 24167 2431
rect 19625 2329 19659 2363
rect 19809 2329 19843 2363
rect 10885 2261 10919 2295
rect 11529 2261 11563 2295
rect 11897 2261 11931 2295
rect 12449 2261 12483 2295
rect 12725 2261 12759 2295
rect 15117 2261 15151 2295
rect 16313 2261 16347 2295
rect 17233 2261 17267 2295
rect 17969 2261 18003 2295
rect 18245 2261 18279 2295
rect 18613 2261 18647 2295
rect 20177 2261 20211 2295
rect 22293 2261 22327 2295
rect 23121 2261 23155 2295
rect 23581 2261 23615 2295
rect 1777 2057 1811 2091
rect 2053 2057 2087 2091
rect 5365 2057 5399 2091
rect 5917 2057 5951 2091
rect 6837 2057 6871 2091
rect 7113 2057 7147 2091
rect 9781 2057 9815 2091
rect 10057 2057 10091 2091
rect 14473 2057 14507 2091
rect 15025 2057 15059 2091
rect 20913 2057 20947 2091
rect 21465 2057 21499 2091
rect 21833 2057 21867 2091
rect 22385 2057 22419 2091
rect 22661 2057 22695 2091
rect 22937 2057 22971 2091
rect 23213 2057 23247 2091
rect 23489 2057 23523 2091
rect 24041 2057 24075 2091
rect 10223 1989 10257 2023
rect 10977 1989 11011 2023
rect 11897 1989 11931 2023
rect 15485 1989 15519 2023
rect 16773 1989 16807 2023
rect 18245 1989 18279 2023
rect 18797 1989 18831 2023
rect 19349 1989 19383 2023
rect 20453 1989 20487 2023
rect 1593 1921 1627 1955
rect 1869 1921 1903 1955
rect 2145 1921 2179 1955
rect 2421 1921 2455 1955
rect 5181 1921 5215 1955
rect 5457 1921 5491 1955
rect 5733 1921 5767 1955
rect 6009 1921 6043 1955
rect 6653 1921 6687 1955
rect 6929 1921 6963 1955
rect 7573 1921 7607 1955
rect 7665 1921 7699 1955
rect 8125 1921 8159 1955
rect 8493 1921 8527 1955
rect 8769 1921 8803 1955
rect 9229 1921 9263 1955
rect 9321 1921 9355 1955
rect 9605 1921 9639 1955
rect 9873 1921 9907 1955
rect 11529 1921 11563 1955
rect 12449 1921 12483 1955
rect 12725 1921 12759 1955
rect 13185 1921 13219 1955
rect 13461 1921 13495 1955
rect 13737 1921 13771 1955
rect 14013 1921 14047 1955
rect 14289 1921 14323 1955
rect 14565 1921 14599 1955
rect 14841 1921 14875 1955
rect 15945 1921 15979 1955
rect 16313 1921 16347 1955
rect 17233 1921 17267 1955
rect 17693 1921 17727 1955
rect 20177 1921 20211 1955
rect 21097 1921 21131 1955
rect 21373 1921 21407 1955
rect 21649 1921 21683 1955
rect 22017 1921 22051 1955
rect 22293 1921 22327 1955
rect 22569 1921 22603 1955
rect 22845 1921 22879 1955
rect 23121 1921 23155 1955
rect 23397 1921 23431 1955
rect 23673 1921 23707 1955
rect 23949 1921 23983 1955
rect 24225 1921 24259 1955
rect 2605 1785 2639 1819
rect 5641 1785 5675 1819
rect 6193 1785 6227 1819
rect 9505 1785 9539 1819
rect 13921 1785 13955 1819
rect 14197 1785 14231 1819
rect 21189 1785 21223 1819
rect 22109 1785 22143 1819
rect 23765 1785 23799 1819
rect 2329 1717 2363 1751
rect 7389 1717 7423 1751
rect 7849 1717 7883 1751
rect 8309 1717 8343 1751
rect 8677 1717 8711 1751
rect 8953 1717 8987 1751
rect 9045 1717 9079 1751
rect 10333 1717 10367 1751
rect 11069 1717 11103 1751
rect 11713 1717 11747 1751
rect 11989 1717 12023 1751
rect 12633 1717 12667 1751
rect 12909 1717 12943 1751
rect 13369 1717 13403 1751
rect 13645 1717 13679 1751
rect 14749 1717 14783 1751
rect 15577 1717 15611 1751
rect 16865 1717 16899 1751
rect 17417 1717 17451 1751
rect 17969 1717 18003 1751
rect 18337 1717 18371 1751
rect 18889 1717 18923 1751
rect 19441 1717 19475 1751
rect 19901 1717 19935 1751
rect 20545 1717 20579 1751
rect 3065 1513 3099 1547
rect 5089 1513 5123 1547
rect 7389 1513 7423 1547
rect 14657 1513 14691 1547
rect 15393 1513 15427 1547
rect 15945 1513 15979 1547
rect 16313 1513 16347 1547
rect 18521 1513 18555 1547
rect 19993 1513 20027 1547
rect 20545 1513 20579 1547
rect 21833 1513 21867 1547
rect 22661 1513 22695 1547
rect 23489 1513 23523 1547
rect 3341 1445 3375 1479
rect 9505 1445 9539 1479
rect 17509 1445 17543 1479
rect 21281 1445 21315 1479
rect 11069 1377 11103 1411
rect 19625 1377 19659 1411
rect 1501 1309 1535 1343
rect 1777 1309 1811 1343
rect 2053 1309 2087 1343
rect 2329 1309 2363 1343
rect 2605 1309 2639 1343
rect 2881 1309 2915 1343
rect 3157 1309 3191 1343
rect 3433 1309 3467 1343
rect 3801 1309 3835 1343
rect 4077 1309 4111 1343
rect 4353 1309 4387 1343
rect 4629 1309 4663 1343
rect 4905 1309 4939 1343
rect 5181 1309 5215 1343
rect 5457 1309 5491 1343
rect 5733 1309 5767 1343
rect 6009 1309 6043 1343
rect 6377 1309 6411 1343
rect 6653 1309 6687 1343
rect 6929 1309 6963 1343
rect 7205 1309 7239 1343
rect 7481 1309 7515 1343
rect 7757 1309 7791 1343
rect 8033 1309 8067 1343
rect 8309 1309 8343 1343
rect 8585 1309 8619 1343
rect 9045 1309 9079 1343
rect 9321 1309 9355 1343
rect 9597 1309 9631 1343
rect 9965 1309 9999 1343
rect 10333 1309 10367 1343
rect 11621 1309 11655 1343
rect 11989 1309 12023 1343
rect 13093 1309 13127 1343
rect 13461 1309 13495 1343
rect 14105 1309 14139 1343
rect 15301 1309 15335 1343
rect 15853 1309 15887 1343
rect 16497 1309 16531 1343
rect 16773 1309 16807 1343
rect 18429 1309 18463 1343
rect 18889 1309 18923 1343
rect 21189 1309 21223 1343
rect 21465 1309 21499 1343
rect 22017 1309 22051 1343
rect 22293 1309 22327 1343
rect 22569 1309 22603 1343
rect 22845 1309 22879 1343
rect 23121 1309 23155 1343
rect 23397 1309 23431 1343
rect 23673 1309 23707 1343
rect 23949 1309 23983 1343
rect 24225 1309 24259 1343
rect 10793 1241 10827 1275
rect 12449 1241 12483 1275
rect 14565 1241 14599 1275
rect 17325 1241 17359 1275
rect 17877 1241 17911 1275
rect 19349 1241 19383 1275
rect 19901 1241 19935 1275
rect 20453 1241 20487 1275
rect 1685 1173 1719 1207
rect 1961 1173 1995 1207
rect 2237 1173 2271 1207
rect 2513 1173 2547 1207
rect 2789 1173 2823 1207
rect 3617 1173 3651 1207
rect 3985 1173 4019 1207
rect 4261 1173 4295 1207
rect 4537 1173 4571 1207
rect 4813 1173 4847 1207
rect 5365 1173 5399 1207
rect 5641 1173 5675 1207
rect 5917 1173 5951 1207
rect 6193 1173 6227 1207
rect 6561 1173 6595 1207
rect 6837 1173 6871 1207
rect 7113 1173 7147 1207
rect 7665 1173 7699 1207
rect 7941 1173 7975 1207
rect 8217 1173 8251 1207
rect 8493 1173 8527 1207
rect 8769 1173 8803 1207
rect 9229 1173 9263 1207
rect 9781 1173 9815 1207
rect 10149 1173 10183 1207
rect 10517 1173 10551 1207
rect 11805 1173 11839 1207
rect 12173 1173 12207 1207
rect 12541 1173 12575 1207
rect 13277 1173 13311 1207
rect 13645 1173 13679 1207
rect 14289 1173 14323 1207
rect 16865 1173 16899 1207
rect 17969 1173 18003 1207
rect 19073 1173 19107 1207
rect 21005 1173 21039 1207
rect 22109 1173 22143 1207
rect 22385 1173 22419 1207
rect 22937 1173 22971 1207
rect 23213 1173 23247 1207
rect 23765 1173 23799 1207
rect 24041 1173 24075 1207
<< metal1 >>
rect 1104 8730 24723 8752
rect 1104 8678 6814 8730
rect 6866 8678 6878 8730
rect 6930 8678 6942 8730
rect 6994 8678 7006 8730
rect 7058 8678 7070 8730
rect 7122 8678 12679 8730
rect 12731 8678 12743 8730
rect 12795 8678 12807 8730
rect 12859 8678 12871 8730
rect 12923 8678 12935 8730
rect 12987 8678 18544 8730
rect 18596 8678 18608 8730
rect 18660 8678 18672 8730
rect 18724 8678 18736 8730
rect 18788 8678 18800 8730
rect 18852 8678 24409 8730
rect 24461 8678 24473 8730
rect 24525 8678 24537 8730
rect 24589 8678 24601 8730
rect 24653 8678 24665 8730
rect 24717 8678 24723 8730
rect 1104 8656 24723 8678
rect 2038 8576 2044 8628
rect 2096 8616 2102 8628
rect 2225 8619 2283 8625
rect 2225 8616 2237 8619
rect 2096 8588 2237 8616
rect 2096 8576 2102 8588
rect 2225 8585 2237 8588
rect 2271 8585 2283 8619
rect 2225 8579 2283 8585
rect 3234 8576 3240 8628
rect 3292 8616 3298 8628
rect 3421 8619 3479 8625
rect 3421 8616 3433 8619
rect 3292 8588 3433 8616
rect 3292 8576 3298 8588
rect 3421 8585 3433 8588
rect 3467 8585 3479 8619
rect 3421 8579 3479 8585
rect 4430 8576 4436 8628
rect 4488 8616 4494 8628
rect 4617 8619 4675 8625
rect 4617 8616 4629 8619
rect 4488 8588 4629 8616
rect 4488 8576 4494 8588
rect 4617 8585 4629 8588
rect 4663 8585 4675 8619
rect 4617 8579 4675 8585
rect 5626 8576 5632 8628
rect 5684 8616 5690 8628
rect 5905 8619 5963 8625
rect 5905 8616 5917 8619
rect 5684 8588 5917 8616
rect 5684 8576 5690 8588
rect 5905 8585 5917 8588
rect 5951 8585 5963 8619
rect 5905 8579 5963 8585
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 7101 8619 7159 8625
rect 7101 8616 7113 8619
rect 6788 8588 7113 8616
rect 6788 8576 6794 8588
rect 7101 8585 7113 8588
rect 7147 8585 7159 8619
rect 7101 8579 7159 8585
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 8297 8619 8355 8625
rect 8297 8616 8309 8619
rect 8076 8588 8309 8616
rect 8076 8576 8082 8588
rect 8297 8585 8309 8588
rect 8343 8585 8355 8619
rect 8297 8579 8355 8585
rect 9214 8576 9220 8628
rect 9272 8616 9278 8628
rect 9493 8619 9551 8625
rect 9493 8616 9505 8619
rect 9272 8588 9505 8616
rect 9272 8576 9278 8588
rect 9493 8585 9505 8588
rect 9539 8585 9551 8619
rect 9493 8579 9551 8585
rect 10410 8576 10416 8628
rect 10468 8616 10474 8628
rect 10689 8619 10747 8625
rect 10689 8616 10701 8619
rect 10468 8588 10701 8616
rect 10468 8576 10474 8588
rect 10689 8585 10701 8588
rect 10735 8585 10747 8619
rect 10689 8579 10747 8585
rect 11606 8576 11612 8628
rect 11664 8616 11670 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11664 8588 11897 8616
rect 11664 8576 11670 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 13078 8576 13084 8628
rect 13136 8576 13142 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 14056 8588 14289 8616
rect 14056 8576 14062 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 15194 8576 15200 8628
rect 15252 8616 15258 8628
rect 15473 8619 15531 8625
rect 15473 8616 15485 8619
rect 15252 8588 15485 8616
rect 15252 8576 15258 8588
rect 15473 8585 15485 8588
rect 15519 8585 15531 8619
rect 15473 8579 15531 8585
rect 17221 8619 17279 8625
rect 17221 8585 17233 8619
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 1394 8508 1400 8560
rect 1452 8508 1458 8560
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 16669 8551 16727 8557
rect 16669 8548 16681 8551
rect 16448 8520 16681 8548
rect 16448 8508 16454 8520
rect 16669 8517 16681 8520
rect 16715 8517 16727 8551
rect 16669 8511 16727 8517
rect 17037 8551 17095 8557
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 17236 8548 17264 8579
rect 17586 8576 17592 8628
rect 17644 8616 17650 8628
rect 17773 8619 17831 8625
rect 17773 8616 17785 8619
rect 17644 8588 17785 8616
rect 17644 8576 17650 8588
rect 17773 8585 17785 8588
rect 17819 8585 17831 8619
rect 17773 8579 17831 8585
rect 18874 8576 18880 8628
rect 18932 8616 18938 8628
rect 19429 8619 19487 8625
rect 19429 8616 19441 8619
rect 18932 8588 19441 8616
rect 18932 8576 18938 8588
rect 19429 8585 19441 8588
rect 19475 8585 19487 8619
rect 19429 8579 19487 8585
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 20165 8619 20223 8625
rect 20165 8616 20177 8619
rect 20036 8588 20177 8616
rect 20036 8576 20042 8588
rect 20165 8585 20177 8588
rect 20211 8585 20223 8619
rect 20165 8579 20223 8585
rect 21174 8576 21180 8628
rect 21232 8616 21238 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 21232 8588 21373 8616
rect 21232 8576 21238 8588
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 22370 8576 22376 8628
rect 22428 8616 22434 8628
rect 22557 8619 22615 8625
rect 22557 8616 22569 8619
rect 22428 8588 22569 8616
rect 22428 8576 22434 8588
rect 22557 8585 22569 8588
rect 22603 8585 22615 8619
rect 22557 8579 22615 8585
rect 23566 8576 23572 8628
rect 23624 8616 23630 8628
rect 23845 8619 23903 8625
rect 23845 8616 23857 8619
rect 23624 8588 23857 8616
rect 23624 8576 23630 8588
rect 23845 8585 23857 8588
rect 23891 8585 23903 8619
rect 23845 8579 23903 8585
rect 24854 8548 24860 8560
rect 17083 8520 17264 8548
rect 17972 8520 24860 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 1762 8440 1768 8492
rect 1820 8440 1826 8492
rect 2406 8440 2412 8492
rect 2464 8440 2470 8492
rect 3602 8440 3608 8492
rect 3660 8440 3666 8492
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 5810 8440 5816 8492
rect 5868 8440 5874 8492
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 8202 8440 8208 8492
rect 8260 8440 8266 8492
rect 9306 8440 9312 8492
rect 9364 8440 9370 8492
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8480 12955 8483
rect 13170 8480 13176 8492
rect 12943 8452 13176 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 14090 8440 14096 8492
rect 14148 8440 14154 8492
rect 15378 8440 15384 8492
rect 15436 8440 15442 8492
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17972 8489 18000 8520
rect 24854 8508 24860 8520
rect 24912 8508 24918 8560
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 19242 8440 19248 8492
rect 19300 8480 19306 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19300 8452 19349 8480
rect 19300 8440 19306 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8449 20407 8483
rect 20349 8443 20407 8449
rect 21545 8483 21603 8489
rect 21545 8449 21557 8483
rect 21591 8480 21603 8483
rect 22002 8480 22008 8492
rect 21591 8452 22008 8480
rect 21591 8449 21603 8452
rect 21545 8443 21603 8449
rect 20364 8412 20392 8443
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 22741 8483 22799 8489
rect 22741 8449 22753 8483
rect 22787 8449 22799 8483
rect 22741 8443 22799 8449
rect 22554 8412 22560 8424
rect 20364 8384 22560 8412
rect 22554 8372 22560 8384
rect 22612 8372 22618 8424
rect 22756 8344 22784 8443
rect 23474 8440 23480 8492
rect 23532 8440 23538 8492
rect 23750 8440 23756 8492
rect 23808 8440 23814 8492
rect 23201 8415 23259 8421
rect 23201 8381 23213 8415
rect 23247 8412 23259 8415
rect 24762 8412 24768 8424
rect 23247 8384 24768 8412
rect 23247 8381 23259 8384
rect 23201 8375 23259 8381
rect 24762 8372 24768 8384
rect 24820 8372 24826 8424
rect 23934 8344 23940 8356
rect 22756 8316 23940 8344
rect 23934 8304 23940 8316
rect 23992 8304 23998 8356
rect 1104 8186 24564 8208
rect 1104 8134 3882 8186
rect 3934 8134 3946 8186
rect 3998 8134 4010 8186
rect 4062 8134 4074 8186
rect 4126 8134 4138 8186
rect 4190 8134 9747 8186
rect 9799 8134 9811 8186
rect 9863 8134 9875 8186
rect 9927 8134 9939 8186
rect 9991 8134 10003 8186
rect 10055 8134 15612 8186
rect 15664 8134 15676 8186
rect 15728 8134 15740 8186
rect 15792 8134 15804 8186
rect 15856 8134 15868 8186
rect 15920 8134 21477 8186
rect 21529 8134 21541 8186
rect 21593 8134 21605 8186
rect 21657 8134 21669 8186
rect 21721 8134 21733 8186
rect 21785 8134 24564 8186
rect 1104 8112 24564 8134
rect 16761 8075 16819 8081
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 17402 8072 17408 8084
rect 16807 8044 17408 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 17402 8032 17408 8044
rect 17460 8032 17466 8084
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 17126 7868 17132 7880
rect 16623 7840 17132 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 1104 7642 24723 7664
rect 1104 7590 6814 7642
rect 6866 7590 6878 7642
rect 6930 7590 6942 7642
rect 6994 7590 7006 7642
rect 7058 7590 7070 7642
rect 7122 7590 12679 7642
rect 12731 7590 12743 7642
rect 12795 7590 12807 7642
rect 12859 7590 12871 7642
rect 12923 7590 12935 7642
rect 12987 7590 18544 7642
rect 18596 7590 18608 7642
rect 18660 7590 18672 7642
rect 18724 7590 18736 7642
rect 18788 7590 18800 7642
rect 18852 7590 24409 7642
rect 24461 7590 24473 7642
rect 24525 7590 24537 7642
rect 24589 7590 24601 7642
rect 24653 7590 24665 7642
rect 24717 7590 24723 7642
rect 1104 7568 24723 7590
rect 1104 7098 24564 7120
rect 1104 7046 3882 7098
rect 3934 7046 3946 7098
rect 3998 7046 4010 7098
rect 4062 7046 4074 7098
rect 4126 7046 4138 7098
rect 4190 7046 9747 7098
rect 9799 7046 9811 7098
rect 9863 7046 9875 7098
rect 9927 7046 9939 7098
rect 9991 7046 10003 7098
rect 10055 7046 15612 7098
rect 15664 7046 15676 7098
rect 15728 7046 15740 7098
rect 15792 7046 15804 7098
rect 15856 7046 15868 7098
rect 15920 7046 21477 7098
rect 21529 7046 21541 7098
rect 21593 7046 21605 7098
rect 21657 7046 21669 7098
rect 21721 7046 21733 7098
rect 21785 7046 24564 7098
rect 1104 7024 24564 7046
rect 1104 6554 24723 6576
rect 1104 6502 6814 6554
rect 6866 6502 6878 6554
rect 6930 6502 6942 6554
rect 6994 6502 7006 6554
rect 7058 6502 7070 6554
rect 7122 6502 12679 6554
rect 12731 6502 12743 6554
rect 12795 6502 12807 6554
rect 12859 6502 12871 6554
rect 12923 6502 12935 6554
rect 12987 6502 18544 6554
rect 18596 6502 18608 6554
rect 18660 6502 18672 6554
rect 18724 6502 18736 6554
rect 18788 6502 18800 6554
rect 18852 6502 24409 6554
rect 24461 6502 24473 6554
rect 24525 6502 24537 6554
rect 24589 6502 24601 6554
rect 24653 6502 24665 6554
rect 24717 6502 24723 6554
rect 1104 6480 24723 6502
rect 1104 6010 24564 6032
rect 1104 5958 3882 6010
rect 3934 5958 3946 6010
rect 3998 5958 4010 6010
rect 4062 5958 4074 6010
rect 4126 5958 4138 6010
rect 4190 5958 9747 6010
rect 9799 5958 9811 6010
rect 9863 5958 9875 6010
rect 9927 5958 9939 6010
rect 9991 5958 10003 6010
rect 10055 5958 15612 6010
rect 15664 5958 15676 6010
rect 15728 5958 15740 6010
rect 15792 5958 15804 6010
rect 15856 5958 15868 6010
rect 15920 5958 21477 6010
rect 21529 5958 21541 6010
rect 21593 5958 21605 6010
rect 21657 5958 21669 6010
rect 21721 5958 21733 6010
rect 21785 5958 24564 6010
rect 1104 5936 24564 5958
rect 1104 5466 24723 5488
rect 1104 5414 6814 5466
rect 6866 5414 6878 5466
rect 6930 5414 6942 5466
rect 6994 5414 7006 5466
rect 7058 5414 7070 5466
rect 7122 5414 12679 5466
rect 12731 5414 12743 5466
rect 12795 5414 12807 5466
rect 12859 5414 12871 5466
rect 12923 5414 12935 5466
rect 12987 5414 18544 5466
rect 18596 5414 18608 5466
rect 18660 5414 18672 5466
rect 18724 5414 18736 5466
rect 18788 5414 18800 5466
rect 18852 5414 24409 5466
rect 24461 5414 24473 5466
rect 24525 5414 24537 5466
rect 24589 5414 24601 5466
rect 24653 5414 24665 5466
rect 24717 5414 24723 5466
rect 1104 5392 24723 5414
rect 1104 4922 24564 4944
rect 1104 4870 3882 4922
rect 3934 4870 3946 4922
rect 3998 4870 4010 4922
rect 4062 4870 4074 4922
rect 4126 4870 4138 4922
rect 4190 4870 9747 4922
rect 9799 4870 9811 4922
rect 9863 4870 9875 4922
rect 9927 4870 9939 4922
rect 9991 4870 10003 4922
rect 10055 4870 15612 4922
rect 15664 4870 15676 4922
rect 15728 4870 15740 4922
rect 15792 4870 15804 4922
rect 15856 4870 15868 4922
rect 15920 4870 21477 4922
rect 21529 4870 21541 4922
rect 21593 4870 21605 4922
rect 21657 4870 21669 4922
rect 21721 4870 21733 4922
rect 21785 4870 24564 4922
rect 1104 4848 24564 4870
rect 1104 4378 24723 4400
rect 1104 4326 6814 4378
rect 6866 4326 6878 4378
rect 6930 4326 6942 4378
rect 6994 4326 7006 4378
rect 7058 4326 7070 4378
rect 7122 4326 12679 4378
rect 12731 4326 12743 4378
rect 12795 4326 12807 4378
rect 12859 4326 12871 4378
rect 12923 4326 12935 4378
rect 12987 4326 18544 4378
rect 18596 4326 18608 4378
rect 18660 4326 18672 4378
rect 18724 4326 18736 4378
rect 18788 4326 18800 4378
rect 18852 4326 24409 4378
rect 24461 4326 24473 4378
rect 24525 4326 24537 4378
rect 24589 4326 24601 4378
rect 24653 4326 24665 4378
rect 24717 4326 24723 4378
rect 1104 4304 24723 4326
rect 9490 4088 9496 4140
rect 9548 4088 9554 4140
rect 10686 4088 10692 4140
rect 10744 4088 10750 4140
rect 11882 4088 11888 4140
rect 11940 4088 11946 4140
rect 13078 4088 13084 4140
rect 13136 4088 13142 4140
rect 19978 4088 19984 4140
rect 20036 4088 20042 4140
rect 24026 4088 24032 4140
rect 24084 4088 24090 4140
rect 22738 4060 22744 4072
rect 10796 4032 22744 4060
rect 10796 3936 10824 4032
rect 22738 4020 22744 4032
rect 22796 4020 22802 4072
rect 19794 3952 19800 4004
rect 19852 3952 19858 4004
rect 9306 3884 9312 3936
rect 9364 3884 9370 3936
rect 10502 3884 10508 3936
rect 10560 3884 10566 3936
rect 10778 3884 10784 3936
rect 10836 3884 10842 3936
rect 11698 3884 11704 3936
rect 11756 3884 11762 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13170 3924 13176 3936
rect 12943 3896 13176 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13170 3884 13176 3896
rect 13228 3884 13234 3936
rect 23474 3884 23480 3936
rect 23532 3924 23538 3936
rect 23845 3927 23903 3933
rect 23845 3924 23857 3927
rect 23532 3896 23857 3924
rect 23532 3884 23538 3896
rect 23845 3893 23857 3896
rect 23891 3893 23903 3927
rect 23845 3887 23903 3893
rect 1104 3834 24564 3856
rect 1104 3782 3882 3834
rect 3934 3782 3946 3834
rect 3998 3782 4010 3834
rect 4062 3782 4074 3834
rect 4126 3782 4138 3834
rect 4190 3782 9747 3834
rect 9799 3782 9811 3834
rect 9863 3782 9875 3834
rect 9927 3782 9939 3834
rect 9991 3782 10003 3834
rect 10055 3782 15612 3834
rect 15664 3782 15676 3834
rect 15728 3782 15740 3834
rect 15792 3782 15804 3834
rect 15856 3782 15868 3834
rect 15920 3782 21477 3834
rect 21529 3782 21541 3834
rect 21593 3782 21605 3834
rect 21657 3782 21669 3834
rect 21721 3782 21733 3834
rect 21785 3782 24564 3834
rect 1104 3760 24564 3782
rect 9490 3680 9496 3732
rect 9548 3680 9554 3732
rect 10597 3723 10655 3729
rect 10597 3689 10609 3723
rect 10643 3720 10655 3723
rect 10686 3720 10692 3732
rect 10643 3692 10692 3720
rect 10643 3689 10655 3692
rect 10597 3683 10655 3689
rect 10686 3680 10692 3692
rect 10744 3680 10750 3732
rect 11793 3723 11851 3729
rect 11793 3689 11805 3723
rect 11839 3720 11851 3723
rect 11882 3720 11888 3732
rect 11839 3692 11888 3720
rect 11839 3689 11851 3692
rect 11793 3683 11851 3689
rect 11882 3680 11888 3692
rect 11940 3680 11946 3732
rect 12989 3723 13047 3729
rect 12989 3689 13001 3723
rect 13035 3720 13047 3723
rect 13078 3720 13084 3732
rect 13035 3692 13084 3720
rect 13035 3689 13047 3692
rect 12989 3683 13047 3689
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 14090 3680 14096 3732
rect 14148 3680 14154 3732
rect 15289 3723 15347 3729
rect 15289 3689 15301 3723
rect 15335 3720 15347 3723
rect 15378 3720 15384 3732
rect 15335 3692 15384 3720
rect 15335 3689 15347 3692
rect 15289 3683 15347 3689
rect 15378 3680 15384 3692
rect 15436 3680 15442 3732
rect 19978 3680 19984 3732
rect 20036 3680 20042 3732
rect 24026 3680 24032 3732
rect 24084 3680 24090 3732
rect 23198 3612 23204 3664
rect 23256 3652 23262 3664
rect 23569 3655 23627 3661
rect 23569 3652 23581 3655
rect 23256 3624 23581 3652
rect 23256 3612 23262 3624
rect 23569 3621 23581 3624
rect 23615 3621 23627 3655
rect 24210 3652 24216 3664
rect 23569 3615 23627 3621
rect 23676 3624 24216 3652
rect 19518 3584 19524 3596
rect 13188 3556 14504 3584
rect 9677 3519 9735 3525
rect 9677 3485 9689 3519
rect 9723 3516 9735 3519
rect 10594 3516 10600 3528
rect 9723 3488 10600 3516
rect 9723 3485 9735 3488
rect 9677 3479 9735 3485
rect 10594 3476 10600 3488
rect 10652 3476 10658 3528
rect 10778 3476 10784 3528
rect 10836 3476 10842 3528
rect 11974 3476 11980 3528
rect 12032 3476 12038 3528
rect 13188 3525 13216 3556
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 13173 3479 13231 3485
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14323 3488 14412 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14384 3389 14412 3488
rect 14476 3448 14504 3556
rect 14568 3556 19524 3584
rect 14568 3525 14596 3556
rect 19518 3544 19524 3556
rect 19576 3544 19582 3596
rect 23676 3584 23704 3624
rect 24210 3612 24216 3624
rect 24268 3612 24274 3664
rect 24302 3584 24308 3596
rect 22066 3556 23704 3584
rect 23768 3556 24308 3584
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 15470 3476 15476 3528
rect 15528 3476 15534 3528
rect 20165 3519 20223 3525
rect 20165 3485 20177 3519
rect 20211 3516 20223 3519
rect 20622 3516 20628 3528
rect 20211 3488 20628 3516
rect 20211 3485 20223 3488
rect 20165 3479 20223 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 22066 3448 22094 3556
rect 23290 3476 23296 3528
rect 23348 3516 23354 3528
rect 23768 3525 23796 3556
rect 24302 3544 24308 3556
rect 24360 3544 24366 3596
rect 23477 3519 23535 3525
rect 23477 3516 23489 3519
rect 23348 3488 23489 3516
rect 23348 3476 23354 3488
rect 23477 3485 23489 3488
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 23753 3519 23811 3525
rect 23753 3485 23765 3519
rect 23799 3485 23811 3519
rect 23753 3479 23811 3485
rect 23845 3519 23903 3525
rect 23845 3485 23857 3519
rect 23891 3485 23903 3519
rect 23845 3479 23903 3485
rect 23860 3448 23888 3479
rect 14476 3420 22094 3448
rect 23492 3420 23888 3448
rect 23492 3392 23520 3420
rect 14369 3383 14427 3389
rect 14369 3349 14381 3383
rect 14415 3349 14427 3383
rect 14369 3343 14427 3349
rect 19886 3340 19892 3392
rect 19944 3380 19950 3392
rect 23293 3383 23351 3389
rect 23293 3380 23305 3383
rect 19944 3352 23305 3380
rect 19944 3340 19950 3352
rect 23293 3349 23305 3352
rect 23339 3349 23351 3383
rect 23293 3343 23351 3349
rect 23474 3340 23480 3392
rect 23532 3340 23538 3392
rect 1104 3290 24723 3312
rect 1104 3238 6814 3290
rect 6866 3238 6878 3290
rect 6930 3238 6942 3290
rect 6994 3238 7006 3290
rect 7058 3238 7070 3290
rect 7122 3238 12679 3290
rect 12731 3238 12743 3290
rect 12795 3238 12807 3290
rect 12859 3238 12871 3290
rect 12923 3238 12935 3290
rect 12987 3238 18544 3290
rect 18596 3238 18608 3290
rect 18660 3238 18672 3290
rect 18724 3238 18736 3290
rect 18788 3238 18800 3290
rect 18852 3238 24409 3290
rect 24461 3238 24473 3290
rect 24525 3238 24537 3290
rect 24589 3238 24601 3290
rect 24653 3238 24665 3290
rect 24717 3238 24723 3290
rect 1104 3216 24723 3238
rect 8113 3179 8171 3185
rect 8113 3145 8125 3179
rect 8159 3176 8171 3179
rect 8202 3176 8208 3188
rect 8159 3148 8208 3176
rect 8159 3145 8171 3148
rect 8113 3139 8171 3145
rect 8202 3136 8208 3148
rect 8260 3136 8266 3188
rect 15381 3179 15439 3185
rect 15381 3145 15393 3179
rect 15427 3176 15439 3179
rect 15470 3176 15476 3188
rect 15427 3148 15476 3176
rect 15427 3145 15439 3148
rect 15381 3139 15439 3145
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 19886 3176 19892 3188
rect 19444 3148 19892 3176
rect 6638 3068 6644 3120
rect 6696 3108 6702 3120
rect 16482 3108 16488 3120
rect 6696 3080 16488 3108
rect 6696 3068 6702 3080
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 15565 3043 15623 3049
rect 9640 3012 14412 3040
rect 9640 3000 9646 3012
rect 14384 2984 14412 3012
rect 15565 3009 15577 3043
rect 15611 3040 15623 3043
rect 19444 3040 19472 3148
rect 19886 3136 19892 3148
rect 19944 3136 19950 3188
rect 22738 3136 22744 3188
rect 22796 3136 22802 3188
rect 23201 3179 23259 3185
rect 23201 3145 23213 3179
rect 23247 3176 23259 3179
rect 23658 3176 23664 3188
rect 23247 3148 23664 3176
rect 23247 3145 23259 3148
rect 23201 3139 23259 3145
rect 23658 3136 23664 3148
rect 23716 3136 23722 3188
rect 19518 3068 19524 3120
rect 19576 3068 19582 3120
rect 25498 3108 25504 3120
rect 23400 3080 25504 3108
rect 15611 3012 19472 3040
rect 15611 3009 15623 3012
rect 15565 3003 15623 3009
rect 9122 2932 9128 2984
rect 9180 2972 9186 2984
rect 12250 2972 12256 2984
rect 9180 2944 12256 2972
rect 9180 2932 9186 2944
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 14366 2932 14372 2984
rect 14424 2932 14430 2984
rect 7834 2864 7840 2916
rect 7892 2904 7898 2916
rect 16666 2904 16672 2916
rect 7892 2876 16672 2904
rect 7892 2864 7898 2876
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 19536 2904 19564 3068
rect 22646 3000 22652 3052
rect 22704 3000 22710 3052
rect 22925 3043 22983 3049
rect 22925 3009 22937 3043
rect 22971 3009 22983 3043
rect 22925 3003 22983 3009
rect 22370 2932 22376 2984
rect 22428 2972 22434 2984
rect 22940 2972 22968 3003
rect 23014 3000 23020 3052
rect 23072 3000 23078 3052
rect 23293 3044 23351 3049
rect 23400 3044 23428 3080
rect 25498 3068 25504 3080
rect 25556 3068 25562 3120
rect 23293 3043 23428 3044
rect 23293 3009 23305 3043
rect 23339 3016 23428 3043
rect 23753 3043 23811 3049
rect 23339 3009 23351 3016
rect 23293 3003 23351 3009
rect 23753 3009 23765 3043
rect 23799 3040 23811 3043
rect 23842 3040 23848 3052
rect 23799 3012 23848 3040
rect 23799 3009 23811 3012
rect 23753 3003 23811 3009
rect 23842 3000 23848 3012
rect 23900 3000 23906 3052
rect 24029 3043 24087 3049
rect 24029 3009 24041 3043
rect 24075 3009 24087 3043
rect 24029 3003 24087 3009
rect 22428 2944 22968 2972
rect 22428 2932 22434 2944
rect 23382 2932 23388 2984
rect 23440 2972 23446 2984
rect 24044 2972 24072 3003
rect 23440 2944 24072 2972
rect 23440 2932 23446 2944
rect 22465 2907 22523 2913
rect 22465 2904 22477 2907
rect 19536 2876 22477 2904
rect 22465 2873 22477 2876
rect 22511 2873 22523 2907
rect 22465 2867 22523 2873
rect 22664 2876 23888 2904
rect 8846 2796 8852 2848
rect 8904 2836 8910 2848
rect 14090 2836 14096 2848
rect 8904 2808 14096 2836
rect 8904 2796 8910 2808
rect 14090 2796 14096 2808
rect 14148 2796 14154 2848
rect 19886 2796 19892 2848
rect 19944 2836 19950 2848
rect 22664 2836 22692 2876
rect 19944 2808 22692 2836
rect 19944 2796 19950 2808
rect 23106 2796 23112 2848
rect 23164 2836 23170 2848
rect 23382 2836 23388 2848
rect 23164 2808 23388 2836
rect 23164 2796 23170 2808
rect 23382 2796 23388 2808
rect 23440 2796 23446 2848
rect 23474 2796 23480 2848
rect 23532 2796 23538 2848
rect 23566 2796 23572 2848
rect 23624 2796 23630 2848
rect 23860 2845 23888 2876
rect 23845 2839 23903 2845
rect 23845 2805 23857 2839
rect 23891 2805 23903 2839
rect 23845 2799 23903 2805
rect 1104 2746 24564 2768
rect 1104 2694 3882 2746
rect 3934 2694 3946 2746
rect 3998 2694 4010 2746
rect 4062 2694 4074 2746
rect 4126 2694 4138 2746
rect 4190 2694 9747 2746
rect 9799 2694 9811 2746
rect 9863 2694 9875 2746
rect 9927 2694 9939 2746
rect 9991 2694 10003 2746
rect 10055 2694 15612 2746
rect 15664 2694 15676 2746
rect 15728 2694 15740 2746
rect 15792 2694 15804 2746
rect 15856 2694 15868 2746
rect 15920 2694 21477 2746
rect 21529 2694 21541 2746
rect 21593 2694 21605 2746
rect 21657 2694 21669 2746
rect 21721 2694 21733 2746
rect 21785 2694 24564 2746
rect 1104 2672 24564 2694
rect 1857 2635 1915 2641
rect 1857 2632 1869 2635
rect 1504 2604 1869 2632
rect 1504 2496 1532 2604
rect 1857 2601 1869 2604
rect 1903 2601 1915 2635
rect 1857 2595 1915 2601
rect 2133 2635 2191 2641
rect 2133 2601 2145 2635
rect 2179 2632 2191 2635
rect 6822 2632 6828 2644
rect 2179 2604 6828 2632
rect 2179 2601 2191 2604
rect 2133 2595 2191 2601
rect 6822 2592 6828 2604
rect 6880 2592 6886 2644
rect 8205 2635 8263 2641
rect 8205 2601 8217 2635
rect 8251 2632 8263 2635
rect 8294 2632 8300 2644
rect 8251 2604 8300 2632
rect 8251 2601 8263 2604
rect 8205 2595 8263 2601
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8938 2592 8944 2644
rect 8996 2632 9002 2644
rect 8996 2604 14780 2632
rect 8996 2592 9002 2604
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 1627 2536 9904 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 5534 2496 5540 2508
rect 1504 2468 5540 2496
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 9582 2496 9588 2508
rect 5644 2468 9588 2496
rect 106 2388 112 2440
rect 164 2428 170 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 164 2400 1409 2428
rect 164 2388 170 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 658 2320 664 2372
rect 716 2360 722 2372
rect 1688 2360 1716 2391
rect 1946 2388 1952 2440
rect 2004 2388 2010 2440
rect 5644 2428 5672 2468
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 9876 2440 9904 2536
rect 10594 2456 10600 2508
rect 10652 2496 10658 2508
rect 14550 2496 14556 2508
rect 10652 2468 14556 2496
rect 10652 2456 10658 2468
rect 14550 2456 14556 2468
rect 14608 2456 14614 2508
rect 14752 2496 14780 2604
rect 14826 2592 14832 2644
rect 14884 2632 14890 2644
rect 14884 2604 18276 2632
rect 14884 2592 14890 2604
rect 16945 2567 17003 2573
rect 16945 2533 16957 2567
rect 16991 2564 17003 2567
rect 17402 2564 17408 2576
rect 16991 2536 17408 2564
rect 16991 2533 17003 2536
rect 16945 2527 17003 2533
rect 17402 2524 17408 2536
rect 17460 2524 17466 2576
rect 17497 2567 17555 2573
rect 17497 2533 17509 2567
rect 17543 2564 17555 2567
rect 18138 2564 18144 2576
rect 17543 2536 18144 2564
rect 17543 2533 17555 2536
rect 17497 2527 17555 2533
rect 18138 2524 18144 2536
rect 18196 2524 18202 2576
rect 18248 2564 18276 2604
rect 19242 2592 19248 2644
rect 19300 2592 19306 2644
rect 23017 2635 23075 2641
rect 23017 2601 23029 2635
rect 23063 2632 23075 2635
rect 23106 2632 23112 2644
rect 23063 2604 23112 2632
rect 23063 2601 23075 2604
rect 23017 2595 23075 2601
rect 23106 2592 23112 2604
rect 23164 2592 23170 2644
rect 23661 2635 23719 2641
rect 23661 2601 23673 2635
rect 23707 2632 23719 2635
rect 23750 2632 23756 2644
rect 23707 2604 23756 2632
rect 23707 2601 23719 2604
rect 23661 2595 23719 2601
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 23860 2604 24164 2632
rect 20806 2564 20812 2576
rect 18248 2536 20812 2564
rect 20806 2524 20812 2536
rect 20864 2524 20870 2576
rect 22189 2567 22247 2573
rect 22189 2533 22201 2567
rect 22235 2564 22247 2567
rect 22554 2564 22560 2576
rect 22235 2536 22560 2564
rect 22235 2533 22247 2536
rect 22189 2527 22247 2533
rect 22554 2524 22560 2536
rect 22612 2524 22618 2576
rect 22741 2567 22799 2573
rect 22741 2533 22753 2567
rect 22787 2564 22799 2567
rect 23860 2564 23888 2604
rect 22787 2536 23888 2564
rect 23937 2567 23995 2573
rect 22787 2533 22799 2536
rect 22741 2527 22799 2533
rect 23937 2533 23949 2567
rect 23983 2533 23995 2567
rect 23937 2527 23995 2533
rect 14752 2468 17080 2496
rect 2056 2400 5672 2428
rect 8389 2431 8447 2437
rect 716 2332 1716 2360
rect 716 2320 722 2332
rect 1854 2320 1860 2372
rect 1912 2360 1918 2372
rect 2056 2360 2084 2400
rect 8389 2397 8401 2431
rect 8435 2428 8447 2431
rect 8846 2428 8852 2440
rect 8435 2400 8852 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8846 2388 8852 2400
rect 8904 2388 8910 2440
rect 9858 2388 9864 2440
rect 9916 2388 9922 2440
rect 10042 2388 10048 2440
rect 10100 2428 10106 2440
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10100 2400 10701 2428
rect 10100 2388 10106 2400
rect 10689 2397 10701 2400
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 11330 2388 11336 2440
rect 11388 2388 11394 2440
rect 11698 2388 11704 2440
rect 11756 2388 11762 2440
rect 12250 2388 12256 2440
rect 12308 2388 12314 2440
rect 12342 2388 12348 2440
rect 12400 2428 12406 2440
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12400 2400 12541 2428
rect 12400 2388 12406 2400
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 12529 2391 12587 2397
rect 13630 2388 13636 2440
rect 13688 2428 13694 2440
rect 14921 2431 14979 2437
rect 14921 2428 14933 2431
rect 13688 2400 14933 2428
rect 13688 2388 13694 2400
rect 14921 2397 14933 2400
rect 14967 2397 14979 2431
rect 14921 2391 14979 2397
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 16117 2431 16175 2437
rect 16117 2428 16129 2431
rect 15988 2400 16129 2428
rect 15988 2388 15994 2400
rect 16117 2397 16129 2400
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 16758 2388 16764 2440
rect 16816 2388 16822 2440
rect 17052 2437 17080 2468
rect 17126 2456 17132 2508
rect 17184 2496 17190 2508
rect 17184 2468 22416 2496
rect 17184 2456 17190 2468
rect 17037 2431 17095 2437
rect 17037 2397 17049 2431
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 1912 2332 2084 2360
rect 1912 2320 1918 2332
rect 8570 2320 8576 2372
rect 8628 2360 8634 2372
rect 17328 2360 17356 2391
rect 17678 2388 17684 2440
rect 17736 2428 17742 2440
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 17736 2400 17785 2428
rect 17736 2388 17742 2400
rect 17773 2397 17785 2400
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2428 18107 2431
rect 18230 2428 18236 2440
rect 18095 2400 18236 2428
rect 18095 2397 18107 2400
rect 18049 2391 18107 2397
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 18417 2431 18475 2437
rect 18417 2397 18429 2431
rect 18463 2428 18475 2431
rect 19058 2428 19064 2440
rect 18463 2400 19064 2428
rect 18463 2397 18475 2400
rect 18417 2391 18475 2397
rect 19058 2388 19064 2400
rect 19116 2388 19122 2440
rect 19429 2431 19487 2437
rect 19429 2397 19441 2431
rect 19475 2428 19487 2431
rect 19886 2428 19892 2440
rect 19475 2400 19892 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 19886 2388 19892 2400
rect 19944 2388 19950 2440
rect 19978 2388 19984 2440
rect 20036 2388 20042 2440
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2428 22063 2431
rect 22051 2400 22324 2428
rect 22051 2397 22063 2400
rect 22005 2391 22063 2397
rect 8628 2332 17356 2360
rect 8628 2320 8634 2332
rect 19610 2320 19616 2372
rect 19668 2320 19674 2372
rect 19797 2363 19855 2369
rect 19797 2329 19809 2363
rect 19843 2360 19855 2363
rect 21818 2360 21824 2372
rect 19843 2332 21824 2360
rect 19843 2329 19855 2332
rect 19797 2323 19855 2329
rect 21818 2320 21824 2332
rect 21876 2320 21882 2372
rect 5718 2252 5724 2304
rect 5776 2292 5782 2304
rect 9214 2292 9220 2304
rect 5776 2264 9220 2292
rect 5776 2252 5782 2264
rect 9214 2252 9220 2264
rect 9272 2252 9278 2304
rect 9398 2252 9404 2304
rect 9456 2292 9462 2304
rect 10226 2292 10232 2304
rect 9456 2264 10232 2292
rect 9456 2252 9462 2264
rect 10226 2252 10232 2264
rect 10284 2252 10290 2304
rect 10870 2252 10876 2304
rect 10928 2252 10934 2304
rect 11514 2252 11520 2304
rect 11572 2252 11578 2304
rect 11882 2252 11888 2304
rect 11940 2252 11946 2304
rect 12434 2252 12440 2304
rect 12492 2252 12498 2304
rect 12713 2295 12771 2301
rect 12713 2261 12725 2295
rect 12759 2292 12771 2295
rect 13078 2292 13084 2304
rect 12759 2264 13084 2292
rect 12759 2261 12771 2264
rect 12713 2255 12771 2261
rect 13078 2252 13084 2264
rect 13136 2252 13142 2304
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 13722 2292 13728 2304
rect 13320 2264 13728 2292
rect 13320 2252 13326 2264
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 15102 2252 15108 2304
rect 15160 2252 15166 2304
rect 16301 2295 16359 2301
rect 16301 2261 16313 2295
rect 16347 2292 16359 2295
rect 17126 2292 17132 2304
rect 16347 2264 17132 2292
rect 16347 2261 16359 2264
rect 16301 2255 16359 2261
rect 17126 2252 17132 2264
rect 17184 2252 17190 2304
rect 17218 2252 17224 2304
rect 17276 2252 17282 2304
rect 17957 2295 18015 2301
rect 17957 2261 17969 2295
rect 18003 2292 18015 2295
rect 18046 2292 18052 2304
rect 18003 2264 18052 2292
rect 18003 2261 18015 2264
rect 17957 2255 18015 2261
rect 18046 2252 18052 2264
rect 18104 2252 18110 2304
rect 18233 2295 18291 2301
rect 18233 2261 18245 2295
rect 18279 2292 18291 2295
rect 18414 2292 18420 2304
rect 18279 2264 18420 2292
rect 18279 2261 18291 2264
rect 18233 2255 18291 2261
rect 18414 2252 18420 2264
rect 18472 2252 18478 2304
rect 18601 2295 18659 2301
rect 18601 2261 18613 2295
rect 18647 2292 18659 2295
rect 19242 2292 19248 2304
rect 18647 2264 19248 2292
rect 18647 2261 18659 2264
rect 18601 2255 18659 2261
rect 19242 2252 19248 2264
rect 19300 2252 19306 2304
rect 20162 2252 20168 2304
rect 20220 2252 20226 2304
rect 22296 2301 22324 2400
rect 22281 2295 22339 2301
rect 22281 2261 22293 2295
rect 22327 2261 22339 2295
rect 22388 2292 22416 2468
rect 23216 2468 23796 2496
rect 22465 2431 22523 2437
rect 22465 2397 22477 2431
rect 22511 2397 22523 2431
rect 22465 2391 22523 2397
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2428 22615 2431
rect 22738 2428 22744 2440
rect 22603 2400 22744 2428
rect 22603 2397 22615 2400
rect 22557 2391 22615 2397
rect 22480 2360 22508 2391
rect 22738 2388 22744 2400
rect 22796 2388 22802 2440
rect 22833 2431 22891 2437
rect 22833 2397 22845 2431
rect 22879 2428 22891 2431
rect 23216 2428 23244 2468
rect 22879 2400 23244 2428
rect 23293 2431 23351 2437
rect 22879 2397 22891 2400
rect 22833 2391 22891 2397
rect 23293 2397 23305 2431
rect 23339 2397 23351 2431
rect 23293 2391 23351 2397
rect 23385 2431 23443 2437
rect 23385 2397 23397 2431
rect 23431 2428 23443 2431
rect 23566 2428 23572 2440
rect 23431 2400 23572 2428
rect 23431 2397 23443 2400
rect 23385 2391 23443 2397
rect 22922 2360 22928 2372
rect 22480 2332 22928 2360
rect 22922 2320 22928 2332
rect 22980 2320 22986 2372
rect 23308 2360 23336 2391
rect 23566 2388 23572 2400
rect 23624 2388 23630 2440
rect 23474 2360 23480 2372
rect 23308 2332 23480 2360
rect 23474 2320 23480 2332
rect 23532 2320 23538 2372
rect 23768 2360 23796 2468
rect 23845 2431 23903 2437
rect 23845 2397 23857 2431
rect 23891 2428 23903 2431
rect 23952 2428 23980 2527
rect 24136 2437 24164 2604
rect 23891 2400 23980 2428
rect 24121 2431 24179 2437
rect 23891 2397 23903 2400
rect 23845 2391 23903 2397
rect 24121 2397 24133 2431
rect 24167 2397 24179 2431
rect 24121 2391 24179 2397
rect 23768 2332 24164 2360
rect 24136 2304 24164 2332
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 22388 2264 23121 2292
rect 22281 2255 22339 2261
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 23569 2295 23627 2301
rect 23569 2261 23581 2295
rect 23615 2292 23627 2295
rect 24026 2292 24032 2304
rect 23615 2264 24032 2292
rect 23615 2261 23627 2264
rect 23569 2255 23627 2261
rect 24026 2252 24032 2264
rect 24084 2252 24090 2304
rect 24118 2252 24124 2304
rect 24176 2252 24182 2304
rect 1104 2202 24723 2224
rect 1104 2150 6814 2202
rect 6866 2150 6878 2202
rect 6930 2150 6942 2202
rect 6994 2150 7006 2202
rect 7058 2150 7070 2202
rect 7122 2150 12679 2202
rect 12731 2150 12743 2202
rect 12795 2150 12807 2202
rect 12859 2150 12871 2202
rect 12923 2150 12935 2202
rect 12987 2150 18544 2202
rect 18596 2150 18608 2202
rect 18660 2150 18672 2202
rect 18724 2150 18736 2202
rect 18788 2150 18800 2202
rect 18852 2150 24409 2202
rect 24461 2150 24473 2202
rect 24525 2150 24537 2202
rect 24589 2150 24601 2202
rect 24653 2150 24665 2202
rect 24717 2150 24723 2202
rect 1104 2128 24723 2150
rect 1765 2091 1823 2097
rect 1765 2057 1777 2091
rect 1811 2088 1823 2091
rect 1854 2088 1860 2100
rect 1811 2060 1860 2088
rect 1811 2057 1823 2060
rect 1765 2051 1823 2057
rect 1854 2048 1860 2060
rect 1912 2048 1918 2100
rect 2041 2091 2099 2097
rect 2041 2057 2053 2091
rect 2087 2057 2099 2091
rect 2041 2051 2099 2057
rect 5353 2091 5411 2097
rect 5353 2057 5365 2091
rect 5399 2088 5411 2091
rect 5718 2088 5724 2100
rect 5399 2060 5724 2088
rect 5399 2057 5411 2060
rect 5353 2051 5411 2057
rect 2056 2020 2084 2051
rect 5718 2048 5724 2060
rect 5776 2048 5782 2100
rect 5810 2048 5816 2100
rect 5868 2088 5874 2100
rect 5905 2091 5963 2097
rect 5905 2088 5917 2091
rect 5868 2060 5917 2088
rect 5868 2048 5874 2060
rect 5905 2057 5917 2060
rect 5951 2057 5963 2091
rect 5905 2051 5963 2057
rect 6822 2048 6828 2100
rect 6880 2048 6886 2100
rect 7101 2091 7159 2097
rect 7101 2057 7113 2091
rect 7147 2088 7159 2091
rect 7190 2088 7196 2100
rect 7147 2060 7196 2088
rect 7147 2057 7159 2060
rect 7101 2051 7159 2057
rect 7190 2048 7196 2060
rect 7248 2048 7254 2100
rect 9674 2088 9680 2100
rect 7300 2060 9680 2088
rect 7300 2020 7328 2060
rect 9674 2048 9680 2060
rect 9732 2048 9738 2100
rect 9769 2091 9827 2097
rect 9769 2057 9781 2091
rect 9815 2057 9827 2091
rect 9769 2051 9827 2057
rect 10045 2091 10103 2097
rect 10045 2057 10057 2091
rect 10091 2088 10103 2091
rect 10091 2060 10548 2088
rect 10091 2057 10103 2060
rect 10045 2051 10103 2057
rect 9398 2020 9404 2032
rect 2056 1992 7328 2020
rect 7944 1992 9404 2020
rect 1578 1912 1584 1964
rect 1636 1912 1642 1964
rect 1857 1955 1915 1961
rect 1857 1921 1869 1955
rect 1903 1921 1915 1955
rect 1857 1915 1915 1921
rect 2133 1955 2191 1961
rect 2133 1921 2145 1955
rect 2179 1921 2191 1955
rect 2133 1915 2191 1921
rect 1210 1844 1216 1896
rect 1268 1884 1274 1896
rect 1872 1884 1900 1915
rect 1268 1856 1900 1884
rect 1268 1844 1274 1856
rect 382 1776 388 1828
rect 440 1816 446 1828
rect 2148 1816 2176 1915
rect 2406 1912 2412 1964
rect 2464 1912 2470 1964
rect 5166 1912 5172 1964
rect 5224 1912 5230 1964
rect 5442 1912 5448 1964
rect 5500 1912 5506 1964
rect 5718 1912 5724 1964
rect 5776 1912 5782 1964
rect 5997 1955 6055 1961
rect 5997 1921 6009 1955
rect 6043 1921 6055 1955
rect 5997 1915 6055 1921
rect 6012 1884 6040 1915
rect 6638 1912 6644 1964
rect 6696 1912 6702 1964
rect 6822 1912 6828 1964
rect 6880 1952 6886 1964
rect 6917 1955 6975 1961
rect 6917 1952 6929 1955
rect 6880 1924 6929 1952
rect 6880 1912 6886 1924
rect 6917 1921 6929 1924
rect 6963 1921 6975 1955
rect 6917 1915 6975 1921
rect 7282 1912 7288 1964
rect 7340 1952 7346 1964
rect 7561 1955 7619 1961
rect 7561 1952 7573 1955
rect 7340 1924 7573 1952
rect 7340 1912 7346 1924
rect 7561 1921 7573 1924
rect 7607 1921 7619 1955
rect 7561 1915 7619 1921
rect 7650 1912 7656 1964
rect 7708 1912 7714 1964
rect 2608 1856 6040 1884
rect 2608 1825 2636 1856
rect 440 1788 2176 1816
rect 2593 1819 2651 1825
rect 440 1776 446 1788
rect 2593 1785 2605 1819
rect 2639 1785 2651 1819
rect 2593 1779 2651 1785
rect 5629 1819 5687 1825
rect 5629 1785 5641 1819
rect 5675 1816 5687 1819
rect 6086 1816 6092 1828
rect 5675 1788 6092 1816
rect 5675 1785 5687 1788
rect 5629 1779 5687 1785
rect 6086 1776 6092 1788
rect 6144 1776 6150 1828
rect 6181 1819 6239 1825
rect 6181 1785 6193 1819
rect 6227 1816 6239 1819
rect 7944 1816 7972 1992
rect 9398 1980 9404 1992
rect 9456 1980 9462 2032
rect 8110 1912 8116 1964
rect 8168 1912 8174 1964
rect 8478 1912 8484 1964
rect 8536 1912 8542 1964
rect 8754 1912 8760 1964
rect 8812 1912 8818 1964
rect 8938 1912 8944 1964
rect 8996 1952 9002 1964
rect 9217 1955 9275 1961
rect 9217 1952 9229 1955
rect 8996 1924 9229 1952
rect 8996 1912 9002 1924
rect 9217 1921 9229 1924
rect 9263 1921 9275 1955
rect 9217 1915 9275 1921
rect 9306 1912 9312 1964
rect 9364 1912 9370 1964
rect 9593 1955 9651 1961
rect 9593 1921 9605 1955
rect 9639 1952 9651 1955
rect 9639 1924 9720 1952
rect 9639 1921 9651 1924
rect 9593 1915 9651 1921
rect 9692 1884 9720 1924
rect 9508 1856 9720 1884
rect 9784 1884 9812 2051
rect 10226 2029 10232 2032
rect 10211 2023 10232 2029
rect 10211 1989 10223 2023
rect 10211 1983 10232 1989
rect 10226 1980 10232 1983
rect 10284 1980 10290 2032
rect 10520 2020 10548 2060
rect 10870 2048 10876 2100
rect 10928 2088 10934 2100
rect 10928 2060 11928 2088
rect 10928 2048 10934 2060
rect 11900 2029 11928 2060
rect 12434 2048 12440 2100
rect 12492 2048 12498 2100
rect 12526 2048 12532 2100
rect 12584 2088 12590 2100
rect 14461 2091 14519 2097
rect 12584 2060 13216 2088
rect 12584 2048 12590 2060
rect 10965 2023 11023 2029
rect 10965 2020 10977 2023
rect 10520 1992 10977 2020
rect 10965 1989 10977 1992
rect 11011 1989 11023 2023
rect 10965 1983 11023 1989
rect 11885 2023 11943 2029
rect 11885 1989 11897 2023
rect 11931 1989 11943 2023
rect 12452 2020 12480 2048
rect 12452 1992 12756 2020
rect 11885 1983 11943 1989
rect 9858 1912 9864 1964
rect 9916 1912 9922 1964
rect 10502 1912 10508 1964
rect 10560 1952 10566 1964
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 10560 1924 11529 1952
rect 10560 1912 10566 1924
rect 11517 1921 11529 1924
rect 11563 1921 11575 1955
rect 11517 1915 11575 1921
rect 12066 1912 12072 1964
rect 12124 1952 12130 1964
rect 12728 1961 12756 1992
rect 13188 1961 13216 2060
rect 14461 2057 14473 2091
rect 14507 2057 14519 2091
rect 14461 2051 14519 2057
rect 14476 2020 14504 2051
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 15013 2091 15071 2097
rect 15013 2088 15025 2091
rect 14608 2060 15025 2088
rect 14608 2048 14614 2060
rect 15013 2057 15025 2060
rect 15059 2057 15071 2091
rect 15013 2051 15071 2057
rect 15102 2048 15108 2100
rect 15160 2088 15166 2100
rect 15160 2060 15516 2088
rect 15160 2048 15166 2060
rect 15378 2020 15384 2032
rect 14476 1992 15384 2020
rect 15378 1980 15384 1992
rect 15436 1980 15442 2032
rect 15488 2029 15516 2060
rect 17218 2048 17224 2100
rect 17276 2048 17282 2100
rect 17402 2048 17408 2100
rect 17460 2088 17466 2100
rect 17460 2060 18368 2088
rect 17460 2048 17466 2060
rect 15473 2023 15531 2029
rect 15473 1989 15485 2023
rect 15519 1989 15531 2023
rect 15473 1983 15531 1989
rect 16666 1980 16672 2032
rect 16724 2020 16730 2032
rect 16761 2023 16819 2029
rect 16761 2020 16773 2023
rect 16724 1992 16773 2020
rect 16724 1980 16730 1992
rect 16761 1989 16773 1992
rect 16807 1989 16819 2023
rect 16761 1983 16819 1989
rect 12437 1955 12495 1961
rect 12437 1952 12449 1955
rect 12124 1924 12449 1952
rect 12124 1912 12130 1924
rect 12437 1921 12449 1924
rect 12483 1921 12495 1955
rect 12437 1915 12495 1921
rect 12713 1955 12771 1961
rect 12713 1921 12725 1955
rect 12759 1921 12771 1955
rect 12713 1915 12771 1921
rect 13173 1955 13231 1961
rect 13173 1921 13185 1955
rect 13219 1921 13231 1955
rect 13173 1915 13231 1921
rect 13446 1912 13452 1964
rect 13504 1912 13510 1964
rect 13630 1912 13636 1964
rect 13688 1912 13694 1964
rect 13722 1912 13728 1964
rect 13780 1912 13786 1964
rect 13998 1912 14004 1964
rect 14056 1912 14062 1964
rect 14274 1912 14280 1964
rect 14332 1912 14338 1964
rect 14366 1912 14372 1964
rect 14424 1952 14430 1964
rect 14553 1955 14611 1961
rect 14553 1952 14565 1955
rect 14424 1924 14565 1952
rect 14424 1912 14430 1924
rect 14553 1921 14565 1924
rect 14599 1921 14611 1955
rect 14553 1915 14611 1921
rect 14829 1955 14887 1961
rect 14829 1921 14841 1955
rect 14875 1921 14887 1955
rect 14829 1915 14887 1921
rect 13354 1884 13360 1896
rect 9784 1856 13360 1884
rect 9398 1816 9404 1828
rect 6227 1788 7972 1816
rect 8312 1788 9404 1816
rect 6227 1785 6239 1788
rect 6181 1779 6239 1785
rect 2317 1751 2375 1757
rect 2317 1717 2329 1751
rect 2363 1748 2375 1751
rect 5994 1748 6000 1760
rect 2363 1720 6000 1748
rect 2363 1717 2375 1720
rect 2317 1711 2375 1717
rect 5994 1708 6000 1720
rect 6052 1708 6058 1760
rect 6638 1708 6644 1760
rect 6696 1748 6702 1760
rect 7377 1751 7435 1757
rect 7377 1748 7389 1751
rect 6696 1720 7389 1748
rect 6696 1708 6702 1720
rect 7377 1717 7389 1720
rect 7423 1717 7435 1751
rect 7377 1711 7435 1717
rect 7837 1751 7895 1757
rect 7837 1717 7849 1751
rect 7883 1748 7895 1751
rect 8202 1748 8208 1760
rect 7883 1720 8208 1748
rect 7883 1717 7895 1720
rect 7837 1711 7895 1717
rect 8202 1708 8208 1720
rect 8260 1708 8266 1760
rect 8312 1757 8340 1788
rect 9398 1776 9404 1788
rect 9456 1776 9462 1828
rect 9508 1825 9536 1856
rect 13354 1844 13360 1856
rect 13412 1844 13418 1896
rect 9493 1819 9551 1825
rect 9493 1785 9505 1819
rect 9539 1785 9551 1819
rect 9493 1779 9551 1785
rect 9674 1776 9680 1828
rect 9732 1816 9738 1828
rect 13648 1816 13676 1912
rect 14844 1884 14872 1915
rect 15562 1912 15568 1964
rect 15620 1952 15626 1964
rect 15933 1955 15991 1961
rect 15933 1952 15945 1955
rect 15620 1924 15945 1952
rect 15620 1912 15626 1924
rect 15933 1921 15945 1924
rect 15979 1921 15991 1955
rect 15933 1915 15991 1921
rect 16298 1912 16304 1964
rect 16356 1912 16362 1964
rect 17236 1961 17264 2048
rect 17954 1980 17960 2032
rect 18012 2020 18018 2032
rect 18233 2023 18291 2029
rect 18233 2020 18245 2023
rect 18012 1992 18245 2020
rect 18012 1980 18018 1992
rect 18233 1989 18245 1992
rect 18279 1989 18291 2023
rect 18340 2020 18368 2060
rect 18414 2048 18420 2100
rect 18472 2088 18478 2100
rect 18472 2060 19380 2088
rect 18472 2048 18478 2060
rect 19352 2029 19380 2060
rect 20162 2048 20168 2100
rect 20220 2048 20226 2100
rect 20901 2091 20959 2097
rect 20901 2057 20913 2091
rect 20947 2057 20959 2091
rect 20901 2051 20959 2057
rect 21453 2091 21511 2097
rect 21453 2057 21465 2091
rect 21499 2057 21511 2091
rect 21453 2051 21511 2057
rect 18785 2023 18843 2029
rect 18785 2020 18797 2023
rect 18340 1992 18797 2020
rect 18233 1983 18291 1989
rect 18785 1989 18797 1992
rect 18831 1989 18843 2023
rect 18785 1983 18843 1989
rect 19337 2023 19395 2029
rect 19337 1989 19349 2023
rect 19383 1989 19395 2023
rect 20180 2020 20208 2048
rect 20441 2023 20499 2029
rect 20441 2020 20453 2023
rect 20180 1992 20453 2020
rect 19337 1983 19395 1989
rect 20441 1989 20453 1992
rect 20487 1989 20499 2023
rect 20441 1983 20499 1989
rect 17221 1955 17279 1961
rect 17221 1921 17233 1955
rect 17267 1921 17279 1955
rect 17221 1915 17279 1921
rect 17681 1955 17739 1961
rect 17681 1921 17693 1955
rect 17727 1921 17739 1955
rect 17681 1915 17739 1921
rect 20165 1955 20223 1961
rect 20165 1921 20177 1955
rect 20211 1952 20223 1955
rect 20916 1952 20944 2051
rect 20211 1924 20944 1952
rect 21085 1955 21143 1961
rect 20211 1921 20223 1924
rect 20165 1915 20223 1921
rect 21085 1921 21097 1955
rect 21131 1921 21143 1955
rect 21085 1915 21143 1921
rect 21361 1955 21419 1961
rect 21361 1921 21373 1955
rect 21407 1952 21419 1955
rect 21468 1952 21496 2051
rect 21542 2048 21548 2100
rect 21600 2088 21606 2100
rect 21821 2091 21879 2097
rect 21821 2088 21833 2091
rect 21600 2060 21833 2088
rect 21600 2048 21606 2060
rect 21821 2057 21833 2060
rect 21867 2057 21879 2091
rect 21821 2051 21879 2057
rect 22002 2048 22008 2100
rect 22060 2088 22066 2100
rect 22373 2091 22431 2097
rect 22373 2088 22385 2091
rect 22060 2060 22385 2088
rect 22060 2048 22066 2060
rect 22373 2057 22385 2060
rect 22419 2057 22431 2091
rect 22373 2051 22431 2057
rect 22554 2048 22560 2100
rect 22612 2048 22618 2100
rect 22646 2048 22652 2100
rect 22704 2048 22710 2100
rect 22925 2091 22983 2097
rect 22925 2057 22937 2091
rect 22971 2057 22983 2091
rect 22925 2051 22983 2057
rect 22186 2020 22192 2032
rect 21652 1992 22192 2020
rect 21652 1961 21680 1992
rect 22186 1980 22192 1992
rect 22244 1980 22250 2032
rect 22572 2020 22600 2048
rect 22572 1992 22784 2020
rect 21407 1924 21496 1952
rect 21637 1955 21695 1961
rect 21407 1921 21419 1924
rect 21361 1915 21419 1921
rect 21637 1921 21649 1955
rect 21683 1921 21695 1955
rect 21637 1915 21695 1921
rect 22005 1955 22063 1961
rect 22005 1921 22017 1955
rect 22051 1952 22063 1955
rect 22051 1924 22140 1952
rect 22051 1921 22063 1924
rect 22005 1915 22063 1921
rect 13924 1856 14872 1884
rect 13924 1825 13952 1856
rect 14918 1844 14924 1896
rect 14976 1884 14982 1896
rect 17696 1884 17724 1915
rect 14976 1856 17724 1884
rect 14976 1844 14982 1856
rect 18046 1844 18052 1896
rect 18104 1884 18110 1896
rect 19610 1884 19616 1896
rect 18104 1856 19616 1884
rect 18104 1844 18110 1856
rect 19610 1844 19616 1856
rect 19668 1844 19674 1896
rect 20714 1844 20720 1896
rect 20772 1884 20778 1896
rect 21100 1884 21128 1915
rect 20772 1856 21128 1884
rect 20772 1844 20778 1856
rect 9732 1788 13676 1816
rect 13909 1819 13967 1825
rect 9732 1776 9738 1788
rect 13909 1785 13921 1819
rect 13955 1785 13967 1819
rect 13909 1779 13967 1785
rect 14185 1819 14243 1825
rect 14185 1785 14197 1819
rect 14231 1816 14243 1819
rect 15194 1816 15200 1828
rect 14231 1788 15200 1816
rect 14231 1785 14243 1788
rect 14185 1779 14243 1785
rect 15194 1776 15200 1788
rect 15252 1776 15258 1828
rect 16666 1776 16672 1828
rect 16724 1816 16730 1828
rect 16724 1788 17448 1816
rect 16724 1776 16730 1788
rect 8297 1751 8355 1757
rect 8297 1717 8309 1751
rect 8343 1717 8355 1751
rect 8297 1711 8355 1717
rect 8570 1708 8576 1760
rect 8628 1748 8634 1760
rect 8665 1751 8723 1757
rect 8665 1748 8677 1751
rect 8628 1720 8677 1748
rect 8628 1708 8634 1720
rect 8665 1717 8677 1720
rect 8711 1717 8723 1751
rect 8665 1711 8723 1717
rect 8846 1708 8852 1760
rect 8904 1748 8910 1760
rect 8941 1751 8999 1757
rect 8941 1748 8953 1751
rect 8904 1720 8953 1748
rect 8904 1708 8910 1720
rect 8941 1717 8953 1720
rect 8987 1717 8999 1751
rect 8941 1711 8999 1717
rect 9030 1708 9036 1760
rect 9088 1708 9094 1760
rect 10318 1708 10324 1760
rect 10376 1708 10382 1760
rect 11054 1708 11060 1760
rect 11112 1708 11118 1760
rect 11698 1708 11704 1760
rect 11756 1708 11762 1760
rect 11790 1708 11796 1760
rect 11848 1748 11854 1760
rect 11977 1751 12035 1757
rect 11977 1748 11989 1751
rect 11848 1720 11989 1748
rect 11848 1708 11854 1720
rect 11977 1717 11989 1720
rect 12023 1717 12035 1751
rect 11977 1711 12035 1717
rect 12618 1708 12624 1760
rect 12676 1708 12682 1760
rect 12894 1708 12900 1760
rect 12952 1708 12958 1760
rect 13357 1751 13415 1757
rect 13357 1717 13369 1751
rect 13403 1748 13415 1751
rect 13538 1748 13544 1760
rect 13403 1720 13544 1748
rect 13403 1717 13415 1720
rect 13357 1711 13415 1717
rect 13538 1708 13544 1720
rect 13596 1708 13602 1760
rect 13630 1708 13636 1760
rect 13688 1708 13694 1760
rect 14737 1751 14795 1757
rect 14737 1717 14749 1751
rect 14783 1748 14795 1751
rect 14918 1748 14924 1760
rect 14783 1720 14924 1748
rect 14783 1717 14795 1720
rect 14737 1711 14795 1717
rect 14918 1708 14924 1720
rect 14976 1708 14982 1760
rect 15286 1708 15292 1760
rect 15344 1748 15350 1760
rect 15565 1751 15623 1757
rect 15565 1748 15577 1751
rect 15344 1720 15577 1748
rect 15344 1708 15350 1720
rect 15565 1717 15577 1720
rect 15611 1717 15623 1751
rect 15565 1711 15623 1717
rect 16390 1708 16396 1760
rect 16448 1748 16454 1760
rect 17420 1757 17448 1788
rect 17494 1776 17500 1828
rect 17552 1816 17558 1828
rect 17552 1788 18920 1816
rect 17552 1776 17558 1788
rect 16853 1751 16911 1757
rect 16853 1748 16865 1751
rect 16448 1720 16865 1748
rect 16448 1708 16454 1720
rect 16853 1717 16865 1720
rect 16899 1717 16911 1751
rect 16853 1711 16911 1717
rect 17405 1751 17463 1757
rect 17405 1717 17417 1751
rect 17451 1717 17463 1751
rect 17405 1711 17463 1717
rect 17586 1708 17592 1760
rect 17644 1748 17650 1760
rect 17957 1751 18015 1757
rect 17957 1748 17969 1751
rect 17644 1720 17969 1748
rect 17644 1708 17650 1720
rect 17957 1717 17969 1720
rect 18003 1717 18015 1751
rect 17957 1711 18015 1717
rect 18046 1708 18052 1760
rect 18104 1748 18110 1760
rect 18892 1757 18920 1788
rect 19150 1776 19156 1828
rect 19208 1816 19214 1828
rect 19208 1788 20576 1816
rect 19208 1776 19214 1788
rect 18325 1751 18383 1757
rect 18325 1748 18337 1751
rect 18104 1720 18337 1748
rect 18104 1708 18110 1720
rect 18325 1717 18337 1720
rect 18371 1717 18383 1751
rect 18325 1711 18383 1717
rect 18877 1751 18935 1757
rect 18877 1717 18889 1751
rect 18923 1717 18935 1751
rect 18877 1711 18935 1717
rect 18966 1708 18972 1760
rect 19024 1748 19030 1760
rect 19429 1751 19487 1757
rect 19429 1748 19441 1751
rect 19024 1720 19441 1748
rect 19024 1708 19030 1720
rect 19429 1717 19441 1720
rect 19475 1717 19487 1751
rect 19429 1711 19487 1717
rect 19886 1708 19892 1760
rect 19944 1708 19950 1760
rect 20548 1757 20576 1788
rect 21174 1776 21180 1828
rect 21232 1776 21238 1828
rect 22112 1825 22140 1924
rect 22278 1912 22284 1964
rect 22336 1912 22342 1964
rect 22557 1955 22615 1961
rect 22557 1921 22569 1955
rect 22603 1952 22615 1955
rect 22646 1952 22652 1964
rect 22603 1924 22652 1952
rect 22603 1921 22615 1924
rect 22557 1915 22615 1921
rect 22646 1912 22652 1924
rect 22704 1912 22710 1964
rect 22756 1884 22784 1992
rect 22833 1955 22891 1961
rect 22833 1921 22845 1955
rect 22879 1952 22891 1955
rect 22940 1952 22968 2051
rect 23198 2048 23204 2100
rect 23256 2048 23262 2100
rect 23477 2091 23535 2097
rect 23477 2057 23489 2091
rect 23523 2088 23535 2091
rect 23934 2088 23940 2100
rect 23523 2060 23940 2088
rect 23523 2057 23535 2060
rect 23477 2051 23535 2057
rect 23934 2048 23940 2060
rect 23992 2048 23998 2100
rect 24029 2091 24087 2097
rect 24029 2057 24041 2091
rect 24075 2088 24087 2091
rect 24210 2088 24216 2100
rect 24075 2060 24216 2088
rect 24075 2057 24087 2060
rect 24029 2051 24087 2057
rect 24210 2048 24216 2060
rect 24268 2048 24274 2100
rect 23014 1980 23020 2032
rect 23072 2020 23078 2032
rect 23072 1992 24256 2020
rect 23072 1980 23078 1992
rect 22879 1924 22968 1952
rect 22879 1921 22891 1924
rect 22833 1915 22891 1921
rect 23106 1912 23112 1964
rect 23164 1912 23170 1964
rect 23382 1912 23388 1964
rect 23440 1912 23446 1964
rect 23661 1955 23719 1961
rect 23661 1921 23673 1955
rect 23707 1921 23719 1955
rect 23661 1915 23719 1921
rect 23676 1884 23704 1915
rect 23750 1912 23756 1964
rect 23808 1952 23814 1964
rect 24228 1961 24256 1992
rect 23937 1955 23995 1961
rect 23937 1952 23949 1955
rect 23808 1924 23949 1952
rect 23808 1912 23814 1924
rect 23937 1921 23949 1924
rect 23983 1921 23995 1955
rect 23937 1915 23995 1921
rect 24213 1955 24271 1961
rect 24213 1921 24225 1955
rect 24259 1921 24271 1955
rect 24213 1915 24271 1921
rect 22756 1856 23704 1884
rect 22097 1819 22155 1825
rect 22097 1785 22109 1819
rect 22143 1785 22155 1819
rect 23198 1816 23204 1828
rect 22097 1779 22155 1785
rect 22664 1788 23204 1816
rect 20533 1751 20591 1757
rect 20533 1717 20545 1751
rect 20579 1717 20591 1751
rect 20533 1711 20591 1717
rect 20806 1708 20812 1760
rect 20864 1748 20870 1760
rect 22664 1748 22692 1788
rect 23198 1776 23204 1788
rect 23256 1776 23262 1828
rect 23566 1776 23572 1828
rect 23624 1816 23630 1828
rect 23753 1819 23811 1825
rect 23753 1816 23765 1819
rect 23624 1788 23765 1816
rect 23624 1776 23630 1788
rect 23753 1785 23765 1788
rect 23799 1785 23811 1819
rect 23753 1779 23811 1785
rect 20864 1720 22692 1748
rect 20864 1708 20870 1720
rect 22738 1708 22744 1760
rect 22796 1748 22802 1760
rect 25222 1748 25228 1760
rect 22796 1720 25228 1748
rect 22796 1708 22802 1720
rect 25222 1708 25228 1720
rect 25280 1708 25286 1760
rect 1104 1658 24564 1680
rect 1104 1606 3882 1658
rect 3934 1606 3946 1658
rect 3998 1606 4010 1658
rect 4062 1606 4074 1658
rect 4126 1606 4138 1658
rect 4190 1606 9747 1658
rect 9799 1606 9811 1658
rect 9863 1606 9875 1658
rect 9927 1606 9939 1658
rect 9991 1606 10003 1658
rect 10055 1606 15612 1658
rect 15664 1606 15676 1658
rect 15728 1606 15740 1658
rect 15792 1606 15804 1658
rect 15856 1606 15868 1658
rect 15920 1606 21477 1658
rect 21529 1606 21541 1658
rect 21593 1606 21605 1658
rect 21657 1606 21669 1658
rect 21721 1606 21733 1658
rect 21785 1606 24564 1658
rect 1104 1584 24564 1606
rect 934 1504 940 1556
rect 992 1544 998 1556
rect 2406 1544 2412 1556
rect 992 1516 2412 1544
rect 992 1504 998 1516
rect 2406 1504 2412 1516
rect 2464 1504 2470 1556
rect 3053 1547 3111 1553
rect 3053 1513 3065 1547
rect 3099 1544 3111 1547
rect 4430 1544 4436 1556
rect 3099 1516 4436 1544
rect 3099 1513 3111 1516
rect 3053 1507 3111 1513
rect 4430 1504 4436 1516
rect 4488 1504 4494 1556
rect 5077 1547 5135 1553
rect 5077 1513 5089 1547
rect 5123 1544 5135 1547
rect 5718 1544 5724 1556
rect 5123 1516 5724 1544
rect 5123 1513 5135 1516
rect 5077 1507 5135 1513
rect 5718 1504 5724 1516
rect 5776 1504 5782 1556
rect 6086 1504 6092 1556
rect 6144 1544 6150 1556
rect 7377 1547 7435 1553
rect 6144 1516 7328 1544
rect 6144 1504 6150 1516
rect 3329 1479 3387 1485
rect 3329 1445 3341 1479
rect 3375 1476 3387 1479
rect 4338 1476 4344 1488
rect 3375 1448 4344 1476
rect 3375 1445 3387 1448
rect 3329 1439 3387 1445
rect 4338 1436 4344 1448
rect 4396 1436 4402 1488
rect 5534 1436 5540 1488
rect 5592 1476 5598 1488
rect 5592 1448 6868 1476
rect 5592 1436 5598 1448
rect 2130 1408 2136 1420
rect 1964 1380 2136 1408
rect 1489 1343 1547 1349
rect 1489 1309 1501 1343
rect 1535 1309 1547 1343
rect 1489 1303 1547 1309
rect 1765 1343 1823 1349
rect 1765 1309 1777 1343
rect 1811 1340 1823 1343
rect 1964 1340 1992 1380
rect 2130 1368 2136 1380
rect 2188 1368 2194 1420
rect 3712 1380 3924 1408
rect 1811 1312 1992 1340
rect 2041 1343 2099 1349
rect 1811 1309 1823 1312
rect 1765 1303 1823 1309
rect 2041 1309 2053 1343
rect 2087 1340 2099 1343
rect 2317 1343 2375 1349
rect 2087 1312 2268 1340
rect 2087 1309 2099 1312
rect 2041 1303 2099 1309
rect 1504 1272 1532 1303
rect 2240 1272 2268 1312
rect 2317 1309 2329 1343
rect 2363 1340 2375 1343
rect 2498 1340 2504 1352
rect 2363 1312 2504 1340
rect 2363 1309 2375 1312
rect 2317 1303 2375 1309
rect 2498 1300 2504 1312
rect 2556 1300 2562 1352
rect 2590 1300 2596 1352
rect 2648 1300 2654 1352
rect 2866 1300 2872 1352
rect 2924 1300 2930 1352
rect 3145 1343 3203 1349
rect 3145 1309 3157 1343
rect 3191 1309 3203 1343
rect 3145 1303 3203 1309
rect 3421 1343 3479 1349
rect 3421 1309 3433 1343
rect 3467 1340 3479 1343
rect 3712 1340 3740 1380
rect 3896 1352 3924 1380
rect 6288 1380 6500 1408
rect 3467 1312 3740 1340
rect 3789 1343 3847 1349
rect 3467 1309 3479 1312
rect 3421 1303 3479 1309
rect 3789 1309 3801 1343
rect 3835 1309 3847 1343
rect 3789 1303 3847 1309
rect 3160 1272 3188 1303
rect 3694 1272 3700 1284
rect 1504 1244 2084 1272
rect 2240 1244 2636 1272
rect 3160 1244 3700 1272
rect 2056 1216 2084 1244
rect 2608 1216 2636 1244
rect 3694 1232 3700 1244
rect 3752 1232 3758 1284
rect 3804 1272 3832 1303
rect 3878 1300 3884 1352
rect 3936 1300 3942 1352
rect 4065 1343 4123 1349
rect 4065 1309 4077 1343
rect 4111 1340 4123 1343
rect 4246 1340 4252 1352
rect 4111 1312 4252 1340
rect 4111 1309 4123 1312
rect 4065 1303 4123 1309
rect 4246 1300 4252 1312
rect 4304 1300 4310 1352
rect 4341 1343 4399 1349
rect 4341 1309 4353 1343
rect 4387 1340 4399 1343
rect 4522 1340 4528 1352
rect 4387 1312 4528 1340
rect 4387 1309 4399 1312
rect 4341 1303 4399 1309
rect 4522 1300 4528 1312
rect 4580 1300 4586 1352
rect 4617 1343 4675 1349
rect 4617 1309 4629 1343
rect 4663 1309 4675 1343
rect 4617 1303 4675 1309
rect 4154 1272 4160 1284
rect 3804 1244 4160 1272
rect 4154 1232 4160 1244
rect 4212 1232 4218 1284
rect 4632 1272 4660 1303
rect 4890 1300 4896 1352
rect 4948 1300 4954 1352
rect 5169 1343 5227 1349
rect 5169 1309 5181 1343
rect 5215 1309 5227 1343
rect 5169 1303 5227 1309
rect 5445 1343 5503 1349
rect 5445 1309 5457 1343
rect 5491 1340 5503 1343
rect 5626 1340 5632 1352
rect 5491 1312 5632 1340
rect 5491 1309 5503 1312
rect 5445 1303 5503 1309
rect 4982 1272 4988 1284
rect 4632 1244 4988 1272
rect 4982 1232 4988 1244
rect 5040 1232 5046 1284
rect 5184 1272 5212 1303
rect 5626 1300 5632 1312
rect 5684 1300 5690 1352
rect 5721 1343 5779 1349
rect 5721 1309 5733 1343
rect 5767 1309 5779 1343
rect 5721 1303 5779 1309
rect 5997 1343 6055 1349
rect 5997 1309 6009 1343
rect 6043 1340 6055 1343
rect 6288 1340 6316 1380
rect 6043 1312 6316 1340
rect 6043 1309 6055 1312
rect 5997 1303 6055 1309
rect 5534 1272 5540 1284
rect 5184 1244 5540 1272
rect 5534 1232 5540 1244
rect 5592 1232 5598 1284
rect 5736 1272 5764 1303
rect 6362 1300 6368 1352
rect 6420 1300 6426 1352
rect 6472 1340 6500 1380
rect 6546 1340 6552 1352
rect 6472 1312 6552 1340
rect 6546 1300 6552 1312
rect 6604 1300 6610 1352
rect 6638 1300 6644 1352
rect 6696 1300 6702 1352
rect 6730 1300 6736 1352
rect 6788 1300 6794 1352
rect 6840 1340 6868 1448
rect 7098 1436 7104 1488
rect 7156 1436 7162 1488
rect 7300 1476 7328 1516
rect 7377 1513 7389 1547
rect 7423 1544 7435 1547
rect 8110 1544 8116 1556
rect 7423 1516 8116 1544
rect 7423 1513 7435 1516
rect 7377 1507 7435 1513
rect 8110 1504 8116 1516
rect 8168 1504 8174 1556
rect 9398 1504 9404 1556
rect 9456 1544 9462 1556
rect 9456 1516 12434 1544
rect 9456 1504 9462 1516
rect 8662 1476 8668 1488
rect 7300 1448 8668 1476
rect 8662 1436 8668 1448
rect 8720 1436 8726 1488
rect 9030 1436 9036 1488
rect 9088 1436 9094 1488
rect 9493 1479 9551 1485
rect 9493 1445 9505 1479
rect 9539 1445 9551 1479
rect 12406 1476 12434 1516
rect 13906 1504 13912 1556
rect 13964 1544 13970 1556
rect 14645 1547 14703 1553
rect 14645 1544 14657 1547
rect 13964 1516 14657 1544
rect 13964 1504 13970 1516
rect 14645 1513 14657 1516
rect 14691 1513 14703 1547
rect 14645 1507 14703 1513
rect 14734 1504 14740 1556
rect 14792 1544 14798 1556
rect 15381 1547 15439 1553
rect 15381 1544 15393 1547
rect 14792 1516 15393 1544
rect 14792 1504 14798 1516
rect 15381 1513 15393 1516
rect 15427 1513 15439 1547
rect 15381 1507 15439 1513
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 14826 1476 14832 1488
rect 12406 1448 14832 1476
rect 9493 1439 9551 1445
rect 7116 1408 7144 1436
rect 9048 1408 9076 1436
rect 7116 1380 7788 1408
rect 6917 1343 6975 1349
rect 6917 1340 6929 1343
rect 6840 1312 6929 1340
rect 6917 1309 6929 1312
rect 6963 1309 6975 1343
rect 6917 1303 6975 1309
rect 7193 1343 7251 1349
rect 7193 1309 7205 1343
rect 7239 1309 7251 1343
rect 7193 1303 7251 1309
rect 6454 1272 6460 1284
rect 5736 1244 6460 1272
rect 6454 1232 6460 1244
rect 6512 1232 6518 1284
rect 1670 1164 1676 1216
rect 1728 1164 1734 1216
rect 1946 1164 1952 1216
rect 2004 1164 2010 1216
rect 2038 1164 2044 1216
rect 2096 1164 2102 1216
rect 2225 1207 2283 1213
rect 2225 1173 2237 1207
rect 2271 1204 2283 1207
rect 2406 1204 2412 1216
rect 2271 1176 2412 1204
rect 2271 1173 2283 1176
rect 2225 1167 2283 1173
rect 2406 1164 2412 1176
rect 2464 1164 2470 1216
rect 2498 1164 2504 1216
rect 2556 1164 2562 1216
rect 2590 1164 2596 1216
rect 2648 1164 2654 1216
rect 2777 1207 2835 1213
rect 2777 1173 2789 1207
rect 2823 1204 2835 1207
rect 3510 1204 3516 1216
rect 2823 1176 3516 1204
rect 2823 1173 2835 1176
rect 2777 1167 2835 1173
rect 3510 1164 3516 1176
rect 3568 1164 3574 1216
rect 3602 1164 3608 1216
rect 3660 1164 3666 1216
rect 3973 1207 4031 1213
rect 3973 1173 3985 1207
rect 4019 1204 4031 1207
rect 4062 1204 4068 1216
rect 4019 1176 4068 1204
rect 4019 1173 4031 1176
rect 3973 1167 4031 1173
rect 4062 1164 4068 1176
rect 4120 1164 4126 1216
rect 4246 1164 4252 1216
rect 4304 1164 4310 1216
rect 4522 1164 4528 1216
rect 4580 1164 4586 1216
rect 4798 1164 4804 1216
rect 4856 1164 4862 1216
rect 5350 1164 5356 1216
rect 5408 1164 5414 1216
rect 5626 1164 5632 1216
rect 5684 1164 5690 1216
rect 5905 1207 5963 1213
rect 5905 1173 5917 1207
rect 5951 1204 5963 1207
rect 6086 1204 6092 1216
rect 5951 1176 6092 1204
rect 5951 1173 5963 1176
rect 5905 1167 5963 1173
rect 6086 1164 6092 1176
rect 6144 1164 6150 1216
rect 6178 1164 6184 1216
rect 6236 1164 6242 1216
rect 6549 1207 6607 1213
rect 6549 1173 6561 1207
rect 6595 1204 6607 1207
rect 6638 1204 6644 1216
rect 6595 1176 6644 1204
rect 6595 1173 6607 1176
rect 6549 1167 6607 1173
rect 6638 1164 6644 1176
rect 6696 1164 6702 1216
rect 6748 1204 6776 1300
rect 7208 1272 7236 1303
rect 7466 1300 7472 1352
rect 7524 1300 7530 1352
rect 7760 1349 7788 1380
rect 8220 1380 9076 1408
rect 9508 1408 9536 1439
rect 14826 1436 14832 1448
rect 14884 1436 14890 1488
rect 14918 1436 14924 1488
rect 14976 1436 14982 1488
rect 15102 1436 15108 1488
rect 15160 1476 15166 1488
rect 15948 1476 15976 1507
rect 16298 1504 16304 1556
rect 16356 1504 16362 1556
rect 16942 1504 16948 1556
rect 17000 1544 17006 1556
rect 18509 1547 18567 1553
rect 18509 1544 18521 1547
rect 17000 1516 18521 1544
rect 17000 1504 17006 1516
rect 18509 1513 18521 1516
rect 18555 1513 18567 1547
rect 18509 1507 18567 1513
rect 19518 1504 19524 1556
rect 19576 1544 19582 1556
rect 19981 1547 20039 1553
rect 19981 1544 19993 1547
rect 19576 1516 19993 1544
rect 19576 1504 19582 1516
rect 19981 1513 19993 1516
rect 20027 1513 20039 1547
rect 19981 1507 20039 1513
rect 20533 1547 20591 1553
rect 20533 1513 20545 1547
rect 20579 1513 20591 1547
rect 20533 1507 20591 1513
rect 15160 1448 15976 1476
rect 15160 1436 15166 1448
rect 16022 1436 16028 1488
rect 16080 1476 16086 1488
rect 17497 1479 17555 1485
rect 17497 1476 17509 1479
rect 16080 1448 17509 1476
rect 16080 1436 16086 1448
rect 17497 1445 17509 1448
rect 17543 1445 17555 1479
rect 17497 1439 17555 1445
rect 18874 1436 18880 1488
rect 18932 1476 18938 1488
rect 20548 1476 20576 1507
rect 21818 1504 21824 1556
rect 21876 1504 21882 1556
rect 22278 1504 22284 1556
rect 22336 1544 22342 1556
rect 22649 1547 22707 1553
rect 22649 1544 22661 1547
rect 22336 1516 22661 1544
rect 22336 1504 22342 1516
rect 22649 1513 22661 1516
rect 22695 1513 22707 1547
rect 22649 1507 22707 1513
rect 22738 1504 22744 1556
rect 22796 1544 22802 1556
rect 23477 1547 23535 1553
rect 23477 1544 23489 1547
rect 22796 1516 23489 1544
rect 22796 1504 22802 1516
rect 23477 1513 23489 1516
rect 23523 1513 23535 1547
rect 23477 1507 23535 1513
rect 18932 1448 20576 1476
rect 21269 1479 21327 1485
rect 18932 1436 18938 1448
rect 21269 1445 21281 1479
rect 21315 1445 21327 1479
rect 21269 1439 21327 1445
rect 9508 1380 10088 1408
rect 7745 1343 7803 1349
rect 7745 1309 7757 1343
rect 7791 1309 7803 1343
rect 7745 1303 7803 1309
rect 7834 1300 7840 1352
rect 7892 1300 7898 1352
rect 8021 1343 8079 1349
rect 8021 1309 8033 1343
rect 8067 1340 8079 1343
rect 8220 1340 8248 1380
rect 8067 1312 8248 1340
rect 8297 1343 8355 1349
rect 8067 1309 8079 1312
rect 8021 1303 8079 1309
rect 8297 1309 8309 1343
rect 8343 1309 8355 1343
rect 8297 1303 8355 1309
rect 7852 1272 7880 1300
rect 8312 1272 8340 1303
rect 8570 1300 8576 1352
rect 8628 1300 8634 1352
rect 8662 1300 8668 1352
rect 8720 1340 8726 1352
rect 9033 1343 9091 1349
rect 9033 1340 9045 1343
rect 8720 1312 9045 1340
rect 8720 1300 8726 1312
rect 9033 1309 9045 1312
rect 9079 1309 9091 1343
rect 9033 1303 9091 1309
rect 9214 1300 9220 1352
rect 9272 1340 9278 1352
rect 9309 1343 9367 1349
rect 9309 1340 9321 1343
rect 9272 1312 9321 1340
rect 9272 1300 9278 1312
rect 9309 1309 9321 1312
rect 9355 1309 9367 1343
rect 9309 1303 9367 1309
rect 9398 1300 9404 1352
rect 9456 1340 9462 1352
rect 9585 1343 9643 1349
rect 9585 1340 9597 1343
rect 9456 1312 9597 1340
rect 9456 1300 9462 1312
rect 9585 1309 9597 1312
rect 9631 1309 9643 1343
rect 9585 1303 9643 1309
rect 9674 1300 9680 1352
rect 9732 1340 9738 1352
rect 9953 1343 10011 1349
rect 9953 1340 9965 1343
rect 9732 1312 9965 1340
rect 9732 1300 9738 1312
rect 9953 1309 9965 1312
rect 9999 1309 10011 1343
rect 10060 1340 10088 1380
rect 11054 1368 11060 1420
rect 11112 1368 11118 1420
rect 14936 1408 14964 1436
rect 14936 1380 16804 1408
rect 10321 1343 10379 1349
rect 10321 1340 10333 1343
rect 10060 1312 10333 1340
rect 9953 1303 10011 1309
rect 10321 1309 10333 1312
rect 10367 1309 10379 1343
rect 10321 1303 10379 1309
rect 11514 1300 11520 1352
rect 11572 1340 11578 1352
rect 11609 1343 11667 1349
rect 11609 1340 11621 1343
rect 11572 1312 11621 1340
rect 11572 1300 11578 1312
rect 11609 1309 11621 1312
rect 11655 1309 11667 1343
rect 11609 1303 11667 1309
rect 11882 1300 11888 1352
rect 11940 1340 11946 1352
rect 11977 1343 12035 1349
rect 11977 1340 11989 1343
rect 11940 1312 11989 1340
rect 11940 1300 11946 1312
rect 11977 1309 11989 1312
rect 12023 1309 12035 1343
rect 11977 1303 12035 1309
rect 12618 1300 12624 1352
rect 12676 1300 12682 1352
rect 13078 1300 13084 1352
rect 13136 1300 13142 1352
rect 13449 1343 13507 1349
rect 13449 1309 13461 1343
rect 13495 1309 13507 1343
rect 13449 1303 13507 1309
rect 9122 1272 9128 1284
rect 7208 1244 7788 1272
rect 7852 1244 8248 1272
rect 8312 1244 9128 1272
rect 7760 1216 7788 1244
rect 6825 1207 6883 1213
rect 6825 1204 6837 1207
rect 6748 1176 6837 1204
rect 6825 1173 6837 1176
rect 6871 1173 6883 1207
rect 6825 1167 6883 1173
rect 7101 1207 7159 1213
rect 7101 1173 7113 1207
rect 7147 1204 7159 1207
rect 7374 1204 7380 1216
rect 7147 1176 7380 1204
rect 7147 1173 7159 1176
rect 7101 1167 7159 1173
rect 7374 1164 7380 1176
rect 7432 1164 7438 1216
rect 7650 1164 7656 1216
rect 7708 1164 7714 1216
rect 7742 1164 7748 1216
rect 7800 1164 7806 1216
rect 7929 1207 7987 1213
rect 7929 1173 7941 1207
rect 7975 1204 7987 1207
rect 8110 1204 8116 1216
rect 7975 1176 8116 1204
rect 7975 1173 7987 1176
rect 7929 1167 7987 1173
rect 8110 1164 8116 1176
rect 8168 1164 8174 1216
rect 8220 1213 8248 1244
rect 9122 1232 9128 1244
rect 9180 1232 9186 1284
rect 10781 1275 10839 1281
rect 10781 1272 10793 1275
rect 9232 1244 10793 1272
rect 8205 1207 8263 1213
rect 8205 1173 8217 1207
rect 8251 1173 8263 1207
rect 8205 1167 8263 1173
rect 8478 1164 8484 1216
rect 8536 1164 8542 1216
rect 8757 1207 8815 1213
rect 8757 1173 8769 1207
rect 8803 1204 8815 1207
rect 9030 1204 9036 1216
rect 8803 1176 9036 1204
rect 8803 1173 8815 1176
rect 8757 1167 8815 1173
rect 9030 1164 9036 1176
rect 9088 1164 9094 1216
rect 9232 1213 9260 1244
rect 10781 1241 10793 1244
rect 10827 1241 10839 1275
rect 10781 1235 10839 1241
rect 11698 1232 11704 1284
rect 11756 1272 11762 1284
rect 12437 1275 12495 1281
rect 12437 1272 12449 1275
rect 11756 1244 12449 1272
rect 11756 1232 11762 1244
rect 12437 1241 12449 1244
rect 12483 1241 12495 1275
rect 12636 1272 12664 1300
rect 13464 1272 13492 1303
rect 13538 1300 13544 1352
rect 13596 1300 13602 1352
rect 13630 1300 13636 1352
rect 13688 1340 13694 1352
rect 14093 1343 14151 1349
rect 14093 1340 14105 1343
rect 13688 1312 14105 1340
rect 13688 1300 13694 1312
rect 14093 1309 14105 1312
rect 14139 1309 14151 1343
rect 14093 1303 14151 1309
rect 15194 1300 15200 1352
rect 15252 1340 15258 1352
rect 15289 1343 15347 1349
rect 15289 1340 15301 1343
rect 15252 1312 15301 1340
rect 15252 1300 15258 1312
rect 15289 1309 15301 1312
rect 15335 1309 15347 1343
rect 15289 1303 15347 1309
rect 15378 1300 15384 1352
rect 15436 1340 15442 1352
rect 15841 1343 15899 1349
rect 15841 1340 15853 1343
rect 15436 1312 15853 1340
rect 15436 1300 15442 1312
rect 15841 1309 15853 1312
rect 15887 1309 15899 1343
rect 15841 1303 15899 1309
rect 16114 1300 16120 1352
rect 16172 1340 16178 1352
rect 16776 1349 16804 1380
rect 17862 1368 17868 1420
rect 17920 1408 17926 1420
rect 19613 1411 19671 1417
rect 19613 1408 19625 1411
rect 17920 1380 19625 1408
rect 17920 1368 17926 1380
rect 19613 1377 19625 1380
rect 19659 1377 19671 1411
rect 19613 1371 19671 1377
rect 16485 1343 16543 1349
rect 16485 1340 16497 1343
rect 16172 1312 16497 1340
rect 16172 1300 16178 1312
rect 16485 1309 16497 1312
rect 16531 1309 16543 1343
rect 16485 1303 16543 1309
rect 16761 1343 16819 1349
rect 16761 1309 16773 1343
rect 16807 1309 16819 1343
rect 16761 1303 16819 1309
rect 16850 1300 16856 1352
rect 16908 1340 16914 1352
rect 16908 1312 17080 1340
rect 16908 1300 16914 1312
rect 12636 1244 13492 1272
rect 13556 1272 13584 1300
rect 14553 1275 14611 1281
rect 14553 1272 14565 1275
rect 13556 1244 14565 1272
rect 12437 1235 12495 1241
rect 14553 1241 14565 1244
rect 14599 1241 14611 1275
rect 14553 1235 14611 1241
rect 16298 1232 16304 1284
rect 16356 1272 16362 1284
rect 17052 1272 17080 1312
rect 17126 1300 17132 1352
rect 17184 1340 17190 1352
rect 17184 1312 17908 1340
rect 17184 1300 17190 1312
rect 17880 1281 17908 1312
rect 18138 1300 18144 1352
rect 18196 1340 18202 1352
rect 18417 1343 18475 1349
rect 18417 1340 18429 1343
rect 18196 1312 18429 1340
rect 18196 1300 18202 1312
rect 18417 1309 18429 1312
rect 18463 1309 18475 1343
rect 18417 1303 18475 1309
rect 18877 1343 18935 1349
rect 18877 1309 18889 1343
rect 18923 1309 18935 1343
rect 18877 1303 18935 1309
rect 17313 1275 17371 1281
rect 17313 1272 17325 1275
rect 16356 1244 16988 1272
rect 17052 1244 17325 1272
rect 16356 1232 16362 1244
rect 9217 1207 9275 1213
rect 9217 1173 9229 1207
rect 9263 1173 9275 1207
rect 9217 1167 9275 1173
rect 9769 1207 9827 1213
rect 9769 1173 9781 1207
rect 9815 1204 9827 1207
rect 10042 1204 10048 1216
rect 9815 1176 10048 1204
rect 9815 1173 9827 1176
rect 9769 1167 9827 1173
rect 10042 1164 10048 1176
rect 10100 1164 10106 1216
rect 10137 1207 10195 1213
rect 10137 1173 10149 1207
rect 10183 1204 10195 1207
rect 10410 1204 10416 1216
rect 10183 1176 10416 1204
rect 10183 1173 10195 1176
rect 10137 1167 10195 1173
rect 10410 1164 10416 1176
rect 10468 1164 10474 1216
rect 10505 1207 10563 1213
rect 10505 1173 10517 1207
rect 10551 1204 10563 1207
rect 11146 1204 11152 1216
rect 10551 1176 11152 1204
rect 10551 1173 10563 1176
rect 10505 1167 10563 1173
rect 11146 1164 11152 1176
rect 11204 1164 11210 1216
rect 11790 1164 11796 1216
rect 11848 1164 11854 1216
rect 12158 1164 12164 1216
rect 12216 1164 12222 1216
rect 12526 1164 12532 1216
rect 12584 1164 12590 1216
rect 13170 1164 13176 1216
rect 13228 1204 13234 1216
rect 13265 1207 13323 1213
rect 13265 1204 13277 1207
rect 13228 1176 13277 1204
rect 13228 1164 13234 1176
rect 13265 1173 13277 1176
rect 13311 1173 13323 1207
rect 13265 1167 13323 1173
rect 13354 1164 13360 1216
rect 13412 1204 13418 1216
rect 13633 1207 13691 1213
rect 13633 1204 13645 1207
rect 13412 1176 13645 1204
rect 13412 1164 13418 1176
rect 13633 1173 13645 1176
rect 13679 1173 13691 1207
rect 13633 1167 13691 1173
rect 13906 1164 13912 1216
rect 13964 1204 13970 1216
rect 14277 1207 14335 1213
rect 14277 1204 14289 1207
rect 13964 1176 14289 1204
rect 13964 1164 13970 1176
rect 14277 1173 14289 1176
rect 14323 1173 14335 1207
rect 14277 1167 14335 1173
rect 15010 1164 15016 1216
rect 15068 1204 15074 1216
rect 16853 1207 16911 1213
rect 16853 1204 16865 1207
rect 15068 1176 16865 1204
rect 15068 1164 15074 1176
rect 16853 1173 16865 1176
rect 16899 1173 16911 1207
rect 16960 1204 16988 1244
rect 17313 1241 17325 1244
rect 17359 1241 17371 1275
rect 17313 1235 17371 1241
rect 17865 1275 17923 1281
rect 17865 1241 17877 1275
rect 17911 1241 17923 1275
rect 17865 1235 17923 1241
rect 18230 1232 18236 1284
rect 18288 1272 18294 1284
rect 18892 1272 18920 1303
rect 19242 1300 19248 1352
rect 19300 1340 19306 1352
rect 19300 1312 19472 1340
rect 19300 1300 19306 1312
rect 19337 1275 19395 1281
rect 19337 1272 19349 1275
rect 18288 1244 18920 1272
rect 19076 1244 19349 1272
rect 18288 1232 18294 1244
rect 19076 1213 19104 1244
rect 19337 1241 19349 1244
rect 19383 1241 19395 1275
rect 19337 1235 19395 1241
rect 17957 1207 18015 1213
rect 17957 1204 17969 1207
rect 16960 1176 17969 1204
rect 16853 1167 16911 1173
rect 17957 1173 17969 1176
rect 18003 1173 18015 1207
rect 17957 1167 18015 1173
rect 19061 1207 19119 1213
rect 19061 1173 19073 1207
rect 19107 1173 19119 1207
rect 19444 1204 19472 1312
rect 19518 1300 19524 1352
rect 19576 1340 19582 1352
rect 21177 1343 21235 1349
rect 19576 1312 20576 1340
rect 19576 1300 19582 1312
rect 19610 1232 19616 1284
rect 19668 1272 19674 1284
rect 19889 1275 19947 1281
rect 19889 1272 19901 1275
rect 19668 1244 19901 1272
rect 19668 1232 19674 1244
rect 19889 1241 19901 1244
rect 19935 1241 19947 1275
rect 19889 1235 19947 1241
rect 20441 1275 20499 1281
rect 20441 1241 20453 1275
rect 20487 1241 20499 1275
rect 20441 1235 20499 1241
rect 20456 1204 20484 1235
rect 19444 1176 20484 1204
rect 20548 1204 20576 1312
rect 21177 1309 21189 1343
rect 21223 1340 21235 1343
rect 21284 1340 21312 1439
rect 22094 1436 22100 1488
rect 22152 1476 22158 1488
rect 23382 1476 23388 1488
rect 22152 1448 23388 1476
rect 22152 1436 22158 1448
rect 23382 1436 23388 1448
rect 23440 1436 23446 1488
rect 23566 1436 23572 1488
rect 23624 1476 23630 1488
rect 24946 1476 24952 1488
rect 23624 1448 24952 1476
rect 23624 1436 23630 1448
rect 24946 1436 24952 1448
rect 25004 1436 25010 1488
rect 21358 1368 21364 1420
rect 21416 1408 21422 1420
rect 21416 1380 22416 1408
rect 21416 1368 21422 1380
rect 21223 1312 21312 1340
rect 21223 1309 21235 1312
rect 21177 1303 21235 1309
rect 21450 1300 21456 1352
rect 21508 1300 21514 1352
rect 21542 1300 21548 1352
rect 21600 1340 21606 1352
rect 22005 1343 22063 1349
rect 22005 1340 22017 1343
rect 21600 1312 22017 1340
rect 21600 1300 21606 1312
rect 22005 1309 22017 1312
rect 22051 1309 22063 1343
rect 22005 1303 22063 1309
rect 22281 1343 22339 1349
rect 22281 1309 22293 1343
rect 22327 1309 22339 1343
rect 22281 1303 22339 1309
rect 20622 1232 20628 1284
rect 20680 1272 20686 1284
rect 20680 1244 21404 1272
rect 20680 1232 20686 1244
rect 20993 1207 21051 1213
rect 20993 1204 21005 1207
rect 20548 1176 21005 1204
rect 19061 1167 19119 1173
rect 20993 1173 21005 1176
rect 21039 1173 21051 1207
rect 21376 1204 21404 1244
rect 21726 1232 21732 1284
rect 21784 1272 21790 1284
rect 22296 1272 22324 1303
rect 21784 1244 22324 1272
rect 22388 1272 22416 1380
rect 22738 1368 22744 1420
rect 22796 1408 22802 1420
rect 23750 1408 23756 1420
rect 22796 1380 23756 1408
rect 22796 1368 22802 1380
rect 23750 1368 23756 1380
rect 23808 1368 23814 1420
rect 22554 1300 22560 1352
rect 22612 1300 22618 1352
rect 22646 1300 22652 1352
rect 22704 1340 22710 1352
rect 22833 1343 22891 1349
rect 22833 1340 22845 1343
rect 22704 1312 22845 1340
rect 22704 1300 22710 1312
rect 22833 1309 22845 1312
rect 22879 1309 22891 1343
rect 22833 1303 22891 1309
rect 23109 1343 23167 1349
rect 23109 1309 23121 1343
rect 23155 1309 23167 1343
rect 23109 1303 23167 1309
rect 23124 1272 23152 1303
rect 23198 1300 23204 1352
rect 23256 1340 23262 1352
rect 23385 1343 23443 1349
rect 23385 1340 23397 1343
rect 23256 1312 23397 1340
rect 23256 1300 23262 1312
rect 23385 1309 23397 1312
rect 23431 1309 23443 1343
rect 23385 1303 23443 1309
rect 23658 1300 23664 1352
rect 23716 1300 23722 1352
rect 23934 1300 23940 1352
rect 23992 1300 23998 1352
rect 24026 1300 24032 1352
rect 24084 1340 24090 1352
rect 24213 1343 24271 1349
rect 24213 1340 24225 1343
rect 24084 1312 24225 1340
rect 24084 1300 24090 1312
rect 24213 1309 24225 1312
rect 24259 1309 24271 1343
rect 24213 1303 24271 1309
rect 24854 1300 24860 1352
rect 24912 1300 24918 1352
rect 22388 1244 23152 1272
rect 21784 1232 21790 1244
rect 22097 1207 22155 1213
rect 22097 1204 22109 1207
rect 21376 1176 22109 1204
rect 20993 1167 21051 1173
rect 22097 1173 22109 1176
rect 22143 1173 22155 1207
rect 22097 1167 22155 1173
rect 22186 1164 22192 1216
rect 22244 1204 22250 1216
rect 22373 1207 22431 1213
rect 22373 1204 22385 1207
rect 22244 1176 22385 1204
rect 22244 1164 22250 1176
rect 22373 1173 22385 1176
rect 22419 1173 22431 1207
rect 22373 1167 22431 1173
rect 22922 1164 22928 1216
rect 22980 1164 22986 1216
rect 23198 1164 23204 1216
rect 23256 1164 23262 1216
rect 23750 1164 23756 1216
rect 23808 1164 23814 1216
rect 24029 1207 24087 1213
rect 24029 1173 24041 1207
rect 24075 1204 24087 1207
rect 24872 1204 24900 1300
rect 24075 1176 24900 1204
rect 24075 1173 24087 1176
rect 24029 1167 24087 1173
rect 1104 1114 24723 1136
rect 1104 1062 6814 1114
rect 6866 1062 6878 1114
rect 6930 1062 6942 1114
rect 6994 1062 7006 1114
rect 7058 1062 7070 1114
rect 7122 1062 12679 1114
rect 12731 1062 12743 1114
rect 12795 1062 12807 1114
rect 12859 1062 12871 1114
rect 12923 1062 12935 1114
rect 12987 1062 18544 1114
rect 18596 1062 18608 1114
rect 18660 1062 18672 1114
rect 18724 1062 18736 1114
rect 18788 1062 18800 1114
rect 18852 1062 24409 1114
rect 24461 1062 24473 1114
rect 24525 1062 24537 1114
rect 24589 1062 24601 1114
rect 24653 1062 24665 1114
rect 24717 1062 24723 1114
rect 1104 1040 24723 1062
rect 2498 960 2504 1012
rect 2556 960 2562 1012
rect 7374 960 7380 1012
rect 7432 960 7438 1012
rect 7650 960 7656 1012
rect 7708 1000 7714 1012
rect 7708 972 12434 1000
rect 7708 960 7714 972
rect 2516 728 2544 960
rect 7392 932 7420 960
rect 9398 932 9404 944
rect 7392 904 9404 932
rect 9398 892 9404 904
rect 9456 892 9462 944
rect 10502 892 10508 944
rect 10560 892 10566 944
rect 4522 824 4528 876
rect 4580 864 4586 876
rect 8018 864 8024 876
rect 4580 836 8024 864
rect 4580 824 4586 836
rect 8018 824 8024 836
rect 8076 824 8082 876
rect 10520 864 10548 892
rect 8128 836 10548 864
rect 12406 864 12434 972
rect 19978 960 19984 1012
rect 20036 1000 20042 1012
rect 21542 1000 21548 1012
rect 20036 972 21548 1000
rect 20036 960 20042 972
rect 21542 960 21548 972
rect 21600 960 21606 1012
rect 22554 1000 22560 1012
rect 22066 972 22560 1000
rect 20530 892 20536 944
rect 20588 932 20594 944
rect 22066 932 22094 972
rect 22554 960 22560 972
rect 22612 960 22618 1012
rect 23750 960 23756 1012
rect 23808 960 23814 1012
rect 23934 960 23940 1012
rect 23992 960 23998 1012
rect 20588 904 22094 932
rect 20588 892 20594 904
rect 16758 864 16764 876
rect 12406 836 16764 864
rect 3602 756 3608 808
rect 3660 796 3666 808
rect 8128 796 8156 836
rect 16758 824 16764 836
rect 16816 824 16822 876
rect 23768 864 23796 960
rect 17052 836 23796 864
rect 3660 768 8156 796
rect 3660 756 3666 768
rect 9030 756 9036 808
rect 9088 796 9094 808
rect 16114 796 16120 808
rect 9088 768 16120 796
rect 9088 756 9094 768
rect 16114 756 16120 768
rect 16172 756 16178 808
rect 2516 700 12434 728
rect 2682 620 2688 672
rect 2740 660 2746 672
rect 3142 660 3148 672
rect 2740 632 3148 660
rect 2740 620 2746 632
rect 3142 620 3148 632
rect 3200 620 3206 672
rect 6362 620 6368 672
rect 6420 660 6426 672
rect 7006 660 7012 672
rect 6420 632 7012 660
rect 6420 620 6426 632
rect 7006 620 7012 632
rect 7064 620 7070 672
rect 7466 620 7472 672
rect 7524 660 7530 672
rect 8110 660 8116 672
rect 7524 632 8116 660
rect 7524 620 7530 632
rect 8110 620 8116 632
rect 8168 620 8174 672
rect 8570 620 8576 672
rect 8628 660 8634 672
rect 9582 660 9588 672
rect 8628 632 9588 660
rect 8628 620 8634 632
rect 9582 620 9588 632
rect 9640 620 9646 672
rect 12066 620 12072 672
rect 12124 620 12130 672
rect 3510 552 3516 604
rect 3568 592 3574 604
rect 12084 592 12112 620
rect 3568 564 12112 592
rect 12406 604 12434 700
rect 14090 688 14096 740
rect 14148 728 14154 740
rect 17052 728 17080 836
rect 21358 756 21364 808
rect 21416 796 21422 808
rect 23106 796 23112 808
rect 21416 768 23112 796
rect 21416 756 21422 768
rect 23106 756 23112 768
rect 23164 756 23170 808
rect 14148 700 17080 728
rect 14148 688 14154 700
rect 21634 688 21640 740
rect 21692 728 21698 740
rect 23952 728 23980 960
rect 21692 700 23980 728
rect 21692 688 21698 700
rect 16482 620 16488 672
rect 16540 660 16546 672
rect 16540 632 18368 660
rect 16540 620 16546 632
rect 12406 564 12440 604
rect 3568 552 3574 564
rect 12434 552 12440 564
rect 12492 552 12498 604
rect 18230 552 18236 604
rect 18288 552 18294 604
rect 6638 484 6644 536
rect 6696 524 6702 536
rect 17678 524 17684 536
rect 6696 496 17684 524
rect 6696 484 6702 496
rect 17678 484 17684 496
rect 17736 484 17742 536
rect 8202 416 8208 468
rect 8260 456 8266 468
rect 18248 456 18276 552
rect 18340 524 18368 632
rect 18414 620 18420 672
rect 18472 660 18478 672
rect 19242 660 19248 672
rect 18472 632 19248 660
rect 18472 620 18478 632
rect 19242 620 19248 632
rect 19300 620 19306 672
rect 20898 620 20904 672
rect 20956 660 20962 672
rect 22646 660 22652 672
rect 20956 632 22652 660
rect 20956 620 20962 632
rect 22646 620 22652 632
rect 22704 620 22710 672
rect 23198 620 23204 672
rect 23256 620 23262 672
rect 20438 552 20444 604
rect 20496 592 20502 604
rect 21726 592 21732 604
rect 20496 564 21732 592
rect 20496 552 20502 564
rect 21726 552 21732 564
rect 21784 552 21790 604
rect 23216 524 23244 620
rect 18340 496 23244 524
rect 8260 428 18276 456
rect 8260 416 8266 428
rect 18874 416 18880 468
rect 18932 416 18938 468
rect 4246 348 4252 400
rect 4304 388 4310 400
rect 8294 388 8300 400
rect 4304 360 8300 388
rect 4304 348 4310 360
rect 8294 348 8300 360
rect 8352 348 8358 400
rect 8478 348 8484 400
rect 8536 388 8542 400
rect 15930 388 15936 400
rect 8536 360 15936 388
rect 8536 348 8542 360
rect 15930 348 15936 360
rect 15988 348 15994 400
rect 2406 280 2412 332
rect 2464 320 2470 332
rect 13446 320 13452 332
rect 2464 292 13452 320
rect 2464 280 2470 292
rect 13446 280 13452 292
rect 13504 280 13510 332
rect 18892 264 18920 416
rect 22738 348 22744 400
rect 22796 388 22802 400
rect 23014 388 23020 400
rect 22796 360 23020 388
rect 22796 348 22802 360
rect 23014 348 23020 360
rect 23072 348 23078 400
rect 1946 212 1952 264
rect 2004 252 2010 264
rect 2004 224 12434 252
rect 2004 212 2010 224
rect 4062 144 4068 196
rect 4120 184 4126 196
rect 9398 184 9404 196
rect 4120 156 9404 184
rect 4120 144 4126 156
rect 9398 144 9404 156
rect 9456 144 9462 196
rect 4982 76 4988 128
rect 5040 116 5046 128
rect 5534 116 5540 128
rect 5040 88 5540 116
rect 5040 76 5046 88
rect 5534 76 5540 88
rect 5592 76 5598 128
rect 12406 116 12434 224
rect 18874 212 18880 264
rect 18932 212 18938 264
rect 13262 116 13268 128
rect 12406 88 13268 116
rect 13262 76 13268 88
rect 13320 76 13326 128
<< via1 >>
rect 6814 8678 6866 8730
rect 6878 8678 6930 8730
rect 6942 8678 6994 8730
rect 7006 8678 7058 8730
rect 7070 8678 7122 8730
rect 12679 8678 12731 8730
rect 12743 8678 12795 8730
rect 12807 8678 12859 8730
rect 12871 8678 12923 8730
rect 12935 8678 12987 8730
rect 18544 8678 18596 8730
rect 18608 8678 18660 8730
rect 18672 8678 18724 8730
rect 18736 8678 18788 8730
rect 18800 8678 18852 8730
rect 24409 8678 24461 8730
rect 24473 8678 24525 8730
rect 24537 8678 24589 8730
rect 24601 8678 24653 8730
rect 24665 8678 24717 8730
rect 2044 8576 2096 8628
rect 3240 8576 3292 8628
rect 4436 8576 4488 8628
rect 5632 8576 5684 8628
rect 6736 8576 6788 8628
rect 8024 8576 8076 8628
rect 9220 8576 9272 8628
rect 10416 8576 10468 8628
rect 11612 8576 11664 8628
rect 13084 8619 13136 8628
rect 13084 8585 13093 8619
rect 13093 8585 13127 8619
rect 13127 8585 13136 8619
rect 13084 8576 13136 8585
rect 14004 8576 14056 8628
rect 15200 8576 15252 8628
rect 1400 8551 1452 8560
rect 1400 8517 1409 8551
rect 1409 8517 1443 8551
rect 1443 8517 1452 8551
rect 1400 8508 1452 8517
rect 16396 8508 16448 8560
rect 17592 8576 17644 8628
rect 18880 8576 18932 8628
rect 19984 8576 20036 8628
rect 21180 8576 21232 8628
rect 22376 8576 22428 8628
rect 23572 8576 23624 8628
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 2412 8483 2464 8492
rect 2412 8449 2421 8483
rect 2421 8449 2455 8483
rect 2455 8449 2464 8483
rect 2412 8440 2464 8449
rect 3608 8483 3660 8492
rect 3608 8449 3617 8483
rect 3617 8449 3651 8483
rect 3651 8449 3660 8483
rect 3608 8440 3660 8449
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5816 8483 5868 8492
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 9312 8483 9364 8492
rect 9312 8449 9321 8483
rect 9321 8449 9355 8483
rect 9355 8449 9364 8483
rect 9312 8440 9364 8449
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 13176 8440 13228 8492
rect 14096 8483 14148 8492
rect 14096 8449 14105 8483
rect 14105 8449 14139 8483
rect 14139 8449 14148 8483
rect 14096 8440 14148 8449
rect 15384 8483 15436 8492
rect 15384 8449 15393 8483
rect 15393 8449 15427 8483
rect 15427 8449 15436 8483
rect 15384 8440 15436 8449
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 24860 8508 24912 8560
rect 19248 8440 19300 8492
rect 22008 8440 22060 8492
rect 22560 8372 22612 8424
rect 23480 8483 23532 8492
rect 23480 8449 23489 8483
rect 23489 8449 23523 8483
rect 23523 8449 23532 8483
rect 23480 8440 23532 8449
rect 23756 8483 23808 8492
rect 23756 8449 23765 8483
rect 23765 8449 23799 8483
rect 23799 8449 23808 8483
rect 23756 8440 23808 8449
rect 24768 8372 24820 8424
rect 23940 8304 23992 8356
rect 3882 8134 3934 8186
rect 3946 8134 3998 8186
rect 4010 8134 4062 8186
rect 4074 8134 4126 8186
rect 4138 8134 4190 8186
rect 9747 8134 9799 8186
rect 9811 8134 9863 8186
rect 9875 8134 9927 8186
rect 9939 8134 9991 8186
rect 10003 8134 10055 8186
rect 15612 8134 15664 8186
rect 15676 8134 15728 8186
rect 15740 8134 15792 8186
rect 15804 8134 15856 8186
rect 15868 8134 15920 8186
rect 21477 8134 21529 8186
rect 21541 8134 21593 8186
rect 21605 8134 21657 8186
rect 21669 8134 21721 8186
rect 21733 8134 21785 8186
rect 17408 8032 17460 8084
rect 17132 7828 17184 7880
rect 6814 7590 6866 7642
rect 6878 7590 6930 7642
rect 6942 7590 6994 7642
rect 7006 7590 7058 7642
rect 7070 7590 7122 7642
rect 12679 7590 12731 7642
rect 12743 7590 12795 7642
rect 12807 7590 12859 7642
rect 12871 7590 12923 7642
rect 12935 7590 12987 7642
rect 18544 7590 18596 7642
rect 18608 7590 18660 7642
rect 18672 7590 18724 7642
rect 18736 7590 18788 7642
rect 18800 7590 18852 7642
rect 24409 7590 24461 7642
rect 24473 7590 24525 7642
rect 24537 7590 24589 7642
rect 24601 7590 24653 7642
rect 24665 7590 24717 7642
rect 3882 7046 3934 7098
rect 3946 7046 3998 7098
rect 4010 7046 4062 7098
rect 4074 7046 4126 7098
rect 4138 7046 4190 7098
rect 9747 7046 9799 7098
rect 9811 7046 9863 7098
rect 9875 7046 9927 7098
rect 9939 7046 9991 7098
rect 10003 7046 10055 7098
rect 15612 7046 15664 7098
rect 15676 7046 15728 7098
rect 15740 7046 15792 7098
rect 15804 7046 15856 7098
rect 15868 7046 15920 7098
rect 21477 7046 21529 7098
rect 21541 7046 21593 7098
rect 21605 7046 21657 7098
rect 21669 7046 21721 7098
rect 21733 7046 21785 7098
rect 6814 6502 6866 6554
rect 6878 6502 6930 6554
rect 6942 6502 6994 6554
rect 7006 6502 7058 6554
rect 7070 6502 7122 6554
rect 12679 6502 12731 6554
rect 12743 6502 12795 6554
rect 12807 6502 12859 6554
rect 12871 6502 12923 6554
rect 12935 6502 12987 6554
rect 18544 6502 18596 6554
rect 18608 6502 18660 6554
rect 18672 6502 18724 6554
rect 18736 6502 18788 6554
rect 18800 6502 18852 6554
rect 24409 6502 24461 6554
rect 24473 6502 24525 6554
rect 24537 6502 24589 6554
rect 24601 6502 24653 6554
rect 24665 6502 24717 6554
rect 3882 5958 3934 6010
rect 3946 5958 3998 6010
rect 4010 5958 4062 6010
rect 4074 5958 4126 6010
rect 4138 5958 4190 6010
rect 9747 5958 9799 6010
rect 9811 5958 9863 6010
rect 9875 5958 9927 6010
rect 9939 5958 9991 6010
rect 10003 5958 10055 6010
rect 15612 5958 15664 6010
rect 15676 5958 15728 6010
rect 15740 5958 15792 6010
rect 15804 5958 15856 6010
rect 15868 5958 15920 6010
rect 21477 5958 21529 6010
rect 21541 5958 21593 6010
rect 21605 5958 21657 6010
rect 21669 5958 21721 6010
rect 21733 5958 21785 6010
rect 6814 5414 6866 5466
rect 6878 5414 6930 5466
rect 6942 5414 6994 5466
rect 7006 5414 7058 5466
rect 7070 5414 7122 5466
rect 12679 5414 12731 5466
rect 12743 5414 12795 5466
rect 12807 5414 12859 5466
rect 12871 5414 12923 5466
rect 12935 5414 12987 5466
rect 18544 5414 18596 5466
rect 18608 5414 18660 5466
rect 18672 5414 18724 5466
rect 18736 5414 18788 5466
rect 18800 5414 18852 5466
rect 24409 5414 24461 5466
rect 24473 5414 24525 5466
rect 24537 5414 24589 5466
rect 24601 5414 24653 5466
rect 24665 5414 24717 5466
rect 3882 4870 3934 4922
rect 3946 4870 3998 4922
rect 4010 4870 4062 4922
rect 4074 4870 4126 4922
rect 4138 4870 4190 4922
rect 9747 4870 9799 4922
rect 9811 4870 9863 4922
rect 9875 4870 9927 4922
rect 9939 4870 9991 4922
rect 10003 4870 10055 4922
rect 15612 4870 15664 4922
rect 15676 4870 15728 4922
rect 15740 4870 15792 4922
rect 15804 4870 15856 4922
rect 15868 4870 15920 4922
rect 21477 4870 21529 4922
rect 21541 4870 21593 4922
rect 21605 4870 21657 4922
rect 21669 4870 21721 4922
rect 21733 4870 21785 4922
rect 6814 4326 6866 4378
rect 6878 4326 6930 4378
rect 6942 4326 6994 4378
rect 7006 4326 7058 4378
rect 7070 4326 7122 4378
rect 12679 4326 12731 4378
rect 12743 4326 12795 4378
rect 12807 4326 12859 4378
rect 12871 4326 12923 4378
rect 12935 4326 12987 4378
rect 18544 4326 18596 4378
rect 18608 4326 18660 4378
rect 18672 4326 18724 4378
rect 18736 4326 18788 4378
rect 18800 4326 18852 4378
rect 24409 4326 24461 4378
rect 24473 4326 24525 4378
rect 24537 4326 24589 4378
rect 24601 4326 24653 4378
rect 24665 4326 24717 4378
rect 9496 4131 9548 4140
rect 9496 4097 9505 4131
rect 9505 4097 9539 4131
rect 9539 4097 9548 4131
rect 9496 4088 9548 4097
rect 10692 4131 10744 4140
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 11888 4131 11940 4140
rect 11888 4097 11897 4131
rect 11897 4097 11931 4131
rect 11931 4097 11940 4131
rect 11888 4088 11940 4097
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 19984 4131 20036 4140
rect 19984 4097 19993 4131
rect 19993 4097 20027 4131
rect 20027 4097 20036 4131
rect 19984 4088 20036 4097
rect 24032 4131 24084 4140
rect 24032 4097 24041 4131
rect 24041 4097 24075 4131
rect 24075 4097 24084 4131
rect 24032 4088 24084 4097
rect 22744 4020 22796 4072
rect 19800 3995 19852 4004
rect 19800 3961 19809 3995
rect 19809 3961 19843 3995
rect 19843 3961 19852 3995
rect 19800 3952 19852 3961
rect 9312 3927 9364 3936
rect 9312 3893 9321 3927
rect 9321 3893 9355 3927
rect 9355 3893 9364 3927
rect 9312 3884 9364 3893
rect 10508 3927 10560 3936
rect 10508 3893 10517 3927
rect 10517 3893 10551 3927
rect 10551 3893 10560 3927
rect 10508 3884 10560 3893
rect 10784 3884 10836 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 13176 3884 13228 3936
rect 23480 3884 23532 3936
rect 3882 3782 3934 3834
rect 3946 3782 3998 3834
rect 4010 3782 4062 3834
rect 4074 3782 4126 3834
rect 4138 3782 4190 3834
rect 9747 3782 9799 3834
rect 9811 3782 9863 3834
rect 9875 3782 9927 3834
rect 9939 3782 9991 3834
rect 10003 3782 10055 3834
rect 15612 3782 15664 3834
rect 15676 3782 15728 3834
rect 15740 3782 15792 3834
rect 15804 3782 15856 3834
rect 15868 3782 15920 3834
rect 21477 3782 21529 3834
rect 21541 3782 21593 3834
rect 21605 3782 21657 3834
rect 21669 3782 21721 3834
rect 21733 3782 21785 3834
rect 9496 3723 9548 3732
rect 9496 3689 9505 3723
rect 9505 3689 9539 3723
rect 9539 3689 9548 3723
rect 9496 3680 9548 3689
rect 10692 3680 10744 3732
rect 11888 3680 11940 3732
rect 13084 3680 13136 3732
rect 14096 3723 14148 3732
rect 14096 3689 14105 3723
rect 14105 3689 14139 3723
rect 14139 3689 14148 3723
rect 14096 3680 14148 3689
rect 15384 3680 15436 3732
rect 19984 3723 20036 3732
rect 19984 3689 19993 3723
rect 19993 3689 20027 3723
rect 20027 3689 20036 3723
rect 19984 3680 20036 3689
rect 24032 3723 24084 3732
rect 24032 3689 24041 3723
rect 24041 3689 24075 3723
rect 24075 3689 24084 3723
rect 24032 3680 24084 3689
rect 23204 3612 23256 3664
rect 10600 3476 10652 3528
rect 10784 3519 10836 3528
rect 10784 3485 10793 3519
rect 10793 3485 10827 3519
rect 10827 3485 10836 3519
rect 10784 3476 10836 3485
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 19524 3544 19576 3596
rect 24216 3612 24268 3664
rect 15476 3519 15528 3528
rect 15476 3485 15485 3519
rect 15485 3485 15519 3519
rect 15519 3485 15528 3519
rect 15476 3476 15528 3485
rect 20628 3476 20680 3528
rect 23296 3476 23348 3528
rect 24308 3544 24360 3596
rect 19892 3340 19944 3392
rect 23480 3340 23532 3392
rect 6814 3238 6866 3290
rect 6878 3238 6930 3290
rect 6942 3238 6994 3290
rect 7006 3238 7058 3290
rect 7070 3238 7122 3290
rect 12679 3238 12731 3290
rect 12743 3238 12795 3290
rect 12807 3238 12859 3290
rect 12871 3238 12923 3290
rect 12935 3238 12987 3290
rect 18544 3238 18596 3290
rect 18608 3238 18660 3290
rect 18672 3238 18724 3290
rect 18736 3238 18788 3290
rect 18800 3238 18852 3290
rect 24409 3238 24461 3290
rect 24473 3238 24525 3290
rect 24537 3238 24589 3290
rect 24601 3238 24653 3290
rect 24665 3238 24717 3290
rect 8208 3136 8260 3188
rect 15476 3136 15528 3188
rect 6644 3068 6696 3120
rect 16488 3068 16540 3120
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 9588 3000 9640 3052
rect 19892 3136 19944 3188
rect 22744 3179 22796 3188
rect 22744 3145 22753 3179
rect 22753 3145 22787 3179
rect 22787 3145 22796 3179
rect 22744 3136 22796 3145
rect 23664 3136 23716 3188
rect 19524 3068 19576 3120
rect 9128 2932 9180 2984
rect 12256 2932 12308 2984
rect 14372 2932 14424 2984
rect 7840 2864 7892 2916
rect 16672 2864 16724 2916
rect 22652 3043 22704 3052
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 22376 2932 22428 2984
rect 23020 3043 23072 3052
rect 23020 3009 23029 3043
rect 23029 3009 23063 3043
rect 23063 3009 23072 3043
rect 23020 3000 23072 3009
rect 25504 3068 25556 3120
rect 23848 3000 23900 3052
rect 23388 2932 23440 2984
rect 8852 2796 8904 2848
rect 14096 2796 14148 2848
rect 19892 2796 19944 2848
rect 23112 2796 23164 2848
rect 23388 2796 23440 2848
rect 23480 2839 23532 2848
rect 23480 2805 23489 2839
rect 23489 2805 23523 2839
rect 23523 2805 23532 2839
rect 23480 2796 23532 2805
rect 23572 2839 23624 2848
rect 23572 2805 23581 2839
rect 23581 2805 23615 2839
rect 23615 2805 23624 2839
rect 23572 2796 23624 2805
rect 3882 2694 3934 2746
rect 3946 2694 3998 2746
rect 4010 2694 4062 2746
rect 4074 2694 4126 2746
rect 4138 2694 4190 2746
rect 9747 2694 9799 2746
rect 9811 2694 9863 2746
rect 9875 2694 9927 2746
rect 9939 2694 9991 2746
rect 10003 2694 10055 2746
rect 15612 2694 15664 2746
rect 15676 2694 15728 2746
rect 15740 2694 15792 2746
rect 15804 2694 15856 2746
rect 15868 2694 15920 2746
rect 21477 2694 21529 2746
rect 21541 2694 21593 2746
rect 21605 2694 21657 2746
rect 21669 2694 21721 2746
rect 21733 2694 21785 2746
rect 6828 2592 6880 2644
rect 8300 2592 8352 2644
rect 8944 2592 8996 2644
rect 5540 2456 5592 2508
rect 112 2388 164 2440
rect 664 2320 716 2372
rect 1952 2431 2004 2440
rect 1952 2397 1961 2431
rect 1961 2397 1995 2431
rect 1995 2397 2004 2431
rect 1952 2388 2004 2397
rect 9588 2456 9640 2508
rect 10600 2456 10652 2508
rect 14556 2456 14608 2508
rect 14832 2592 14884 2644
rect 17408 2524 17460 2576
rect 18144 2524 18196 2576
rect 19248 2635 19300 2644
rect 19248 2601 19257 2635
rect 19257 2601 19291 2635
rect 19291 2601 19300 2635
rect 19248 2592 19300 2601
rect 23112 2592 23164 2644
rect 23756 2592 23808 2644
rect 20812 2524 20864 2576
rect 22560 2524 22612 2576
rect 1860 2320 1912 2372
rect 8852 2388 8904 2440
rect 9864 2388 9916 2440
rect 10048 2388 10100 2440
rect 11336 2431 11388 2440
rect 11336 2397 11345 2431
rect 11345 2397 11379 2431
rect 11379 2397 11388 2431
rect 11336 2388 11388 2397
rect 11704 2431 11756 2440
rect 11704 2397 11713 2431
rect 11713 2397 11747 2431
rect 11747 2397 11756 2431
rect 11704 2388 11756 2397
rect 12256 2431 12308 2440
rect 12256 2397 12265 2431
rect 12265 2397 12299 2431
rect 12299 2397 12308 2431
rect 12256 2388 12308 2397
rect 12348 2388 12400 2440
rect 13636 2388 13688 2440
rect 15936 2388 15988 2440
rect 16764 2431 16816 2440
rect 16764 2397 16773 2431
rect 16773 2397 16807 2431
rect 16807 2397 16816 2431
rect 16764 2388 16816 2397
rect 17132 2456 17184 2508
rect 8576 2320 8628 2372
rect 17684 2388 17736 2440
rect 18236 2388 18288 2440
rect 19064 2388 19116 2440
rect 19892 2388 19944 2440
rect 19984 2431 20036 2440
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 19616 2363 19668 2372
rect 19616 2329 19625 2363
rect 19625 2329 19659 2363
rect 19659 2329 19668 2363
rect 19616 2320 19668 2329
rect 21824 2320 21876 2372
rect 5724 2252 5776 2304
rect 9220 2252 9272 2304
rect 9404 2252 9456 2304
rect 10232 2252 10284 2304
rect 10876 2295 10928 2304
rect 10876 2261 10885 2295
rect 10885 2261 10919 2295
rect 10919 2261 10928 2295
rect 10876 2252 10928 2261
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 12440 2295 12492 2304
rect 12440 2261 12449 2295
rect 12449 2261 12483 2295
rect 12483 2261 12492 2295
rect 12440 2252 12492 2261
rect 13084 2252 13136 2304
rect 13268 2252 13320 2304
rect 13728 2252 13780 2304
rect 15108 2295 15160 2304
rect 15108 2261 15117 2295
rect 15117 2261 15151 2295
rect 15151 2261 15160 2295
rect 15108 2252 15160 2261
rect 17132 2252 17184 2304
rect 17224 2295 17276 2304
rect 17224 2261 17233 2295
rect 17233 2261 17267 2295
rect 17267 2261 17276 2295
rect 17224 2252 17276 2261
rect 18052 2252 18104 2304
rect 18420 2252 18472 2304
rect 19248 2252 19300 2304
rect 20168 2295 20220 2304
rect 20168 2261 20177 2295
rect 20177 2261 20211 2295
rect 20211 2261 20220 2295
rect 20168 2252 20220 2261
rect 22744 2388 22796 2440
rect 22928 2320 22980 2372
rect 23572 2388 23624 2440
rect 23480 2320 23532 2372
rect 24032 2252 24084 2304
rect 24124 2252 24176 2304
rect 6814 2150 6866 2202
rect 6878 2150 6930 2202
rect 6942 2150 6994 2202
rect 7006 2150 7058 2202
rect 7070 2150 7122 2202
rect 12679 2150 12731 2202
rect 12743 2150 12795 2202
rect 12807 2150 12859 2202
rect 12871 2150 12923 2202
rect 12935 2150 12987 2202
rect 18544 2150 18596 2202
rect 18608 2150 18660 2202
rect 18672 2150 18724 2202
rect 18736 2150 18788 2202
rect 18800 2150 18852 2202
rect 24409 2150 24461 2202
rect 24473 2150 24525 2202
rect 24537 2150 24589 2202
rect 24601 2150 24653 2202
rect 24665 2150 24717 2202
rect 1860 2048 1912 2100
rect 5724 2048 5776 2100
rect 5816 2048 5868 2100
rect 6828 2091 6880 2100
rect 6828 2057 6837 2091
rect 6837 2057 6871 2091
rect 6871 2057 6880 2091
rect 6828 2048 6880 2057
rect 7196 2048 7248 2100
rect 9680 2048 9732 2100
rect 1584 1955 1636 1964
rect 1584 1921 1593 1955
rect 1593 1921 1627 1955
rect 1627 1921 1636 1955
rect 1584 1912 1636 1921
rect 1216 1844 1268 1896
rect 388 1776 440 1828
rect 2412 1955 2464 1964
rect 2412 1921 2421 1955
rect 2421 1921 2455 1955
rect 2455 1921 2464 1955
rect 2412 1912 2464 1921
rect 5172 1955 5224 1964
rect 5172 1921 5181 1955
rect 5181 1921 5215 1955
rect 5215 1921 5224 1955
rect 5172 1912 5224 1921
rect 5448 1955 5500 1964
rect 5448 1921 5457 1955
rect 5457 1921 5491 1955
rect 5491 1921 5500 1955
rect 5448 1912 5500 1921
rect 5724 1955 5776 1964
rect 5724 1921 5733 1955
rect 5733 1921 5767 1955
rect 5767 1921 5776 1955
rect 5724 1912 5776 1921
rect 6644 1955 6696 1964
rect 6644 1921 6653 1955
rect 6653 1921 6687 1955
rect 6687 1921 6696 1955
rect 6644 1912 6696 1921
rect 6828 1912 6880 1964
rect 7288 1912 7340 1964
rect 7656 1955 7708 1964
rect 7656 1921 7665 1955
rect 7665 1921 7699 1955
rect 7699 1921 7708 1955
rect 7656 1912 7708 1921
rect 6092 1776 6144 1828
rect 9404 1980 9456 2032
rect 8116 1955 8168 1964
rect 8116 1921 8125 1955
rect 8125 1921 8159 1955
rect 8159 1921 8168 1955
rect 8116 1912 8168 1921
rect 8484 1955 8536 1964
rect 8484 1921 8493 1955
rect 8493 1921 8527 1955
rect 8527 1921 8536 1955
rect 8484 1912 8536 1921
rect 8760 1955 8812 1964
rect 8760 1921 8769 1955
rect 8769 1921 8803 1955
rect 8803 1921 8812 1955
rect 8760 1912 8812 1921
rect 8944 1912 8996 1964
rect 9312 1955 9364 1964
rect 9312 1921 9321 1955
rect 9321 1921 9355 1955
rect 9355 1921 9364 1955
rect 9312 1912 9364 1921
rect 10232 2023 10284 2032
rect 10232 1989 10257 2023
rect 10257 1989 10284 2023
rect 10232 1980 10284 1989
rect 10876 2048 10928 2100
rect 12440 2048 12492 2100
rect 12532 2048 12584 2100
rect 9864 1955 9916 1964
rect 9864 1921 9873 1955
rect 9873 1921 9907 1955
rect 9907 1921 9916 1955
rect 9864 1912 9916 1921
rect 10508 1912 10560 1964
rect 12072 1912 12124 1964
rect 14556 2048 14608 2100
rect 15108 2048 15160 2100
rect 15384 1980 15436 2032
rect 17224 2048 17276 2100
rect 17408 2048 17460 2100
rect 16672 1980 16724 2032
rect 13452 1955 13504 1964
rect 13452 1921 13461 1955
rect 13461 1921 13495 1955
rect 13495 1921 13504 1955
rect 13452 1912 13504 1921
rect 13636 1912 13688 1964
rect 13728 1955 13780 1964
rect 13728 1921 13737 1955
rect 13737 1921 13771 1955
rect 13771 1921 13780 1955
rect 13728 1912 13780 1921
rect 14004 1955 14056 1964
rect 14004 1921 14013 1955
rect 14013 1921 14047 1955
rect 14047 1921 14056 1955
rect 14004 1912 14056 1921
rect 14280 1955 14332 1964
rect 14280 1921 14289 1955
rect 14289 1921 14323 1955
rect 14323 1921 14332 1955
rect 14280 1912 14332 1921
rect 14372 1912 14424 1964
rect 6000 1708 6052 1760
rect 6644 1708 6696 1760
rect 8208 1708 8260 1760
rect 9404 1776 9456 1828
rect 13360 1844 13412 1896
rect 9680 1776 9732 1828
rect 15568 1912 15620 1964
rect 16304 1955 16356 1964
rect 16304 1921 16313 1955
rect 16313 1921 16347 1955
rect 16347 1921 16356 1955
rect 16304 1912 16356 1921
rect 17960 1980 18012 2032
rect 18420 2048 18472 2100
rect 20168 2048 20220 2100
rect 21548 2048 21600 2100
rect 22008 2048 22060 2100
rect 22560 2048 22612 2100
rect 22652 2091 22704 2100
rect 22652 2057 22661 2091
rect 22661 2057 22695 2091
rect 22695 2057 22704 2091
rect 22652 2048 22704 2057
rect 22192 1980 22244 2032
rect 14924 1844 14976 1896
rect 18052 1844 18104 1896
rect 19616 1844 19668 1896
rect 20720 1844 20772 1896
rect 15200 1776 15252 1828
rect 16672 1776 16724 1828
rect 8576 1708 8628 1760
rect 8852 1708 8904 1760
rect 9036 1751 9088 1760
rect 9036 1717 9045 1751
rect 9045 1717 9079 1751
rect 9079 1717 9088 1751
rect 9036 1708 9088 1717
rect 10324 1751 10376 1760
rect 10324 1717 10333 1751
rect 10333 1717 10367 1751
rect 10367 1717 10376 1751
rect 10324 1708 10376 1717
rect 11060 1751 11112 1760
rect 11060 1717 11069 1751
rect 11069 1717 11103 1751
rect 11103 1717 11112 1751
rect 11060 1708 11112 1717
rect 11704 1751 11756 1760
rect 11704 1717 11713 1751
rect 11713 1717 11747 1751
rect 11747 1717 11756 1751
rect 11704 1708 11756 1717
rect 11796 1708 11848 1760
rect 12624 1751 12676 1760
rect 12624 1717 12633 1751
rect 12633 1717 12667 1751
rect 12667 1717 12676 1751
rect 12624 1708 12676 1717
rect 12900 1751 12952 1760
rect 12900 1717 12909 1751
rect 12909 1717 12943 1751
rect 12943 1717 12952 1751
rect 12900 1708 12952 1717
rect 13544 1708 13596 1760
rect 13636 1751 13688 1760
rect 13636 1717 13645 1751
rect 13645 1717 13679 1751
rect 13679 1717 13688 1751
rect 13636 1708 13688 1717
rect 14924 1708 14976 1760
rect 15292 1708 15344 1760
rect 16396 1708 16448 1760
rect 17500 1776 17552 1828
rect 17592 1708 17644 1760
rect 18052 1708 18104 1760
rect 19156 1776 19208 1828
rect 18972 1708 19024 1760
rect 19892 1751 19944 1760
rect 19892 1717 19901 1751
rect 19901 1717 19935 1751
rect 19935 1717 19944 1751
rect 19892 1708 19944 1717
rect 21180 1819 21232 1828
rect 21180 1785 21189 1819
rect 21189 1785 21223 1819
rect 21223 1785 21232 1819
rect 21180 1776 21232 1785
rect 22284 1955 22336 1964
rect 22284 1921 22293 1955
rect 22293 1921 22327 1955
rect 22327 1921 22336 1955
rect 22284 1912 22336 1921
rect 22652 1912 22704 1964
rect 23204 2091 23256 2100
rect 23204 2057 23213 2091
rect 23213 2057 23247 2091
rect 23247 2057 23256 2091
rect 23204 2048 23256 2057
rect 23940 2048 23992 2100
rect 24216 2048 24268 2100
rect 23020 1980 23072 2032
rect 23112 1955 23164 1964
rect 23112 1921 23121 1955
rect 23121 1921 23155 1955
rect 23155 1921 23164 1955
rect 23112 1912 23164 1921
rect 23388 1955 23440 1964
rect 23388 1921 23397 1955
rect 23397 1921 23431 1955
rect 23431 1921 23440 1955
rect 23388 1912 23440 1921
rect 23756 1912 23808 1964
rect 20812 1708 20864 1760
rect 23204 1776 23256 1828
rect 23572 1776 23624 1828
rect 22744 1708 22796 1760
rect 25228 1708 25280 1760
rect 3882 1606 3934 1658
rect 3946 1606 3998 1658
rect 4010 1606 4062 1658
rect 4074 1606 4126 1658
rect 4138 1606 4190 1658
rect 9747 1606 9799 1658
rect 9811 1606 9863 1658
rect 9875 1606 9927 1658
rect 9939 1606 9991 1658
rect 10003 1606 10055 1658
rect 15612 1606 15664 1658
rect 15676 1606 15728 1658
rect 15740 1606 15792 1658
rect 15804 1606 15856 1658
rect 15868 1606 15920 1658
rect 21477 1606 21529 1658
rect 21541 1606 21593 1658
rect 21605 1606 21657 1658
rect 21669 1606 21721 1658
rect 21733 1606 21785 1658
rect 940 1504 992 1556
rect 2412 1504 2464 1556
rect 4436 1504 4488 1556
rect 5724 1504 5776 1556
rect 6092 1504 6144 1556
rect 4344 1436 4396 1488
rect 5540 1436 5592 1488
rect 2136 1368 2188 1420
rect 2504 1300 2556 1352
rect 2596 1343 2648 1352
rect 2596 1309 2605 1343
rect 2605 1309 2639 1343
rect 2639 1309 2648 1343
rect 2596 1300 2648 1309
rect 2872 1343 2924 1352
rect 2872 1309 2881 1343
rect 2881 1309 2915 1343
rect 2915 1309 2924 1343
rect 2872 1300 2924 1309
rect 3700 1232 3752 1284
rect 3884 1300 3936 1352
rect 4252 1300 4304 1352
rect 4528 1300 4580 1352
rect 4160 1232 4212 1284
rect 4896 1343 4948 1352
rect 4896 1309 4905 1343
rect 4905 1309 4939 1343
rect 4939 1309 4948 1343
rect 4896 1300 4948 1309
rect 4988 1232 5040 1284
rect 5632 1300 5684 1352
rect 5540 1232 5592 1284
rect 6368 1343 6420 1352
rect 6368 1309 6377 1343
rect 6377 1309 6411 1343
rect 6411 1309 6420 1343
rect 6368 1300 6420 1309
rect 6552 1300 6604 1352
rect 6644 1343 6696 1352
rect 6644 1309 6653 1343
rect 6653 1309 6687 1343
rect 6687 1309 6696 1343
rect 6644 1300 6696 1309
rect 6736 1300 6788 1352
rect 7104 1436 7156 1488
rect 8116 1504 8168 1556
rect 9404 1504 9456 1556
rect 8668 1436 8720 1488
rect 9036 1436 9088 1488
rect 13912 1504 13964 1556
rect 14740 1504 14792 1556
rect 6460 1232 6512 1284
rect 1676 1207 1728 1216
rect 1676 1173 1685 1207
rect 1685 1173 1719 1207
rect 1719 1173 1728 1207
rect 1676 1164 1728 1173
rect 1952 1207 2004 1216
rect 1952 1173 1961 1207
rect 1961 1173 1995 1207
rect 1995 1173 2004 1207
rect 1952 1164 2004 1173
rect 2044 1164 2096 1216
rect 2412 1164 2464 1216
rect 2504 1207 2556 1216
rect 2504 1173 2513 1207
rect 2513 1173 2547 1207
rect 2547 1173 2556 1207
rect 2504 1164 2556 1173
rect 2596 1164 2648 1216
rect 3516 1164 3568 1216
rect 3608 1207 3660 1216
rect 3608 1173 3617 1207
rect 3617 1173 3651 1207
rect 3651 1173 3660 1207
rect 3608 1164 3660 1173
rect 4068 1164 4120 1216
rect 4252 1207 4304 1216
rect 4252 1173 4261 1207
rect 4261 1173 4295 1207
rect 4295 1173 4304 1207
rect 4252 1164 4304 1173
rect 4528 1207 4580 1216
rect 4528 1173 4537 1207
rect 4537 1173 4571 1207
rect 4571 1173 4580 1207
rect 4528 1164 4580 1173
rect 4804 1207 4856 1216
rect 4804 1173 4813 1207
rect 4813 1173 4847 1207
rect 4847 1173 4856 1207
rect 4804 1164 4856 1173
rect 5356 1207 5408 1216
rect 5356 1173 5365 1207
rect 5365 1173 5399 1207
rect 5399 1173 5408 1207
rect 5356 1164 5408 1173
rect 5632 1207 5684 1216
rect 5632 1173 5641 1207
rect 5641 1173 5675 1207
rect 5675 1173 5684 1207
rect 5632 1164 5684 1173
rect 6092 1164 6144 1216
rect 6184 1207 6236 1216
rect 6184 1173 6193 1207
rect 6193 1173 6227 1207
rect 6227 1173 6236 1207
rect 6184 1164 6236 1173
rect 6644 1164 6696 1216
rect 7472 1343 7524 1352
rect 7472 1309 7481 1343
rect 7481 1309 7515 1343
rect 7515 1309 7524 1343
rect 7472 1300 7524 1309
rect 14832 1436 14884 1488
rect 14924 1436 14976 1488
rect 15108 1436 15160 1488
rect 16304 1547 16356 1556
rect 16304 1513 16313 1547
rect 16313 1513 16347 1547
rect 16347 1513 16356 1547
rect 16304 1504 16356 1513
rect 16948 1504 17000 1556
rect 19524 1504 19576 1556
rect 16028 1436 16080 1488
rect 18880 1436 18932 1488
rect 21824 1547 21876 1556
rect 21824 1513 21833 1547
rect 21833 1513 21867 1547
rect 21867 1513 21876 1547
rect 21824 1504 21876 1513
rect 22284 1504 22336 1556
rect 22744 1504 22796 1556
rect 7840 1300 7892 1352
rect 8576 1343 8628 1352
rect 8576 1309 8585 1343
rect 8585 1309 8619 1343
rect 8619 1309 8628 1343
rect 8576 1300 8628 1309
rect 8668 1300 8720 1352
rect 9220 1300 9272 1352
rect 9404 1300 9456 1352
rect 9680 1300 9732 1352
rect 11060 1411 11112 1420
rect 11060 1377 11069 1411
rect 11069 1377 11103 1411
rect 11103 1377 11112 1411
rect 11060 1368 11112 1377
rect 11520 1300 11572 1352
rect 11888 1300 11940 1352
rect 12624 1300 12676 1352
rect 13084 1343 13136 1352
rect 13084 1309 13093 1343
rect 13093 1309 13127 1343
rect 13127 1309 13136 1343
rect 13084 1300 13136 1309
rect 7380 1164 7432 1216
rect 7656 1207 7708 1216
rect 7656 1173 7665 1207
rect 7665 1173 7699 1207
rect 7699 1173 7708 1207
rect 7656 1164 7708 1173
rect 7748 1164 7800 1216
rect 8116 1164 8168 1216
rect 9128 1232 9180 1284
rect 8484 1207 8536 1216
rect 8484 1173 8493 1207
rect 8493 1173 8527 1207
rect 8527 1173 8536 1207
rect 8484 1164 8536 1173
rect 9036 1164 9088 1216
rect 11704 1232 11756 1284
rect 13544 1300 13596 1352
rect 13636 1300 13688 1352
rect 15200 1300 15252 1352
rect 15384 1300 15436 1352
rect 16120 1300 16172 1352
rect 17868 1368 17920 1420
rect 16856 1300 16908 1352
rect 16304 1232 16356 1284
rect 17132 1300 17184 1352
rect 18144 1300 18196 1352
rect 10048 1164 10100 1216
rect 10416 1164 10468 1216
rect 11152 1164 11204 1216
rect 11796 1207 11848 1216
rect 11796 1173 11805 1207
rect 11805 1173 11839 1207
rect 11839 1173 11848 1207
rect 11796 1164 11848 1173
rect 12164 1207 12216 1216
rect 12164 1173 12173 1207
rect 12173 1173 12207 1207
rect 12207 1173 12216 1207
rect 12164 1164 12216 1173
rect 12532 1207 12584 1216
rect 12532 1173 12541 1207
rect 12541 1173 12575 1207
rect 12575 1173 12584 1207
rect 12532 1164 12584 1173
rect 13176 1164 13228 1216
rect 13360 1164 13412 1216
rect 13912 1164 13964 1216
rect 15016 1164 15068 1216
rect 18236 1232 18288 1284
rect 19248 1300 19300 1352
rect 19524 1300 19576 1352
rect 19616 1232 19668 1284
rect 22100 1436 22152 1488
rect 23388 1436 23440 1488
rect 23572 1436 23624 1488
rect 24952 1436 25004 1488
rect 21364 1368 21416 1420
rect 21456 1343 21508 1352
rect 21456 1309 21465 1343
rect 21465 1309 21499 1343
rect 21499 1309 21508 1343
rect 21456 1300 21508 1309
rect 21548 1300 21600 1352
rect 20628 1232 20680 1284
rect 21732 1232 21784 1284
rect 22744 1368 22796 1420
rect 23756 1368 23808 1420
rect 22560 1343 22612 1352
rect 22560 1309 22569 1343
rect 22569 1309 22603 1343
rect 22603 1309 22612 1343
rect 22560 1300 22612 1309
rect 22652 1300 22704 1352
rect 23204 1300 23256 1352
rect 23664 1343 23716 1352
rect 23664 1309 23673 1343
rect 23673 1309 23707 1343
rect 23707 1309 23716 1343
rect 23664 1300 23716 1309
rect 23940 1343 23992 1352
rect 23940 1309 23949 1343
rect 23949 1309 23983 1343
rect 23983 1309 23992 1343
rect 23940 1300 23992 1309
rect 24032 1300 24084 1352
rect 24860 1300 24912 1352
rect 22192 1164 22244 1216
rect 22928 1207 22980 1216
rect 22928 1173 22937 1207
rect 22937 1173 22971 1207
rect 22971 1173 22980 1207
rect 22928 1164 22980 1173
rect 23204 1207 23256 1216
rect 23204 1173 23213 1207
rect 23213 1173 23247 1207
rect 23247 1173 23256 1207
rect 23204 1164 23256 1173
rect 23756 1207 23808 1216
rect 23756 1173 23765 1207
rect 23765 1173 23799 1207
rect 23799 1173 23808 1207
rect 23756 1164 23808 1173
rect 6814 1062 6866 1114
rect 6878 1062 6930 1114
rect 6942 1062 6994 1114
rect 7006 1062 7058 1114
rect 7070 1062 7122 1114
rect 12679 1062 12731 1114
rect 12743 1062 12795 1114
rect 12807 1062 12859 1114
rect 12871 1062 12923 1114
rect 12935 1062 12987 1114
rect 18544 1062 18596 1114
rect 18608 1062 18660 1114
rect 18672 1062 18724 1114
rect 18736 1062 18788 1114
rect 18800 1062 18852 1114
rect 24409 1062 24461 1114
rect 24473 1062 24525 1114
rect 24537 1062 24589 1114
rect 24601 1062 24653 1114
rect 24665 1062 24717 1114
rect 2504 960 2556 1012
rect 7380 960 7432 1012
rect 7656 960 7708 1012
rect 9404 892 9456 944
rect 10508 892 10560 944
rect 4528 824 4580 876
rect 8024 824 8076 876
rect 19984 960 20036 1012
rect 21548 960 21600 1012
rect 20536 892 20588 944
rect 22560 960 22612 1012
rect 23756 960 23808 1012
rect 23940 960 23992 1012
rect 3608 756 3660 808
rect 16764 824 16816 876
rect 9036 756 9088 808
rect 16120 756 16172 808
rect 2688 620 2740 672
rect 3148 620 3200 672
rect 6368 620 6420 672
rect 7012 620 7064 672
rect 7472 620 7524 672
rect 8116 620 8168 672
rect 8576 620 8628 672
rect 9588 620 9640 672
rect 12072 620 12124 672
rect 3516 552 3568 604
rect 14096 688 14148 740
rect 21364 756 21416 808
rect 23112 756 23164 808
rect 21640 688 21692 740
rect 16488 620 16540 672
rect 12440 552 12492 604
rect 18236 552 18288 604
rect 6644 484 6696 536
rect 17684 484 17736 536
rect 8208 416 8260 468
rect 18420 620 18472 672
rect 19248 620 19300 672
rect 20904 620 20956 672
rect 22652 620 22704 672
rect 23204 620 23256 672
rect 20444 552 20496 604
rect 21732 552 21784 604
rect 18880 416 18932 468
rect 4252 348 4304 400
rect 8300 348 8352 400
rect 8484 348 8536 400
rect 15936 348 15988 400
rect 2412 280 2464 332
rect 13452 280 13504 332
rect 22744 348 22796 400
rect 23020 348 23072 400
rect 1952 212 2004 264
rect 4068 144 4120 196
rect 9404 144 9456 196
rect 4988 76 5040 128
rect 5540 76 5592 128
rect 18880 212 18932 264
rect 13268 76 13320 128
<< metal2 >>
rect 846 9840 902 10300
rect 952 9846 1440 9874
rect 860 9738 888 9840
rect 952 9738 980 9846
rect 860 9710 980 9738
rect 1412 8566 1440 9846
rect 2042 9840 2098 10300
rect 3238 9840 3294 10300
rect 4434 9840 4490 10300
rect 5630 9840 5686 10300
rect 6826 9840 6882 10300
rect 8022 9840 8078 10300
rect 9218 9840 9274 10300
rect 10414 9840 10470 10300
rect 11610 9840 11666 10300
rect 12806 9840 12862 10300
rect 12912 9846 13124 9874
rect 2056 8634 2084 9840
rect 3252 8634 3280 9840
rect 4448 8634 4476 9840
rect 5644 8634 5672 9840
rect 6840 9194 6868 9840
rect 6748 9166 6868 9194
rect 6748 8634 6776 9166
rect 6814 8732 7122 8741
rect 6814 8730 6820 8732
rect 6876 8730 6900 8732
rect 6956 8730 6980 8732
rect 7036 8730 7060 8732
rect 7116 8730 7122 8732
rect 6876 8678 6878 8730
rect 7058 8678 7060 8730
rect 6814 8676 6820 8678
rect 6876 8676 6900 8678
rect 6956 8676 6980 8678
rect 7036 8676 7060 8678
rect 7116 8676 7122 8678
rect 6814 8667 7122 8676
rect 8036 8634 8064 9840
rect 9232 8634 9260 9840
rect 10428 8634 10456 9840
rect 11624 8634 11652 9840
rect 12820 9738 12848 9840
rect 12912 9738 12940 9846
rect 12820 9710 12940 9738
rect 12679 8732 12987 8741
rect 12679 8730 12685 8732
rect 12741 8730 12765 8732
rect 12821 8730 12845 8732
rect 12901 8730 12925 8732
rect 12981 8730 12987 8732
rect 12741 8678 12743 8730
rect 12923 8678 12925 8730
rect 12679 8676 12685 8678
rect 12741 8676 12765 8678
rect 12821 8676 12845 8678
rect 12901 8676 12925 8678
rect 12981 8676 12987 8678
rect 12679 8667 12987 8676
rect 13096 8634 13124 9846
rect 14002 9840 14058 10300
rect 15198 9840 15254 10300
rect 16394 9840 16450 10300
rect 17590 9840 17646 10300
rect 18786 9840 18842 10300
rect 19982 9840 20038 10300
rect 21178 9840 21234 10300
rect 22374 9840 22430 10300
rect 23570 9840 23626 10300
rect 24766 9840 24822 10300
rect 14016 8634 14044 9840
rect 15212 8634 15240 9840
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 3240 8628 3292 8634
rect 3240 8570 3292 8576
rect 4436 8628 4488 8634
rect 4436 8570 4488 8576
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 11612 8628 11664 8634
rect 11612 8570 11664 8576
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 16408 8566 16436 9840
rect 17604 8634 17632 9840
rect 18800 9058 18828 9840
rect 18800 9030 18920 9058
rect 18544 8732 18852 8741
rect 18544 8730 18550 8732
rect 18606 8730 18630 8732
rect 18686 8730 18710 8732
rect 18766 8730 18790 8732
rect 18846 8730 18852 8732
rect 18606 8678 18608 8730
rect 18788 8678 18790 8730
rect 18544 8676 18550 8678
rect 18606 8676 18630 8678
rect 18686 8676 18710 8678
rect 18766 8676 18790 8678
rect 18846 8676 18852 8678
rect 18544 8667 18852 8676
rect 18892 8634 18920 9030
rect 19996 8634 20024 9840
rect 21192 8634 21220 9840
rect 22388 8634 22416 9840
rect 23584 8634 23612 9840
rect 24409 8732 24717 8741
rect 24409 8730 24415 8732
rect 24471 8730 24495 8732
rect 24551 8730 24575 8732
rect 24631 8730 24655 8732
rect 24711 8730 24717 8732
rect 24471 8678 24473 8730
rect 24653 8678 24655 8730
rect 24409 8676 24415 8678
rect 24471 8676 24495 8678
rect 24551 8676 24575 8678
rect 24631 8676 24655 8678
rect 24711 8676 24717 8678
rect 24409 8667 24717 8676
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 18880 8628 18932 8634
rect 18880 8570 18932 8576
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 1400 8560 1452 8566
rect 1400 8502 1452 8508
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 14096 8492 14148 8498
rect 14096 8434 14148 8440
rect 15384 8492 15436 8498
rect 15384 8434 15436 8440
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 19248 8492 19300 8498
rect 19248 8434 19300 8440
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 112 2440 164 2446
rect 1780 2417 1808 8434
rect 2424 4049 2452 8434
rect 2410 4040 2466 4049
rect 2410 3975 2466 3984
rect 1952 2440 2004 2446
rect 112 2382 164 2388
rect 1766 2408 1822 2417
rect 124 160 152 2382
rect 664 2372 716 2378
rect 1952 2382 2004 2388
rect 1766 2343 1822 2352
rect 1860 2372 1912 2378
rect 664 2314 716 2320
rect 1860 2314 1912 2320
rect 388 1828 440 1834
rect 388 1770 440 1776
rect 400 160 428 1770
rect 676 160 704 2314
rect 1872 2106 1900 2314
rect 1860 2100 1912 2106
rect 1860 2042 1912 2048
rect 1584 1964 1636 1970
rect 1504 1924 1584 1952
rect 1216 1896 1268 1902
rect 1216 1838 1268 1844
rect 940 1556 992 1562
rect 940 1498 992 1504
rect 952 160 980 1498
rect 1228 160 1256 1838
rect 1504 160 1532 1924
rect 1584 1906 1636 1912
rect 1964 1306 1992 2382
rect 2412 1964 2464 1970
rect 2412 1906 2464 1912
rect 2424 1562 2452 1906
rect 3620 1873 3648 8434
rect 3882 8188 4190 8197
rect 3882 8186 3888 8188
rect 3944 8186 3968 8188
rect 4024 8186 4048 8188
rect 4104 8186 4128 8188
rect 4184 8186 4190 8188
rect 3944 8134 3946 8186
rect 4126 8134 4128 8186
rect 3882 8132 3888 8134
rect 3944 8132 3968 8134
rect 4024 8132 4048 8134
rect 4104 8132 4128 8134
rect 4184 8132 4190 8134
rect 3882 8123 4190 8132
rect 3882 7100 4190 7109
rect 3882 7098 3888 7100
rect 3944 7098 3968 7100
rect 4024 7098 4048 7100
rect 4104 7098 4128 7100
rect 4184 7098 4190 7100
rect 3944 7046 3946 7098
rect 4126 7046 4128 7098
rect 3882 7044 3888 7046
rect 3944 7044 3968 7046
rect 4024 7044 4048 7046
rect 4104 7044 4128 7046
rect 4184 7044 4190 7046
rect 3882 7035 4190 7044
rect 3882 6012 4190 6021
rect 3882 6010 3888 6012
rect 3944 6010 3968 6012
rect 4024 6010 4048 6012
rect 4104 6010 4128 6012
rect 4184 6010 4190 6012
rect 3944 5958 3946 6010
rect 4126 5958 4128 6010
rect 3882 5956 3888 5958
rect 3944 5956 3968 5958
rect 4024 5956 4048 5958
rect 4104 5956 4128 5958
rect 4184 5956 4190 5958
rect 3882 5947 4190 5956
rect 3882 4924 4190 4933
rect 3882 4922 3888 4924
rect 3944 4922 3968 4924
rect 4024 4922 4048 4924
rect 4104 4922 4128 4924
rect 4184 4922 4190 4924
rect 3944 4870 3946 4922
rect 4126 4870 4128 4922
rect 3882 4868 3888 4870
rect 3944 4868 3968 4870
rect 4024 4868 4048 4870
rect 4104 4868 4128 4870
rect 4184 4868 4190 4870
rect 3882 4859 4190 4868
rect 3882 3836 4190 3845
rect 3882 3834 3888 3836
rect 3944 3834 3968 3836
rect 4024 3834 4048 3836
rect 4104 3834 4128 3836
rect 4184 3834 4190 3836
rect 3944 3782 3946 3834
rect 4126 3782 4128 3834
rect 3882 3780 3888 3782
rect 3944 3780 3968 3782
rect 4024 3780 4048 3782
rect 4104 3780 4128 3782
rect 4184 3780 4190 3782
rect 3882 3771 4190 3780
rect 4434 3088 4490 3097
rect 4434 3023 4490 3032
rect 3882 2748 4190 2757
rect 3882 2746 3888 2748
rect 3944 2746 3968 2748
rect 4024 2746 4048 2748
rect 4104 2746 4128 2748
rect 4184 2746 4190 2748
rect 3944 2694 3946 2746
rect 4126 2694 4128 2746
rect 3882 2692 3888 2694
rect 3944 2692 3968 2694
rect 4024 2692 4048 2694
rect 4104 2692 4128 2694
rect 4184 2692 4190 2694
rect 3882 2683 4190 2692
rect 3606 1864 3662 1873
rect 3606 1799 3662 1808
rect 3882 1660 4190 1669
rect 3882 1658 3888 1660
rect 3944 1658 3968 1660
rect 4024 1658 4048 1660
rect 4104 1658 4128 1660
rect 4184 1658 4190 1660
rect 3944 1606 3946 1658
rect 4126 1606 4128 1658
rect 3882 1604 3888 1606
rect 3944 1604 3968 1606
rect 4024 1604 4048 1606
rect 4104 1604 4128 1606
rect 4184 1604 4190 1606
rect 3882 1595 4190 1604
rect 4342 1592 4398 1601
rect 2412 1556 2464 1562
rect 4448 1562 4476 3023
rect 4816 2009 4844 8434
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 4802 2000 4858 2009
rect 4802 1935 4858 1944
rect 5172 1964 5224 1970
rect 5172 1906 5224 1912
rect 5448 1964 5500 1970
rect 5448 1906 5500 1912
rect 4342 1527 4398 1536
rect 4436 1556 4488 1562
rect 2412 1498 2464 1504
rect 4356 1494 4384 1527
rect 4436 1498 4488 1504
rect 4344 1488 4396 1494
rect 2136 1420 2188 1426
rect 2136 1362 2188 1368
rect 2516 1414 2820 1442
rect 4344 1430 4396 1436
rect 4894 1456 4950 1465
rect 1780 1278 1992 1306
rect 1676 1216 1728 1222
rect 1676 1158 1728 1164
rect 1688 377 1716 1158
rect 1674 368 1730 377
rect 1674 303 1730 312
rect 1780 160 1808 1278
rect 1952 1216 2004 1222
rect 1952 1158 2004 1164
rect 2044 1216 2096 1222
rect 2044 1158 2096 1164
rect 1964 270 1992 1158
rect 1952 264 2004 270
rect 1952 206 2004 212
rect 2056 160 2084 1158
rect 2148 762 2176 1362
rect 2516 1358 2544 1414
rect 2504 1352 2556 1358
rect 2504 1294 2556 1300
rect 2596 1352 2648 1358
rect 2648 1300 2728 1306
rect 2596 1294 2728 1300
rect 2608 1278 2728 1294
rect 2412 1216 2464 1222
rect 2412 1158 2464 1164
rect 2504 1216 2556 1222
rect 2504 1158 2556 1164
rect 2596 1216 2648 1222
rect 2596 1158 2648 1164
rect 2148 734 2360 762
rect 2332 160 2360 734
rect 2424 338 2452 1158
rect 2516 1018 2544 1158
rect 2504 1012 2556 1018
rect 2504 954 2556 960
rect 2412 332 2464 338
rect 2412 274 2464 280
rect 2608 160 2636 1158
rect 2700 678 2728 1278
rect 2792 762 2820 1414
rect 4894 1391 4950 1400
rect 4908 1358 4936 1391
rect 2872 1352 2924 1358
rect 3884 1352 3936 1358
rect 2924 1312 3464 1340
rect 2872 1294 2924 1300
rect 2792 734 2912 762
rect 2688 672 2740 678
rect 2688 614 2740 620
rect 2884 160 2912 734
rect 3148 672 3200 678
rect 3148 614 3200 620
rect 3160 160 3188 614
rect 3436 160 3464 1312
rect 3884 1294 3936 1300
rect 4252 1352 4304 1358
rect 4528 1352 4580 1358
rect 4304 1312 4384 1340
rect 4252 1294 4304 1300
rect 3700 1284 3752 1290
rect 3700 1226 3752 1232
rect 3516 1216 3568 1222
rect 3516 1158 3568 1164
rect 3608 1216 3660 1222
rect 3608 1158 3660 1164
rect 3528 610 3556 1158
rect 3620 814 3648 1158
rect 3608 808 3660 814
rect 3608 750 3660 756
rect 3516 604 3568 610
rect 3516 546 3568 552
rect 3712 160 3740 1226
rect 110 -300 166 160
rect 386 -300 442 160
rect 662 -300 718 160
rect 938 -300 994 160
rect 1214 -300 1270 160
rect 1490 -300 1546 160
rect 1766 -300 1822 160
rect 2042 -300 2098 160
rect 2318 -300 2374 160
rect 2594 -300 2650 160
rect 2870 -300 2926 160
rect 3146 -300 3202 160
rect 3422 -300 3478 160
rect 3698 -300 3754 160
rect 3896 82 3924 1294
rect 4160 1284 4212 1290
rect 4160 1226 4212 1232
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 4080 202 4108 1158
rect 4068 196 4120 202
rect 3974 82 4030 160
rect 4068 138 4120 144
rect 3896 54 4030 82
rect 4172 82 4200 1226
rect 4252 1216 4304 1222
rect 4252 1158 4304 1164
rect 4264 406 4292 1158
rect 4252 400 4304 406
rect 4252 342 4304 348
rect 4250 82 4306 160
rect 4172 54 4306 82
rect 4356 82 4384 1312
rect 4896 1352 4948 1358
rect 4580 1312 4660 1340
rect 4528 1294 4580 1300
rect 4528 1216 4580 1222
rect 4528 1158 4580 1164
rect 4540 882 4568 1158
rect 4528 876 4580 882
rect 4528 818 4580 824
rect 4526 82 4582 160
rect 4356 54 4582 82
rect 4632 82 4660 1312
rect 4896 1294 4948 1300
rect 4988 1284 5040 1290
rect 4988 1226 5040 1232
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4816 649 4844 1158
rect 4802 640 4858 649
rect 4802 575 4858 584
rect 4802 82 4858 160
rect 5000 134 5028 1226
rect 4632 54 4858 82
rect 4988 128 5040 134
rect 4988 70 5040 76
rect 5078 82 5134 160
rect 5184 82 5212 1906
rect 5356 1216 5408 1222
rect 5356 1158 5408 1164
rect 5368 921 5396 1158
rect 5354 912 5410 921
rect 5354 847 5410 856
rect 3974 -300 4030 54
rect 4250 -300 4306 54
rect 4526 -300 4582 54
rect 4802 -300 4858 54
rect 5078 54 5212 82
rect 5354 82 5410 160
rect 5460 82 5488 1906
rect 5552 1494 5580 2450
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 5736 2106 5764 2246
rect 5828 2106 5856 8434
rect 7024 7834 7052 8434
rect 7024 7806 7236 7834
rect 6814 7644 7122 7653
rect 6814 7642 6820 7644
rect 6876 7642 6900 7644
rect 6956 7642 6980 7644
rect 7036 7642 7060 7644
rect 7116 7642 7122 7644
rect 6876 7590 6878 7642
rect 7058 7590 7060 7642
rect 6814 7588 6820 7590
rect 6876 7588 6900 7590
rect 6956 7588 6980 7590
rect 7036 7588 7060 7590
rect 7116 7588 7122 7590
rect 6814 7579 7122 7588
rect 6814 6556 7122 6565
rect 6814 6554 6820 6556
rect 6876 6554 6900 6556
rect 6956 6554 6980 6556
rect 7036 6554 7060 6556
rect 7116 6554 7122 6556
rect 6876 6502 6878 6554
rect 7058 6502 7060 6554
rect 6814 6500 6820 6502
rect 6876 6500 6900 6502
rect 6956 6500 6980 6502
rect 7036 6500 7060 6502
rect 7116 6500 7122 6502
rect 6814 6491 7122 6500
rect 6814 5468 7122 5477
rect 6814 5466 6820 5468
rect 6876 5466 6900 5468
rect 6956 5466 6980 5468
rect 7036 5466 7060 5468
rect 7116 5466 7122 5468
rect 6876 5414 6878 5466
rect 7058 5414 7060 5466
rect 6814 5412 6820 5414
rect 6876 5412 6900 5414
rect 6956 5412 6980 5414
rect 7036 5412 7060 5414
rect 7116 5412 7122 5414
rect 6814 5403 7122 5412
rect 6814 4380 7122 4389
rect 6814 4378 6820 4380
rect 6876 4378 6900 4380
rect 6956 4378 6980 4380
rect 7036 4378 7060 4380
rect 7116 4378 7122 4380
rect 6876 4326 6878 4378
rect 7058 4326 7060 4378
rect 6814 4324 6820 4326
rect 6876 4324 6900 4326
rect 6956 4324 6980 4326
rect 7036 4324 7060 4326
rect 7116 4324 7122 4326
rect 6814 4315 7122 4324
rect 6814 3292 7122 3301
rect 6814 3290 6820 3292
rect 6876 3290 6900 3292
rect 6956 3290 6980 3292
rect 7036 3290 7060 3292
rect 7116 3290 7122 3292
rect 6876 3238 6878 3290
rect 7058 3238 7060 3290
rect 6814 3236 6820 3238
rect 6876 3236 6900 3238
rect 6956 3236 6980 3238
rect 7036 3236 7060 3238
rect 7116 3236 7122 3238
rect 6814 3227 7122 3236
rect 6644 3120 6696 3126
rect 6644 3062 6696 3068
rect 5724 2100 5776 2106
rect 5724 2042 5776 2048
rect 5816 2100 5868 2106
rect 5816 2042 5868 2048
rect 6656 1970 6684 3062
rect 6826 2952 6882 2961
rect 6748 2910 6826 2938
rect 5724 1964 5776 1970
rect 5724 1906 5776 1912
rect 6644 1964 6696 1970
rect 6644 1906 6696 1912
rect 5736 1562 5764 1906
rect 6092 1828 6144 1834
rect 6092 1770 6144 1776
rect 6000 1760 6052 1766
rect 5998 1728 6000 1737
rect 6052 1728 6054 1737
rect 5998 1663 6054 1672
rect 6104 1562 6132 1770
rect 6644 1760 6696 1766
rect 6644 1702 6696 1708
rect 5724 1556 5776 1562
rect 5724 1498 5776 1504
rect 6092 1556 6144 1562
rect 6092 1498 6144 1504
rect 5540 1488 5592 1494
rect 5540 1430 5592 1436
rect 6656 1358 6684 1702
rect 6748 1358 6776 2910
rect 6826 2887 6882 2896
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6840 2553 6868 2586
rect 6826 2544 6882 2553
rect 6826 2479 6882 2488
rect 6814 2204 7122 2213
rect 6814 2202 6820 2204
rect 6876 2202 6900 2204
rect 6956 2202 6980 2204
rect 7036 2202 7060 2204
rect 7116 2202 7122 2204
rect 6876 2150 6878 2202
rect 7058 2150 7060 2202
rect 6814 2148 6820 2150
rect 6876 2148 6900 2150
rect 6956 2148 6980 2150
rect 7036 2148 7060 2150
rect 7116 2148 7122 2150
rect 6814 2139 7122 2148
rect 7208 2106 7236 7806
rect 8220 3194 8248 8434
rect 9324 3942 9352 8434
rect 9747 8188 10055 8197
rect 9747 8186 9753 8188
rect 9809 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10055 8188
rect 9809 8134 9811 8186
rect 9991 8134 9993 8186
rect 9747 8132 9753 8134
rect 9809 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10055 8134
rect 9747 8123 10055 8132
rect 9747 7100 10055 7109
rect 9747 7098 9753 7100
rect 9809 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10055 7100
rect 9809 7046 9811 7098
rect 9991 7046 9993 7098
rect 9747 7044 9753 7046
rect 9809 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10055 7046
rect 9747 7035 10055 7044
rect 9747 6012 10055 6021
rect 9747 6010 9753 6012
rect 9809 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10055 6012
rect 9809 5958 9811 6010
rect 9991 5958 9993 6010
rect 9747 5956 9753 5958
rect 9809 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10055 5958
rect 9747 5947 10055 5956
rect 9747 4924 10055 4933
rect 9747 4922 9753 4924
rect 9809 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10055 4924
rect 9809 4870 9811 4922
rect 9991 4870 9993 4922
rect 9747 4868 9753 4870
rect 9809 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10055 4870
rect 9747 4859 10055 4868
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9312 3936 9364 3942
rect 9312 3878 9364 3884
rect 9508 3738 9536 4082
rect 10520 3942 10548 8434
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 9747 3836 10055 3845
rect 9747 3834 9753 3836
rect 9809 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10055 3836
rect 9809 3782 9811 3834
rect 9991 3782 9993 3834
rect 9747 3780 9753 3782
rect 9809 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10055 3782
rect 9747 3771 10055 3780
rect 10704 3738 10732 4082
rect 11716 3942 11744 8434
rect 12679 7644 12987 7653
rect 12679 7642 12685 7644
rect 12741 7642 12765 7644
rect 12821 7642 12845 7644
rect 12901 7642 12925 7644
rect 12981 7642 12987 7644
rect 12741 7590 12743 7642
rect 12923 7590 12925 7642
rect 12679 7588 12685 7590
rect 12741 7588 12765 7590
rect 12821 7588 12845 7590
rect 12901 7588 12925 7590
rect 12981 7588 12987 7590
rect 12679 7579 12987 7588
rect 12679 6556 12987 6565
rect 12679 6554 12685 6556
rect 12741 6554 12765 6556
rect 12821 6554 12845 6556
rect 12901 6554 12925 6556
rect 12981 6554 12987 6556
rect 12741 6502 12743 6554
rect 12923 6502 12925 6554
rect 12679 6500 12685 6502
rect 12741 6500 12765 6502
rect 12821 6500 12845 6502
rect 12901 6500 12925 6502
rect 12981 6500 12987 6502
rect 12679 6491 12987 6500
rect 12679 5468 12987 5477
rect 12679 5466 12685 5468
rect 12741 5466 12765 5468
rect 12821 5466 12845 5468
rect 12901 5466 12925 5468
rect 12981 5466 12987 5468
rect 12741 5414 12743 5466
rect 12923 5414 12925 5466
rect 12679 5412 12685 5414
rect 12741 5412 12765 5414
rect 12821 5412 12845 5414
rect 12901 5412 12925 5414
rect 12981 5412 12987 5414
rect 12679 5403 12987 5412
rect 12679 4380 12987 4389
rect 12679 4378 12685 4380
rect 12741 4378 12765 4380
rect 12821 4378 12845 4380
rect 12901 4378 12925 4380
rect 12981 4378 12987 4380
rect 12741 4326 12743 4378
rect 12923 4326 12925 4378
rect 12679 4324 12685 4326
rect 12741 4324 12765 4326
rect 12821 4324 12845 4326
rect 12901 4324 12925 4326
rect 12981 4324 12987 4326
rect 12679 4315 12987 4324
rect 11888 4140 11940 4146
rect 11888 4082 11940 4088
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10796 3534 10824 3878
rect 11900 3738 11928 4082
rect 13096 3738 13124 4082
rect 13188 3942 13216 8434
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 14108 3738 14136 8434
rect 15396 3738 15424 8434
rect 15612 8188 15920 8197
rect 15612 8186 15618 8188
rect 15674 8186 15698 8188
rect 15754 8186 15778 8188
rect 15834 8186 15858 8188
rect 15914 8186 15920 8188
rect 15674 8134 15676 8186
rect 15856 8134 15858 8186
rect 15612 8132 15618 8134
rect 15674 8132 15698 8134
rect 15754 8132 15778 8134
rect 15834 8132 15858 8134
rect 15914 8132 15920 8134
rect 15612 8123 15920 8132
rect 17420 8090 17448 8434
rect 17408 8084 17460 8090
rect 17408 8026 17460 8032
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 15612 7100 15920 7109
rect 15612 7098 15618 7100
rect 15674 7098 15698 7100
rect 15754 7098 15778 7100
rect 15834 7098 15858 7100
rect 15914 7098 15920 7100
rect 15674 7046 15676 7098
rect 15856 7046 15858 7098
rect 15612 7044 15618 7046
rect 15674 7044 15698 7046
rect 15754 7044 15778 7046
rect 15834 7044 15858 7046
rect 15914 7044 15920 7046
rect 15612 7035 15920 7044
rect 15612 6012 15920 6021
rect 15612 6010 15618 6012
rect 15674 6010 15698 6012
rect 15754 6010 15778 6012
rect 15834 6010 15858 6012
rect 15914 6010 15920 6012
rect 15674 5958 15676 6010
rect 15856 5958 15858 6010
rect 15612 5956 15618 5958
rect 15674 5956 15698 5958
rect 15754 5956 15778 5958
rect 15834 5956 15858 5958
rect 15914 5956 15920 5958
rect 15612 5947 15920 5956
rect 15612 4924 15920 4933
rect 15612 4922 15618 4924
rect 15674 4922 15698 4924
rect 15754 4922 15778 4924
rect 15834 4922 15858 4924
rect 15914 4922 15920 4924
rect 15674 4870 15676 4922
rect 15856 4870 15858 4922
rect 15612 4868 15618 4870
rect 15674 4868 15698 4870
rect 15754 4868 15778 4870
rect 15834 4868 15858 4870
rect 15914 4868 15920 4870
rect 15612 4859 15920 4868
rect 15612 3836 15920 3845
rect 15612 3834 15618 3836
rect 15674 3834 15698 3836
rect 15754 3834 15778 3836
rect 15834 3834 15858 3836
rect 15914 3834 15920 3836
rect 15674 3782 15676 3834
rect 15856 3782 15858 3834
rect 15612 3780 15618 3782
rect 15674 3780 15698 3782
rect 15754 3780 15778 3782
rect 15834 3780 15858 3782
rect 15914 3780 15920 3782
rect 15612 3771 15920 3780
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 14096 3732 14148 3738
rect 14096 3674 14148 3680
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 7840 2916 7892 2922
rect 7840 2858 7892 2864
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 6840 1970 6868 2042
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 7288 1964 7340 1970
rect 7656 1964 7708 1970
rect 7288 1906 7340 1912
rect 7576 1924 7656 1952
rect 7102 1728 7158 1737
rect 7102 1663 7158 1672
rect 7116 1494 7144 1663
rect 7104 1488 7156 1494
rect 7104 1430 7156 1436
rect 5632 1352 5684 1358
rect 6368 1352 6420 1358
rect 5684 1312 6040 1340
rect 5632 1294 5684 1300
rect 5540 1284 5592 1290
rect 5540 1226 5592 1232
rect 5552 218 5580 1226
rect 5632 1216 5684 1222
rect 5632 1158 5684 1164
rect 5644 513 5672 1158
rect 5630 504 5686 513
rect 5630 439 5686 448
rect 5552 190 5764 218
rect 5354 54 5488 82
rect 5540 128 5592 134
rect 5630 82 5686 160
rect 5592 76 5686 82
rect 5540 70 5686 76
rect 5552 54 5686 70
rect 5736 82 5764 190
rect 5906 82 5962 160
rect 5736 54 5962 82
rect 6012 82 6040 1312
rect 6368 1294 6420 1300
rect 6552 1352 6604 1358
rect 6552 1294 6604 1300
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 6092 1216 6144 1222
rect 6092 1158 6144 1164
rect 6184 1216 6236 1222
rect 6184 1158 6236 1164
rect 6104 241 6132 1158
rect 6196 785 6224 1158
rect 6182 776 6238 785
rect 6182 711 6238 720
rect 6380 678 6408 1294
rect 6460 1284 6512 1290
rect 6460 1226 6512 1232
rect 6368 672 6420 678
rect 6368 614 6420 620
rect 6090 232 6146 241
rect 6090 167 6146 176
rect 6472 160 6500 1226
rect 6182 82 6238 160
rect 6012 54 6238 82
rect 5078 -300 5134 54
rect 5354 -300 5410 54
rect 5630 -300 5686 54
rect 5906 -300 5962 54
rect 6182 -300 6238 54
rect 6458 -300 6514 160
rect 6564 82 6592 1294
rect 6644 1216 6696 1222
rect 6644 1158 6696 1164
rect 6656 542 6684 1158
rect 6814 1116 7122 1125
rect 6814 1114 6820 1116
rect 6876 1114 6900 1116
rect 6956 1114 6980 1116
rect 7036 1114 7060 1116
rect 7116 1114 7122 1116
rect 6876 1062 6878 1114
rect 7058 1062 7060 1114
rect 6814 1060 6820 1062
rect 6876 1060 6900 1062
rect 6956 1060 6980 1062
rect 7036 1060 7060 1062
rect 7116 1060 7122 1062
rect 6814 1051 7122 1060
rect 7012 672 7064 678
rect 7012 614 7064 620
rect 6644 536 6696 542
rect 6644 478 6696 484
rect 7024 160 7052 614
rect 7300 160 7328 1906
rect 7472 1352 7524 1358
rect 7472 1294 7524 1300
rect 7380 1216 7432 1222
rect 7380 1158 7432 1164
rect 7392 1018 7420 1158
rect 7380 1012 7432 1018
rect 7380 954 7432 960
rect 7484 678 7512 1294
rect 7472 672 7524 678
rect 7472 614 7524 620
rect 7576 160 7604 1924
rect 7656 1906 7708 1912
rect 7852 1358 7880 2858
rect 8312 2650 8340 2994
rect 9128 2984 9180 2990
rect 9128 2926 9180 2932
rect 8852 2848 8904 2854
rect 8852 2790 8904 2796
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8864 2446 8892 2790
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 8852 2440 8904 2446
rect 8852 2382 8904 2388
rect 8576 2372 8628 2378
rect 8576 2314 8628 2320
rect 8206 2272 8262 2281
rect 8036 2230 8206 2258
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 7656 1216 7708 1222
rect 7656 1158 7708 1164
rect 7748 1216 7800 1222
rect 7748 1158 7800 1164
rect 7668 1018 7696 1158
rect 7656 1012 7708 1018
rect 7656 954 7708 960
rect 6734 82 6790 160
rect 6564 54 6790 82
rect 6734 -300 6790 54
rect 7010 -300 7066 160
rect 7286 -300 7342 160
rect 7562 -300 7618 160
rect 7760 82 7788 1158
rect 8036 882 8064 2230
rect 8206 2207 8262 2216
rect 8116 1964 8168 1970
rect 8484 1964 8536 1970
rect 8116 1906 8168 1912
rect 8404 1924 8484 1952
rect 8128 1562 8156 1906
rect 8208 1760 8260 1766
rect 8208 1702 8260 1708
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 8116 1216 8168 1222
rect 8114 1184 8116 1193
rect 8168 1184 8170 1193
rect 8114 1119 8170 1128
rect 8024 876 8076 882
rect 8024 818 8076 824
rect 8116 672 8168 678
rect 8116 614 8168 620
rect 8128 160 8156 614
rect 8220 474 8248 1702
rect 8298 1320 8354 1329
rect 8298 1255 8354 1264
rect 8208 468 8260 474
rect 8208 410 8260 416
rect 8312 406 8340 1255
rect 8300 400 8352 406
rect 8300 342 8352 348
rect 8404 160 8432 1924
rect 8484 1906 8536 1912
rect 8588 1766 8616 2314
rect 8956 2122 8984 2586
rect 8864 2094 8984 2122
rect 8760 1964 8812 1970
rect 8760 1906 8812 1912
rect 8576 1760 8628 1766
rect 8576 1702 8628 1708
rect 8668 1488 8720 1494
rect 8668 1430 8720 1436
rect 8680 1358 8708 1430
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 8484 1216 8536 1222
rect 8484 1158 8536 1164
rect 8496 406 8524 1158
rect 8588 678 8616 1294
rect 8576 672 8628 678
rect 8576 614 8628 620
rect 8484 400 8536 406
rect 8484 342 8536 348
rect 7838 82 7894 160
rect 7760 54 7894 82
rect 7838 -300 7894 54
rect 8114 -300 8170 160
rect 8390 -300 8446 160
rect 8666 82 8722 160
rect 8772 82 8800 1906
rect 8864 1766 8892 2094
rect 8944 1964 8996 1970
rect 8944 1906 8996 1912
rect 8852 1760 8904 1766
rect 8852 1702 8904 1708
rect 8956 160 8984 1906
rect 9036 1760 9088 1766
rect 9036 1702 9088 1708
rect 9048 1494 9076 1702
rect 9140 1601 9168 2926
rect 9600 2514 9628 2994
rect 9747 2748 10055 2757
rect 9747 2746 9753 2748
rect 9809 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10055 2748
rect 9809 2694 9811 2746
rect 9991 2694 9993 2746
rect 9747 2692 9753 2694
rect 9809 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10055 2694
rect 9747 2683 10055 2692
rect 10612 2514 10640 3470
rect 11992 2553 12020 3470
rect 12679 3292 12987 3301
rect 12679 3290 12685 3292
rect 12741 3290 12765 3292
rect 12821 3290 12845 3292
rect 12901 3290 12925 3292
rect 12981 3290 12987 3292
rect 12741 3238 12743 3290
rect 12923 3238 12925 3290
rect 12679 3236 12685 3238
rect 12741 3236 12765 3238
rect 12821 3236 12845 3238
rect 12901 3236 12925 3238
rect 12981 3236 12987 3238
rect 12679 3227 12987 3236
rect 15488 3194 15516 3470
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 16488 3120 16540 3126
rect 12346 3088 12402 3097
rect 16488 3062 16540 3068
rect 12346 3023 12402 3032
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 11978 2544 12034 2553
rect 9588 2508 9640 2514
rect 9588 2450 9640 2456
rect 10600 2508 10652 2514
rect 11978 2479 12034 2488
rect 10600 2450 10652 2456
rect 12268 2446 12296 2926
rect 12360 2446 12388 3023
rect 14372 2984 14424 2990
rect 14372 2926 14424 2932
rect 14096 2848 14148 2854
rect 14096 2790 14148 2796
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 11336 2440 11388 2446
rect 11336 2382 11388 2388
rect 11704 2440 11756 2446
rect 11704 2382 11756 2388
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9404 2304 9456 2310
rect 9404 2246 9456 2252
rect 9126 1592 9182 1601
rect 9126 1527 9182 1536
rect 9036 1488 9088 1494
rect 9036 1430 9088 1436
rect 9232 1358 9260 2246
rect 9416 2038 9444 2246
rect 9586 2136 9642 2145
rect 9586 2071 9642 2080
rect 9680 2100 9732 2106
rect 9404 2032 9456 2038
rect 9404 1974 9456 1980
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 9220 1352 9272 1358
rect 9220 1294 9272 1300
rect 9128 1284 9180 1290
rect 9128 1226 9180 1232
rect 9036 1216 9088 1222
rect 9036 1158 9088 1164
rect 9048 814 9076 1158
rect 9036 808 9088 814
rect 9036 750 9088 756
rect 9140 660 9168 1226
rect 9140 632 9260 660
rect 9232 160 9260 632
rect 8666 54 8800 82
rect 8666 -300 8722 54
rect 8942 -300 8998 160
rect 9218 -300 9274 160
rect 9324 82 9352 1906
rect 9404 1828 9456 1834
rect 9404 1770 9456 1776
rect 9416 1562 9444 1770
rect 9404 1556 9456 1562
rect 9404 1498 9456 1504
rect 9404 1352 9456 1358
rect 9404 1294 9456 1300
rect 9416 950 9444 1294
rect 9404 944 9456 950
rect 9404 886 9456 892
rect 9600 762 9628 2071
rect 9680 2042 9732 2048
rect 9692 1834 9720 2042
rect 9876 1970 9904 2382
rect 10060 2281 10088 2382
rect 10232 2304 10284 2310
rect 10046 2272 10102 2281
rect 10232 2246 10284 2252
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10046 2207 10102 2216
rect 10244 2038 10272 2246
rect 10888 2106 10916 2246
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10232 2032 10284 2038
rect 10232 1974 10284 1980
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 10508 1964 10560 1970
rect 10508 1906 10560 1912
rect 9680 1828 9732 1834
rect 9680 1770 9732 1776
rect 10324 1760 10376 1766
rect 10152 1720 10324 1748
rect 9747 1660 10055 1669
rect 9747 1658 9753 1660
rect 9809 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10055 1660
rect 9809 1606 9811 1658
rect 9991 1606 9993 1658
rect 9747 1604 9753 1606
rect 9809 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10055 1606
rect 9747 1595 10055 1604
rect 9680 1352 9732 1358
rect 10152 1306 10180 1720
rect 10324 1702 10376 1708
rect 9680 1294 9732 1300
rect 9692 1193 9720 1294
rect 9968 1278 10180 1306
rect 9678 1184 9734 1193
rect 9678 1119 9734 1128
rect 9416 734 9628 762
rect 9416 202 9444 734
rect 9588 672 9640 678
rect 9588 614 9640 620
rect 9404 196 9456 202
rect 9404 138 9456 144
rect 9494 82 9550 160
rect 9324 54 9550 82
rect 9600 82 9628 614
rect 9770 82 9826 160
rect 9600 54 9826 82
rect 9968 82 9996 1278
rect 10048 1216 10100 1222
rect 10416 1216 10468 1222
rect 10100 1176 10364 1204
rect 10048 1158 10100 1164
rect 10336 160 10364 1176
rect 10416 1158 10468 1164
rect 10046 82 10102 160
rect 9968 54 10102 82
rect 9494 -300 9550 54
rect 9770 -300 9826 54
rect 10046 -300 10102 54
rect 10322 -300 10378 160
rect 10428 82 10456 1158
rect 10520 950 10548 1906
rect 11060 1760 11112 1766
rect 10980 1720 11060 1748
rect 10508 944 10560 950
rect 10508 886 10560 892
rect 10598 82 10654 160
rect 10428 54 10654 82
rect 10598 -300 10654 54
rect 10874 82 10930 160
rect 10980 82 11008 1720
rect 11060 1702 11112 1708
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 10874 54 11008 82
rect 11072 82 11100 1362
rect 11348 1329 11376 2382
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11532 1358 11560 2246
rect 11716 2145 11744 2382
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 13084 2304 13136 2310
rect 13084 2246 13136 2252
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 11702 2136 11758 2145
rect 11702 2071 11758 2080
rect 11624 1822 11836 1850
rect 11520 1352 11572 1358
rect 11334 1320 11390 1329
rect 11520 1294 11572 1300
rect 11334 1255 11390 1264
rect 11152 1216 11204 1222
rect 11204 1176 11284 1204
rect 11152 1158 11204 1164
rect 11150 82 11206 160
rect 11072 54 11206 82
rect 11256 82 11284 1176
rect 11624 898 11652 1822
rect 11808 1766 11836 1822
rect 11704 1760 11756 1766
rect 11704 1702 11756 1708
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11716 1290 11744 1702
rect 11900 1358 11928 2246
rect 12452 2106 12480 2246
rect 12679 2204 12987 2213
rect 12679 2202 12685 2204
rect 12741 2202 12765 2204
rect 12821 2202 12845 2204
rect 12901 2202 12925 2204
rect 12981 2202 12987 2204
rect 12741 2150 12743 2202
rect 12923 2150 12925 2202
rect 12679 2148 12685 2150
rect 12741 2148 12765 2150
rect 12821 2148 12845 2150
rect 12901 2148 12925 2150
rect 12981 2148 12987 2150
rect 12679 2139 12987 2148
rect 12440 2100 12492 2106
rect 12440 2042 12492 2048
rect 12532 2100 12584 2106
rect 12532 2042 12584 2048
rect 12072 1964 12124 1970
rect 12072 1906 12124 1912
rect 11888 1352 11940 1358
rect 11888 1294 11940 1300
rect 11704 1284 11756 1290
rect 11704 1226 11756 1232
rect 11796 1216 11848 1222
rect 11848 1176 12020 1204
rect 11796 1158 11848 1164
rect 11624 870 11744 898
rect 11716 160 11744 870
rect 11992 160 12020 1176
rect 12084 678 12112 1906
rect 12544 1306 12572 2042
rect 12624 1760 12676 1766
rect 12624 1702 12676 1708
rect 12900 1760 12952 1766
rect 12900 1702 12952 1708
rect 12636 1358 12664 1702
rect 12452 1278 12572 1306
rect 12624 1352 12676 1358
rect 12624 1294 12676 1300
rect 12164 1216 12216 1222
rect 12216 1176 12296 1204
rect 12164 1158 12216 1164
rect 12072 672 12124 678
rect 12072 614 12124 620
rect 12268 160 12296 1176
rect 12452 610 12480 1278
rect 12532 1216 12584 1222
rect 12912 1204 12940 1702
rect 13096 1358 13124 2246
rect 13084 1352 13136 1358
rect 13084 1294 13136 1300
rect 13176 1216 13228 1222
rect 12912 1176 13124 1204
rect 12532 1158 12584 1164
rect 12440 604 12492 610
rect 12440 546 12492 552
rect 12544 160 12572 1158
rect 12679 1116 12987 1125
rect 12679 1114 12685 1116
rect 12741 1114 12765 1116
rect 12821 1114 12845 1116
rect 12901 1114 12925 1116
rect 12981 1114 12987 1116
rect 12741 1062 12743 1114
rect 12923 1062 12925 1114
rect 12679 1060 12685 1062
rect 12741 1060 12765 1062
rect 12821 1060 12845 1062
rect 12901 1060 12925 1062
rect 12981 1060 12987 1062
rect 12679 1051 12987 1060
rect 13096 490 13124 1176
rect 13176 1158 13228 1164
rect 13004 462 13124 490
rect 11426 82 11482 160
rect 11256 54 11482 82
rect 10874 -300 10930 54
rect 11150 -300 11206 54
rect 11426 -300 11482 54
rect 11702 -300 11758 160
rect 11978 -300 12034 160
rect 12254 -300 12310 160
rect 12530 -300 12586 160
rect 12806 82 12862 160
rect 13004 82 13032 462
rect 13188 354 13216 1158
rect 13096 326 13216 354
rect 13096 160 13124 326
rect 12806 54 13032 82
rect 12806 -300 12862 54
rect 13082 -300 13138 160
rect 13280 134 13308 2246
rect 13648 1970 13676 2382
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13740 1970 13768 2246
rect 13452 1964 13504 1970
rect 13452 1906 13504 1912
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 13728 1964 13780 1970
rect 13728 1906 13780 1912
rect 14004 1964 14056 1970
rect 14004 1906 14056 1912
rect 13360 1896 13412 1902
rect 13360 1838 13412 1844
rect 13372 1465 13400 1838
rect 13358 1456 13414 1465
rect 13358 1391 13414 1400
rect 13360 1216 13412 1222
rect 13360 1158 13412 1164
rect 13372 160 13400 1158
rect 13464 338 13492 1906
rect 13544 1760 13596 1766
rect 13544 1702 13596 1708
rect 13636 1760 13688 1766
rect 13636 1702 13688 1708
rect 13556 1358 13584 1702
rect 13648 1358 13676 1702
rect 13912 1556 13964 1562
rect 13740 1516 13912 1544
rect 13544 1352 13596 1358
rect 13544 1294 13596 1300
rect 13636 1352 13688 1358
rect 13636 1294 13688 1300
rect 13452 332 13504 338
rect 13452 274 13504 280
rect 13268 128 13320 134
rect 13268 70 13320 76
rect 13358 -300 13414 160
rect 13634 82 13690 160
rect 13740 82 13768 1516
rect 13912 1498 13964 1504
rect 13912 1216 13964 1222
rect 13912 1158 13964 1164
rect 13924 160 13952 1158
rect 14016 377 14044 1906
rect 14108 746 14136 2790
rect 14278 2680 14334 2689
rect 14278 2615 14334 2624
rect 14292 1970 14320 2615
rect 14384 1970 14412 2926
rect 15612 2748 15920 2757
rect 15612 2746 15618 2748
rect 15674 2746 15698 2748
rect 15754 2746 15778 2748
rect 15834 2746 15858 2748
rect 15914 2746 15920 2748
rect 15674 2694 15676 2746
rect 15856 2694 15858 2746
rect 15612 2692 15618 2694
rect 15674 2692 15698 2694
rect 15754 2692 15778 2694
rect 15834 2692 15858 2694
rect 15914 2692 15920 2694
rect 15612 2683 15920 2692
rect 14568 2650 14872 2666
rect 14568 2644 14884 2650
rect 14568 2638 14832 2644
rect 14568 2514 14596 2638
rect 14832 2586 14884 2592
rect 14556 2508 14608 2514
rect 14556 2450 14608 2456
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15120 2106 15148 2246
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 15108 2100 15160 2106
rect 15108 2042 15160 2048
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 14096 740 14148 746
rect 14096 682 14148 688
rect 14002 368 14058 377
rect 14002 303 14058 312
rect 14568 218 14596 2042
rect 15384 2032 15436 2038
rect 15384 1974 15436 1980
rect 14924 1896 14976 1902
rect 14844 1844 14924 1850
rect 14844 1838 14976 1844
rect 14844 1822 14964 1838
rect 15200 1828 15252 1834
rect 14740 1556 14792 1562
rect 14384 190 14596 218
rect 14660 1516 14740 1544
rect 13634 54 13768 82
rect 13634 -300 13690 54
rect 13910 -300 13966 160
rect 14186 82 14242 160
rect 14384 82 14412 190
rect 14186 54 14412 82
rect 14462 82 14518 160
rect 14660 82 14688 1516
rect 14740 1498 14792 1504
rect 14844 1494 14872 1822
rect 15200 1770 15252 1776
rect 14924 1760 14976 1766
rect 14924 1702 14976 1708
rect 14936 1494 14964 1702
rect 14832 1488 14884 1494
rect 14832 1430 14884 1436
rect 14924 1488 14976 1494
rect 14924 1430 14976 1436
rect 15108 1488 15160 1494
rect 15108 1430 15160 1436
rect 15120 1306 15148 1430
rect 15212 1358 15240 1770
rect 15292 1760 15344 1766
rect 15292 1702 15344 1708
rect 14936 1278 15148 1306
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 14462 54 14688 82
rect 14738 82 14794 160
rect 14936 82 14964 1278
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 15028 160 15056 1158
rect 15304 160 15332 1702
rect 15396 1358 15424 1974
rect 15568 1964 15620 1970
rect 15488 1924 15568 1952
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 14738 54 14964 82
rect 14186 -300 14242 54
rect 14462 -300 14518 54
rect 14738 -300 14794 54
rect 15014 -300 15070 160
rect 15290 -300 15346 160
rect 15488 82 15516 1924
rect 15568 1906 15620 1912
rect 15612 1660 15920 1669
rect 15612 1658 15618 1660
rect 15674 1658 15698 1660
rect 15754 1658 15778 1660
rect 15834 1658 15858 1660
rect 15914 1658 15920 1660
rect 15674 1606 15676 1658
rect 15856 1606 15858 1658
rect 15612 1604 15618 1606
rect 15674 1604 15698 1606
rect 15754 1604 15778 1606
rect 15834 1604 15858 1606
rect 15914 1604 15920 1606
rect 15612 1595 15920 1604
rect 15948 406 15976 2382
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16316 1562 16344 1906
rect 16396 1760 16448 1766
rect 16396 1702 16448 1708
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 16028 1488 16080 1494
rect 16028 1430 16080 1436
rect 15936 400 15988 406
rect 15936 342 15988 348
rect 15566 82 15622 160
rect 15488 54 15622 82
rect 15566 -300 15622 54
rect 15842 82 15898 160
rect 16040 82 16068 1430
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16132 814 16160 1294
rect 16304 1284 16356 1290
rect 16304 1226 16356 1232
rect 16120 808 16172 814
rect 16120 750 16172 756
rect 16316 626 16344 1226
rect 16132 598 16344 626
rect 16132 160 16160 598
rect 16408 160 16436 1702
rect 16500 1442 16528 3062
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16684 2038 16712 2858
rect 17144 2514 17172 7822
rect 18544 7644 18852 7653
rect 18544 7642 18550 7644
rect 18606 7642 18630 7644
rect 18686 7642 18710 7644
rect 18766 7642 18790 7644
rect 18846 7642 18852 7644
rect 18606 7590 18608 7642
rect 18788 7590 18790 7642
rect 18544 7588 18550 7590
rect 18606 7588 18630 7590
rect 18686 7588 18710 7590
rect 18766 7588 18790 7590
rect 18846 7588 18852 7590
rect 18544 7579 18852 7588
rect 18544 6556 18852 6565
rect 18544 6554 18550 6556
rect 18606 6554 18630 6556
rect 18686 6554 18710 6556
rect 18766 6554 18790 6556
rect 18846 6554 18852 6556
rect 18606 6502 18608 6554
rect 18788 6502 18790 6554
rect 18544 6500 18550 6502
rect 18606 6500 18630 6502
rect 18686 6500 18710 6502
rect 18766 6500 18790 6502
rect 18846 6500 18852 6502
rect 18544 6491 18852 6500
rect 18544 5468 18852 5477
rect 18544 5466 18550 5468
rect 18606 5466 18630 5468
rect 18686 5466 18710 5468
rect 18766 5466 18790 5468
rect 18846 5466 18852 5468
rect 18606 5414 18608 5466
rect 18788 5414 18790 5466
rect 18544 5412 18550 5414
rect 18606 5412 18630 5414
rect 18686 5412 18710 5414
rect 18766 5412 18790 5414
rect 18846 5412 18852 5414
rect 18544 5403 18852 5412
rect 18544 4380 18852 4389
rect 18544 4378 18550 4380
rect 18606 4378 18630 4380
rect 18686 4378 18710 4380
rect 18766 4378 18790 4380
rect 18846 4378 18852 4380
rect 18606 4326 18608 4378
rect 18788 4326 18790 4378
rect 18544 4324 18550 4326
rect 18606 4324 18630 4326
rect 18686 4324 18710 4326
rect 18766 4324 18790 4326
rect 18846 4324 18852 4326
rect 18544 4315 18852 4324
rect 18544 3292 18852 3301
rect 18544 3290 18550 3292
rect 18606 3290 18630 3292
rect 18686 3290 18710 3292
rect 18766 3290 18790 3292
rect 18846 3290 18852 3292
rect 18606 3238 18608 3290
rect 18788 3238 18790 3290
rect 18544 3236 18550 3238
rect 18606 3236 18630 3238
rect 18686 3236 18710 3238
rect 18766 3236 18790 3238
rect 18846 3236 18852 3238
rect 18544 3227 18852 3236
rect 17958 2952 18014 2961
rect 17958 2887 18014 2896
rect 17408 2576 17460 2582
rect 17408 2518 17460 2524
rect 17132 2508 17184 2514
rect 17132 2450 17184 2456
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16672 2032 16724 2038
rect 16672 1974 16724 1980
rect 16672 1828 16724 1834
rect 16672 1770 16724 1776
rect 16500 1414 16620 1442
rect 16592 898 16620 1414
rect 16500 870 16620 898
rect 16500 678 16528 870
rect 16488 672 16540 678
rect 16488 614 16540 620
rect 16684 160 16712 1770
rect 16776 882 16804 2382
rect 17132 2304 17184 2310
rect 17132 2246 17184 2252
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 16948 1556 17000 1562
rect 16948 1498 17000 1504
rect 16854 1456 16910 1465
rect 16854 1391 16910 1400
rect 16868 1358 16896 1391
rect 16856 1352 16908 1358
rect 16856 1294 16908 1300
rect 16764 876 16816 882
rect 16764 818 16816 824
rect 16960 160 16988 1498
rect 17144 1358 17172 2246
rect 17236 2106 17264 2246
rect 17420 2106 17448 2518
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 17224 2100 17276 2106
rect 17224 2042 17276 2048
rect 17408 2100 17460 2106
rect 17408 2042 17460 2048
rect 17500 1828 17552 1834
rect 17236 1788 17500 1816
rect 17132 1352 17184 1358
rect 17132 1294 17184 1300
rect 17236 160 17264 1788
rect 17500 1770 17552 1776
rect 17592 1760 17644 1766
rect 17592 1702 17644 1708
rect 17604 898 17632 1702
rect 17512 870 17632 898
rect 17512 160 17540 870
rect 17696 542 17724 2382
rect 17972 2038 18000 2887
rect 19260 2650 19288 8434
rect 21477 8188 21785 8197
rect 21477 8186 21483 8188
rect 21539 8186 21563 8188
rect 21619 8186 21643 8188
rect 21699 8186 21723 8188
rect 21779 8186 21785 8188
rect 21539 8134 21541 8186
rect 21721 8134 21723 8186
rect 21477 8132 21483 8134
rect 21539 8132 21563 8134
rect 21619 8132 21643 8134
rect 21699 8132 21723 8134
rect 21779 8132 21785 8134
rect 21477 8123 21785 8132
rect 21477 7100 21785 7109
rect 21477 7098 21483 7100
rect 21539 7098 21563 7100
rect 21619 7098 21643 7100
rect 21699 7098 21723 7100
rect 21779 7098 21785 7100
rect 21539 7046 21541 7098
rect 21721 7046 21723 7098
rect 21477 7044 21483 7046
rect 21539 7044 21563 7046
rect 21619 7044 21643 7046
rect 21699 7044 21723 7046
rect 21779 7044 21785 7046
rect 21477 7035 21785 7044
rect 21477 6012 21785 6021
rect 21477 6010 21483 6012
rect 21539 6010 21563 6012
rect 21619 6010 21643 6012
rect 21699 6010 21723 6012
rect 21779 6010 21785 6012
rect 21539 5958 21541 6010
rect 21721 5958 21723 6010
rect 21477 5956 21483 5958
rect 21539 5956 21563 5958
rect 21619 5956 21643 5958
rect 21699 5956 21723 5958
rect 21779 5956 21785 5958
rect 21477 5947 21785 5956
rect 21477 4924 21785 4933
rect 21477 4922 21483 4924
rect 21539 4922 21563 4924
rect 21619 4922 21643 4924
rect 21699 4922 21723 4924
rect 21779 4922 21785 4924
rect 21539 4870 21541 4922
rect 21721 4870 21723 4922
rect 21477 4868 21483 4870
rect 21539 4868 21563 4870
rect 21619 4868 21643 4870
rect 21699 4868 21723 4870
rect 21779 4868 21785 4870
rect 21477 4859 21785 4868
rect 19984 4140 20036 4146
rect 19984 4082 20036 4088
rect 19798 4040 19854 4049
rect 19798 3975 19800 3984
rect 19852 3975 19854 3984
rect 19800 3946 19852 3952
rect 19996 3738 20024 4082
rect 21477 3836 21785 3845
rect 21477 3834 21483 3836
rect 21539 3834 21563 3836
rect 21619 3834 21643 3836
rect 21699 3834 21723 3836
rect 21779 3834 21785 3836
rect 21539 3782 21541 3834
rect 21721 3782 21723 3834
rect 21477 3780 21483 3782
rect 21539 3780 21563 3782
rect 21619 3780 21643 3782
rect 21699 3780 21723 3782
rect 21779 3780 21785 3782
rect 21477 3771 21785 3780
rect 19984 3732 20036 3738
rect 19984 3674 20036 3680
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 19536 3126 19564 3538
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 19892 3392 19944 3398
rect 19892 3334 19944 3340
rect 19904 3194 19932 3334
rect 19892 3188 19944 3194
rect 19892 3130 19944 3136
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19892 2848 19944 2854
rect 19892 2790 19944 2796
rect 19248 2644 19300 2650
rect 19248 2586 19300 2592
rect 18144 2576 18196 2582
rect 18144 2518 18196 2524
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 17960 2032 18012 2038
rect 17960 1974 18012 1980
rect 18064 1902 18092 2246
rect 18052 1896 18104 1902
rect 18052 1838 18104 1844
rect 18052 1760 18104 1766
rect 18052 1702 18104 1708
rect 17868 1420 17920 1426
rect 17788 1380 17868 1408
rect 17684 536 17736 542
rect 17684 478 17736 484
rect 17788 160 17816 1380
rect 17868 1362 17920 1368
rect 18064 160 18092 1702
rect 18156 1358 18184 2518
rect 19904 2446 19932 2790
rect 18236 2440 18288 2446
rect 19064 2440 19116 2446
rect 18288 2400 18368 2428
rect 18236 2382 18288 2388
rect 18340 1578 18368 2400
rect 19892 2440 19944 2446
rect 19064 2382 19116 2388
rect 19614 2408 19670 2417
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18432 2106 18460 2246
rect 18544 2204 18852 2213
rect 18544 2202 18550 2204
rect 18606 2202 18630 2204
rect 18686 2202 18710 2204
rect 18766 2202 18790 2204
rect 18846 2202 18852 2204
rect 18606 2150 18608 2202
rect 18788 2150 18790 2202
rect 18544 2148 18550 2150
rect 18606 2148 18630 2150
rect 18686 2148 18710 2150
rect 18766 2148 18790 2150
rect 18846 2148 18852 2150
rect 18544 2139 18852 2148
rect 18420 2100 18472 2106
rect 18420 2042 18472 2048
rect 18972 1760 19024 1766
rect 18972 1702 19024 1708
rect 18340 1550 18460 1578
rect 18144 1352 18196 1358
rect 18144 1294 18196 1300
rect 18236 1284 18288 1290
rect 18236 1226 18288 1232
rect 18248 610 18276 1226
rect 18432 785 18460 1550
rect 18880 1488 18932 1494
rect 18880 1430 18932 1436
rect 18544 1116 18852 1125
rect 18544 1114 18550 1116
rect 18606 1114 18630 1116
rect 18686 1114 18710 1116
rect 18766 1114 18790 1116
rect 18846 1114 18852 1116
rect 18606 1062 18608 1114
rect 18788 1062 18790 1114
rect 18544 1060 18550 1062
rect 18606 1060 18630 1062
rect 18686 1060 18710 1062
rect 18766 1060 18790 1062
rect 18846 1060 18852 1062
rect 18544 1051 18852 1060
rect 18418 776 18474 785
rect 18418 711 18474 720
rect 18420 672 18472 678
rect 18340 620 18420 626
rect 18340 614 18472 620
rect 18236 604 18288 610
rect 18236 546 18288 552
rect 18340 598 18460 614
rect 18340 160 18368 598
rect 18892 474 18920 1430
rect 18880 468 18932 474
rect 18880 410 18932 416
rect 18984 354 19012 1702
rect 18800 326 19012 354
rect 15842 54 16068 82
rect 15842 -300 15898 54
rect 16118 -300 16174 160
rect 16394 -300 16450 160
rect 16670 -300 16726 160
rect 16946 -300 17002 160
rect 17222 -300 17278 160
rect 17498 -300 17554 160
rect 17774 -300 17830 160
rect 18050 -300 18106 160
rect 18326 -300 18382 160
rect 18602 82 18658 160
rect 18800 82 18828 326
rect 18880 264 18932 270
rect 19076 241 19104 2382
rect 19892 2382 19944 2388
rect 19984 2440 20036 2446
rect 20036 2400 20116 2428
rect 19984 2382 20036 2388
rect 19614 2343 19616 2352
rect 19668 2343 19670 2352
rect 19616 2314 19668 2320
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19156 1828 19208 1834
rect 19156 1770 19208 1776
rect 18880 206 18932 212
rect 19062 232 19118 241
rect 18892 160 18920 206
rect 19062 167 19118 176
rect 19168 160 19196 1770
rect 19260 1358 19288 2246
rect 19616 1896 19668 1902
rect 19616 1838 19668 1844
rect 19524 1556 19576 1562
rect 19352 1516 19524 1544
rect 19248 1352 19300 1358
rect 19248 1294 19300 1300
rect 19352 1204 19380 1516
rect 19524 1498 19576 1504
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 19536 1204 19564 1294
rect 19628 1290 19656 1838
rect 19892 1760 19944 1766
rect 19892 1702 19944 1708
rect 19616 1284 19668 1290
rect 19616 1226 19668 1232
rect 19260 1176 19380 1204
rect 19444 1176 19564 1204
rect 19260 678 19288 1176
rect 19248 672 19300 678
rect 19248 614 19300 620
rect 19444 160 19472 1176
rect 18602 54 18828 82
rect 18602 -300 18658 54
rect 18878 -300 18934 160
rect 19154 -300 19210 160
rect 19430 -300 19486 160
rect 19706 82 19762 160
rect 19904 82 19932 1702
rect 19984 1012 20036 1018
rect 19984 954 20036 960
rect 19996 160 20024 954
rect 20088 649 20116 2400
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 20180 2106 20208 2246
rect 20168 2100 20220 2106
rect 20168 2042 20220 2048
rect 20640 1290 20668 3470
rect 21477 2748 21785 2757
rect 21477 2746 21483 2748
rect 21539 2746 21563 2748
rect 21619 2746 21643 2748
rect 21699 2746 21723 2748
rect 21779 2746 21785 2748
rect 21539 2694 21541 2746
rect 21721 2694 21723 2746
rect 21477 2692 21483 2694
rect 21539 2692 21563 2694
rect 21619 2692 21643 2694
rect 21699 2692 21723 2694
rect 21779 2692 21785 2694
rect 21477 2683 21785 2692
rect 20812 2576 20864 2582
rect 20812 2518 20864 2524
rect 20720 1896 20772 1902
rect 20720 1838 20772 1844
rect 20628 1284 20680 1290
rect 20628 1226 20680 1232
rect 20536 944 20588 950
rect 20536 886 20588 892
rect 20074 640 20130 649
rect 20074 575 20130 584
rect 20444 604 20496 610
rect 20444 546 20496 552
rect 19706 54 19932 82
rect 19706 -300 19762 54
rect 19982 -300 20038 160
rect 20258 82 20314 160
rect 20456 82 20484 546
rect 20548 160 20576 886
rect 20732 785 20760 1838
rect 20824 1766 20852 2518
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 21548 2100 21600 2106
rect 21548 2042 21600 2048
rect 21560 2009 21588 2042
rect 21546 2000 21602 2009
rect 21546 1935 21602 1944
rect 21178 1864 21234 1873
rect 21178 1799 21180 1808
rect 21232 1799 21234 1808
rect 21180 1770 21232 1776
rect 20812 1760 20864 1766
rect 20812 1702 20864 1708
rect 21477 1660 21785 1669
rect 21477 1658 21483 1660
rect 21539 1658 21563 1660
rect 21619 1658 21643 1660
rect 21699 1658 21723 1660
rect 21779 1658 21785 1660
rect 21539 1606 21541 1658
rect 21721 1606 21723 1658
rect 21477 1604 21483 1606
rect 21539 1604 21563 1606
rect 21619 1604 21643 1606
rect 21699 1604 21723 1606
rect 21779 1604 21785 1606
rect 21477 1595 21785 1604
rect 21836 1562 21864 2314
rect 22020 2106 22048 8434
rect 22560 8424 22612 8430
rect 22560 8366 22612 8372
rect 22376 2984 22428 2990
rect 22376 2926 22428 2932
rect 22008 2100 22060 2106
rect 22008 2042 22060 2048
rect 22192 2032 22244 2038
rect 22192 1974 22244 1980
rect 21824 1556 21876 1562
rect 21824 1498 21876 1504
rect 22100 1488 22152 1494
rect 22020 1436 22100 1442
rect 22020 1430 22152 1436
rect 21364 1420 21416 1426
rect 21100 1380 21364 1408
rect 20718 776 20774 785
rect 20718 711 20774 720
rect 20904 672 20956 678
rect 20904 614 20956 620
rect 20916 354 20944 614
rect 20824 326 20944 354
rect 20824 160 20852 326
rect 21100 160 21128 1380
rect 21364 1362 21416 1368
rect 22020 1414 22140 1430
rect 21456 1352 21508 1358
rect 21456 1294 21508 1300
rect 21548 1352 21600 1358
rect 21548 1294 21600 1300
rect 21468 921 21496 1294
rect 21560 1018 21588 1294
rect 21732 1284 21784 1290
rect 21732 1226 21784 1232
rect 21548 1012 21600 1018
rect 21548 954 21600 960
rect 21454 912 21510 921
rect 21454 847 21510 856
rect 21364 808 21416 814
rect 21364 750 21416 756
rect 21376 160 21404 750
rect 21640 740 21692 746
rect 21640 682 21692 688
rect 21652 160 21680 682
rect 21744 610 21772 1226
rect 21732 604 21784 610
rect 21732 546 21784 552
rect 20258 54 20484 82
rect 20258 -300 20314 54
rect 20534 -300 20590 160
rect 20810 -300 20866 160
rect 21086 -300 21142 160
rect 21362 -300 21418 160
rect 21638 -300 21694 160
rect 21914 82 21970 160
rect 22020 82 22048 1414
rect 22204 1222 22232 1974
rect 22284 1964 22336 1970
rect 22284 1906 22336 1912
rect 22296 1562 22324 1906
rect 22284 1556 22336 1562
rect 22284 1498 22336 1504
rect 22192 1216 22244 1222
rect 22192 1158 22244 1164
rect 21914 54 22048 82
rect 22190 82 22246 160
rect 22388 82 22416 2926
rect 22572 2774 22600 8366
rect 22744 4072 22796 4078
rect 22744 4014 22796 4020
rect 22756 3194 22784 4014
rect 23492 3942 23520 8434
rect 23480 3936 23532 3942
rect 23480 3878 23532 3884
rect 23204 3664 23256 3670
rect 23204 3606 23256 3612
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 23020 3052 23072 3058
rect 23020 2994 23072 3000
rect 22664 2938 22692 2994
rect 22664 2910 22876 2938
rect 22572 2746 22692 2774
rect 22560 2576 22612 2582
rect 22560 2518 22612 2524
rect 22572 2106 22600 2518
rect 22664 2106 22692 2746
rect 22744 2440 22796 2446
rect 22744 2382 22796 2388
rect 22560 2100 22612 2106
rect 22560 2042 22612 2048
rect 22652 2100 22704 2106
rect 22652 2042 22704 2048
rect 22652 1964 22704 1970
rect 22652 1906 22704 1912
rect 22664 1578 22692 1906
rect 22756 1766 22784 2382
rect 22744 1760 22796 1766
rect 22744 1702 22796 1708
rect 22664 1562 22784 1578
rect 22664 1556 22796 1562
rect 22664 1550 22744 1556
rect 22744 1498 22796 1504
rect 22744 1420 22796 1426
rect 22744 1362 22796 1368
rect 22560 1352 22612 1358
rect 22560 1294 22612 1300
rect 22652 1352 22704 1358
rect 22652 1294 22704 1300
rect 22572 1018 22600 1294
rect 22560 1012 22612 1018
rect 22560 954 22612 960
rect 22664 678 22692 1294
rect 22652 672 22704 678
rect 22652 614 22704 620
rect 22756 490 22784 1362
rect 22480 462 22784 490
rect 22480 160 22508 462
rect 22744 400 22796 406
rect 22744 342 22796 348
rect 22756 160 22784 342
rect 22190 54 22416 82
rect 21914 -300 21970 54
rect 22190 -300 22246 54
rect 22466 -300 22522 160
rect 22742 -300 22798 160
rect 22848 82 22876 2910
rect 23032 2417 23060 2994
rect 23112 2848 23164 2854
rect 23112 2790 23164 2796
rect 23124 2650 23152 2790
rect 23112 2644 23164 2650
rect 23112 2586 23164 2592
rect 23018 2408 23074 2417
rect 22928 2372 22980 2378
rect 23216 2360 23244 3606
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23018 2343 23074 2352
rect 22928 2314 22980 2320
rect 23124 2332 23244 2360
rect 22940 1737 22968 2314
rect 23020 2032 23072 2038
rect 23020 1974 23072 1980
rect 22926 1728 22982 1737
rect 22926 1663 22982 1672
rect 22928 1216 22980 1222
rect 22928 1158 22980 1164
rect 22940 377 22968 1158
rect 23032 406 23060 1974
rect 23124 1970 23152 2332
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 23112 1964 23164 1970
rect 23112 1906 23164 1912
rect 23216 1834 23244 2042
rect 23204 1828 23256 1834
rect 23204 1770 23256 1776
rect 23204 1352 23256 1358
rect 23124 1300 23204 1306
rect 23124 1294 23256 1300
rect 23124 1278 23244 1294
rect 23124 814 23152 1278
rect 23204 1216 23256 1222
rect 23204 1158 23256 1164
rect 23112 808 23164 814
rect 23112 750 23164 756
rect 23216 678 23244 1158
rect 23204 672 23256 678
rect 23204 614 23256 620
rect 23020 400 23072 406
rect 22926 368 22982 377
rect 23020 342 23072 348
rect 22926 303 22982 312
rect 23308 160 23336 3470
rect 23480 3392 23532 3398
rect 23480 3334 23532 3340
rect 23388 2984 23440 2990
rect 23388 2926 23440 2932
rect 23400 2854 23428 2926
rect 23492 2854 23520 3334
rect 23664 3188 23716 3194
rect 23664 3130 23716 3136
rect 23388 2848 23440 2854
rect 23388 2790 23440 2796
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23572 2848 23624 2854
rect 23572 2790 23624 2796
rect 23584 2446 23612 2790
rect 23572 2440 23624 2446
rect 23572 2382 23624 2388
rect 23480 2372 23532 2378
rect 23480 2314 23532 2320
rect 23388 1964 23440 1970
rect 23388 1906 23440 1912
rect 23400 1494 23428 1906
rect 23388 1488 23440 1494
rect 23388 1430 23440 1436
rect 23018 82 23074 160
rect 22848 54 23074 82
rect 23018 -300 23074 54
rect 23294 -300 23350 160
rect 23492 82 23520 2314
rect 23570 2272 23626 2281
rect 23570 2207 23626 2216
rect 23584 1834 23612 2207
rect 23572 1828 23624 1834
rect 23572 1770 23624 1776
rect 23570 1728 23626 1737
rect 23570 1663 23626 1672
rect 23584 1494 23612 1663
rect 23572 1488 23624 1494
rect 23572 1430 23624 1436
rect 23676 1358 23704 3130
rect 23768 2650 23796 8434
rect 24780 8430 24808 9840
rect 24860 8560 24912 8566
rect 24860 8502 24912 8508
rect 24768 8424 24820 8430
rect 24768 8366 24820 8372
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23848 3052 23900 3058
rect 23848 2994 23900 3000
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23756 1964 23808 1970
rect 23756 1906 23808 1912
rect 23768 1426 23796 1906
rect 23756 1420 23808 1426
rect 23756 1362 23808 1368
rect 23664 1352 23716 1358
rect 23664 1294 23716 1300
rect 23756 1216 23808 1222
rect 23756 1158 23808 1164
rect 23768 1018 23796 1158
rect 23756 1012 23808 1018
rect 23756 954 23808 960
rect 23860 160 23888 2994
rect 23952 2106 23980 8298
rect 24409 7644 24717 7653
rect 24409 7642 24415 7644
rect 24471 7642 24495 7644
rect 24551 7642 24575 7644
rect 24631 7642 24655 7644
rect 24711 7642 24717 7644
rect 24471 7590 24473 7642
rect 24653 7590 24655 7642
rect 24409 7588 24415 7590
rect 24471 7588 24495 7590
rect 24551 7588 24575 7590
rect 24631 7588 24655 7590
rect 24711 7588 24717 7590
rect 24409 7579 24717 7588
rect 24409 6556 24717 6565
rect 24409 6554 24415 6556
rect 24471 6554 24495 6556
rect 24551 6554 24575 6556
rect 24631 6554 24655 6556
rect 24711 6554 24717 6556
rect 24471 6502 24473 6554
rect 24653 6502 24655 6554
rect 24409 6500 24415 6502
rect 24471 6500 24495 6502
rect 24551 6500 24575 6502
rect 24631 6500 24655 6502
rect 24711 6500 24717 6502
rect 24409 6491 24717 6500
rect 24409 5468 24717 5477
rect 24409 5466 24415 5468
rect 24471 5466 24495 5468
rect 24551 5466 24575 5468
rect 24631 5466 24655 5468
rect 24711 5466 24717 5468
rect 24471 5414 24473 5466
rect 24653 5414 24655 5466
rect 24409 5412 24415 5414
rect 24471 5412 24495 5414
rect 24551 5412 24575 5414
rect 24631 5412 24655 5414
rect 24711 5412 24717 5414
rect 24409 5403 24717 5412
rect 24409 4380 24717 4389
rect 24409 4378 24415 4380
rect 24471 4378 24495 4380
rect 24551 4378 24575 4380
rect 24631 4378 24655 4380
rect 24711 4378 24717 4380
rect 24471 4326 24473 4378
rect 24653 4326 24655 4378
rect 24409 4324 24415 4326
rect 24471 4324 24495 4326
rect 24551 4324 24575 4326
rect 24631 4324 24655 4326
rect 24711 4324 24717 4326
rect 24409 4315 24717 4324
rect 24032 4140 24084 4146
rect 24032 4082 24084 4088
rect 24044 3738 24072 4082
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 24216 3664 24268 3670
rect 24216 3606 24268 3612
rect 24032 2304 24084 2310
rect 24032 2246 24084 2252
rect 24124 2304 24176 2310
rect 24124 2246 24176 2252
rect 23940 2100 23992 2106
rect 23940 2042 23992 2048
rect 24044 1358 24072 2246
rect 23940 1352 23992 1358
rect 23940 1294 23992 1300
rect 24032 1352 24084 1358
rect 24032 1294 24084 1300
rect 23952 1018 23980 1294
rect 23940 1012 23992 1018
rect 23940 954 23992 960
rect 24136 160 24164 2246
rect 24228 2106 24256 3606
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 24216 2100 24268 2106
rect 24216 2042 24268 2048
rect 23570 82 23626 160
rect 23492 54 23626 82
rect 23570 -300 23626 54
rect 23846 -300 23902 160
rect 24122 -300 24178 160
rect 24320 82 24348 3538
rect 24409 3292 24717 3301
rect 24409 3290 24415 3292
rect 24471 3290 24495 3292
rect 24551 3290 24575 3292
rect 24631 3290 24655 3292
rect 24711 3290 24717 3292
rect 24471 3238 24473 3290
rect 24653 3238 24655 3290
rect 24409 3236 24415 3238
rect 24471 3236 24495 3238
rect 24551 3236 24575 3238
rect 24631 3236 24655 3238
rect 24711 3236 24717 3238
rect 24409 3227 24717 3236
rect 24674 2408 24730 2417
rect 24730 2366 24808 2394
rect 24674 2343 24730 2352
rect 24409 2204 24717 2213
rect 24409 2202 24415 2204
rect 24471 2202 24495 2204
rect 24551 2202 24575 2204
rect 24631 2202 24655 2204
rect 24711 2202 24717 2204
rect 24471 2150 24473 2202
rect 24653 2150 24655 2202
rect 24409 2148 24415 2150
rect 24471 2148 24495 2150
rect 24551 2148 24575 2150
rect 24631 2148 24655 2150
rect 24711 2148 24717 2150
rect 24409 2139 24717 2148
rect 24409 1116 24717 1125
rect 24409 1114 24415 1116
rect 24471 1114 24495 1116
rect 24551 1114 24575 1116
rect 24631 1114 24655 1116
rect 24711 1114 24717 1116
rect 24471 1062 24473 1114
rect 24653 1062 24655 1114
rect 24409 1060 24415 1062
rect 24471 1060 24495 1062
rect 24551 1060 24575 1062
rect 24631 1060 24655 1062
rect 24711 1060 24717 1062
rect 24409 1051 24717 1060
rect 24398 82 24454 160
rect 24320 54 24454 82
rect 24398 -300 24454 54
rect 24674 82 24730 160
rect 24780 82 24808 2366
rect 24872 1358 24900 8502
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 25228 1760 25280 1766
rect 25228 1702 25280 1708
rect 24952 1488 25004 1494
rect 24952 1430 25004 1436
rect 24860 1352 24912 1358
rect 24860 1294 24912 1300
rect 24964 160 24992 1430
rect 25240 160 25268 1702
rect 25516 160 25544 3062
rect 24674 54 24808 82
rect 24674 -300 24730 54
rect 24950 -300 25006 160
rect 25226 -300 25282 160
rect 25502 -300 25558 160
<< via2 >>
rect 6820 8730 6876 8732
rect 6900 8730 6956 8732
rect 6980 8730 7036 8732
rect 7060 8730 7116 8732
rect 6820 8678 6866 8730
rect 6866 8678 6876 8730
rect 6900 8678 6930 8730
rect 6930 8678 6942 8730
rect 6942 8678 6956 8730
rect 6980 8678 6994 8730
rect 6994 8678 7006 8730
rect 7006 8678 7036 8730
rect 7060 8678 7070 8730
rect 7070 8678 7116 8730
rect 6820 8676 6876 8678
rect 6900 8676 6956 8678
rect 6980 8676 7036 8678
rect 7060 8676 7116 8678
rect 12685 8730 12741 8732
rect 12765 8730 12821 8732
rect 12845 8730 12901 8732
rect 12925 8730 12981 8732
rect 12685 8678 12731 8730
rect 12731 8678 12741 8730
rect 12765 8678 12795 8730
rect 12795 8678 12807 8730
rect 12807 8678 12821 8730
rect 12845 8678 12859 8730
rect 12859 8678 12871 8730
rect 12871 8678 12901 8730
rect 12925 8678 12935 8730
rect 12935 8678 12981 8730
rect 12685 8676 12741 8678
rect 12765 8676 12821 8678
rect 12845 8676 12901 8678
rect 12925 8676 12981 8678
rect 18550 8730 18606 8732
rect 18630 8730 18686 8732
rect 18710 8730 18766 8732
rect 18790 8730 18846 8732
rect 18550 8678 18596 8730
rect 18596 8678 18606 8730
rect 18630 8678 18660 8730
rect 18660 8678 18672 8730
rect 18672 8678 18686 8730
rect 18710 8678 18724 8730
rect 18724 8678 18736 8730
rect 18736 8678 18766 8730
rect 18790 8678 18800 8730
rect 18800 8678 18846 8730
rect 18550 8676 18606 8678
rect 18630 8676 18686 8678
rect 18710 8676 18766 8678
rect 18790 8676 18846 8678
rect 24415 8730 24471 8732
rect 24495 8730 24551 8732
rect 24575 8730 24631 8732
rect 24655 8730 24711 8732
rect 24415 8678 24461 8730
rect 24461 8678 24471 8730
rect 24495 8678 24525 8730
rect 24525 8678 24537 8730
rect 24537 8678 24551 8730
rect 24575 8678 24589 8730
rect 24589 8678 24601 8730
rect 24601 8678 24631 8730
rect 24655 8678 24665 8730
rect 24665 8678 24711 8730
rect 24415 8676 24471 8678
rect 24495 8676 24551 8678
rect 24575 8676 24631 8678
rect 24655 8676 24711 8678
rect 2410 3984 2466 4040
rect 1766 2352 1822 2408
rect 3888 8186 3944 8188
rect 3968 8186 4024 8188
rect 4048 8186 4104 8188
rect 4128 8186 4184 8188
rect 3888 8134 3934 8186
rect 3934 8134 3944 8186
rect 3968 8134 3998 8186
rect 3998 8134 4010 8186
rect 4010 8134 4024 8186
rect 4048 8134 4062 8186
rect 4062 8134 4074 8186
rect 4074 8134 4104 8186
rect 4128 8134 4138 8186
rect 4138 8134 4184 8186
rect 3888 8132 3944 8134
rect 3968 8132 4024 8134
rect 4048 8132 4104 8134
rect 4128 8132 4184 8134
rect 3888 7098 3944 7100
rect 3968 7098 4024 7100
rect 4048 7098 4104 7100
rect 4128 7098 4184 7100
rect 3888 7046 3934 7098
rect 3934 7046 3944 7098
rect 3968 7046 3998 7098
rect 3998 7046 4010 7098
rect 4010 7046 4024 7098
rect 4048 7046 4062 7098
rect 4062 7046 4074 7098
rect 4074 7046 4104 7098
rect 4128 7046 4138 7098
rect 4138 7046 4184 7098
rect 3888 7044 3944 7046
rect 3968 7044 4024 7046
rect 4048 7044 4104 7046
rect 4128 7044 4184 7046
rect 3888 6010 3944 6012
rect 3968 6010 4024 6012
rect 4048 6010 4104 6012
rect 4128 6010 4184 6012
rect 3888 5958 3934 6010
rect 3934 5958 3944 6010
rect 3968 5958 3998 6010
rect 3998 5958 4010 6010
rect 4010 5958 4024 6010
rect 4048 5958 4062 6010
rect 4062 5958 4074 6010
rect 4074 5958 4104 6010
rect 4128 5958 4138 6010
rect 4138 5958 4184 6010
rect 3888 5956 3944 5958
rect 3968 5956 4024 5958
rect 4048 5956 4104 5958
rect 4128 5956 4184 5958
rect 3888 4922 3944 4924
rect 3968 4922 4024 4924
rect 4048 4922 4104 4924
rect 4128 4922 4184 4924
rect 3888 4870 3934 4922
rect 3934 4870 3944 4922
rect 3968 4870 3998 4922
rect 3998 4870 4010 4922
rect 4010 4870 4024 4922
rect 4048 4870 4062 4922
rect 4062 4870 4074 4922
rect 4074 4870 4104 4922
rect 4128 4870 4138 4922
rect 4138 4870 4184 4922
rect 3888 4868 3944 4870
rect 3968 4868 4024 4870
rect 4048 4868 4104 4870
rect 4128 4868 4184 4870
rect 3888 3834 3944 3836
rect 3968 3834 4024 3836
rect 4048 3834 4104 3836
rect 4128 3834 4184 3836
rect 3888 3782 3934 3834
rect 3934 3782 3944 3834
rect 3968 3782 3998 3834
rect 3998 3782 4010 3834
rect 4010 3782 4024 3834
rect 4048 3782 4062 3834
rect 4062 3782 4074 3834
rect 4074 3782 4104 3834
rect 4128 3782 4138 3834
rect 4138 3782 4184 3834
rect 3888 3780 3944 3782
rect 3968 3780 4024 3782
rect 4048 3780 4104 3782
rect 4128 3780 4184 3782
rect 4434 3032 4490 3088
rect 3888 2746 3944 2748
rect 3968 2746 4024 2748
rect 4048 2746 4104 2748
rect 4128 2746 4184 2748
rect 3888 2694 3934 2746
rect 3934 2694 3944 2746
rect 3968 2694 3998 2746
rect 3998 2694 4010 2746
rect 4010 2694 4024 2746
rect 4048 2694 4062 2746
rect 4062 2694 4074 2746
rect 4074 2694 4104 2746
rect 4128 2694 4138 2746
rect 4138 2694 4184 2746
rect 3888 2692 3944 2694
rect 3968 2692 4024 2694
rect 4048 2692 4104 2694
rect 4128 2692 4184 2694
rect 3606 1808 3662 1864
rect 3888 1658 3944 1660
rect 3968 1658 4024 1660
rect 4048 1658 4104 1660
rect 4128 1658 4184 1660
rect 3888 1606 3934 1658
rect 3934 1606 3944 1658
rect 3968 1606 3998 1658
rect 3998 1606 4010 1658
rect 4010 1606 4024 1658
rect 4048 1606 4062 1658
rect 4062 1606 4074 1658
rect 4074 1606 4104 1658
rect 4128 1606 4138 1658
rect 4138 1606 4184 1658
rect 3888 1604 3944 1606
rect 3968 1604 4024 1606
rect 4048 1604 4104 1606
rect 4128 1604 4184 1606
rect 4342 1536 4398 1592
rect 4802 1944 4858 2000
rect 1674 312 1730 368
rect 4894 1400 4950 1456
rect 4802 584 4858 640
rect 5354 856 5410 912
rect 6820 7642 6876 7644
rect 6900 7642 6956 7644
rect 6980 7642 7036 7644
rect 7060 7642 7116 7644
rect 6820 7590 6866 7642
rect 6866 7590 6876 7642
rect 6900 7590 6930 7642
rect 6930 7590 6942 7642
rect 6942 7590 6956 7642
rect 6980 7590 6994 7642
rect 6994 7590 7006 7642
rect 7006 7590 7036 7642
rect 7060 7590 7070 7642
rect 7070 7590 7116 7642
rect 6820 7588 6876 7590
rect 6900 7588 6956 7590
rect 6980 7588 7036 7590
rect 7060 7588 7116 7590
rect 6820 6554 6876 6556
rect 6900 6554 6956 6556
rect 6980 6554 7036 6556
rect 7060 6554 7116 6556
rect 6820 6502 6866 6554
rect 6866 6502 6876 6554
rect 6900 6502 6930 6554
rect 6930 6502 6942 6554
rect 6942 6502 6956 6554
rect 6980 6502 6994 6554
rect 6994 6502 7006 6554
rect 7006 6502 7036 6554
rect 7060 6502 7070 6554
rect 7070 6502 7116 6554
rect 6820 6500 6876 6502
rect 6900 6500 6956 6502
rect 6980 6500 7036 6502
rect 7060 6500 7116 6502
rect 6820 5466 6876 5468
rect 6900 5466 6956 5468
rect 6980 5466 7036 5468
rect 7060 5466 7116 5468
rect 6820 5414 6866 5466
rect 6866 5414 6876 5466
rect 6900 5414 6930 5466
rect 6930 5414 6942 5466
rect 6942 5414 6956 5466
rect 6980 5414 6994 5466
rect 6994 5414 7006 5466
rect 7006 5414 7036 5466
rect 7060 5414 7070 5466
rect 7070 5414 7116 5466
rect 6820 5412 6876 5414
rect 6900 5412 6956 5414
rect 6980 5412 7036 5414
rect 7060 5412 7116 5414
rect 6820 4378 6876 4380
rect 6900 4378 6956 4380
rect 6980 4378 7036 4380
rect 7060 4378 7116 4380
rect 6820 4326 6866 4378
rect 6866 4326 6876 4378
rect 6900 4326 6930 4378
rect 6930 4326 6942 4378
rect 6942 4326 6956 4378
rect 6980 4326 6994 4378
rect 6994 4326 7006 4378
rect 7006 4326 7036 4378
rect 7060 4326 7070 4378
rect 7070 4326 7116 4378
rect 6820 4324 6876 4326
rect 6900 4324 6956 4326
rect 6980 4324 7036 4326
rect 7060 4324 7116 4326
rect 6820 3290 6876 3292
rect 6900 3290 6956 3292
rect 6980 3290 7036 3292
rect 7060 3290 7116 3292
rect 6820 3238 6866 3290
rect 6866 3238 6876 3290
rect 6900 3238 6930 3290
rect 6930 3238 6942 3290
rect 6942 3238 6956 3290
rect 6980 3238 6994 3290
rect 6994 3238 7006 3290
rect 7006 3238 7036 3290
rect 7060 3238 7070 3290
rect 7070 3238 7116 3290
rect 6820 3236 6876 3238
rect 6900 3236 6956 3238
rect 6980 3236 7036 3238
rect 7060 3236 7116 3238
rect 5998 1708 6000 1728
rect 6000 1708 6052 1728
rect 6052 1708 6054 1728
rect 5998 1672 6054 1708
rect 6826 2896 6882 2952
rect 6826 2488 6882 2544
rect 6820 2202 6876 2204
rect 6900 2202 6956 2204
rect 6980 2202 7036 2204
rect 7060 2202 7116 2204
rect 6820 2150 6866 2202
rect 6866 2150 6876 2202
rect 6900 2150 6930 2202
rect 6930 2150 6942 2202
rect 6942 2150 6956 2202
rect 6980 2150 6994 2202
rect 6994 2150 7006 2202
rect 7006 2150 7036 2202
rect 7060 2150 7070 2202
rect 7070 2150 7116 2202
rect 6820 2148 6876 2150
rect 6900 2148 6956 2150
rect 6980 2148 7036 2150
rect 7060 2148 7116 2150
rect 9753 8186 9809 8188
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 9753 8134 9799 8186
rect 9799 8134 9809 8186
rect 9833 8134 9863 8186
rect 9863 8134 9875 8186
rect 9875 8134 9889 8186
rect 9913 8134 9927 8186
rect 9927 8134 9939 8186
rect 9939 8134 9969 8186
rect 9993 8134 10003 8186
rect 10003 8134 10049 8186
rect 9753 8132 9809 8134
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 9753 7098 9809 7100
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 9753 7046 9799 7098
rect 9799 7046 9809 7098
rect 9833 7046 9863 7098
rect 9863 7046 9875 7098
rect 9875 7046 9889 7098
rect 9913 7046 9927 7098
rect 9927 7046 9939 7098
rect 9939 7046 9969 7098
rect 9993 7046 10003 7098
rect 10003 7046 10049 7098
rect 9753 7044 9809 7046
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 9753 6010 9809 6012
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 9753 5958 9799 6010
rect 9799 5958 9809 6010
rect 9833 5958 9863 6010
rect 9863 5958 9875 6010
rect 9875 5958 9889 6010
rect 9913 5958 9927 6010
rect 9927 5958 9939 6010
rect 9939 5958 9969 6010
rect 9993 5958 10003 6010
rect 10003 5958 10049 6010
rect 9753 5956 9809 5958
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 9753 4922 9809 4924
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 9753 4870 9799 4922
rect 9799 4870 9809 4922
rect 9833 4870 9863 4922
rect 9863 4870 9875 4922
rect 9875 4870 9889 4922
rect 9913 4870 9927 4922
rect 9927 4870 9939 4922
rect 9939 4870 9969 4922
rect 9993 4870 10003 4922
rect 10003 4870 10049 4922
rect 9753 4868 9809 4870
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 9753 3834 9809 3836
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 9753 3782 9799 3834
rect 9799 3782 9809 3834
rect 9833 3782 9863 3834
rect 9863 3782 9875 3834
rect 9875 3782 9889 3834
rect 9913 3782 9927 3834
rect 9927 3782 9939 3834
rect 9939 3782 9969 3834
rect 9993 3782 10003 3834
rect 10003 3782 10049 3834
rect 9753 3780 9809 3782
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 12685 7642 12741 7644
rect 12765 7642 12821 7644
rect 12845 7642 12901 7644
rect 12925 7642 12981 7644
rect 12685 7590 12731 7642
rect 12731 7590 12741 7642
rect 12765 7590 12795 7642
rect 12795 7590 12807 7642
rect 12807 7590 12821 7642
rect 12845 7590 12859 7642
rect 12859 7590 12871 7642
rect 12871 7590 12901 7642
rect 12925 7590 12935 7642
rect 12935 7590 12981 7642
rect 12685 7588 12741 7590
rect 12765 7588 12821 7590
rect 12845 7588 12901 7590
rect 12925 7588 12981 7590
rect 12685 6554 12741 6556
rect 12765 6554 12821 6556
rect 12845 6554 12901 6556
rect 12925 6554 12981 6556
rect 12685 6502 12731 6554
rect 12731 6502 12741 6554
rect 12765 6502 12795 6554
rect 12795 6502 12807 6554
rect 12807 6502 12821 6554
rect 12845 6502 12859 6554
rect 12859 6502 12871 6554
rect 12871 6502 12901 6554
rect 12925 6502 12935 6554
rect 12935 6502 12981 6554
rect 12685 6500 12741 6502
rect 12765 6500 12821 6502
rect 12845 6500 12901 6502
rect 12925 6500 12981 6502
rect 12685 5466 12741 5468
rect 12765 5466 12821 5468
rect 12845 5466 12901 5468
rect 12925 5466 12981 5468
rect 12685 5414 12731 5466
rect 12731 5414 12741 5466
rect 12765 5414 12795 5466
rect 12795 5414 12807 5466
rect 12807 5414 12821 5466
rect 12845 5414 12859 5466
rect 12859 5414 12871 5466
rect 12871 5414 12901 5466
rect 12925 5414 12935 5466
rect 12935 5414 12981 5466
rect 12685 5412 12741 5414
rect 12765 5412 12821 5414
rect 12845 5412 12901 5414
rect 12925 5412 12981 5414
rect 12685 4378 12741 4380
rect 12765 4378 12821 4380
rect 12845 4378 12901 4380
rect 12925 4378 12981 4380
rect 12685 4326 12731 4378
rect 12731 4326 12741 4378
rect 12765 4326 12795 4378
rect 12795 4326 12807 4378
rect 12807 4326 12821 4378
rect 12845 4326 12859 4378
rect 12859 4326 12871 4378
rect 12871 4326 12901 4378
rect 12925 4326 12935 4378
rect 12935 4326 12981 4378
rect 12685 4324 12741 4326
rect 12765 4324 12821 4326
rect 12845 4324 12901 4326
rect 12925 4324 12981 4326
rect 15618 8186 15674 8188
rect 15698 8186 15754 8188
rect 15778 8186 15834 8188
rect 15858 8186 15914 8188
rect 15618 8134 15664 8186
rect 15664 8134 15674 8186
rect 15698 8134 15728 8186
rect 15728 8134 15740 8186
rect 15740 8134 15754 8186
rect 15778 8134 15792 8186
rect 15792 8134 15804 8186
rect 15804 8134 15834 8186
rect 15858 8134 15868 8186
rect 15868 8134 15914 8186
rect 15618 8132 15674 8134
rect 15698 8132 15754 8134
rect 15778 8132 15834 8134
rect 15858 8132 15914 8134
rect 15618 7098 15674 7100
rect 15698 7098 15754 7100
rect 15778 7098 15834 7100
rect 15858 7098 15914 7100
rect 15618 7046 15664 7098
rect 15664 7046 15674 7098
rect 15698 7046 15728 7098
rect 15728 7046 15740 7098
rect 15740 7046 15754 7098
rect 15778 7046 15792 7098
rect 15792 7046 15804 7098
rect 15804 7046 15834 7098
rect 15858 7046 15868 7098
rect 15868 7046 15914 7098
rect 15618 7044 15674 7046
rect 15698 7044 15754 7046
rect 15778 7044 15834 7046
rect 15858 7044 15914 7046
rect 15618 6010 15674 6012
rect 15698 6010 15754 6012
rect 15778 6010 15834 6012
rect 15858 6010 15914 6012
rect 15618 5958 15664 6010
rect 15664 5958 15674 6010
rect 15698 5958 15728 6010
rect 15728 5958 15740 6010
rect 15740 5958 15754 6010
rect 15778 5958 15792 6010
rect 15792 5958 15804 6010
rect 15804 5958 15834 6010
rect 15858 5958 15868 6010
rect 15868 5958 15914 6010
rect 15618 5956 15674 5958
rect 15698 5956 15754 5958
rect 15778 5956 15834 5958
rect 15858 5956 15914 5958
rect 15618 4922 15674 4924
rect 15698 4922 15754 4924
rect 15778 4922 15834 4924
rect 15858 4922 15914 4924
rect 15618 4870 15664 4922
rect 15664 4870 15674 4922
rect 15698 4870 15728 4922
rect 15728 4870 15740 4922
rect 15740 4870 15754 4922
rect 15778 4870 15792 4922
rect 15792 4870 15804 4922
rect 15804 4870 15834 4922
rect 15858 4870 15868 4922
rect 15868 4870 15914 4922
rect 15618 4868 15674 4870
rect 15698 4868 15754 4870
rect 15778 4868 15834 4870
rect 15858 4868 15914 4870
rect 15618 3834 15674 3836
rect 15698 3834 15754 3836
rect 15778 3834 15834 3836
rect 15858 3834 15914 3836
rect 15618 3782 15664 3834
rect 15664 3782 15674 3834
rect 15698 3782 15728 3834
rect 15728 3782 15740 3834
rect 15740 3782 15754 3834
rect 15778 3782 15792 3834
rect 15792 3782 15804 3834
rect 15804 3782 15834 3834
rect 15858 3782 15868 3834
rect 15868 3782 15914 3834
rect 15618 3780 15674 3782
rect 15698 3780 15754 3782
rect 15778 3780 15834 3782
rect 15858 3780 15914 3782
rect 7102 1672 7158 1728
rect 5630 448 5686 504
rect 6182 720 6238 776
rect 6090 176 6146 232
rect 6820 1114 6876 1116
rect 6900 1114 6956 1116
rect 6980 1114 7036 1116
rect 7060 1114 7116 1116
rect 6820 1062 6866 1114
rect 6866 1062 6876 1114
rect 6900 1062 6930 1114
rect 6930 1062 6942 1114
rect 6942 1062 6956 1114
rect 6980 1062 6994 1114
rect 6994 1062 7006 1114
rect 7006 1062 7036 1114
rect 7060 1062 7070 1114
rect 7070 1062 7116 1114
rect 6820 1060 6876 1062
rect 6900 1060 6956 1062
rect 6980 1060 7036 1062
rect 7060 1060 7116 1062
rect 8206 2216 8262 2272
rect 8114 1164 8116 1184
rect 8116 1164 8168 1184
rect 8168 1164 8170 1184
rect 8114 1128 8170 1164
rect 8298 1264 8354 1320
rect 9753 2746 9809 2748
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 9753 2694 9799 2746
rect 9799 2694 9809 2746
rect 9833 2694 9863 2746
rect 9863 2694 9875 2746
rect 9875 2694 9889 2746
rect 9913 2694 9927 2746
rect 9927 2694 9939 2746
rect 9939 2694 9969 2746
rect 9993 2694 10003 2746
rect 10003 2694 10049 2746
rect 9753 2692 9809 2694
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 12685 3290 12741 3292
rect 12765 3290 12821 3292
rect 12845 3290 12901 3292
rect 12925 3290 12981 3292
rect 12685 3238 12731 3290
rect 12731 3238 12741 3290
rect 12765 3238 12795 3290
rect 12795 3238 12807 3290
rect 12807 3238 12821 3290
rect 12845 3238 12859 3290
rect 12859 3238 12871 3290
rect 12871 3238 12901 3290
rect 12925 3238 12935 3290
rect 12935 3238 12981 3290
rect 12685 3236 12741 3238
rect 12765 3236 12821 3238
rect 12845 3236 12901 3238
rect 12925 3236 12981 3238
rect 12346 3032 12402 3088
rect 11978 2488 12034 2544
rect 9126 1536 9182 1592
rect 9586 2080 9642 2136
rect 10046 2216 10102 2272
rect 9753 1658 9809 1660
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 9753 1606 9799 1658
rect 9799 1606 9809 1658
rect 9833 1606 9863 1658
rect 9863 1606 9875 1658
rect 9875 1606 9889 1658
rect 9913 1606 9927 1658
rect 9927 1606 9939 1658
rect 9939 1606 9969 1658
rect 9993 1606 10003 1658
rect 10003 1606 10049 1658
rect 9753 1604 9809 1606
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 9678 1128 9734 1184
rect 11702 2080 11758 2136
rect 11334 1264 11390 1320
rect 12685 2202 12741 2204
rect 12765 2202 12821 2204
rect 12845 2202 12901 2204
rect 12925 2202 12981 2204
rect 12685 2150 12731 2202
rect 12731 2150 12741 2202
rect 12765 2150 12795 2202
rect 12795 2150 12807 2202
rect 12807 2150 12821 2202
rect 12845 2150 12859 2202
rect 12859 2150 12871 2202
rect 12871 2150 12901 2202
rect 12925 2150 12935 2202
rect 12935 2150 12981 2202
rect 12685 2148 12741 2150
rect 12765 2148 12821 2150
rect 12845 2148 12901 2150
rect 12925 2148 12981 2150
rect 12685 1114 12741 1116
rect 12765 1114 12821 1116
rect 12845 1114 12901 1116
rect 12925 1114 12981 1116
rect 12685 1062 12731 1114
rect 12731 1062 12741 1114
rect 12765 1062 12795 1114
rect 12795 1062 12807 1114
rect 12807 1062 12821 1114
rect 12845 1062 12859 1114
rect 12859 1062 12871 1114
rect 12871 1062 12901 1114
rect 12925 1062 12935 1114
rect 12935 1062 12981 1114
rect 12685 1060 12741 1062
rect 12765 1060 12821 1062
rect 12845 1060 12901 1062
rect 12925 1060 12981 1062
rect 13358 1400 13414 1456
rect 14278 2624 14334 2680
rect 15618 2746 15674 2748
rect 15698 2746 15754 2748
rect 15778 2746 15834 2748
rect 15858 2746 15914 2748
rect 15618 2694 15664 2746
rect 15664 2694 15674 2746
rect 15698 2694 15728 2746
rect 15728 2694 15740 2746
rect 15740 2694 15754 2746
rect 15778 2694 15792 2746
rect 15792 2694 15804 2746
rect 15804 2694 15834 2746
rect 15858 2694 15868 2746
rect 15868 2694 15914 2746
rect 15618 2692 15674 2694
rect 15698 2692 15754 2694
rect 15778 2692 15834 2694
rect 15858 2692 15914 2694
rect 14002 312 14058 368
rect 15618 1658 15674 1660
rect 15698 1658 15754 1660
rect 15778 1658 15834 1660
rect 15858 1658 15914 1660
rect 15618 1606 15664 1658
rect 15664 1606 15674 1658
rect 15698 1606 15728 1658
rect 15728 1606 15740 1658
rect 15740 1606 15754 1658
rect 15778 1606 15792 1658
rect 15792 1606 15804 1658
rect 15804 1606 15834 1658
rect 15858 1606 15868 1658
rect 15868 1606 15914 1658
rect 15618 1604 15674 1606
rect 15698 1604 15754 1606
rect 15778 1604 15834 1606
rect 15858 1604 15914 1606
rect 18550 7642 18606 7644
rect 18630 7642 18686 7644
rect 18710 7642 18766 7644
rect 18790 7642 18846 7644
rect 18550 7590 18596 7642
rect 18596 7590 18606 7642
rect 18630 7590 18660 7642
rect 18660 7590 18672 7642
rect 18672 7590 18686 7642
rect 18710 7590 18724 7642
rect 18724 7590 18736 7642
rect 18736 7590 18766 7642
rect 18790 7590 18800 7642
rect 18800 7590 18846 7642
rect 18550 7588 18606 7590
rect 18630 7588 18686 7590
rect 18710 7588 18766 7590
rect 18790 7588 18846 7590
rect 18550 6554 18606 6556
rect 18630 6554 18686 6556
rect 18710 6554 18766 6556
rect 18790 6554 18846 6556
rect 18550 6502 18596 6554
rect 18596 6502 18606 6554
rect 18630 6502 18660 6554
rect 18660 6502 18672 6554
rect 18672 6502 18686 6554
rect 18710 6502 18724 6554
rect 18724 6502 18736 6554
rect 18736 6502 18766 6554
rect 18790 6502 18800 6554
rect 18800 6502 18846 6554
rect 18550 6500 18606 6502
rect 18630 6500 18686 6502
rect 18710 6500 18766 6502
rect 18790 6500 18846 6502
rect 18550 5466 18606 5468
rect 18630 5466 18686 5468
rect 18710 5466 18766 5468
rect 18790 5466 18846 5468
rect 18550 5414 18596 5466
rect 18596 5414 18606 5466
rect 18630 5414 18660 5466
rect 18660 5414 18672 5466
rect 18672 5414 18686 5466
rect 18710 5414 18724 5466
rect 18724 5414 18736 5466
rect 18736 5414 18766 5466
rect 18790 5414 18800 5466
rect 18800 5414 18846 5466
rect 18550 5412 18606 5414
rect 18630 5412 18686 5414
rect 18710 5412 18766 5414
rect 18790 5412 18846 5414
rect 18550 4378 18606 4380
rect 18630 4378 18686 4380
rect 18710 4378 18766 4380
rect 18790 4378 18846 4380
rect 18550 4326 18596 4378
rect 18596 4326 18606 4378
rect 18630 4326 18660 4378
rect 18660 4326 18672 4378
rect 18672 4326 18686 4378
rect 18710 4326 18724 4378
rect 18724 4326 18736 4378
rect 18736 4326 18766 4378
rect 18790 4326 18800 4378
rect 18800 4326 18846 4378
rect 18550 4324 18606 4326
rect 18630 4324 18686 4326
rect 18710 4324 18766 4326
rect 18790 4324 18846 4326
rect 18550 3290 18606 3292
rect 18630 3290 18686 3292
rect 18710 3290 18766 3292
rect 18790 3290 18846 3292
rect 18550 3238 18596 3290
rect 18596 3238 18606 3290
rect 18630 3238 18660 3290
rect 18660 3238 18672 3290
rect 18672 3238 18686 3290
rect 18710 3238 18724 3290
rect 18724 3238 18736 3290
rect 18736 3238 18766 3290
rect 18790 3238 18800 3290
rect 18800 3238 18846 3290
rect 18550 3236 18606 3238
rect 18630 3236 18686 3238
rect 18710 3236 18766 3238
rect 18790 3236 18846 3238
rect 17958 2896 18014 2952
rect 16854 1400 16910 1456
rect 21483 8186 21539 8188
rect 21563 8186 21619 8188
rect 21643 8186 21699 8188
rect 21723 8186 21779 8188
rect 21483 8134 21529 8186
rect 21529 8134 21539 8186
rect 21563 8134 21593 8186
rect 21593 8134 21605 8186
rect 21605 8134 21619 8186
rect 21643 8134 21657 8186
rect 21657 8134 21669 8186
rect 21669 8134 21699 8186
rect 21723 8134 21733 8186
rect 21733 8134 21779 8186
rect 21483 8132 21539 8134
rect 21563 8132 21619 8134
rect 21643 8132 21699 8134
rect 21723 8132 21779 8134
rect 21483 7098 21539 7100
rect 21563 7098 21619 7100
rect 21643 7098 21699 7100
rect 21723 7098 21779 7100
rect 21483 7046 21529 7098
rect 21529 7046 21539 7098
rect 21563 7046 21593 7098
rect 21593 7046 21605 7098
rect 21605 7046 21619 7098
rect 21643 7046 21657 7098
rect 21657 7046 21669 7098
rect 21669 7046 21699 7098
rect 21723 7046 21733 7098
rect 21733 7046 21779 7098
rect 21483 7044 21539 7046
rect 21563 7044 21619 7046
rect 21643 7044 21699 7046
rect 21723 7044 21779 7046
rect 21483 6010 21539 6012
rect 21563 6010 21619 6012
rect 21643 6010 21699 6012
rect 21723 6010 21779 6012
rect 21483 5958 21529 6010
rect 21529 5958 21539 6010
rect 21563 5958 21593 6010
rect 21593 5958 21605 6010
rect 21605 5958 21619 6010
rect 21643 5958 21657 6010
rect 21657 5958 21669 6010
rect 21669 5958 21699 6010
rect 21723 5958 21733 6010
rect 21733 5958 21779 6010
rect 21483 5956 21539 5958
rect 21563 5956 21619 5958
rect 21643 5956 21699 5958
rect 21723 5956 21779 5958
rect 21483 4922 21539 4924
rect 21563 4922 21619 4924
rect 21643 4922 21699 4924
rect 21723 4922 21779 4924
rect 21483 4870 21529 4922
rect 21529 4870 21539 4922
rect 21563 4870 21593 4922
rect 21593 4870 21605 4922
rect 21605 4870 21619 4922
rect 21643 4870 21657 4922
rect 21657 4870 21669 4922
rect 21669 4870 21699 4922
rect 21723 4870 21733 4922
rect 21733 4870 21779 4922
rect 21483 4868 21539 4870
rect 21563 4868 21619 4870
rect 21643 4868 21699 4870
rect 21723 4868 21779 4870
rect 19798 4004 19854 4040
rect 19798 3984 19800 4004
rect 19800 3984 19852 4004
rect 19852 3984 19854 4004
rect 21483 3834 21539 3836
rect 21563 3834 21619 3836
rect 21643 3834 21699 3836
rect 21723 3834 21779 3836
rect 21483 3782 21529 3834
rect 21529 3782 21539 3834
rect 21563 3782 21593 3834
rect 21593 3782 21605 3834
rect 21605 3782 21619 3834
rect 21643 3782 21657 3834
rect 21657 3782 21669 3834
rect 21669 3782 21699 3834
rect 21723 3782 21733 3834
rect 21733 3782 21779 3834
rect 21483 3780 21539 3782
rect 21563 3780 21619 3782
rect 21643 3780 21699 3782
rect 21723 3780 21779 3782
rect 18550 2202 18606 2204
rect 18630 2202 18686 2204
rect 18710 2202 18766 2204
rect 18790 2202 18846 2204
rect 18550 2150 18596 2202
rect 18596 2150 18606 2202
rect 18630 2150 18660 2202
rect 18660 2150 18672 2202
rect 18672 2150 18686 2202
rect 18710 2150 18724 2202
rect 18724 2150 18736 2202
rect 18736 2150 18766 2202
rect 18790 2150 18800 2202
rect 18800 2150 18846 2202
rect 18550 2148 18606 2150
rect 18630 2148 18686 2150
rect 18710 2148 18766 2150
rect 18790 2148 18846 2150
rect 18550 1114 18606 1116
rect 18630 1114 18686 1116
rect 18710 1114 18766 1116
rect 18790 1114 18846 1116
rect 18550 1062 18596 1114
rect 18596 1062 18606 1114
rect 18630 1062 18660 1114
rect 18660 1062 18672 1114
rect 18672 1062 18686 1114
rect 18710 1062 18724 1114
rect 18724 1062 18736 1114
rect 18736 1062 18766 1114
rect 18790 1062 18800 1114
rect 18800 1062 18846 1114
rect 18550 1060 18606 1062
rect 18630 1060 18686 1062
rect 18710 1060 18766 1062
rect 18790 1060 18846 1062
rect 18418 720 18474 776
rect 19614 2372 19670 2408
rect 19614 2352 19616 2372
rect 19616 2352 19668 2372
rect 19668 2352 19670 2372
rect 19062 176 19118 232
rect 21483 2746 21539 2748
rect 21563 2746 21619 2748
rect 21643 2746 21699 2748
rect 21723 2746 21779 2748
rect 21483 2694 21529 2746
rect 21529 2694 21539 2746
rect 21563 2694 21593 2746
rect 21593 2694 21605 2746
rect 21605 2694 21619 2746
rect 21643 2694 21657 2746
rect 21657 2694 21669 2746
rect 21669 2694 21699 2746
rect 21723 2694 21733 2746
rect 21733 2694 21779 2746
rect 21483 2692 21539 2694
rect 21563 2692 21619 2694
rect 21643 2692 21699 2694
rect 21723 2692 21779 2694
rect 20074 584 20130 640
rect 21546 1944 21602 2000
rect 21178 1828 21234 1864
rect 21178 1808 21180 1828
rect 21180 1808 21232 1828
rect 21232 1808 21234 1828
rect 21483 1658 21539 1660
rect 21563 1658 21619 1660
rect 21643 1658 21699 1660
rect 21723 1658 21779 1660
rect 21483 1606 21529 1658
rect 21529 1606 21539 1658
rect 21563 1606 21593 1658
rect 21593 1606 21605 1658
rect 21605 1606 21619 1658
rect 21643 1606 21657 1658
rect 21657 1606 21669 1658
rect 21669 1606 21699 1658
rect 21723 1606 21733 1658
rect 21733 1606 21779 1658
rect 21483 1604 21539 1606
rect 21563 1604 21619 1606
rect 21643 1604 21699 1606
rect 21723 1604 21779 1606
rect 20718 720 20774 776
rect 21454 856 21510 912
rect 23018 2352 23074 2408
rect 22926 1672 22982 1728
rect 22926 312 22982 368
rect 23570 2216 23626 2272
rect 23570 1672 23626 1728
rect 24415 7642 24471 7644
rect 24495 7642 24551 7644
rect 24575 7642 24631 7644
rect 24655 7642 24711 7644
rect 24415 7590 24461 7642
rect 24461 7590 24471 7642
rect 24495 7590 24525 7642
rect 24525 7590 24537 7642
rect 24537 7590 24551 7642
rect 24575 7590 24589 7642
rect 24589 7590 24601 7642
rect 24601 7590 24631 7642
rect 24655 7590 24665 7642
rect 24665 7590 24711 7642
rect 24415 7588 24471 7590
rect 24495 7588 24551 7590
rect 24575 7588 24631 7590
rect 24655 7588 24711 7590
rect 24415 6554 24471 6556
rect 24495 6554 24551 6556
rect 24575 6554 24631 6556
rect 24655 6554 24711 6556
rect 24415 6502 24461 6554
rect 24461 6502 24471 6554
rect 24495 6502 24525 6554
rect 24525 6502 24537 6554
rect 24537 6502 24551 6554
rect 24575 6502 24589 6554
rect 24589 6502 24601 6554
rect 24601 6502 24631 6554
rect 24655 6502 24665 6554
rect 24665 6502 24711 6554
rect 24415 6500 24471 6502
rect 24495 6500 24551 6502
rect 24575 6500 24631 6502
rect 24655 6500 24711 6502
rect 24415 5466 24471 5468
rect 24495 5466 24551 5468
rect 24575 5466 24631 5468
rect 24655 5466 24711 5468
rect 24415 5414 24461 5466
rect 24461 5414 24471 5466
rect 24495 5414 24525 5466
rect 24525 5414 24537 5466
rect 24537 5414 24551 5466
rect 24575 5414 24589 5466
rect 24589 5414 24601 5466
rect 24601 5414 24631 5466
rect 24655 5414 24665 5466
rect 24665 5414 24711 5466
rect 24415 5412 24471 5414
rect 24495 5412 24551 5414
rect 24575 5412 24631 5414
rect 24655 5412 24711 5414
rect 24415 4378 24471 4380
rect 24495 4378 24551 4380
rect 24575 4378 24631 4380
rect 24655 4378 24711 4380
rect 24415 4326 24461 4378
rect 24461 4326 24471 4378
rect 24495 4326 24525 4378
rect 24525 4326 24537 4378
rect 24537 4326 24551 4378
rect 24575 4326 24589 4378
rect 24589 4326 24601 4378
rect 24601 4326 24631 4378
rect 24655 4326 24665 4378
rect 24665 4326 24711 4378
rect 24415 4324 24471 4326
rect 24495 4324 24551 4326
rect 24575 4324 24631 4326
rect 24655 4324 24711 4326
rect 24415 3290 24471 3292
rect 24495 3290 24551 3292
rect 24575 3290 24631 3292
rect 24655 3290 24711 3292
rect 24415 3238 24461 3290
rect 24461 3238 24471 3290
rect 24495 3238 24525 3290
rect 24525 3238 24537 3290
rect 24537 3238 24551 3290
rect 24575 3238 24589 3290
rect 24589 3238 24601 3290
rect 24601 3238 24631 3290
rect 24655 3238 24665 3290
rect 24665 3238 24711 3290
rect 24415 3236 24471 3238
rect 24495 3236 24551 3238
rect 24575 3236 24631 3238
rect 24655 3236 24711 3238
rect 24674 2352 24730 2408
rect 24415 2202 24471 2204
rect 24495 2202 24551 2204
rect 24575 2202 24631 2204
rect 24655 2202 24711 2204
rect 24415 2150 24461 2202
rect 24461 2150 24471 2202
rect 24495 2150 24525 2202
rect 24525 2150 24537 2202
rect 24537 2150 24551 2202
rect 24575 2150 24589 2202
rect 24589 2150 24601 2202
rect 24601 2150 24631 2202
rect 24655 2150 24665 2202
rect 24665 2150 24711 2202
rect 24415 2148 24471 2150
rect 24495 2148 24551 2150
rect 24575 2148 24631 2150
rect 24655 2148 24711 2150
rect 24415 1114 24471 1116
rect 24495 1114 24551 1116
rect 24575 1114 24631 1116
rect 24655 1114 24711 1116
rect 24415 1062 24461 1114
rect 24461 1062 24471 1114
rect 24495 1062 24525 1114
rect 24525 1062 24537 1114
rect 24537 1062 24551 1114
rect 24575 1062 24589 1114
rect 24589 1062 24601 1114
rect 24601 1062 24631 1114
rect 24655 1062 24665 1114
rect 24665 1062 24711 1114
rect 24415 1060 24471 1062
rect 24495 1060 24551 1062
rect 24575 1060 24631 1062
rect 24655 1060 24711 1062
<< metal3 >>
rect 6810 8736 7126 8737
rect 6810 8672 6816 8736
rect 6880 8672 6896 8736
rect 6960 8672 6976 8736
rect 7040 8672 7056 8736
rect 7120 8672 7126 8736
rect 6810 8671 7126 8672
rect 12675 8736 12991 8737
rect 12675 8672 12681 8736
rect 12745 8672 12761 8736
rect 12825 8672 12841 8736
rect 12905 8672 12921 8736
rect 12985 8672 12991 8736
rect 12675 8671 12991 8672
rect 18540 8736 18856 8737
rect 18540 8672 18546 8736
rect 18610 8672 18626 8736
rect 18690 8672 18706 8736
rect 18770 8672 18786 8736
rect 18850 8672 18856 8736
rect 18540 8671 18856 8672
rect 24405 8736 24721 8737
rect 24405 8672 24411 8736
rect 24475 8672 24491 8736
rect 24555 8672 24571 8736
rect 24635 8672 24651 8736
rect 24715 8672 24721 8736
rect 24405 8671 24721 8672
rect 3878 8192 4194 8193
rect 3878 8128 3884 8192
rect 3948 8128 3964 8192
rect 4028 8128 4044 8192
rect 4108 8128 4124 8192
rect 4188 8128 4194 8192
rect 3878 8127 4194 8128
rect 9743 8192 10059 8193
rect 9743 8128 9749 8192
rect 9813 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10059 8192
rect 9743 8127 10059 8128
rect 15608 8192 15924 8193
rect 15608 8128 15614 8192
rect 15678 8128 15694 8192
rect 15758 8128 15774 8192
rect 15838 8128 15854 8192
rect 15918 8128 15924 8192
rect 15608 8127 15924 8128
rect 21473 8192 21789 8193
rect 21473 8128 21479 8192
rect 21543 8128 21559 8192
rect 21623 8128 21639 8192
rect 21703 8128 21719 8192
rect 21783 8128 21789 8192
rect 21473 8127 21789 8128
rect 6810 7648 7126 7649
rect 6810 7584 6816 7648
rect 6880 7584 6896 7648
rect 6960 7584 6976 7648
rect 7040 7584 7056 7648
rect 7120 7584 7126 7648
rect 6810 7583 7126 7584
rect 12675 7648 12991 7649
rect 12675 7584 12681 7648
rect 12745 7584 12761 7648
rect 12825 7584 12841 7648
rect 12905 7584 12921 7648
rect 12985 7584 12991 7648
rect 12675 7583 12991 7584
rect 18540 7648 18856 7649
rect 18540 7584 18546 7648
rect 18610 7584 18626 7648
rect 18690 7584 18706 7648
rect 18770 7584 18786 7648
rect 18850 7584 18856 7648
rect 18540 7583 18856 7584
rect 24405 7648 24721 7649
rect 24405 7584 24411 7648
rect 24475 7584 24491 7648
rect 24555 7584 24571 7648
rect 24635 7584 24651 7648
rect 24715 7584 24721 7648
rect 24405 7583 24721 7584
rect 3878 7104 4194 7105
rect 3878 7040 3884 7104
rect 3948 7040 3964 7104
rect 4028 7040 4044 7104
rect 4108 7040 4124 7104
rect 4188 7040 4194 7104
rect 3878 7039 4194 7040
rect 9743 7104 10059 7105
rect 9743 7040 9749 7104
rect 9813 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10059 7104
rect 9743 7039 10059 7040
rect 15608 7104 15924 7105
rect 15608 7040 15614 7104
rect 15678 7040 15694 7104
rect 15758 7040 15774 7104
rect 15838 7040 15854 7104
rect 15918 7040 15924 7104
rect 15608 7039 15924 7040
rect 21473 7104 21789 7105
rect 21473 7040 21479 7104
rect 21543 7040 21559 7104
rect 21623 7040 21639 7104
rect 21703 7040 21719 7104
rect 21783 7040 21789 7104
rect 21473 7039 21789 7040
rect 6810 6560 7126 6561
rect 6810 6496 6816 6560
rect 6880 6496 6896 6560
rect 6960 6496 6976 6560
rect 7040 6496 7056 6560
rect 7120 6496 7126 6560
rect 6810 6495 7126 6496
rect 12675 6560 12991 6561
rect 12675 6496 12681 6560
rect 12745 6496 12761 6560
rect 12825 6496 12841 6560
rect 12905 6496 12921 6560
rect 12985 6496 12991 6560
rect 12675 6495 12991 6496
rect 18540 6560 18856 6561
rect 18540 6496 18546 6560
rect 18610 6496 18626 6560
rect 18690 6496 18706 6560
rect 18770 6496 18786 6560
rect 18850 6496 18856 6560
rect 18540 6495 18856 6496
rect 24405 6560 24721 6561
rect 24405 6496 24411 6560
rect 24475 6496 24491 6560
rect 24555 6496 24571 6560
rect 24635 6496 24651 6560
rect 24715 6496 24721 6560
rect 24405 6495 24721 6496
rect 3878 6016 4194 6017
rect 3878 5952 3884 6016
rect 3948 5952 3964 6016
rect 4028 5952 4044 6016
rect 4108 5952 4124 6016
rect 4188 5952 4194 6016
rect 3878 5951 4194 5952
rect 9743 6016 10059 6017
rect 9743 5952 9749 6016
rect 9813 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10059 6016
rect 9743 5951 10059 5952
rect 15608 6016 15924 6017
rect 15608 5952 15614 6016
rect 15678 5952 15694 6016
rect 15758 5952 15774 6016
rect 15838 5952 15854 6016
rect 15918 5952 15924 6016
rect 15608 5951 15924 5952
rect 21473 6016 21789 6017
rect 21473 5952 21479 6016
rect 21543 5952 21559 6016
rect 21623 5952 21639 6016
rect 21703 5952 21719 6016
rect 21783 5952 21789 6016
rect 21473 5951 21789 5952
rect 6810 5472 7126 5473
rect 6810 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6976 5472
rect 7040 5408 7056 5472
rect 7120 5408 7126 5472
rect 6810 5407 7126 5408
rect 12675 5472 12991 5473
rect 12675 5408 12681 5472
rect 12745 5408 12761 5472
rect 12825 5408 12841 5472
rect 12905 5408 12921 5472
rect 12985 5408 12991 5472
rect 12675 5407 12991 5408
rect 18540 5472 18856 5473
rect 18540 5408 18546 5472
rect 18610 5408 18626 5472
rect 18690 5408 18706 5472
rect 18770 5408 18786 5472
rect 18850 5408 18856 5472
rect 18540 5407 18856 5408
rect 24405 5472 24721 5473
rect 24405 5408 24411 5472
rect 24475 5408 24491 5472
rect 24555 5408 24571 5472
rect 24635 5408 24651 5472
rect 24715 5408 24721 5472
rect 24405 5407 24721 5408
rect 3878 4928 4194 4929
rect 3878 4864 3884 4928
rect 3948 4864 3964 4928
rect 4028 4864 4044 4928
rect 4108 4864 4124 4928
rect 4188 4864 4194 4928
rect 3878 4863 4194 4864
rect 9743 4928 10059 4929
rect 9743 4864 9749 4928
rect 9813 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10059 4928
rect 9743 4863 10059 4864
rect 15608 4928 15924 4929
rect 15608 4864 15614 4928
rect 15678 4864 15694 4928
rect 15758 4864 15774 4928
rect 15838 4864 15854 4928
rect 15918 4864 15924 4928
rect 15608 4863 15924 4864
rect 21473 4928 21789 4929
rect 21473 4864 21479 4928
rect 21543 4864 21559 4928
rect 21623 4864 21639 4928
rect 21703 4864 21719 4928
rect 21783 4864 21789 4928
rect 21473 4863 21789 4864
rect 6810 4384 7126 4385
rect 6810 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6976 4384
rect 7040 4320 7056 4384
rect 7120 4320 7126 4384
rect 6810 4319 7126 4320
rect 12675 4384 12991 4385
rect 12675 4320 12681 4384
rect 12745 4320 12761 4384
rect 12825 4320 12841 4384
rect 12905 4320 12921 4384
rect 12985 4320 12991 4384
rect 12675 4319 12991 4320
rect 18540 4384 18856 4385
rect 18540 4320 18546 4384
rect 18610 4320 18626 4384
rect 18690 4320 18706 4384
rect 18770 4320 18786 4384
rect 18850 4320 18856 4384
rect 18540 4319 18856 4320
rect 24405 4384 24721 4385
rect 24405 4320 24411 4384
rect 24475 4320 24491 4384
rect 24555 4320 24571 4384
rect 24635 4320 24651 4384
rect 24715 4320 24721 4384
rect 24405 4319 24721 4320
rect 2405 4042 2471 4045
rect 19793 4042 19859 4045
rect 2405 4040 19859 4042
rect 2405 3984 2410 4040
rect 2466 3984 19798 4040
rect 19854 3984 19859 4040
rect 2405 3982 19859 3984
rect 2405 3979 2471 3982
rect 19793 3979 19859 3982
rect 3878 3840 4194 3841
rect 3878 3776 3884 3840
rect 3948 3776 3964 3840
rect 4028 3776 4044 3840
rect 4108 3776 4124 3840
rect 4188 3776 4194 3840
rect 3878 3775 4194 3776
rect 9743 3840 10059 3841
rect 9743 3776 9749 3840
rect 9813 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10059 3840
rect 9743 3775 10059 3776
rect 15608 3840 15924 3841
rect 15608 3776 15614 3840
rect 15678 3776 15694 3840
rect 15758 3776 15774 3840
rect 15838 3776 15854 3840
rect 15918 3776 15924 3840
rect 15608 3775 15924 3776
rect 21473 3840 21789 3841
rect 21473 3776 21479 3840
rect 21543 3776 21559 3840
rect 21623 3776 21639 3840
rect 21703 3776 21719 3840
rect 21783 3776 21789 3840
rect 21473 3775 21789 3776
rect 6810 3296 7126 3297
rect 6810 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6976 3296
rect 7040 3232 7056 3296
rect 7120 3232 7126 3296
rect 6810 3231 7126 3232
rect 12675 3296 12991 3297
rect 12675 3232 12681 3296
rect 12745 3232 12761 3296
rect 12825 3232 12841 3296
rect 12905 3232 12921 3296
rect 12985 3232 12991 3296
rect 12675 3231 12991 3232
rect 18540 3296 18856 3297
rect 18540 3232 18546 3296
rect 18610 3232 18626 3296
rect 18690 3232 18706 3296
rect 18770 3232 18786 3296
rect 18850 3232 18856 3296
rect 18540 3231 18856 3232
rect 24405 3296 24721 3297
rect 24405 3232 24411 3296
rect 24475 3232 24491 3296
rect 24555 3232 24571 3296
rect 24635 3232 24651 3296
rect 24715 3232 24721 3296
rect 24405 3231 24721 3232
rect 4429 3090 4495 3093
rect 12341 3090 12407 3093
rect 4429 3088 12407 3090
rect 4429 3032 4434 3088
rect 4490 3032 12346 3088
rect 12402 3032 12407 3088
rect 4429 3030 12407 3032
rect 4429 3027 4495 3030
rect 12341 3027 12407 3030
rect 6821 2954 6887 2957
rect 17953 2954 18019 2957
rect 6821 2952 18019 2954
rect 6821 2896 6826 2952
rect 6882 2896 17958 2952
rect 18014 2896 18019 2952
rect 6821 2894 18019 2896
rect 6821 2891 6887 2894
rect 17953 2891 18019 2894
rect 3878 2752 4194 2753
rect 3878 2688 3884 2752
rect 3948 2688 3964 2752
rect 4028 2688 4044 2752
rect 4108 2688 4124 2752
rect 4188 2688 4194 2752
rect 3878 2687 4194 2688
rect 9743 2752 10059 2753
rect 9743 2688 9749 2752
rect 9813 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10059 2752
rect 9743 2687 10059 2688
rect 15608 2752 15924 2753
rect 15608 2688 15614 2752
rect 15678 2688 15694 2752
rect 15758 2688 15774 2752
rect 15838 2688 15854 2752
rect 15918 2688 15924 2752
rect 15608 2687 15924 2688
rect 21473 2752 21789 2753
rect 21473 2688 21479 2752
rect 21543 2688 21559 2752
rect 21623 2688 21639 2752
rect 21703 2688 21719 2752
rect 21783 2688 21789 2752
rect 21473 2687 21789 2688
rect 14273 2682 14339 2685
rect 11286 2680 14339 2682
rect 11286 2624 14278 2680
rect 14334 2624 14339 2680
rect 11286 2622 14339 2624
rect 6821 2546 6887 2549
rect 11286 2546 11346 2622
rect 14273 2619 14339 2622
rect 6821 2544 11346 2546
rect 6821 2488 6826 2544
rect 6882 2488 11346 2544
rect 6821 2486 11346 2488
rect 11973 2546 12039 2549
rect 11973 2544 22110 2546
rect 11973 2488 11978 2544
rect 12034 2488 22110 2544
rect 11973 2486 22110 2488
rect 6821 2483 6887 2486
rect 11973 2483 12039 2486
rect 1761 2410 1827 2413
rect 19609 2410 19675 2413
rect 1761 2408 19675 2410
rect 1761 2352 1766 2408
rect 1822 2352 19614 2408
rect 19670 2352 19675 2408
rect 1761 2350 19675 2352
rect 1761 2347 1827 2350
rect 19609 2347 19675 2350
rect 8201 2274 8267 2277
rect 10041 2274 10107 2277
rect 8201 2272 10107 2274
rect 8201 2216 8206 2272
rect 8262 2216 10046 2272
rect 10102 2216 10107 2272
rect 8201 2214 10107 2216
rect 22050 2274 22110 2486
rect 23013 2410 23079 2413
rect 24669 2410 24735 2413
rect 23013 2408 24735 2410
rect 23013 2352 23018 2408
rect 23074 2352 24674 2408
rect 24730 2352 24735 2408
rect 23013 2350 24735 2352
rect 23013 2347 23079 2350
rect 24669 2347 24735 2350
rect 23565 2274 23631 2277
rect 22050 2272 23631 2274
rect 22050 2216 23570 2272
rect 23626 2216 23631 2272
rect 22050 2214 23631 2216
rect 8201 2211 8267 2214
rect 10041 2211 10107 2214
rect 23565 2211 23631 2214
rect 6810 2208 7126 2209
rect 6810 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6976 2208
rect 7040 2144 7056 2208
rect 7120 2144 7126 2208
rect 6810 2143 7126 2144
rect 12675 2208 12991 2209
rect 12675 2144 12681 2208
rect 12745 2144 12761 2208
rect 12825 2144 12841 2208
rect 12905 2144 12921 2208
rect 12985 2144 12991 2208
rect 12675 2143 12991 2144
rect 18540 2208 18856 2209
rect 18540 2144 18546 2208
rect 18610 2144 18626 2208
rect 18690 2144 18706 2208
rect 18770 2144 18786 2208
rect 18850 2144 18856 2208
rect 18540 2143 18856 2144
rect 24405 2208 24721 2209
rect 24405 2144 24411 2208
rect 24475 2144 24491 2208
rect 24555 2144 24571 2208
rect 24635 2144 24651 2208
rect 24715 2144 24721 2208
rect 24405 2143 24721 2144
rect 9581 2138 9647 2141
rect 11697 2138 11763 2141
rect 9581 2136 11763 2138
rect 9581 2080 9586 2136
rect 9642 2080 11702 2136
rect 11758 2080 11763 2136
rect 9581 2078 11763 2080
rect 9581 2075 9647 2078
rect 11697 2075 11763 2078
rect 4797 2002 4863 2005
rect 21541 2002 21607 2005
rect 4797 2000 21607 2002
rect 4797 1944 4802 2000
rect 4858 1944 21546 2000
rect 21602 1944 21607 2000
rect 4797 1942 21607 1944
rect 4797 1939 4863 1942
rect 21541 1939 21607 1942
rect 3601 1866 3667 1869
rect 21173 1866 21239 1869
rect 3601 1864 21239 1866
rect 3601 1808 3606 1864
rect 3662 1808 21178 1864
rect 21234 1808 21239 1864
rect 3601 1806 21239 1808
rect 3601 1803 3667 1806
rect 21173 1803 21239 1806
rect 5993 1730 6059 1733
rect 7097 1730 7163 1733
rect 13670 1730 13676 1732
rect 5993 1728 7163 1730
rect 5993 1672 5998 1728
rect 6054 1672 7102 1728
rect 7158 1672 7163 1728
rect 5993 1670 7163 1672
rect 5993 1667 6059 1670
rect 7097 1667 7163 1670
rect 12390 1670 13676 1730
rect 3878 1664 4194 1665
rect 3878 1600 3884 1664
rect 3948 1600 3964 1664
rect 4028 1600 4044 1664
rect 4108 1600 4124 1664
rect 4188 1600 4194 1664
rect 3878 1599 4194 1600
rect 9743 1664 10059 1665
rect 9743 1600 9749 1664
rect 9813 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10059 1664
rect 9743 1599 10059 1600
rect 4337 1594 4403 1597
rect 9121 1594 9187 1597
rect 4337 1592 9187 1594
rect 4337 1536 4342 1592
rect 4398 1536 9126 1592
rect 9182 1536 9187 1592
rect 4337 1534 9187 1536
rect 4337 1531 4403 1534
rect 9121 1531 9187 1534
rect 4889 1458 4955 1461
rect 12390 1458 12450 1670
rect 13670 1668 13676 1670
rect 13740 1668 13746 1732
rect 22921 1730 22987 1733
rect 23565 1730 23631 1733
rect 22921 1728 23631 1730
rect 22921 1672 22926 1728
rect 22982 1672 23570 1728
rect 23626 1672 23631 1728
rect 22921 1670 23631 1672
rect 22921 1667 22987 1670
rect 23565 1667 23631 1670
rect 15608 1664 15924 1665
rect 15608 1600 15614 1664
rect 15678 1600 15694 1664
rect 15758 1600 15774 1664
rect 15838 1600 15854 1664
rect 15918 1600 15924 1664
rect 15608 1599 15924 1600
rect 21473 1664 21789 1665
rect 21473 1600 21479 1664
rect 21543 1600 21559 1664
rect 21623 1600 21639 1664
rect 21703 1600 21719 1664
rect 21783 1600 21789 1664
rect 21473 1599 21789 1600
rect 4889 1456 12450 1458
rect 4889 1400 4894 1456
rect 4950 1400 12450 1456
rect 4889 1398 12450 1400
rect 13353 1458 13419 1461
rect 16849 1458 16915 1461
rect 13353 1456 16915 1458
rect 13353 1400 13358 1456
rect 13414 1400 16854 1456
rect 16910 1400 16915 1456
rect 13353 1398 16915 1400
rect 4889 1395 4955 1398
rect 13353 1395 13419 1398
rect 16849 1395 16915 1398
rect 8293 1322 8359 1325
rect 11329 1322 11395 1325
rect 8293 1320 11395 1322
rect 8293 1264 8298 1320
rect 8354 1264 11334 1320
rect 11390 1264 11395 1320
rect 8293 1262 11395 1264
rect 8293 1259 8359 1262
rect 11329 1259 11395 1262
rect 8109 1186 8175 1189
rect 9673 1186 9739 1189
rect 8109 1184 9739 1186
rect 8109 1128 8114 1184
rect 8170 1128 9678 1184
rect 9734 1128 9739 1184
rect 8109 1126 9739 1128
rect 8109 1123 8175 1126
rect 9673 1123 9739 1126
rect 6810 1120 7126 1121
rect 6810 1056 6816 1120
rect 6880 1056 6896 1120
rect 6960 1056 6976 1120
rect 7040 1056 7056 1120
rect 7120 1056 7126 1120
rect 6810 1055 7126 1056
rect 12675 1120 12991 1121
rect 12675 1056 12681 1120
rect 12745 1056 12761 1120
rect 12825 1056 12841 1120
rect 12905 1056 12921 1120
rect 12985 1056 12991 1120
rect 12675 1055 12991 1056
rect 18540 1120 18856 1121
rect 18540 1056 18546 1120
rect 18610 1056 18626 1120
rect 18690 1056 18706 1120
rect 18770 1056 18786 1120
rect 18850 1056 18856 1120
rect 18540 1055 18856 1056
rect 24405 1120 24721 1121
rect 24405 1056 24411 1120
rect 24475 1056 24491 1120
rect 24555 1056 24571 1120
rect 24635 1056 24651 1120
rect 24715 1056 24721 1120
rect 24405 1055 24721 1056
rect 5349 914 5415 917
rect 21449 914 21515 917
rect 5349 912 21515 914
rect 5349 856 5354 912
rect 5410 856 21454 912
rect 21510 856 21515 912
rect 5349 854 21515 856
rect 5349 851 5415 854
rect 21449 851 21515 854
rect 6177 778 6243 781
rect 18413 778 18479 781
rect 20713 778 20779 781
rect 6177 776 18479 778
rect 6177 720 6182 776
rect 6238 720 18418 776
rect 18474 720 18479 776
rect 6177 718 18479 720
rect 6177 715 6243 718
rect 18413 715 18479 718
rect 18646 776 20779 778
rect 18646 720 20718 776
rect 20774 720 20779 776
rect 18646 718 20779 720
rect 4797 642 4863 645
rect 18646 642 18706 718
rect 20713 715 20779 718
rect 20069 642 20135 645
rect 4797 640 18706 642
rect 4797 584 4802 640
rect 4858 584 18706 640
rect 4797 582 18706 584
rect 18830 640 20135 642
rect 18830 584 20074 640
rect 20130 584 20135 640
rect 18830 582 20135 584
rect 4797 579 4863 582
rect 5625 506 5691 509
rect 18830 506 18890 582
rect 20069 579 20135 582
rect 5625 504 18890 506
rect 5625 448 5630 504
rect 5686 448 18890 504
rect 5625 446 18890 448
rect 5625 443 5691 446
rect 1669 370 1735 373
rect 13997 370 14063 373
rect 22921 370 22987 373
rect 1669 368 14063 370
rect 1669 312 1674 368
rect 1730 312 14002 368
rect 14058 312 14063 368
rect 1669 310 14063 312
rect 1669 307 1735 310
rect 13997 307 14063 310
rect 22050 368 22987 370
rect 22050 312 22926 368
rect 22982 312 22987 368
rect 22050 310 22987 312
rect 6085 234 6151 237
rect 19057 234 19123 237
rect 6085 232 19123 234
rect 6085 176 6090 232
rect 6146 176 19062 232
rect 19118 176 19123 232
rect 6085 174 19123 176
rect 6085 171 6151 174
rect 19057 171 19123 174
rect 13670 36 13676 100
rect 13740 98 13746 100
rect 22050 98 22110 310
rect 22921 307 22987 310
rect 13740 38 22110 98
rect 13740 36 13746 38
<< via3 >>
rect 6816 8732 6880 8736
rect 6816 8676 6820 8732
rect 6820 8676 6876 8732
rect 6876 8676 6880 8732
rect 6816 8672 6880 8676
rect 6896 8732 6960 8736
rect 6896 8676 6900 8732
rect 6900 8676 6956 8732
rect 6956 8676 6960 8732
rect 6896 8672 6960 8676
rect 6976 8732 7040 8736
rect 6976 8676 6980 8732
rect 6980 8676 7036 8732
rect 7036 8676 7040 8732
rect 6976 8672 7040 8676
rect 7056 8732 7120 8736
rect 7056 8676 7060 8732
rect 7060 8676 7116 8732
rect 7116 8676 7120 8732
rect 7056 8672 7120 8676
rect 12681 8732 12745 8736
rect 12681 8676 12685 8732
rect 12685 8676 12741 8732
rect 12741 8676 12745 8732
rect 12681 8672 12745 8676
rect 12761 8732 12825 8736
rect 12761 8676 12765 8732
rect 12765 8676 12821 8732
rect 12821 8676 12825 8732
rect 12761 8672 12825 8676
rect 12841 8732 12905 8736
rect 12841 8676 12845 8732
rect 12845 8676 12901 8732
rect 12901 8676 12905 8732
rect 12841 8672 12905 8676
rect 12921 8732 12985 8736
rect 12921 8676 12925 8732
rect 12925 8676 12981 8732
rect 12981 8676 12985 8732
rect 12921 8672 12985 8676
rect 18546 8732 18610 8736
rect 18546 8676 18550 8732
rect 18550 8676 18606 8732
rect 18606 8676 18610 8732
rect 18546 8672 18610 8676
rect 18626 8732 18690 8736
rect 18626 8676 18630 8732
rect 18630 8676 18686 8732
rect 18686 8676 18690 8732
rect 18626 8672 18690 8676
rect 18706 8732 18770 8736
rect 18706 8676 18710 8732
rect 18710 8676 18766 8732
rect 18766 8676 18770 8732
rect 18706 8672 18770 8676
rect 18786 8732 18850 8736
rect 18786 8676 18790 8732
rect 18790 8676 18846 8732
rect 18846 8676 18850 8732
rect 18786 8672 18850 8676
rect 24411 8732 24475 8736
rect 24411 8676 24415 8732
rect 24415 8676 24471 8732
rect 24471 8676 24475 8732
rect 24411 8672 24475 8676
rect 24491 8732 24555 8736
rect 24491 8676 24495 8732
rect 24495 8676 24551 8732
rect 24551 8676 24555 8732
rect 24491 8672 24555 8676
rect 24571 8732 24635 8736
rect 24571 8676 24575 8732
rect 24575 8676 24631 8732
rect 24631 8676 24635 8732
rect 24571 8672 24635 8676
rect 24651 8732 24715 8736
rect 24651 8676 24655 8732
rect 24655 8676 24711 8732
rect 24711 8676 24715 8732
rect 24651 8672 24715 8676
rect 3884 8188 3948 8192
rect 3884 8132 3888 8188
rect 3888 8132 3944 8188
rect 3944 8132 3948 8188
rect 3884 8128 3948 8132
rect 3964 8188 4028 8192
rect 3964 8132 3968 8188
rect 3968 8132 4024 8188
rect 4024 8132 4028 8188
rect 3964 8128 4028 8132
rect 4044 8188 4108 8192
rect 4044 8132 4048 8188
rect 4048 8132 4104 8188
rect 4104 8132 4108 8188
rect 4044 8128 4108 8132
rect 4124 8188 4188 8192
rect 4124 8132 4128 8188
rect 4128 8132 4184 8188
rect 4184 8132 4188 8188
rect 4124 8128 4188 8132
rect 9749 8188 9813 8192
rect 9749 8132 9753 8188
rect 9753 8132 9809 8188
rect 9809 8132 9813 8188
rect 9749 8128 9813 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 15614 8188 15678 8192
rect 15614 8132 15618 8188
rect 15618 8132 15674 8188
rect 15674 8132 15678 8188
rect 15614 8128 15678 8132
rect 15694 8188 15758 8192
rect 15694 8132 15698 8188
rect 15698 8132 15754 8188
rect 15754 8132 15758 8188
rect 15694 8128 15758 8132
rect 15774 8188 15838 8192
rect 15774 8132 15778 8188
rect 15778 8132 15834 8188
rect 15834 8132 15838 8188
rect 15774 8128 15838 8132
rect 15854 8188 15918 8192
rect 15854 8132 15858 8188
rect 15858 8132 15914 8188
rect 15914 8132 15918 8188
rect 15854 8128 15918 8132
rect 21479 8188 21543 8192
rect 21479 8132 21483 8188
rect 21483 8132 21539 8188
rect 21539 8132 21543 8188
rect 21479 8128 21543 8132
rect 21559 8188 21623 8192
rect 21559 8132 21563 8188
rect 21563 8132 21619 8188
rect 21619 8132 21623 8188
rect 21559 8128 21623 8132
rect 21639 8188 21703 8192
rect 21639 8132 21643 8188
rect 21643 8132 21699 8188
rect 21699 8132 21703 8188
rect 21639 8128 21703 8132
rect 21719 8188 21783 8192
rect 21719 8132 21723 8188
rect 21723 8132 21779 8188
rect 21779 8132 21783 8188
rect 21719 8128 21783 8132
rect 6816 7644 6880 7648
rect 6816 7588 6820 7644
rect 6820 7588 6876 7644
rect 6876 7588 6880 7644
rect 6816 7584 6880 7588
rect 6896 7644 6960 7648
rect 6896 7588 6900 7644
rect 6900 7588 6956 7644
rect 6956 7588 6960 7644
rect 6896 7584 6960 7588
rect 6976 7644 7040 7648
rect 6976 7588 6980 7644
rect 6980 7588 7036 7644
rect 7036 7588 7040 7644
rect 6976 7584 7040 7588
rect 7056 7644 7120 7648
rect 7056 7588 7060 7644
rect 7060 7588 7116 7644
rect 7116 7588 7120 7644
rect 7056 7584 7120 7588
rect 12681 7644 12745 7648
rect 12681 7588 12685 7644
rect 12685 7588 12741 7644
rect 12741 7588 12745 7644
rect 12681 7584 12745 7588
rect 12761 7644 12825 7648
rect 12761 7588 12765 7644
rect 12765 7588 12821 7644
rect 12821 7588 12825 7644
rect 12761 7584 12825 7588
rect 12841 7644 12905 7648
rect 12841 7588 12845 7644
rect 12845 7588 12901 7644
rect 12901 7588 12905 7644
rect 12841 7584 12905 7588
rect 12921 7644 12985 7648
rect 12921 7588 12925 7644
rect 12925 7588 12981 7644
rect 12981 7588 12985 7644
rect 12921 7584 12985 7588
rect 18546 7644 18610 7648
rect 18546 7588 18550 7644
rect 18550 7588 18606 7644
rect 18606 7588 18610 7644
rect 18546 7584 18610 7588
rect 18626 7644 18690 7648
rect 18626 7588 18630 7644
rect 18630 7588 18686 7644
rect 18686 7588 18690 7644
rect 18626 7584 18690 7588
rect 18706 7644 18770 7648
rect 18706 7588 18710 7644
rect 18710 7588 18766 7644
rect 18766 7588 18770 7644
rect 18706 7584 18770 7588
rect 18786 7644 18850 7648
rect 18786 7588 18790 7644
rect 18790 7588 18846 7644
rect 18846 7588 18850 7644
rect 18786 7584 18850 7588
rect 24411 7644 24475 7648
rect 24411 7588 24415 7644
rect 24415 7588 24471 7644
rect 24471 7588 24475 7644
rect 24411 7584 24475 7588
rect 24491 7644 24555 7648
rect 24491 7588 24495 7644
rect 24495 7588 24551 7644
rect 24551 7588 24555 7644
rect 24491 7584 24555 7588
rect 24571 7644 24635 7648
rect 24571 7588 24575 7644
rect 24575 7588 24631 7644
rect 24631 7588 24635 7644
rect 24571 7584 24635 7588
rect 24651 7644 24715 7648
rect 24651 7588 24655 7644
rect 24655 7588 24711 7644
rect 24711 7588 24715 7644
rect 24651 7584 24715 7588
rect 3884 7100 3948 7104
rect 3884 7044 3888 7100
rect 3888 7044 3944 7100
rect 3944 7044 3948 7100
rect 3884 7040 3948 7044
rect 3964 7100 4028 7104
rect 3964 7044 3968 7100
rect 3968 7044 4024 7100
rect 4024 7044 4028 7100
rect 3964 7040 4028 7044
rect 4044 7100 4108 7104
rect 4044 7044 4048 7100
rect 4048 7044 4104 7100
rect 4104 7044 4108 7100
rect 4044 7040 4108 7044
rect 4124 7100 4188 7104
rect 4124 7044 4128 7100
rect 4128 7044 4184 7100
rect 4184 7044 4188 7100
rect 4124 7040 4188 7044
rect 9749 7100 9813 7104
rect 9749 7044 9753 7100
rect 9753 7044 9809 7100
rect 9809 7044 9813 7100
rect 9749 7040 9813 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 15614 7100 15678 7104
rect 15614 7044 15618 7100
rect 15618 7044 15674 7100
rect 15674 7044 15678 7100
rect 15614 7040 15678 7044
rect 15694 7100 15758 7104
rect 15694 7044 15698 7100
rect 15698 7044 15754 7100
rect 15754 7044 15758 7100
rect 15694 7040 15758 7044
rect 15774 7100 15838 7104
rect 15774 7044 15778 7100
rect 15778 7044 15834 7100
rect 15834 7044 15838 7100
rect 15774 7040 15838 7044
rect 15854 7100 15918 7104
rect 15854 7044 15858 7100
rect 15858 7044 15914 7100
rect 15914 7044 15918 7100
rect 15854 7040 15918 7044
rect 21479 7100 21543 7104
rect 21479 7044 21483 7100
rect 21483 7044 21539 7100
rect 21539 7044 21543 7100
rect 21479 7040 21543 7044
rect 21559 7100 21623 7104
rect 21559 7044 21563 7100
rect 21563 7044 21619 7100
rect 21619 7044 21623 7100
rect 21559 7040 21623 7044
rect 21639 7100 21703 7104
rect 21639 7044 21643 7100
rect 21643 7044 21699 7100
rect 21699 7044 21703 7100
rect 21639 7040 21703 7044
rect 21719 7100 21783 7104
rect 21719 7044 21723 7100
rect 21723 7044 21779 7100
rect 21779 7044 21783 7100
rect 21719 7040 21783 7044
rect 6816 6556 6880 6560
rect 6816 6500 6820 6556
rect 6820 6500 6876 6556
rect 6876 6500 6880 6556
rect 6816 6496 6880 6500
rect 6896 6556 6960 6560
rect 6896 6500 6900 6556
rect 6900 6500 6956 6556
rect 6956 6500 6960 6556
rect 6896 6496 6960 6500
rect 6976 6556 7040 6560
rect 6976 6500 6980 6556
rect 6980 6500 7036 6556
rect 7036 6500 7040 6556
rect 6976 6496 7040 6500
rect 7056 6556 7120 6560
rect 7056 6500 7060 6556
rect 7060 6500 7116 6556
rect 7116 6500 7120 6556
rect 7056 6496 7120 6500
rect 12681 6556 12745 6560
rect 12681 6500 12685 6556
rect 12685 6500 12741 6556
rect 12741 6500 12745 6556
rect 12681 6496 12745 6500
rect 12761 6556 12825 6560
rect 12761 6500 12765 6556
rect 12765 6500 12821 6556
rect 12821 6500 12825 6556
rect 12761 6496 12825 6500
rect 12841 6556 12905 6560
rect 12841 6500 12845 6556
rect 12845 6500 12901 6556
rect 12901 6500 12905 6556
rect 12841 6496 12905 6500
rect 12921 6556 12985 6560
rect 12921 6500 12925 6556
rect 12925 6500 12981 6556
rect 12981 6500 12985 6556
rect 12921 6496 12985 6500
rect 18546 6556 18610 6560
rect 18546 6500 18550 6556
rect 18550 6500 18606 6556
rect 18606 6500 18610 6556
rect 18546 6496 18610 6500
rect 18626 6556 18690 6560
rect 18626 6500 18630 6556
rect 18630 6500 18686 6556
rect 18686 6500 18690 6556
rect 18626 6496 18690 6500
rect 18706 6556 18770 6560
rect 18706 6500 18710 6556
rect 18710 6500 18766 6556
rect 18766 6500 18770 6556
rect 18706 6496 18770 6500
rect 18786 6556 18850 6560
rect 18786 6500 18790 6556
rect 18790 6500 18846 6556
rect 18846 6500 18850 6556
rect 18786 6496 18850 6500
rect 24411 6556 24475 6560
rect 24411 6500 24415 6556
rect 24415 6500 24471 6556
rect 24471 6500 24475 6556
rect 24411 6496 24475 6500
rect 24491 6556 24555 6560
rect 24491 6500 24495 6556
rect 24495 6500 24551 6556
rect 24551 6500 24555 6556
rect 24491 6496 24555 6500
rect 24571 6556 24635 6560
rect 24571 6500 24575 6556
rect 24575 6500 24631 6556
rect 24631 6500 24635 6556
rect 24571 6496 24635 6500
rect 24651 6556 24715 6560
rect 24651 6500 24655 6556
rect 24655 6500 24711 6556
rect 24711 6500 24715 6556
rect 24651 6496 24715 6500
rect 3884 6012 3948 6016
rect 3884 5956 3888 6012
rect 3888 5956 3944 6012
rect 3944 5956 3948 6012
rect 3884 5952 3948 5956
rect 3964 6012 4028 6016
rect 3964 5956 3968 6012
rect 3968 5956 4024 6012
rect 4024 5956 4028 6012
rect 3964 5952 4028 5956
rect 4044 6012 4108 6016
rect 4044 5956 4048 6012
rect 4048 5956 4104 6012
rect 4104 5956 4108 6012
rect 4044 5952 4108 5956
rect 4124 6012 4188 6016
rect 4124 5956 4128 6012
rect 4128 5956 4184 6012
rect 4184 5956 4188 6012
rect 4124 5952 4188 5956
rect 9749 6012 9813 6016
rect 9749 5956 9753 6012
rect 9753 5956 9809 6012
rect 9809 5956 9813 6012
rect 9749 5952 9813 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 15614 6012 15678 6016
rect 15614 5956 15618 6012
rect 15618 5956 15674 6012
rect 15674 5956 15678 6012
rect 15614 5952 15678 5956
rect 15694 6012 15758 6016
rect 15694 5956 15698 6012
rect 15698 5956 15754 6012
rect 15754 5956 15758 6012
rect 15694 5952 15758 5956
rect 15774 6012 15838 6016
rect 15774 5956 15778 6012
rect 15778 5956 15834 6012
rect 15834 5956 15838 6012
rect 15774 5952 15838 5956
rect 15854 6012 15918 6016
rect 15854 5956 15858 6012
rect 15858 5956 15914 6012
rect 15914 5956 15918 6012
rect 15854 5952 15918 5956
rect 21479 6012 21543 6016
rect 21479 5956 21483 6012
rect 21483 5956 21539 6012
rect 21539 5956 21543 6012
rect 21479 5952 21543 5956
rect 21559 6012 21623 6016
rect 21559 5956 21563 6012
rect 21563 5956 21619 6012
rect 21619 5956 21623 6012
rect 21559 5952 21623 5956
rect 21639 6012 21703 6016
rect 21639 5956 21643 6012
rect 21643 5956 21699 6012
rect 21699 5956 21703 6012
rect 21639 5952 21703 5956
rect 21719 6012 21783 6016
rect 21719 5956 21723 6012
rect 21723 5956 21779 6012
rect 21779 5956 21783 6012
rect 21719 5952 21783 5956
rect 6816 5468 6880 5472
rect 6816 5412 6820 5468
rect 6820 5412 6876 5468
rect 6876 5412 6880 5468
rect 6816 5408 6880 5412
rect 6896 5468 6960 5472
rect 6896 5412 6900 5468
rect 6900 5412 6956 5468
rect 6956 5412 6960 5468
rect 6896 5408 6960 5412
rect 6976 5468 7040 5472
rect 6976 5412 6980 5468
rect 6980 5412 7036 5468
rect 7036 5412 7040 5468
rect 6976 5408 7040 5412
rect 7056 5468 7120 5472
rect 7056 5412 7060 5468
rect 7060 5412 7116 5468
rect 7116 5412 7120 5468
rect 7056 5408 7120 5412
rect 12681 5468 12745 5472
rect 12681 5412 12685 5468
rect 12685 5412 12741 5468
rect 12741 5412 12745 5468
rect 12681 5408 12745 5412
rect 12761 5468 12825 5472
rect 12761 5412 12765 5468
rect 12765 5412 12821 5468
rect 12821 5412 12825 5468
rect 12761 5408 12825 5412
rect 12841 5468 12905 5472
rect 12841 5412 12845 5468
rect 12845 5412 12901 5468
rect 12901 5412 12905 5468
rect 12841 5408 12905 5412
rect 12921 5468 12985 5472
rect 12921 5412 12925 5468
rect 12925 5412 12981 5468
rect 12981 5412 12985 5468
rect 12921 5408 12985 5412
rect 18546 5468 18610 5472
rect 18546 5412 18550 5468
rect 18550 5412 18606 5468
rect 18606 5412 18610 5468
rect 18546 5408 18610 5412
rect 18626 5468 18690 5472
rect 18626 5412 18630 5468
rect 18630 5412 18686 5468
rect 18686 5412 18690 5468
rect 18626 5408 18690 5412
rect 18706 5468 18770 5472
rect 18706 5412 18710 5468
rect 18710 5412 18766 5468
rect 18766 5412 18770 5468
rect 18706 5408 18770 5412
rect 18786 5468 18850 5472
rect 18786 5412 18790 5468
rect 18790 5412 18846 5468
rect 18846 5412 18850 5468
rect 18786 5408 18850 5412
rect 24411 5468 24475 5472
rect 24411 5412 24415 5468
rect 24415 5412 24471 5468
rect 24471 5412 24475 5468
rect 24411 5408 24475 5412
rect 24491 5468 24555 5472
rect 24491 5412 24495 5468
rect 24495 5412 24551 5468
rect 24551 5412 24555 5468
rect 24491 5408 24555 5412
rect 24571 5468 24635 5472
rect 24571 5412 24575 5468
rect 24575 5412 24631 5468
rect 24631 5412 24635 5468
rect 24571 5408 24635 5412
rect 24651 5468 24715 5472
rect 24651 5412 24655 5468
rect 24655 5412 24711 5468
rect 24711 5412 24715 5468
rect 24651 5408 24715 5412
rect 3884 4924 3948 4928
rect 3884 4868 3888 4924
rect 3888 4868 3944 4924
rect 3944 4868 3948 4924
rect 3884 4864 3948 4868
rect 3964 4924 4028 4928
rect 3964 4868 3968 4924
rect 3968 4868 4024 4924
rect 4024 4868 4028 4924
rect 3964 4864 4028 4868
rect 4044 4924 4108 4928
rect 4044 4868 4048 4924
rect 4048 4868 4104 4924
rect 4104 4868 4108 4924
rect 4044 4864 4108 4868
rect 4124 4924 4188 4928
rect 4124 4868 4128 4924
rect 4128 4868 4184 4924
rect 4184 4868 4188 4924
rect 4124 4864 4188 4868
rect 9749 4924 9813 4928
rect 9749 4868 9753 4924
rect 9753 4868 9809 4924
rect 9809 4868 9813 4924
rect 9749 4864 9813 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 15614 4924 15678 4928
rect 15614 4868 15618 4924
rect 15618 4868 15674 4924
rect 15674 4868 15678 4924
rect 15614 4864 15678 4868
rect 15694 4924 15758 4928
rect 15694 4868 15698 4924
rect 15698 4868 15754 4924
rect 15754 4868 15758 4924
rect 15694 4864 15758 4868
rect 15774 4924 15838 4928
rect 15774 4868 15778 4924
rect 15778 4868 15834 4924
rect 15834 4868 15838 4924
rect 15774 4864 15838 4868
rect 15854 4924 15918 4928
rect 15854 4868 15858 4924
rect 15858 4868 15914 4924
rect 15914 4868 15918 4924
rect 15854 4864 15918 4868
rect 21479 4924 21543 4928
rect 21479 4868 21483 4924
rect 21483 4868 21539 4924
rect 21539 4868 21543 4924
rect 21479 4864 21543 4868
rect 21559 4924 21623 4928
rect 21559 4868 21563 4924
rect 21563 4868 21619 4924
rect 21619 4868 21623 4924
rect 21559 4864 21623 4868
rect 21639 4924 21703 4928
rect 21639 4868 21643 4924
rect 21643 4868 21699 4924
rect 21699 4868 21703 4924
rect 21639 4864 21703 4868
rect 21719 4924 21783 4928
rect 21719 4868 21723 4924
rect 21723 4868 21779 4924
rect 21779 4868 21783 4924
rect 21719 4864 21783 4868
rect 6816 4380 6880 4384
rect 6816 4324 6820 4380
rect 6820 4324 6876 4380
rect 6876 4324 6880 4380
rect 6816 4320 6880 4324
rect 6896 4380 6960 4384
rect 6896 4324 6900 4380
rect 6900 4324 6956 4380
rect 6956 4324 6960 4380
rect 6896 4320 6960 4324
rect 6976 4380 7040 4384
rect 6976 4324 6980 4380
rect 6980 4324 7036 4380
rect 7036 4324 7040 4380
rect 6976 4320 7040 4324
rect 7056 4380 7120 4384
rect 7056 4324 7060 4380
rect 7060 4324 7116 4380
rect 7116 4324 7120 4380
rect 7056 4320 7120 4324
rect 12681 4380 12745 4384
rect 12681 4324 12685 4380
rect 12685 4324 12741 4380
rect 12741 4324 12745 4380
rect 12681 4320 12745 4324
rect 12761 4380 12825 4384
rect 12761 4324 12765 4380
rect 12765 4324 12821 4380
rect 12821 4324 12825 4380
rect 12761 4320 12825 4324
rect 12841 4380 12905 4384
rect 12841 4324 12845 4380
rect 12845 4324 12901 4380
rect 12901 4324 12905 4380
rect 12841 4320 12905 4324
rect 12921 4380 12985 4384
rect 12921 4324 12925 4380
rect 12925 4324 12981 4380
rect 12981 4324 12985 4380
rect 12921 4320 12985 4324
rect 18546 4380 18610 4384
rect 18546 4324 18550 4380
rect 18550 4324 18606 4380
rect 18606 4324 18610 4380
rect 18546 4320 18610 4324
rect 18626 4380 18690 4384
rect 18626 4324 18630 4380
rect 18630 4324 18686 4380
rect 18686 4324 18690 4380
rect 18626 4320 18690 4324
rect 18706 4380 18770 4384
rect 18706 4324 18710 4380
rect 18710 4324 18766 4380
rect 18766 4324 18770 4380
rect 18706 4320 18770 4324
rect 18786 4380 18850 4384
rect 18786 4324 18790 4380
rect 18790 4324 18846 4380
rect 18846 4324 18850 4380
rect 18786 4320 18850 4324
rect 24411 4380 24475 4384
rect 24411 4324 24415 4380
rect 24415 4324 24471 4380
rect 24471 4324 24475 4380
rect 24411 4320 24475 4324
rect 24491 4380 24555 4384
rect 24491 4324 24495 4380
rect 24495 4324 24551 4380
rect 24551 4324 24555 4380
rect 24491 4320 24555 4324
rect 24571 4380 24635 4384
rect 24571 4324 24575 4380
rect 24575 4324 24631 4380
rect 24631 4324 24635 4380
rect 24571 4320 24635 4324
rect 24651 4380 24715 4384
rect 24651 4324 24655 4380
rect 24655 4324 24711 4380
rect 24711 4324 24715 4380
rect 24651 4320 24715 4324
rect 3884 3836 3948 3840
rect 3884 3780 3888 3836
rect 3888 3780 3944 3836
rect 3944 3780 3948 3836
rect 3884 3776 3948 3780
rect 3964 3836 4028 3840
rect 3964 3780 3968 3836
rect 3968 3780 4024 3836
rect 4024 3780 4028 3836
rect 3964 3776 4028 3780
rect 4044 3836 4108 3840
rect 4044 3780 4048 3836
rect 4048 3780 4104 3836
rect 4104 3780 4108 3836
rect 4044 3776 4108 3780
rect 4124 3836 4188 3840
rect 4124 3780 4128 3836
rect 4128 3780 4184 3836
rect 4184 3780 4188 3836
rect 4124 3776 4188 3780
rect 9749 3836 9813 3840
rect 9749 3780 9753 3836
rect 9753 3780 9809 3836
rect 9809 3780 9813 3836
rect 9749 3776 9813 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 15614 3836 15678 3840
rect 15614 3780 15618 3836
rect 15618 3780 15674 3836
rect 15674 3780 15678 3836
rect 15614 3776 15678 3780
rect 15694 3836 15758 3840
rect 15694 3780 15698 3836
rect 15698 3780 15754 3836
rect 15754 3780 15758 3836
rect 15694 3776 15758 3780
rect 15774 3836 15838 3840
rect 15774 3780 15778 3836
rect 15778 3780 15834 3836
rect 15834 3780 15838 3836
rect 15774 3776 15838 3780
rect 15854 3836 15918 3840
rect 15854 3780 15858 3836
rect 15858 3780 15914 3836
rect 15914 3780 15918 3836
rect 15854 3776 15918 3780
rect 21479 3836 21543 3840
rect 21479 3780 21483 3836
rect 21483 3780 21539 3836
rect 21539 3780 21543 3836
rect 21479 3776 21543 3780
rect 21559 3836 21623 3840
rect 21559 3780 21563 3836
rect 21563 3780 21619 3836
rect 21619 3780 21623 3836
rect 21559 3776 21623 3780
rect 21639 3836 21703 3840
rect 21639 3780 21643 3836
rect 21643 3780 21699 3836
rect 21699 3780 21703 3836
rect 21639 3776 21703 3780
rect 21719 3836 21783 3840
rect 21719 3780 21723 3836
rect 21723 3780 21779 3836
rect 21779 3780 21783 3836
rect 21719 3776 21783 3780
rect 6816 3292 6880 3296
rect 6816 3236 6820 3292
rect 6820 3236 6876 3292
rect 6876 3236 6880 3292
rect 6816 3232 6880 3236
rect 6896 3292 6960 3296
rect 6896 3236 6900 3292
rect 6900 3236 6956 3292
rect 6956 3236 6960 3292
rect 6896 3232 6960 3236
rect 6976 3292 7040 3296
rect 6976 3236 6980 3292
rect 6980 3236 7036 3292
rect 7036 3236 7040 3292
rect 6976 3232 7040 3236
rect 7056 3292 7120 3296
rect 7056 3236 7060 3292
rect 7060 3236 7116 3292
rect 7116 3236 7120 3292
rect 7056 3232 7120 3236
rect 12681 3292 12745 3296
rect 12681 3236 12685 3292
rect 12685 3236 12741 3292
rect 12741 3236 12745 3292
rect 12681 3232 12745 3236
rect 12761 3292 12825 3296
rect 12761 3236 12765 3292
rect 12765 3236 12821 3292
rect 12821 3236 12825 3292
rect 12761 3232 12825 3236
rect 12841 3292 12905 3296
rect 12841 3236 12845 3292
rect 12845 3236 12901 3292
rect 12901 3236 12905 3292
rect 12841 3232 12905 3236
rect 12921 3292 12985 3296
rect 12921 3236 12925 3292
rect 12925 3236 12981 3292
rect 12981 3236 12985 3292
rect 12921 3232 12985 3236
rect 18546 3292 18610 3296
rect 18546 3236 18550 3292
rect 18550 3236 18606 3292
rect 18606 3236 18610 3292
rect 18546 3232 18610 3236
rect 18626 3292 18690 3296
rect 18626 3236 18630 3292
rect 18630 3236 18686 3292
rect 18686 3236 18690 3292
rect 18626 3232 18690 3236
rect 18706 3292 18770 3296
rect 18706 3236 18710 3292
rect 18710 3236 18766 3292
rect 18766 3236 18770 3292
rect 18706 3232 18770 3236
rect 18786 3292 18850 3296
rect 18786 3236 18790 3292
rect 18790 3236 18846 3292
rect 18846 3236 18850 3292
rect 18786 3232 18850 3236
rect 24411 3292 24475 3296
rect 24411 3236 24415 3292
rect 24415 3236 24471 3292
rect 24471 3236 24475 3292
rect 24411 3232 24475 3236
rect 24491 3292 24555 3296
rect 24491 3236 24495 3292
rect 24495 3236 24551 3292
rect 24551 3236 24555 3292
rect 24491 3232 24555 3236
rect 24571 3292 24635 3296
rect 24571 3236 24575 3292
rect 24575 3236 24631 3292
rect 24631 3236 24635 3292
rect 24571 3232 24635 3236
rect 24651 3292 24715 3296
rect 24651 3236 24655 3292
rect 24655 3236 24711 3292
rect 24711 3236 24715 3292
rect 24651 3232 24715 3236
rect 3884 2748 3948 2752
rect 3884 2692 3888 2748
rect 3888 2692 3944 2748
rect 3944 2692 3948 2748
rect 3884 2688 3948 2692
rect 3964 2748 4028 2752
rect 3964 2692 3968 2748
rect 3968 2692 4024 2748
rect 4024 2692 4028 2748
rect 3964 2688 4028 2692
rect 4044 2748 4108 2752
rect 4044 2692 4048 2748
rect 4048 2692 4104 2748
rect 4104 2692 4108 2748
rect 4044 2688 4108 2692
rect 4124 2748 4188 2752
rect 4124 2692 4128 2748
rect 4128 2692 4184 2748
rect 4184 2692 4188 2748
rect 4124 2688 4188 2692
rect 9749 2748 9813 2752
rect 9749 2692 9753 2748
rect 9753 2692 9809 2748
rect 9809 2692 9813 2748
rect 9749 2688 9813 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 15614 2748 15678 2752
rect 15614 2692 15618 2748
rect 15618 2692 15674 2748
rect 15674 2692 15678 2748
rect 15614 2688 15678 2692
rect 15694 2748 15758 2752
rect 15694 2692 15698 2748
rect 15698 2692 15754 2748
rect 15754 2692 15758 2748
rect 15694 2688 15758 2692
rect 15774 2748 15838 2752
rect 15774 2692 15778 2748
rect 15778 2692 15834 2748
rect 15834 2692 15838 2748
rect 15774 2688 15838 2692
rect 15854 2748 15918 2752
rect 15854 2692 15858 2748
rect 15858 2692 15914 2748
rect 15914 2692 15918 2748
rect 15854 2688 15918 2692
rect 21479 2748 21543 2752
rect 21479 2692 21483 2748
rect 21483 2692 21539 2748
rect 21539 2692 21543 2748
rect 21479 2688 21543 2692
rect 21559 2748 21623 2752
rect 21559 2692 21563 2748
rect 21563 2692 21619 2748
rect 21619 2692 21623 2748
rect 21559 2688 21623 2692
rect 21639 2748 21703 2752
rect 21639 2692 21643 2748
rect 21643 2692 21699 2748
rect 21699 2692 21703 2748
rect 21639 2688 21703 2692
rect 21719 2748 21783 2752
rect 21719 2692 21723 2748
rect 21723 2692 21779 2748
rect 21779 2692 21783 2748
rect 21719 2688 21783 2692
rect 6816 2204 6880 2208
rect 6816 2148 6820 2204
rect 6820 2148 6876 2204
rect 6876 2148 6880 2204
rect 6816 2144 6880 2148
rect 6896 2204 6960 2208
rect 6896 2148 6900 2204
rect 6900 2148 6956 2204
rect 6956 2148 6960 2204
rect 6896 2144 6960 2148
rect 6976 2204 7040 2208
rect 6976 2148 6980 2204
rect 6980 2148 7036 2204
rect 7036 2148 7040 2204
rect 6976 2144 7040 2148
rect 7056 2204 7120 2208
rect 7056 2148 7060 2204
rect 7060 2148 7116 2204
rect 7116 2148 7120 2204
rect 7056 2144 7120 2148
rect 12681 2204 12745 2208
rect 12681 2148 12685 2204
rect 12685 2148 12741 2204
rect 12741 2148 12745 2204
rect 12681 2144 12745 2148
rect 12761 2204 12825 2208
rect 12761 2148 12765 2204
rect 12765 2148 12821 2204
rect 12821 2148 12825 2204
rect 12761 2144 12825 2148
rect 12841 2204 12905 2208
rect 12841 2148 12845 2204
rect 12845 2148 12901 2204
rect 12901 2148 12905 2204
rect 12841 2144 12905 2148
rect 12921 2204 12985 2208
rect 12921 2148 12925 2204
rect 12925 2148 12981 2204
rect 12981 2148 12985 2204
rect 12921 2144 12985 2148
rect 18546 2204 18610 2208
rect 18546 2148 18550 2204
rect 18550 2148 18606 2204
rect 18606 2148 18610 2204
rect 18546 2144 18610 2148
rect 18626 2204 18690 2208
rect 18626 2148 18630 2204
rect 18630 2148 18686 2204
rect 18686 2148 18690 2204
rect 18626 2144 18690 2148
rect 18706 2204 18770 2208
rect 18706 2148 18710 2204
rect 18710 2148 18766 2204
rect 18766 2148 18770 2204
rect 18706 2144 18770 2148
rect 18786 2204 18850 2208
rect 18786 2148 18790 2204
rect 18790 2148 18846 2204
rect 18846 2148 18850 2204
rect 18786 2144 18850 2148
rect 24411 2204 24475 2208
rect 24411 2148 24415 2204
rect 24415 2148 24471 2204
rect 24471 2148 24475 2204
rect 24411 2144 24475 2148
rect 24491 2204 24555 2208
rect 24491 2148 24495 2204
rect 24495 2148 24551 2204
rect 24551 2148 24555 2204
rect 24491 2144 24555 2148
rect 24571 2204 24635 2208
rect 24571 2148 24575 2204
rect 24575 2148 24631 2204
rect 24631 2148 24635 2204
rect 24571 2144 24635 2148
rect 24651 2204 24715 2208
rect 24651 2148 24655 2204
rect 24655 2148 24711 2204
rect 24711 2148 24715 2204
rect 24651 2144 24715 2148
rect 3884 1660 3948 1664
rect 3884 1604 3888 1660
rect 3888 1604 3944 1660
rect 3944 1604 3948 1660
rect 3884 1600 3948 1604
rect 3964 1660 4028 1664
rect 3964 1604 3968 1660
rect 3968 1604 4024 1660
rect 4024 1604 4028 1660
rect 3964 1600 4028 1604
rect 4044 1660 4108 1664
rect 4044 1604 4048 1660
rect 4048 1604 4104 1660
rect 4104 1604 4108 1660
rect 4044 1600 4108 1604
rect 4124 1660 4188 1664
rect 4124 1604 4128 1660
rect 4128 1604 4184 1660
rect 4184 1604 4188 1660
rect 4124 1600 4188 1604
rect 9749 1660 9813 1664
rect 9749 1604 9753 1660
rect 9753 1604 9809 1660
rect 9809 1604 9813 1660
rect 9749 1600 9813 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 13676 1668 13740 1732
rect 15614 1660 15678 1664
rect 15614 1604 15618 1660
rect 15618 1604 15674 1660
rect 15674 1604 15678 1660
rect 15614 1600 15678 1604
rect 15694 1660 15758 1664
rect 15694 1604 15698 1660
rect 15698 1604 15754 1660
rect 15754 1604 15758 1660
rect 15694 1600 15758 1604
rect 15774 1660 15838 1664
rect 15774 1604 15778 1660
rect 15778 1604 15834 1660
rect 15834 1604 15838 1660
rect 15774 1600 15838 1604
rect 15854 1660 15918 1664
rect 15854 1604 15858 1660
rect 15858 1604 15914 1660
rect 15914 1604 15918 1660
rect 15854 1600 15918 1604
rect 21479 1660 21543 1664
rect 21479 1604 21483 1660
rect 21483 1604 21539 1660
rect 21539 1604 21543 1660
rect 21479 1600 21543 1604
rect 21559 1660 21623 1664
rect 21559 1604 21563 1660
rect 21563 1604 21619 1660
rect 21619 1604 21623 1660
rect 21559 1600 21623 1604
rect 21639 1660 21703 1664
rect 21639 1604 21643 1660
rect 21643 1604 21699 1660
rect 21699 1604 21703 1660
rect 21639 1600 21703 1604
rect 21719 1660 21783 1664
rect 21719 1604 21723 1660
rect 21723 1604 21779 1660
rect 21779 1604 21783 1660
rect 21719 1600 21783 1604
rect 6816 1116 6880 1120
rect 6816 1060 6820 1116
rect 6820 1060 6876 1116
rect 6876 1060 6880 1116
rect 6816 1056 6880 1060
rect 6896 1116 6960 1120
rect 6896 1060 6900 1116
rect 6900 1060 6956 1116
rect 6956 1060 6960 1116
rect 6896 1056 6960 1060
rect 6976 1116 7040 1120
rect 6976 1060 6980 1116
rect 6980 1060 7036 1116
rect 7036 1060 7040 1116
rect 6976 1056 7040 1060
rect 7056 1116 7120 1120
rect 7056 1060 7060 1116
rect 7060 1060 7116 1116
rect 7116 1060 7120 1116
rect 7056 1056 7120 1060
rect 12681 1116 12745 1120
rect 12681 1060 12685 1116
rect 12685 1060 12741 1116
rect 12741 1060 12745 1116
rect 12681 1056 12745 1060
rect 12761 1116 12825 1120
rect 12761 1060 12765 1116
rect 12765 1060 12821 1116
rect 12821 1060 12825 1116
rect 12761 1056 12825 1060
rect 12841 1116 12905 1120
rect 12841 1060 12845 1116
rect 12845 1060 12901 1116
rect 12901 1060 12905 1116
rect 12841 1056 12905 1060
rect 12921 1116 12985 1120
rect 12921 1060 12925 1116
rect 12925 1060 12981 1116
rect 12981 1060 12985 1116
rect 12921 1056 12985 1060
rect 18546 1116 18610 1120
rect 18546 1060 18550 1116
rect 18550 1060 18606 1116
rect 18606 1060 18610 1116
rect 18546 1056 18610 1060
rect 18626 1116 18690 1120
rect 18626 1060 18630 1116
rect 18630 1060 18686 1116
rect 18686 1060 18690 1116
rect 18626 1056 18690 1060
rect 18706 1116 18770 1120
rect 18706 1060 18710 1116
rect 18710 1060 18766 1116
rect 18766 1060 18770 1116
rect 18706 1056 18770 1060
rect 18786 1116 18850 1120
rect 18786 1060 18790 1116
rect 18790 1060 18846 1116
rect 18846 1060 18850 1116
rect 18786 1056 18850 1060
rect 24411 1116 24475 1120
rect 24411 1060 24415 1116
rect 24415 1060 24471 1116
rect 24471 1060 24475 1116
rect 24411 1056 24475 1060
rect 24491 1116 24555 1120
rect 24491 1060 24495 1116
rect 24495 1060 24551 1116
rect 24551 1060 24555 1116
rect 24491 1056 24555 1060
rect 24571 1116 24635 1120
rect 24571 1060 24575 1116
rect 24575 1060 24631 1116
rect 24631 1060 24635 1116
rect 24571 1056 24635 1060
rect 24651 1116 24715 1120
rect 24651 1060 24655 1116
rect 24655 1060 24711 1116
rect 24711 1060 24715 1116
rect 24651 1056 24715 1060
rect 13676 36 13740 100
<< metal4 >>
rect 3876 8192 4196 8752
rect 3876 8128 3884 8192
rect 3948 8128 3964 8192
rect 4028 8128 4044 8192
rect 4108 8128 4124 8192
rect 4188 8128 4196 8192
rect 3876 7104 4196 8128
rect 3876 7040 3884 7104
rect 3948 7040 3964 7104
rect 4028 7040 4044 7104
rect 4108 7040 4124 7104
rect 4188 7040 4196 7104
rect 3876 6016 4196 7040
rect 3876 5952 3884 6016
rect 3948 5952 3964 6016
rect 4028 5952 4044 6016
rect 4108 5952 4124 6016
rect 4188 5952 4196 6016
rect 3876 4928 4196 5952
rect 3876 4864 3884 4928
rect 3948 4864 3964 4928
rect 4028 4864 4044 4928
rect 4108 4864 4124 4928
rect 4188 4864 4196 4928
rect 3876 3840 4196 4864
rect 3876 3776 3884 3840
rect 3948 3776 3964 3840
rect 4028 3776 4044 3840
rect 4108 3776 4124 3840
rect 4188 3776 4196 3840
rect 3876 2752 4196 3776
rect 3876 2688 3884 2752
rect 3948 2688 3964 2752
rect 4028 2688 4044 2752
rect 4108 2688 4124 2752
rect 4188 2688 4196 2752
rect 3876 1664 4196 2688
rect 3876 1600 3884 1664
rect 3948 1600 3964 1664
rect 4028 1600 4044 1664
rect 4108 1600 4124 1664
rect 4188 1600 4196 1664
rect 3876 1040 4196 1600
rect 6808 8736 7128 8752
rect 6808 8672 6816 8736
rect 6880 8672 6896 8736
rect 6960 8672 6976 8736
rect 7040 8672 7056 8736
rect 7120 8672 7128 8736
rect 6808 7648 7128 8672
rect 6808 7584 6816 7648
rect 6880 7584 6896 7648
rect 6960 7584 6976 7648
rect 7040 7584 7056 7648
rect 7120 7584 7128 7648
rect 6808 6560 7128 7584
rect 6808 6496 6816 6560
rect 6880 6496 6896 6560
rect 6960 6496 6976 6560
rect 7040 6496 7056 6560
rect 7120 6496 7128 6560
rect 6808 5472 7128 6496
rect 6808 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6976 5472
rect 7040 5408 7056 5472
rect 7120 5408 7128 5472
rect 6808 4384 7128 5408
rect 6808 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6976 4384
rect 7040 4320 7056 4384
rect 7120 4320 7128 4384
rect 6808 3296 7128 4320
rect 6808 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6976 3296
rect 7040 3232 7056 3296
rect 7120 3232 7128 3296
rect 6808 2208 7128 3232
rect 6808 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6976 2208
rect 7040 2144 7056 2208
rect 7120 2144 7128 2208
rect 6808 1120 7128 2144
rect 6808 1056 6816 1120
rect 6880 1056 6896 1120
rect 6960 1056 6976 1120
rect 7040 1056 7056 1120
rect 7120 1056 7128 1120
rect 6808 1040 7128 1056
rect 9741 8192 10061 8752
rect 9741 8128 9749 8192
rect 9813 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10061 8192
rect 9741 7104 10061 8128
rect 9741 7040 9749 7104
rect 9813 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10061 7104
rect 9741 6016 10061 7040
rect 9741 5952 9749 6016
rect 9813 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10061 6016
rect 9741 4928 10061 5952
rect 9741 4864 9749 4928
rect 9813 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10061 4928
rect 9741 3840 10061 4864
rect 9741 3776 9749 3840
rect 9813 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10061 3840
rect 9741 2752 10061 3776
rect 9741 2688 9749 2752
rect 9813 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10061 2752
rect 9741 1664 10061 2688
rect 9741 1600 9749 1664
rect 9813 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10061 1664
rect 9741 1040 10061 1600
rect 12673 8736 12993 8752
rect 12673 8672 12681 8736
rect 12745 8672 12761 8736
rect 12825 8672 12841 8736
rect 12905 8672 12921 8736
rect 12985 8672 12993 8736
rect 12673 7648 12993 8672
rect 12673 7584 12681 7648
rect 12745 7584 12761 7648
rect 12825 7584 12841 7648
rect 12905 7584 12921 7648
rect 12985 7584 12993 7648
rect 12673 6560 12993 7584
rect 12673 6496 12681 6560
rect 12745 6496 12761 6560
rect 12825 6496 12841 6560
rect 12905 6496 12921 6560
rect 12985 6496 12993 6560
rect 12673 5472 12993 6496
rect 12673 5408 12681 5472
rect 12745 5408 12761 5472
rect 12825 5408 12841 5472
rect 12905 5408 12921 5472
rect 12985 5408 12993 5472
rect 12673 4384 12993 5408
rect 12673 4320 12681 4384
rect 12745 4320 12761 4384
rect 12825 4320 12841 4384
rect 12905 4320 12921 4384
rect 12985 4320 12993 4384
rect 12673 3296 12993 4320
rect 12673 3232 12681 3296
rect 12745 3232 12761 3296
rect 12825 3232 12841 3296
rect 12905 3232 12921 3296
rect 12985 3232 12993 3296
rect 12673 2208 12993 3232
rect 12673 2144 12681 2208
rect 12745 2144 12761 2208
rect 12825 2144 12841 2208
rect 12905 2144 12921 2208
rect 12985 2144 12993 2208
rect 12673 1120 12993 2144
rect 15606 8192 15926 8752
rect 15606 8128 15614 8192
rect 15678 8128 15694 8192
rect 15758 8128 15774 8192
rect 15838 8128 15854 8192
rect 15918 8128 15926 8192
rect 15606 7104 15926 8128
rect 15606 7040 15614 7104
rect 15678 7040 15694 7104
rect 15758 7040 15774 7104
rect 15838 7040 15854 7104
rect 15918 7040 15926 7104
rect 15606 6016 15926 7040
rect 15606 5952 15614 6016
rect 15678 5952 15694 6016
rect 15758 5952 15774 6016
rect 15838 5952 15854 6016
rect 15918 5952 15926 6016
rect 15606 4928 15926 5952
rect 15606 4864 15614 4928
rect 15678 4864 15694 4928
rect 15758 4864 15774 4928
rect 15838 4864 15854 4928
rect 15918 4864 15926 4928
rect 15606 3840 15926 4864
rect 15606 3776 15614 3840
rect 15678 3776 15694 3840
rect 15758 3776 15774 3840
rect 15838 3776 15854 3840
rect 15918 3776 15926 3840
rect 15606 2752 15926 3776
rect 15606 2688 15614 2752
rect 15678 2688 15694 2752
rect 15758 2688 15774 2752
rect 15838 2688 15854 2752
rect 15918 2688 15926 2752
rect 13675 1732 13741 1733
rect 13675 1668 13676 1732
rect 13740 1668 13741 1732
rect 13675 1667 13741 1668
rect 12673 1056 12681 1120
rect 12745 1056 12761 1120
rect 12825 1056 12841 1120
rect 12905 1056 12921 1120
rect 12985 1056 12993 1120
rect 12673 1040 12993 1056
rect 13678 101 13738 1667
rect 15606 1664 15926 2688
rect 15606 1600 15614 1664
rect 15678 1600 15694 1664
rect 15758 1600 15774 1664
rect 15838 1600 15854 1664
rect 15918 1600 15926 1664
rect 15606 1040 15926 1600
rect 18538 8736 18858 8752
rect 18538 8672 18546 8736
rect 18610 8672 18626 8736
rect 18690 8672 18706 8736
rect 18770 8672 18786 8736
rect 18850 8672 18858 8736
rect 18538 7648 18858 8672
rect 18538 7584 18546 7648
rect 18610 7584 18626 7648
rect 18690 7584 18706 7648
rect 18770 7584 18786 7648
rect 18850 7584 18858 7648
rect 18538 6560 18858 7584
rect 18538 6496 18546 6560
rect 18610 6496 18626 6560
rect 18690 6496 18706 6560
rect 18770 6496 18786 6560
rect 18850 6496 18858 6560
rect 18538 5472 18858 6496
rect 18538 5408 18546 5472
rect 18610 5408 18626 5472
rect 18690 5408 18706 5472
rect 18770 5408 18786 5472
rect 18850 5408 18858 5472
rect 18538 4384 18858 5408
rect 18538 4320 18546 4384
rect 18610 4320 18626 4384
rect 18690 4320 18706 4384
rect 18770 4320 18786 4384
rect 18850 4320 18858 4384
rect 18538 3296 18858 4320
rect 18538 3232 18546 3296
rect 18610 3232 18626 3296
rect 18690 3232 18706 3296
rect 18770 3232 18786 3296
rect 18850 3232 18858 3296
rect 18538 2208 18858 3232
rect 18538 2144 18546 2208
rect 18610 2144 18626 2208
rect 18690 2144 18706 2208
rect 18770 2144 18786 2208
rect 18850 2144 18858 2208
rect 18538 1120 18858 2144
rect 18538 1056 18546 1120
rect 18610 1056 18626 1120
rect 18690 1056 18706 1120
rect 18770 1056 18786 1120
rect 18850 1056 18858 1120
rect 18538 1040 18858 1056
rect 21471 8192 21791 8752
rect 21471 8128 21479 8192
rect 21543 8128 21559 8192
rect 21623 8128 21639 8192
rect 21703 8128 21719 8192
rect 21783 8128 21791 8192
rect 21471 7104 21791 8128
rect 21471 7040 21479 7104
rect 21543 7040 21559 7104
rect 21623 7040 21639 7104
rect 21703 7040 21719 7104
rect 21783 7040 21791 7104
rect 21471 6016 21791 7040
rect 21471 5952 21479 6016
rect 21543 5952 21559 6016
rect 21623 5952 21639 6016
rect 21703 5952 21719 6016
rect 21783 5952 21791 6016
rect 21471 4928 21791 5952
rect 21471 4864 21479 4928
rect 21543 4864 21559 4928
rect 21623 4864 21639 4928
rect 21703 4864 21719 4928
rect 21783 4864 21791 4928
rect 21471 3840 21791 4864
rect 21471 3776 21479 3840
rect 21543 3776 21559 3840
rect 21623 3776 21639 3840
rect 21703 3776 21719 3840
rect 21783 3776 21791 3840
rect 21471 2752 21791 3776
rect 21471 2688 21479 2752
rect 21543 2688 21559 2752
rect 21623 2688 21639 2752
rect 21703 2688 21719 2752
rect 21783 2688 21791 2752
rect 21471 1664 21791 2688
rect 21471 1600 21479 1664
rect 21543 1600 21559 1664
rect 21623 1600 21639 1664
rect 21703 1600 21719 1664
rect 21783 1600 21791 1664
rect 21471 1040 21791 1600
rect 24403 8736 24723 8752
rect 24403 8672 24411 8736
rect 24475 8672 24491 8736
rect 24555 8672 24571 8736
rect 24635 8672 24651 8736
rect 24715 8672 24723 8736
rect 24403 7648 24723 8672
rect 24403 7584 24411 7648
rect 24475 7584 24491 7648
rect 24555 7584 24571 7648
rect 24635 7584 24651 7648
rect 24715 7584 24723 7648
rect 24403 6560 24723 7584
rect 24403 6496 24411 6560
rect 24475 6496 24491 6560
rect 24555 6496 24571 6560
rect 24635 6496 24651 6560
rect 24715 6496 24723 6560
rect 24403 5472 24723 6496
rect 24403 5408 24411 5472
rect 24475 5408 24491 5472
rect 24555 5408 24571 5472
rect 24635 5408 24651 5472
rect 24715 5408 24723 5472
rect 24403 4384 24723 5408
rect 24403 4320 24411 4384
rect 24475 4320 24491 4384
rect 24555 4320 24571 4384
rect 24635 4320 24651 4384
rect 24715 4320 24723 4384
rect 24403 3296 24723 4320
rect 24403 3232 24411 3296
rect 24475 3232 24491 3296
rect 24555 3232 24571 3296
rect 24635 3232 24651 3296
rect 24715 3232 24723 3296
rect 24403 2208 24723 3232
rect 24403 2144 24411 2208
rect 24475 2144 24491 2208
rect 24555 2144 24571 2208
rect 24635 2144 24651 2208
rect 24715 2144 24723 2208
rect 24403 1120 24723 2144
rect 24403 1056 24411 1120
rect 24475 1056 24491 1120
rect 24555 1056 24571 1120
rect 24635 1056 24651 1120
rect 24715 1056 24723 1120
rect 24403 1040 24723 1056
rect 13675 100 13741 101
rect 13675 36 13676 100
rect 13740 36 13741 100
rect 13675 35 13741 36
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_128
timestamp 1688980957
transform 1 0 12880 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1688980957
transform 1 0 13800 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp 1688980957
transform 1 0 21528 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_17 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2668 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_29
timestamp 1688980957
transform 1 0 3772 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_41 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4876 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_66
timestamp 1688980957
transform 1 0 7176 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_74
timestamp 1688980957
transform 1 0 7912 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_79
timestamp 1688980957
transform 1 0 8372 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_104
timestamp 1688980957
transform 1 0 10672 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_122
timestamp 1688980957
transform 1 0 12328 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_130
timestamp 1688980957
transform 1 0 13064 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_153
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_12
timestamp 1688980957
transform 1 0 2208 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_24 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_80
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_103
timestamp 1688980957
transform 1 0 10580 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_107
timestamp 1688980957
transform 1 0 10948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_114
timestamp 1688980957
transform 1 0 11592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_118
timestamp 1688980957
transform 1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_127
timestamp 1688980957
transform 1 0 12788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_161
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_166
timestamp 1688980957
transform 1 0 16376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_179
timestamp 1688980957
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_187
timestamp 1688980957
transform 1 0 18308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_191
timestamp 1688980957
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_200
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_208
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_220
timestamp 1688980957
transform 1 0 21344 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_226
timestamp 1688980957
transform 1 0 21896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_75
timestamp 1688980957
transform 1 0 8004 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_79
timestamp 1688980957
transform 1 0 8372 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_91
timestamp 1688980957
transform 1 0 9476 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_103
timestamp 1688980957
transform 1 0 10580 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_158
timestamp 1688980957
transform 1 0 15640 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1688980957
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_231
timestamp 1688980957
transform 1 0 22356 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_250
timestamp 1688980957
transform 1 0 24104 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_94
timestamp 1688980957
transform 1 0 9752 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_102
timestamp 1688980957
transform 1 0 10488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_106
timestamp 1688980957
transform 1 0 10856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_114
timestamp 1688980957
transform 1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_119
timestamp 1688980957
transform 1 0 12052 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_127
timestamp 1688980957
transform 1 0 12788 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_132
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_147
timestamp 1688980957
transform 1 0 14628 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_157
timestamp 1688980957
transform 1 0 15548 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_169
timestamp 1688980957
transform 1 0 16652 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1688980957
transform 1 0 17756 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_208
timestamp 1688980957
transform 1 0 20240 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_220
timestamp 1688980957
transform 1 0 21344 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_232
timestamp 1688980957
transform 1 0 22448 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_240
timestamp 1688980957
transform 1 0 23184 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_92
timestamp 1688980957
transform 1 0 9568 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_100
timestamp 1688980957
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_118
timestamp 1688980957
transform 1 0 11960 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_126
timestamp 1688980957
transform 1 0 12696 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_131
timestamp 1688980957
transform 1 0 13156 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_143
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_155
timestamp 1688980957
transform 1 0 15364 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_201
timestamp 1688980957
transform 1 0 19596 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_206
timestamp 1688980957
transform 1 0 20056 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_218
timestamp 1688980957
transform 1 0 21160 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_245
timestamp 1688980957
transform 1 0 23644 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_250
timestamp 1688980957
transform 1 0 24104 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_171
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_183
timestamp 1688980957
transform 1 0 17940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_23
timestamp 1688980957
transform 1 0 3220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_41
timestamp 1688980957
transform 1 0 4876 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_49
timestamp 1688980957
transform 1 0 5612 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_75
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_82
timestamp 1688980957
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_101
timestamp 1688980957
transform 1 0 10396 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_106
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_119
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_127
timestamp 1688980957
transform 1 0 12788 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_132
timestamp 1688980957
transform 1 0 13248 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_145
timestamp 1688980957
transform 1 0 14444 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_153
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_160
timestamp 1688980957
transform 1 0 15824 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_178
timestamp 1688980957
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_184
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_203
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_210
timestamp 1688980957
transform 1 0 20424 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_218
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_231
timestamp 1688980957
transform 1 0 22356 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_236
timestamp 1688980957
transform 1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_251
timestamp 1688980957
transform 1 0 24196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1688980957
transform -1 0 23368 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 23092 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 23552 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform -1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform -1 0 23184 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform -1 0 23460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform -1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform -1 0 23460 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform -1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform -1 0 24012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform -1 0 24288 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform -1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform -1 0 2392 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform -1 0 2668 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 2852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input26
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 1688980957
transform 1 0 3404 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform -1 0 4048 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform -1 0 4324 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform -1 0 4600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform -1 0 5428 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform -1 0 5704 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 1564 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 1748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 2024 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 2300 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 4600 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform -1 0 8740 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform -1 0 9016 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 9016 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform -1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform -1 0 9568 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform -1 0 8832 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input49
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input50
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 7360 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input54
timestamp 1688980957
transform 1 0 7636 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform -1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input56
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__00_
timestamp 1688980957
transform -1 0 6256 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__01_
timestamp 1688980957
transform -1 0 7176 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__02_
timestamp 1688980957
transform -1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__03_
timestamp 1688980957
transform -1 0 10120 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__04_
timestamp 1688980957
transform -1 0 12696 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__05_
timestamp 1688980957
transform -1 0 13432 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__06_
timestamp 1688980957
transform -1 0 13708 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__07_
timestamp 1688980957
transform -1 0 13984 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__08_
timestamp 1688980957
transform -1 0 14260 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__09_
timestamp 1688980957
transform -1 0 14536 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__10_
timestamp 1688980957
transform -1 0 14812 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__11_
timestamp 1688980957
transform -1 0 15180 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__12_
timestamp 1688980957
transform -1 0 9292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__13_
timestamp 1688980957
transform -1 0 9568 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__14_
timestamp 1688980957
transform -1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__15_
timestamp 1688980957
transform -1 0 11592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__16_
timestamp 1688980957
transform -1 0 11960 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__17_
timestamp 1688980957
transform -1 0 11776 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__18_
timestamp 1688980957
transform -1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__19_
timestamp 1688980957
transform -1 0 12788 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__20_
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__21_
timestamp 1688980957
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__22_
timestamp 1688980957
transform -1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__23_
timestamp 1688980957
transform -1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__24_
timestamp 1688980957
transform -1 0 18676 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__25_
timestamp 1688980957
transform -1 0 20240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__26_
timestamp 1688980957
transform 1 0 21252 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__27_
timestamp 1688980957
transform 1 0 20884 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__28_
timestamp 1688980957
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix__29_
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__30_
timestamp 1688980957
transform -1 0 17296 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__31_
timestamp 1688980957
transform -1 0 17572 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__32_
timestamp 1688980957
transform -1 0 17020 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__33_
timestamp 1688980957
transform -1 0 8372 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_N_term_RAM_IO_switch_matrix__34_
timestamp 1688980957
transform -1 0 19136 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_N_term_RAM_IO_switch_matrix__35_
timestamp 1688980957
transform 1 0 6624 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 2484 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output60 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform -1 0 17204 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1688980957
transform -1 0 18032 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1688980957
transform -1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1688980957
transform -1 0 21620 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1688980957
transform -1 0 22816 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 23644 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform -1 0 23644 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1688980957
transform -1 0 3680 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1688980957
transform -1 0 4876 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1688980957
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 6900 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 8096 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1688980957
transform 1 0 9292 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1688980957
transform 1 0 11684 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 10120 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 14444 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 15364 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 10672 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 10304 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 11776 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1688980957
transform 1 0 11592 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1688980957
transform 1 0 11960 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 12696 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1688980957
transform 1 0 13064 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform -1 0 16468 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 19780 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 19228 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output102
timestamp 1688980957
transform 1 0 20332 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1688980957
transform -1 0 21252 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform -1 0 20332 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1688980957
transform 1 0 17204 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 18308 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 18676 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 17572 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform 1 0 18124 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output114
timestamp 1688980957
transform -1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24564 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24564 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 24564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 19964 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 22080 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform -1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform -1 0 6900 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 9476 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 11776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 12972 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 15364 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform -1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform -1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 22908 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 23460 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform -1 0 22264 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 23920 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform -1 0 24104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform -1 0 20056 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform -1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform -1 0 22080 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform -1 0 5980 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform -1 0 7176 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 11684 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 12880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 15272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform -1 0 24288 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 22632 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 22356 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 23460 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 23828 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 20258 -300 20314 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 23018 -300 23074 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 23294 -300 23350 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 23570 -300 23626 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 23846 -300 23902 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 24122 -300 24178 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 24398 -300 24454 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 24674 -300 24730 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 24950 -300 25006 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 25226 -300 25282 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 25502 -300 25558 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 20534 -300 20590 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 20810 -300 20866 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 21086 -300 21142 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 21362 -300 21418 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 21638 -300 21694 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 21914 -300 21970 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 22190 -300 22246 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 22466 -300 22522 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 22742 -300 22798 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 2042 9840 2098 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 14002 9840 14058 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 15198 9840 15254 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 16394 9840 16450 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 17590 9840 17646 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 18786 9840 18842 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 19982 9840 20038 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 21178 9840 21234 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 22374 9840 22430 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 23570 9840 23626 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 24766 9840 24822 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 3238 9840 3294 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 4434 9840 4490 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 5630 9840 5686 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 6826 9840 6882 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 8022 9840 8078 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 9218 9840 9274 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 10414 9840 10470 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 11610 9840 11666 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 12806 9840 12862 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 110 -300 166 160 0 FreeSans 224 90 0 0 N1END[0]
port 40 nsew signal input
flabel metal2 s 386 -300 442 160 0 FreeSans 224 90 0 0 N1END[1]
port 41 nsew signal input
flabel metal2 s 662 -300 718 160 0 FreeSans 224 90 0 0 N1END[2]
port 42 nsew signal input
flabel metal2 s 938 -300 994 160 0 FreeSans 224 90 0 0 N1END[3]
port 43 nsew signal input
flabel metal2 s 3422 -300 3478 160 0 FreeSans 224 90 0 0 N2END[0]
port 44 nsew signal input
flabel metal2 s 3698 -300 3754 160 0 FreeSans 224 90 0 0 N2END[1]
port 45 nsew signal input
flabel metal2 s 3974 -300 4030 160 0 FreeSans 224 90 0 0 N2END[2]
port 46 nsew signal input
flabel metal2 s 4250 -300 4306 160 0 FreeSans 224 90 0 0 N2END[3]
port 47 nsew signal input
flabel metal2 s 4526 -300 4582 160 0 FreeSans 224 90 0 0 N2END[4]
port 48 nsew signal input
flabel metal2 s 4802 -300 4858 160 0 FreeSans 224 90 0 0 N2END[5]
port 49 nsew signal input
flabel metal2 s 5078 -300 5134 160 0 FreeSans 224 90 0 0 N2END[6]
port 50 nsew signal input
flabel metal2 s 5354 -300 5410 160 0 FreeSans 224 90 0 0 N2END[7]
port 51 nsew signal input
flabel metal2 s 1214 -300 1270 160 0 FreeSans 224 90 0 0 N2MID[0]
port 52 nsew signal input
flabel metal2 s 1490 -300 1546 160 0 FreeSans 224 90 0 0 N2MID[1]
port 53 nsew signal input
flabel metal2 s 1766 -300 1822 160 0 FreeSans 224 90 0 0 N2MID[2]
port 54 nsew signal input
flabel metal2 s 2042 -300 2098 160 0 FreeSans 224 90 0 0 N2MID[3]
port 55 nsew signal input
flabel metal2 s 2318 -300 2374 160 0 FreeSans 224 90 0 0 N2MID[4]
port 56 nsew signal input
flabel metal2 s 2594 -300 2650 160 0 FreeSans 224 90 0 0 N2MID[5]
port 57 nsew signal input
flabel metal2 s 2870 -300 2926 160 0 FreeSans 224 90 0 0 N2MID[6]
port 58 nsew signal input
flabel metal2 s 3146 -300 3202 160 0 FreeSans 224 90 0 0 N2MID[7]
port 59 nsew signal input
flabel metal2 s 5630 -300 5686 160 0 FreeSans 224 90 0 0 N4END[0]
port 60 nsew signal input
flabel metal2 s 8390 -300 8446 160 0 FreeSans 224 90 0 0 N4END[10]
port 61 nsew signal input
flabel metal2 s 8666 -300 8722 160 0 FreeSans 224 90 0 0 N4END[11]
port 62 nsew signal input
flabel metal2 s 8942 -300 8998 160 0 FreeSans 224 90 0 0 N4END[12]
port 63 nsew signal input
flabel metal2 s 9218 -300 9274 160 0 FreeSans 224 90 0 0 N4END[13]
port 64 nsew signal input
flabel metal2 s 9494 -300 9550 160 0 FreeSans 224 90 0 0 N4END[14]
port 65 nsew signal input
flabel metal2 s 9770 -300 9826 160 0 FreeSans 224 90 0 0 N4END[15]
port 66 nsew signal input
flabel metal2 s 5906 -300 5962 160 0 FreeSans 224 90 0 0 N4END[1]
port 67 nsew signal input
flabel metal2 s 6182 -300 6238 160 0 FreeSans 224 90 0 0 N4END[2]
port 68 nsew signal input
flabel metal2 s 6458 -300 6514 160 0 FreeSans 224 90 0 0 N4END[3]
port 69 nsew signal input
flabel metal2 s 6734 -300 6790 160 0 FreeSans 224 90 0 0 N4END[4]
port 70 nsew signal input
flabel metal2 s 7010 -300 7066 160 0 FreeSans 224 90 0 0 N4END[5]
port 71 nsew signal input
flabel metal2 s 7286 -300 7342 160 0 FreeSans 224 90 0 0 N4END[6]
port 72 nsew signal input
flabel metal2 s 7562 -300 7618 160 0 FreeSans 224 90 0 0 N4END[7]
port 73 nsew signal input
flabel metal2 s 7838 -300 7894 160 0 FreeSans 224 90 0 0 N4END[8]
port 74 nsew signal input
flabel metal2 s 8114 -300 8170 160 0 FreeSans 224 90 0 0 N4END[9]
port 75 nsew signal input
flabel metal2 s 10046 -300 10102 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 76 nsew signal tristate
flabel metal2 s 10322 -300 10378 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 77 nsew signal tristate
flabel metal2 s 10598 -300 10654 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 78 nsew signal tristate
flabel metal2 s 10874 -300 10930 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 79 nsew signal tristate
flabel metal2 s 13358 -300 13414 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 80 nsew signal tristate
flabel metal2 s 13634 -300 13690 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 81 nsew signal tristate
flabel metal2 s 13910 -300 13966 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 82 nsew signal tristate
flabel metal2 s 14186 -300 14242 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 83 nsew signal tristate
flabel metal2 s 14462 -300 14518 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 84 nsew signal tristate
flabel metal2 s 14738 -300 14794 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 85 nsew signal tristate
flabel metal2 s 15014 -300 15070 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 86 nsew signal tristate
flabel metal2 s 15290 -300 15346 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 87 nsew signal tristate
flabel metal2 s 11150 -300 11206 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 88 nsew signal tristate
flabel metal2 s 11426 -300 11482 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 89 nsew signal tristate
flabel metal2 s 11702 -300 11758 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 90 nsew signal tristate
flabel metal2 s 11978 -300 12034 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 91 nsew signal tristate
flabel metal2 s 12254 -300 12310 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 92 nsew signal tristate
flabel metal2 s 12530 -300 12586 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 93 nsew signal tristate
flabel metal2 s 12806 -300 12862 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 94 nsew signal tristate
flabel metal2 s 13082 -300 13138 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 95 nsew signal tristate
flabel metal2 s 15566 -300 15622 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 96 nsew signal tristate
flabel metal2 s 18326 -300 18382 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 97 nsew signal tristate
flabel metal2 s 18602 -300 18658 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 98 nsew signal tristate
flabel metal2 s 18878 -300 18934 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 99 nsew signal tristate
flabel metal2 s 19154 -300 19210 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 100 nsew signal tristate
flabel metal2 s 19430 -300 19486 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 101 nsew signal tristate
flabel metal2 s 19706 -300 19762 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 102 nsew signal tristate
flabel metal2 s 15842 -300 15898 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 103 nsew signal tristate
flabel metal2 s 16118 -300 16174 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 104 nsew signal tristate
flabel metal2 s 16394 -300 16450 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 105 nsew signal tristate
flabel metal2 s 16670 -300 16726 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 106 nsew signal tristate
flabel metal2 s 16946 -300 17002 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 107 nsew signal tristate
flabel metal2 s 17222 -300 17278 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 108 nsew signal tristate
flabel metal2 s 17498 -300 17554 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 109 nsew signal tristate
flabel metal2 s 17774 -300 17830 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 110 nsew signal tristate
flabel metal2 s 18050 -300 18106 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 111 nsew signal tristate
flabel metal2 s 19982 -300 20038 160 0 FreeSans 224 90 0 0 UserCLK
port 112 nsew signal input
flabel metal2 s 846 9840 902 10300 0 FreeSans 224 90 0 0 UserCLKo
port 113 nsew signal tristate
flabel metal4 s 6808 1040 7128 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 12673 1040 12993 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 18538 1040 18858 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 24403 1040 24723 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 3876 1040 4196 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 9741 1040 10061 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 15606 1040 15926 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 21471 1040 21791 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
rlabel via1 12913 8704 12913 8704 0 VGND
rlabel metal1 12834 8160 12834 8160 0 VPWR
rlabel metal2 20385 68 20385 68 0 FrameStrobe[0]
rlabel metal2 22947 68 22947 68 0 FrameStrobe[10]
rlabel metal1 23414 3502 23414 3502 0 FrameStrobe[11]
rlabel metal2 23545 68 23545 68 0 FrameStrobe[12]
rlabel metal1 23828 3026 23828 3026 0 FrameStrobe[13]
rlabel metal2 24150 1180 24150 1180 0 FrameStrobe[14]
rlabel metal2 24373 68 24373 68 0 FrameStrobe[15]
rlabel metal2 24755 68 24755 68 0 FrameStrobe[16]
rlabel metal2 24978 772 24978 772 0 FrameStrobe[17]
rlabel metal2 25254 908 25254 908 0 FrameStrobe[18]
rlabel metal2 25530 1588 25530 1588 0 FrameStrobe[19]
rlabel metal2 20562 500 20562 500 0 FrameStrobe[1]
rlabel metal2 20838 211 20838 211 0 FrameStrobe[2]
rlabel metal2 21114 738 21114 738 0 FrameStrobe[3]
rlabel metal2 21390 432 21390 432 0 FrameStrobe[4]
rlabel metal2 21666 398 21666 398 0 FrameStrobe[5]
rlabel metal2 21995 68 21995 68 0 FrameStrobe[6]
rlabel metal2 22317 68 22317 68 0 FrameStrobe[7]
rlabel metal2 22494 279 22494 279 0 FrameStrobe[8]
rlabel metal2 22770 228 22770 228 0 FrameStrobe[9]
rlabel metal1 2162 8602 2162 8602 0 FrameStrobe_O[0]
rlabel metal1 14168 8602 14168 8602 0 FrameStrobe_O[10]
rlabel metal2 15226 9224 15226 9224 0 FrameStrobe_O[11]
rlabel metal2 16422 9190 16422 9190 0 FrameStrobe_O[12]
rlabel metal1 17710 8602 17710 8602 0 FrameStrobe_O[13]
rlabel metal2 18814 9445 18814 9445 0 FrameStrobe_O[14]
rlabel metal1 20102 8602 20102 8602 0 FrameStrobe_O[15]
rlabel metal1 21298 8602 21298 8602 0 FrameStrobe_O[16]
rlabel metal1 22494 8602 22494 8602 0 FrameStrobe_O[17]
rlabel metal2 23598 9224 23598 9224 0 FrameStrobe_O[18]
rlabel metal1 24012 8398 24012 8398 0 FrameStrobe_O[19]
rlabel metal1 3358 8602 3358 8602 0 FrameStrobe_O[1]
rlabel metal1 4554 8602 4554 8602 0 FrameStrobe_O[2]
rlabel metal2 5658 9224 5658 9224 0 FrameStrobe_O[3]
rlabel metal2 6854 9513 6854 9513 0 FrameStrobe_O[4]
rlabel metal2 8050 9224 8050 9224 0 FrameStrobe_O[5]
rlabel metal1 9384 8602 9384 8602 0 FrameStrobe_O[6]
rlabel metal1 10580 8602 10580 8602 0 FrameStrobe_O[7]
rlabel metal1 11776 8602 11776 8602 0 FrameStrobe_O[8]
rlabel metal2 13110 9231 13110 9231 0 FrameStrobe_O[9]
rlabel metal2 20010 3910 20010 3910 0 FrameStrobe_O_i\[0\]
rlabel metal1 14352 3502 14352 3502 0 FrameStrobe_O_i\[10\]
rlabel metal1 15456 3162 15456 3162 0 FrameStrobe_O_i\[11\]
rlabel metal1 17112 8058 17112 8058 0 FrameStrobe_O_i\[12\]
rlabel metal1 24150 1326 24150 1326 0 FrameStrobe_O_i\[13\]
rlabel metal1 19688 2414 19688 2414 0 FrameStrobe_O_i\[14\]
rlabel metal1 22908 1938 22908 1938 0 FrameStrobe_O_i\[15\]
rlabel metal1 23138 1530 23138 1530 0 FrameStrobe_O_i\[16\]
rlabel metal1 23690 1904 23690 1904 0 FrameStrobe_O_i\[17\]
rlabel metal1 23920 2414 23920 2414 0 FrameStrobe_O_i\[18\]
rlabel metal2 24058 3910 24058 3910 0 FrameStrobe_O_i\[19\]
rlabel metal1 21436 1938 21436 1938 0 FrameStrobe_O_i\[1\]
rlabel metal1 22126 1870 22126 1870 0 FrameStrobe_O_i\[2\]
rlabel metal1 5428 1530 5428 1530 0 FrameStrobe_O_i\[3\]
rlabel metal1 6900 1938 6900 1938 0 FrameStrobe_O_i\[4\]
rlabel metal1 8280 2618 8280 2618 0 FrameStrobe_O_i\[5\]
rlabel metal2 9522 3910 9522 3910 0 FrameStrobe_O_i\[6\]
rlabel metal1 10672 3706 10672 3706 0 FrameStrobe_O_i\[7\]
rlabel metal1 11868 3706 11868 3706 0 FrameStrobe_O_i\[8\]
rlabel metal1 13064 3706 13064 3706 0 FrameStrobe_O_i\[9\]
rlabel metal2 138 1248 138 1248 0 N1END[0]
rlabel metal2 414 942 414 942 0 N1END[1]
rlabel metal2 690 1214 690 1214 0 N1END[2]
rlabel metal2 966 806 966 806 0 N1END[3]
rlabel metal2 3450 704 3450 704 0 N2END[0]
rlabel metal2 3726 670 3726 670 0 N2END[1]
rlabel metal2 3949 68 3949 68 0 N2END[2]
rlabel metal2 4225 68 4225 68 0 N2END[3]
rlabel metal2 4455 68 4455 68 0 N2END[4]
rlabel metal2 4731 68 4731 68 0 N2END[5]
rlabel metal2 5159 68 5159 68 0 N2END[6]
rlabel metal2 5435 68 5435 68 0 N2END[7]
rlabel metal2 1242 976 1242 976 0 N2MID[0]
rlabel metal2 1518 1010 1518 1010 0 N2MID[1]
rlabel metal2 1794 687 1794 687 0 N2MID[2]
rlabel metal2 2070 636 2070 636 0 N2MID[3]
rlabel metal2 2346 415 2346 415 0 N2MID[4]
rlabel metal2 2622 636 2622 636 0 N2MID[5]
rlabel metal2 2530 1377 2530 1377 0 N2MID[6]
rlabel metal2 2714 969 2714 969 0 N2MID[7]
rlabel metal2 5605 68 5605 68 0 N4END[0]
rlabel metal2 8418 1010 8418 1010 0 N4END[10]
rlabel metal2 8747 68 8747 68 0 N4END[11]
rlabel metal2 8970 1010 8970 1010 0 N4END[12]
rlabel metal2 9246 364 9246 364 0 N4END[13]
rlabel metal2 9423 68 9423 68 0 N4END[14]
rlabel metal2 9699 68 9699 68 0 N4END[15]
rlabel metal2 5835 68 5835 68 0 N4END[1]
rlabel metal2 6111 68 6111 68 0 N4END[2]
rlabel metal2 6486 670 6486 670 0 N4END[3]
rlabel metal2 6663 68 6663 68 0 N4END[4]
rlabel metal2 7038 364 7038 364 0 N4END[5]
rlabel metal2 7314 1010 7314 1010 0 N4END[6]
rlabel metal2 7590 1010 7590 1010 0 N4END[7]
rlabel metal2 7813 68 7813 68 0 N4END[8]
rlabel metal2 8142 364 8142 364 0 N4END[9]
rlabel metal2 10021 68 10021 68 0 S1BEG[0]
rlabel metal2 10350 636 10350 636 0 S1BEG[1]
rlabel metal2 10527 68 10527 68 0 S1BEG[2]
rlabel metal2 10955 68 10955 68 0 S1BEG[3]
rlabel metal2 13386 636 13386 636 0 S2BEG[0]
rlabel metal2 13715 68 13715 68 0 S2BEG[1]
rlabel metal2 13938 636 13938 636 0 S2BEG[2]
rlabel metal2 14313 68 14313 68 0 S2BEG[3]
rlabel metal2 14589 68 14589 68 0 S2BEG[4]
rlabel metal2 14865 68 14865 68 0 S2BEG[5]
rlabel metal2 15042 636 15042 636 0 S2BEG[6]
rlabel metal2 15318 908 15318 908 0 S2BEG[7]
rlabel metal2 11125 68 11125 68 0 S2BEGb[0]
rlabel metal2 11355 68 11355 68 0 S2BEGb[1]
rlabel metal2 11730 483 11730 483 0 S2BEGb[2]
rlabel metal2 12006 636 12006 636 0 S2BEGb[3]
rlabel metal2 12282 636 12282 636 0 S2BEGb[4]
rlabel metal2 12558 636 12558 636 0 S2BEGb[5]
rlabel metal2 12933 68 12933 68 0 S2BEGb[6]
rlabel metal2 13110 211 13110 211 0 S2BEGb[7]
rlabel metal2 15541 68 15541 68 0 S4BEG[0]
rlabel metal2 18354 347 18354 347 0 S4BEG[10]
rlabel metal2 18729 68 18729 68 0 S4BEG[11]
rlabel metal2 18906 160 18906 160 0 S4BEG[12]
rlabel metal2 19182 942 19182 942 0 S4BEG[13]
rlabel metal2 19458 636 19458 636 0 S4BEG[14]
rlabel metal2 19833 68 19833 68 0 S4BEG[15]
rlabel metal2 15969 68 15969 68 0 S4BEG[1]
rlabel metal2 16146 347 16146 347 0 S4BEG[2]
rlabel metal2 16422 908 16422 908 0 S4BEG[3]
rlabel metal2 16698 942 16698 942 0 S4BEG[4]
rlabel metal2 16974 806 16974 806 0 S4BEG[5]
rlabel metal2 17250 942 17250 942 0 S4BEG[6]
rlabel metal2 17526 483 17526 483 0 S4BEG[7]
rlabel metal2 17802 738 17802 738 0 S4BEG[8]
rlabel metal2 18078 908 18078 908 0 S4BEG[9]
rlabel metal2 20010 534 20010 534 0 UserCLK
rlabel metal2 874 9785 874 9785 0 UserCLKo
rlabel metal1 20424 3502 20424 3502 0 net1
rlabel metal1 24150 2516 24150 2516 0 net10
rlabel metal1 19366 2040 19366 2040 0 net100
rlabel metal1 20470 1224 20470 1224 0 net101
rlabel metal1 20332 2006 20332 2006 0 net102
rlabel metal1 21252 1326 21252 1326 0 net103
rlabel metal1 20562 1938 20562 1938 0 net104
rlabel metal1 17204 1258 17204 1258 0 net105
rlabel metal1 17894 1292 17894 1292 0 net106
rlabel metal1 12282 2890 12282 2890 0 net107
rlabel metal1 17250 2006 17250 2006 0 net108
rlabel metal1 18308 1326 18308 1326 0 net109
rlabel metal2 23506 3094 23506 3094 0 net11
rlabel metal1 18584 2006 18584 2006 0 net110
rlabel metal2 14858 1649 14858 1649 0 net111
rlabel metal1 19228 1258 19228 1258 0 net112
rlabel metal2 6808 2924 6808 2924 0 net113
rlabel metal2 1794 5423 1794 5423 0 net114
rlabel metal1 21666 1972 21666 1972 0 net12
rlabel metal1 22494 1530 22494 1530 0 net13
rlabel metal4 13708 884 13708 884 0 net14
rlabel metal1 11592 3094 11592 3094 0 net15
rlabel metal1 11500 2822 11500 2822 0 net16
rlabel metal1 10166 3502 10166 3502 0 net17
rlabel metal1 10810 3978 10810 3978 0 net18
rlabel metal2 12006 3009 12006 3009 0 net19
rlabel metal1 19550 2992 19550 2992 0 net2
rlabel metal1 14490 3502 14490 3502 0 net20
rlabel metal1 9890 2482 9890 2482 0 net21
rlabel metal1 7774 1360 7774 1360 0 net22
rlabel metal1 1518 2550 1518 2550 0 net23
rlabel metal1 2622 1836 2622 1836 0 net24
rlabel metal3 8418 3060 8418 3060 0 net25
rlabel metal1 3864 1462 3864 1462 0 net26
rlabel metal2 3634 986 3634 986 0 net27
rlabel metal1 4048 1190 4048 1190 0 net28
rlabel metal2 4278 782 4278 782 0 net29
rlabel metal1 19458 3094 19458 3094 0 net3
rlabel metal2 4554 1020 4554 1020 0 net30
rlabel metal1 9292 1326 9292 1326 0 net31
rlabel metal1 8878 1326 8878 1326 0 net32
rlabel metal1 2070 2040 2070 2040 0 net33
rlabel metal1 1840 2074 1840 2074 0 net34
rlabel metal2 6854 2567 6854 2567 0 net35
rlabel metal2 1702 765 1702 765 0 net36
rlabel metal2 13294 1190 13294 1190 0 net37
rlabel metal2 13478 1122 13478 1122 0 net38
rlabel metal1 2530 850 2530 850 0 net39
rlabel metal1 16882 7854 16882 7854 0 net4
rlabel metal1 3174 1190 3174 1190 0 net40
rlabel metal3 18676 680 18676 680 0 net41
rlabel metal1 17342 2380 17342 2380 0 net42
rlabel metal1 8924 1734 8924 1734 0 net43
rlabel metal1 8142 1326 8142 1326 0 net44
rlabel metal2 15962 1394 15962 1394 0 net45
rlabel metal1 9664 1938 9664 1938 0 net46
rlabel metal2 16146 1054 16146 1054 0 net47
rlabel metal2 21482 1105 21482 1105 0 net48
rlabel metal3 18860 544 18860 544 0 net49
rlabel metal1 23506 2414 23506 2414 0 net5
rlabel metal2 19090 1309 19090 1309 0 net50
rlabel metal2 18446 1156 18446 1156 0 net51
rlabel metal2 17710 1462 17710 1462 0 net52
rlabel metal2 6670 1530 6670 1530 0 net53
rlabel metal1 18262 510 18262 510 0 net54
rlabel metal1 7774 1530 7774 1530 0 net55
rlabel metal2 16790 1632 16790 1632 0 net56
rlabel metal2 21850 1938 21850 1938 0 net57
rlabel via2 19826 3995 19826 3995 0 net58
rlabel metal2 14122 6086 14122 6086 0 net59
rlabel metal1 23092 2618 23092 2618 0 net6
rlabel metal1 15364 3706 15364 3706 0 net60
rlabel metal1 17158 8534 17158 8534 0 net61
rlabel metal1 17986 8500 17986 8500 0 net62
rlabel metal1 19320 8466 19320 8466 0 net63
rlabel metal1 20378 8432 20378 8432 0 net64
rlabel metal1 21804 8466 21804 8466 0 net65
rlabel metal1 23736 2074 23736 2074 0 net66
rlabel metal1 23736 2618 23736 2618 0 net67
rlabel metal1 23690 3910 23690 3910 0 net68
rlabel via2 21206 1819 21206 1819 0 net69
rlabel metal2 23184 2346 23184 2346 0 net7
rlabel metal2 21574 2023 21574 2023 0 net70
rlabel metal1 5888 2074 5888 2074 0 net71
rlabel metal2 7130 7820 7130 7820 0 net72
rlabel metal1 8188 3162 8188 3162 0 net73
rlabel metal2 9338 6188 9338 6188 0 net74
rlabel metal2 10534 6188 10534 6188 0 net75
rlabel metal2 11730 6188 11730 6188 0 net76
rlabel metal1 13064 3910 13064 3910 0 net77
rlabel metal1 7958 1904 7958 1904 0 net78
rlabel metal1 9522 1326 9522 1326 0 net79
rlabel metal1 23460 3162 23460 3162 0 net8
rlabel metal1 9844 1326 9844 1326 0 net80
rlabel metal1 10764 2006 10764 2006 0 net81
rlabel metal1 13478 1292 13478 1292 0 net82
rlabel metal1 14076 1258 14076 1258 0 net83
rlabel metal1 13892 1326 13892 1326 0 net84
rlabel metal1 14858 1904 14858 1904 0 net85
rlabel metal1 15272 1326 15272 1326 0 net86
rlabel metal1 15640 1326 15640 1326 0 net87
rlabel metal1 16790 1360 16790 1360 0 net88
rlabel metal1 15502 2040 15502 2040 0 net89
rlabel metal1 22310 2346 22310 2346 0 net9
rlabel metal1 10028 1258 10028 1258 0 net90
rlabel metal1 10212 1326 10212 1326 0 net91
rlabel metal1 11914 2040 11914 2040 0 net92
rlabel metal1 11592 1326 11592 1326 0 net93
rlabel metal1 11960 1326 11960 1326 0 net94
rlabel metal2 11730 1496 11730 1496 0 net95
rlabel metal1 12742 1972 12742 1972 0 net96
rlabel metal2 13110 1802 13110 1802 0 net97
rlabel metal2 16330 1734 16330 1734 0 net98
rlabel metal1 19780 1258 19780 1258 0 net99
<< properties >>
string FIXED_BBOX 0 0 25700 10000
<< end >>
