// This is the unpowered netlist.
module RAM_IO (Config_accessC_bit0,
    Config_accessC_bit1,
    Config_accessC_bit2,
    Config_accessC_bit3,
    FAB2RAM_A0_O0,
    FAB2RAM_A0_O1,
    FAB2RAM_A0_O2,
    FAB2RAM_A0_O3,
    FAB2RAM_A1_O0,
    FAB2RAM_A1_O1,
    FAB2RAM_A1_O2,
    FAB2RAM_A1_O3,
    FAB2RAM_C_O0,
    FAB2RAM_C_O1,
    FAB2RAM_C_O2,
    FAB2RAM_C_O3,
    FAB2RAM_D0_O0,
    FAB2RAM_D0_O1,
    FAB2RAM_D0_O2,
    FAB2RAM_D0_O3,
    FAB2RAM_D1_O0,
    FAB2RAM_D1_O1,
    FAB2RAM_D1_O2,
    FAB2RAM_D1_O3,
    FAB2RAM_D2_O0,
    FAB2RAM_D2_O1,
    FAB2RAM_D2_O2,
    FAB2RAM_D2_O3,
    FAB2RAM_D3_O0,
    FAB2RAM_D3_O1,
    FAB2RAM_D3_O2,
    FAB2RAM_D3_O3,
    RAM2FAB_D0_I0,
    RAM2FAB_D0_I1,
    RAM2FAB_D0_I2,
    RAM2FAB_D0_I3,
    RAM2FAB_D1_I0,
    RAM2FAB_D1_I1,
    RAM2FAB_D1_I2,
    RAM2FAB_D1_I3,
    RAM2FAB_D2_I0,
    RAM2FAB_D2_I1,
    RAM2FAB_D2_I2,
    RAM2FAB_D2_I3,
    RAM2FAB_D3_I0,
    RAM2FAB_D3_I1,
    RAM2FAB_D3_I2,
    RAM2FAB_D3_I3,
    UserCLK,
    UserCLKo,
    E1END,
    E2END,
    E2MID,
    E6END,
    EE4END,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1BEG,
    N1END,
    N2BEG,
    N2BEGb,
    N2END,
    N2MID,
    N4BEG,
    N4END,
    S1BEG,
    S1END,
    S2BEG,
    S2BEGb,
    S2END,
    S2MID,
    S4BEG,
    S4END,
    W1BEG,
    W2BEG,
    W2BEGb,
    W6BEG,
    WW4BEG);
 output Config_accessC_bit0;
 output Config_accessC_bit1;
 output Config_accessC_bit2;
 output Config_accessC_bit3;
 output FAB2RAM_A0_O0;
 output FAB2RAM_A0_O1;
 output FAB2RAM_A0_O2;
 output FAB2RAM_A0_O3;
 output FAB2RAM_A1_O0;
 output FAB2RAM_A1_O1;
 output FAB2RAM_A1_O2;
 output FAB2RAM_A1_O3;
 output FAB2RAM_C_O0;
 output FAB2RAM_C_O1;
 output FAB2RAM_C_O2;
 output FAB2RAM_C_O3;
 output FAB2RAM_D0_O0;
 output FAB2RAM_D0_O1;
 output FAB2RAM_D0_O2;
 output FAB2RAM_D0_O3;
 output FAB2RAM_D1_O0;
 output FAB2RAM_D1_O1;
 output FAB2RAM_D1_O2;
 output FAB2RAM_D1_O3;
 output FAB2RAM_D2_O0;
 output FAB2RAM_D2_O1;
 output FAB2RAM_D2_O2;
 output FAB2RAM_D2_O3;
 output FAB2RAM_D3_O0;
 output FAB2RAM_D3_O1;
 output FAB2RAM_D3_O2;
 output FAB2RAM_D3_O3;
 input RAM2FAB_D0_I0;
 input RAM2FAB_D0_I1;
 input RAM2FAB_D0_I2;
 input RAM2FAB_D0_I3;
 input RAM2FAB_D1_I0;
 input RAM2FAB_D1_I1;
 input RAM2FAB_D1_I2;
 input RAM2FAB_D1_I3;
 input RAM2FAB_D2_I0;
 input RAM2FAB_D2_I1;
 input RAM2FAB_D2_I2;
 input RAM2FAB_D2_I3;
 input RAM2FAB_D3_I0;
 input RAM2FAB_D3_I1;
 input RAM2FAB_D3_I2;
 input RAM2FAB_D3_I3;
 input UserCLK;
 output UserCLKo;
 input [3:0] E1END;
 input [7:0] E2END;
 input [7:0] E2MID;
 input [11:0] E6END;
 input [15:0] EE4END;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 output [3:0] N1BEG;
 input [3:0] N1END;
 output [7:0] N2BEG;
 output [7:0] N2BEGb;
 input [7:0] N2END;
 input [7:0] N2MID;
 output [15:0] N4BEG;
 input [15:0] N4END;
 output [3:0] S1BEG;
 input [3:0] S1END;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 input [7:0] S2END;
 input [7:0] S2MID;
 output [15:0] S4BEG;
 input [15:0] S4END;
 output [3:0] W1BEG;
 output [7:0] W2BEG;
 output [7:0] W2BEGb;
 output [11:0] W6BEG;
 output [15:0] WW4BEG;

 wire \ConfigBits[0] ;
 wire \ConfigBits[100] ;
 wire \ConfigBits[101] ;
 wire \ConfigBits[102] ;
 wire \ConfigBits[103] ;
 wire \ConfigBits[104] ;
 wire \ConfigBits[105] ;
 wire \ConfigBits[106] ;
 wire \ConfigBits[107] ;
 wire \ConfigBits[108] ;
 wire \ConfigBits[109] ;
 wire \ConfigBits[10] ;
 wire \ConfigBits[110] ;
 wire \ConfigBits[111] ;
 wire \ConfigBits[112] ;
 wire \ConfigBits[113] ;
 wire \ConfigBits[114] ;
 wire \ConfigBits[115] ;
 wire \ConfigBits[116] ;
 wire \ConfigBits[117] ;
 wire \ConfigBits[118] ;
 wire \ConfigBits[119] ;
 wire \ConfigBits[11] ;
 wire \ConfigBits[120] ;
 wire \ConfigBits[121] ;
 wire \ConfigBits[122] ;
 wire \ConfigBits[123] ;
 wire \ConfigBits[124] ;
 wire \ConfigBits[125] ;
 wire \ConfigBits[126] ;
 wire \ConfigBits[127] ;
 wire \ConfigBits[128] ;
 wire \ConfigBits[129] ;
 wire \ConfigBits[12] ;
 wire \ConfigBits[130] ;
 wire \ConfigBits[131] ;
 wire \ConfigBits[132] ;
 wire \ConfigBits[133] ;
 wire \ConfigBits[134] ;
 wire \ConfigBits[135] ;
 wire \ConfigBits[136] ;
 wire \ConfigBits[137] ;
 wire \ConfigBits[138] ;
 wire \ConfigBits[139] ;
 wire \ConfigBits[13] ;
 wire \ConfigBits[140] ;
 wire \ConfigBits[141] ;
 wire \ConfigBits[142] ;
 wire \ConfigBits[143] ;
 wire \ConfigBits[144] ;
 wire \ConfigBits[145] ;
 wire \ConfigBits[146] ;
 wire \ConfigBits[147] ;
 wire \ConfigBits[148] ;
 wire \ConfigBits[149] ;
 wire \ConfigBits[14] ;
 wire \ConfigBits[150] ;
 wire \ConfigBits[151] ;
 wire \ConfigBits[152] ;
 wire \ConfigBits[153] ;
 wire \ConfigBits[154] ;
 wire \ConfigBits[155] ;
 wire \ConfigBits[156] ;
 wire \ConfigBits[157] ;
 wire \ConfigBits[158] ;
 wire \ConfigBits[159] ;
 wire \ConfigBits[15] ;
 wire \ConfigBits[160] ;
 wire \ConfigBits[161] ;
 wire \ConfigBits[162] ;
 wire \ConfigBits[163] ;
 wire \ConfigBits[164] ;
 wire \ConfigBits[165] ;
 wire \ConfigBits[166] ;
 wire \ConfigBits[167] ;
 wire \ConfigBits[168] ;
 wire \ConfigBits[169] ;
 wire \ConfigBits[16] ;
 wire \ConfigBits[170] ;
 wire \ConfigBits[171] ;
 wire \ConfigBits[172] ;
 wire \ConfigBits[173] ;
 wire \ConfigBits[174] ;
 wire \ConfigBits[175] ;
 wire \ConfigBits[176] ;
 wire \ConfigBits[177] ;
 wire \ConfigBits[178] ;
 wire \ConfigBits[179] ;
 wire \ConfigBits[17] ;
 wire \ConfigBits[180] ;
 wire \ConfigBits[181] ;
 wire \ConfigBits[182] ;
 wire \ConfigBits[183] ;
 wire \ConfigBits[184] ;
 wire \ConfigBits[185] ;
 wire \ConfigBits[186] ;
 wire \ConfigBits[187] ;
 wire \ConfigBits[188] ;
 wire \ConfigBits[189] ;
 wire \ConfigBits[18] ;
 wire \ConfigBits[190] ;
 wire \ConfigBits[191] ;
 wire \ConfigBits[192] ;
 wire \ConfigBits[193] ;
 wire \ConfigBits[194] ;
 wire \ConfigBits[195] ;
 wire \ConfigBits[196] ;
 wire \ConfigBits[197] ;
 wire \ConfigBits[198] ;
 wire \ConfigBits[199] ;
 wire \ConfigBits[19] ;
 wire \ConfigBits[1] ;
 wire \ConfigBits[200] ;
 wire \ConfigBits[201] ;
 wire \ConfigBits[202] ;
 wire \ConfigBits[203] ;
 wire \ConfigBits[204] ;
 wire \ConfigBits[205] ;
 wire \ConfigBits[206] ;
 wire \ConfigBits[207] ;
 wire \ConfigBits[208] ;
 wire \ConfigBits[209] ;
 wire \ConfigBits[20] ;
 wire \ConfigBits[210] ;
 wire \ConfigBits[211] ;
 wire \ConfigBits[212] ;
 wire \ConfigBits[213] ;
 wire \ConfigBits[214] ;
 wire \ConfigBits[215] ;
 wire \ConfigBits[216] ;
 wire \ConfigBits[217] ;
 wire \ConfigBits[218] ;
 wire \ConfigBits[219] ;
 wire \ConfigBits[21] ;
 wire \ConfigBits[220] ;
 wire \ConfigBits[221] ;
 wire \ConfigBits[222] ;
 wire \ConfigBits[223] ;
 wire \ConfigBits[224] ;
 wire \ConfigBits[225] ;
 wire \ConfigBits[226] ;
 wire \ConfigBits[227] ;
 wire \ConfigBits[228] ;
 wire \ConfigBits[229] ;
 wire \ConfigBits[22] ;
 wire \ConfigBits[230] ;
 wire \ConfigBits[231] ;
 wire \ConfigBits[232] ;
 wire \ConfigBits[233] ;
 wire \ConfigBits[234] ;
 wire \ConfigBits[235] ;
 wire \ConfigBits[236] ;
 wire \ConfigBits[237] ;
 wire \ConfigBits[238] ;
 wire \ConfigBits[239] ;
 wire \ConfigBits[23] ;
 wire \ConfigBits[240] ;
 wire \ConfigBits[241] ;
 wire \ConfigBits[242] ;
 wire \ConfigBits[243] ;
 wire \ConfigBits[244] ;
 wire \ConfigBits[245] ;
 wire \ConfigBits[246] ;
 wire \ConfigBits[247] ;
 wire \ConfigBits[248] ;
 wire \ConfigBits[249] ;
 wire \ConfigBits[24] ;
 wire \ConfigBits[250] ;
 wire \ConfigBits[251] ;
 wire \ConfigBits[252] ;
 wire \ConfigBits[253] ;
 wire \ConfigBits[254] ;
 wire \ConfigBits[255] ;
 wire \ConfigBits[256] ;
 wire \ConfigBits[257] ;
 wire \ConfigBits[258] ;
 wire \ConfigBits[259] ;
 wire \ConfigBits[25] ;
 wire \ConfigBits[260] ;
 wire \ConfigBits[261] ;
 wire \ConfigBits[262] ;
 wire \ConfigBits[263] ;
 wire \ConfigBits[264] ;
 wire \ConfigBits[265] ;
 wire \ConfigBits[266] ;
 wire \ConfigBits[267] ;
 wire \ConfigBits[268] ;
 wire \ConfigBits[269] ;
 wire \ConfigBits[26] ;
 wire \ConfigBits[270] ;
 wire \ConfigBits[271] ;
 wire \ConfigBits[272] ;
 wire \ConfigBits[273] ;
 wire \ConfigBits[274] ;
 wire \ConfigBits[275] ;
 wire \ConfigBits[276] ;
 wire \ConfigBits[277] ;
 wire \ConfigBits[278] ;
 wire \ConfigBits[279] ;
 wire \ConfigBits[27] ;
 wire \ConfigBits[280] ;
 wire \ConfigBits[281] ;
 wire \ConfigBits[282] ;
 wire \ConfigBits[283] ;
 wire \ConfigBits[284] ;
 wire \ConfigBits[285] ;
 wire \ConfigBits[286] ;
 wire \ConfigBits[287] ;
 wire \ConfigBits[288] ;
 wire \ConfigBits[289] ;
 wire \ConfigBits[28] ;
 wire \ConfigBits[290] ;
 wire \ConfigBits[291] ;
 wire \ConfigBits[292] ;
 wire \ConfigBits[293] ;
 wire \ConfigBits[294] ;
 wire \ConfigBits[295] ;
 wire \ConfigBits[296] ;
 wire \ConfigBits[297] ;
 wire \ConfigBits[298] ;
 wire \ConfigBits[299] ;
 wire \ConfigBits[29] ;
 wire \ConfigBits[2] ;
 wire \ConfigBits[300] ;
 wire \ConfigBits[301] ;
 wire \ConfigBits[302] ;
 wire \ConfigBits[303] ;
 wire \ConfigBits[304] ;
 wire \ConfigBits[305] ;
 wire \ConfigBits[306] ;
 wire \ConfigBits[307] ;
 wire \ConfigBits[308] ;
 wire \ConfigBits[309] ;
 wire \ConfigBits[30] ;
 wire \ConfigBits[310] ;
 wire \ConfigBits[311] ;
 wire \ConfigBits[312] ;
 wire \ConfigBits[313] ;
 wire \ConfigBits[314] ;
 wire \ConfigBits[315] ;
 wire \ConfigBits[316] ;
 wire \ConfigBits[317] ;
 wire \ConfigBits[318] ;
 wire \ConfigBits[319] ;
 wire \ConfigBits[31] ;
 wire \ConfigBits[320] ;
 wire \ConfigBits[321] ;
 wire \ConfigBits[322] ;
 wire \ConfigBits[323] ;
 wire \ConfigBits[324] ;
 wire \ConfigBits[325] ;
 wire \ConfigBits[326] ;
 wire \ConfigBits[327] ;
 wire \ConfigBits[32] ;
 wire \ConfigBits[33] ;
 wire \ConfigBits[34] ;
 wire \ConfigBits[35] ;
 wire \ConfigBits[36] ;
 wire \ConfigBits[37] ;
 wire \ConfigBits[38] ;
 wire \ConfigBits[39] ;
 wire \ConfigBits[3] ;
 wire \ConfigBits[40] ;
 wire \ConfigBits[41] ;
 wire \ConfigBits[42] ;
 wire \ConfigBits[43] ;
 wire \ConfigBits[44] ;
 wire \ConfigBits[45] ;
 wire \ConfigBits[46] ;
 wire \ConfigBits[47] ;
 wire \ConfigBits[48] ;
 wire \ConfigBits[49] ;
 wire \ConfigBits[4] ;
 wire \ConfigBits[50] ;
 wire \ConfigBits[51] ;
 wire \ConfigBits[52] ;
 wire \ConfigBits[53] ;
 wire \ConfigBits[54] ;
 wire \ConfigBits[55] ;
 wire \ConfigBits[56] ;
 wire \ConfigBits[57] ;
 wire \ConfigBits[58] ;
 wire \ConfigBits[59] ;
 wire \ConfigBits[5] ;
 wire \ConfigBits[60] ;
 wire \ConfigBits[61] ;
 wire \ConfigBits[62] ;
 wire \ConfigBits[63] ;
 wire \ConfigBits[64] ;
 wire \ConfigBits[65] ;
 wire \ConfigBits[66] ;
 wire \ConfigBits[67] ;
 wire \ConfigBits[68] ;
 wire \ConfigBits[69] ;
 wire \ConfigBits[6] ;
 wire \ConfigBits[70] ;
 wire \ConfigBits[71] ;
 wire \ConfigBits[72] ;
 wire \ConfigBits[73] ;
 wire \ConfigBits[74] ;
 wire \ConfigBits[75] ;
 wire \ConfigBits[76] ;
 wire \ConfigBits[77] ;
 wire \ConfigBits[78] ;
 wire \ConfigBits[79] ;
 wire \ConfigBits[7] ;
 wire \ConfigBits[80] ;
 wire \ConfigBits[81] ;
 wire \ConfigBits[82] ;
 wire \ConfigBits[83] ;
 wire \ConfigBits[84] ;
 wire \ConfigBits[85] ;
 wire \ConfigBits[86] ;
 wire \ConfigBits[87] ;
 wire \ConfigBits[88] ;
 wire \ConfigBits[89] ;
 wire \ConfigBits[8] ;
 wire \ConfigBits[90] ;
 wire \ConfigBits[91] ;
 wire \ConfigBits[92] ;
 wire \ConfigBits[93] ;
 wire \ConfigBits[94] ;
 wire \ConfigBits[95] ;
 wire \ConfigBits[96] ;
 wire \ConfigBits[97] ;
 wire \ConfigBits[98] ;
 wire \ConfigBits[99] ;
 wire \ConfigBits[9] ;
 wire \ConfigBits_N[0] ;
 wire \ConfigBits_N[100] ;
 wire \ConfigBits_N[101] ;
 wire \ConfigBits_N[102] ;
 wire \ConfigBits_N[103] ;
 wire \ConfigBits_N[104] ;
 wire \ConfigBits_N[105] ;
 wire \ConfigBits_N[106] ;
 wire \ConfigBits_N[107] ;
 wire \ConfigBits_N[108] ;
 wire \ConfigBits_N[109] ;
 wire \ConfigBits_N[10] ;
 wire \ConfigBits_N[110] ;
 wire \ConfigBits_N[111] ;
 wire \ConfigBits_N[112] ;
 wire \ConfigBits_N[113] ;
 wire \ConfigBits_N[114] ;
 wire \ConfigBits_N[115] ;
 wire \ConfigBits_N[116] ;
 wire \ConfigBits_N[117] ;
 wire \ConfigBits_N[118] ;
 wire \ConfigBits_N[119] ;
 wire \ConfigBits_N[11] ;
 wire \ConfigBits_N[120] ;
 wire \ConfigBits_N[121] ;
 wire \ConfigBits_N[122] ;
 wire \ConfigBits_N[123] ;
 wire \ConfigBits_N[124] ;
 wire \ConfigBits_N[125] ;
 wire \ConfigBits_N[126] ;
 wire \ConfigBits_N[127] ;
 wire \ConfigBits_N[128] ;
 wire \ConfigBits_N[129] ;
 wire \ConfigBits_N[12] ;
 wire \ConfigBits_N[130] ;
 wire \ConfigBits_N[131] ;
 wire \ConfigBits_N[132] ;
 wire \ConfigBits_N[133] ;
 wire \ConfigBits_N[134] ;
 wire \ConfigBits_N[135] ;
 wire \ConfigBits_N[136] ;
 wire \ConfigBits_N[137] ;
 wire \ConfigBits_N[138] ;
 wire \ConfigBits_N[139] ;
 wire \ConfigBits_N[13] ;
 wire \ConfigBits_N[140] ;
 wire \ConfigBits_N[141] ;
 wire \ConfigBits_N[142] ;
 wire \ConfigBits_N[143] ;
 wire \ConfigBits_N[144] ;
 wire \ConfigBits_N[145] ;
 wire \ConfigBits_N[146] ;
 wire \ConfigBits_N[147] ;
 wire \ConfigBits_N[148] ;
 wire \ConfigBits_N[149] ;
 wire \ConfigBits_N[14] ;
 wire \ConfigBits_N[150] ;
 wire \ConfigBits_N[151] ;
 wire \ConfigBits_N[152] ;
 wire \ConfigBits_N[153] ;
 wire \ConfigBits_N[154] ;
 wire \ConfigBits_N[155] ;
 wire \ConfigBits_N[156] ;
 wire \ConfigBits_N[157] ;
 wire \ConfigBits_N[158] ;
 wire \ConfigBits_N[159] ;
 wire \ConfigBits_N[15] ;
 wire \ConfigBits_N[160] ;
 wire \ConfigBits_N[161] ;
 wire \ConfigBits_N[162] ;
 wire \ConfigBits_N[163] ;
 wire \ConfigBits_N[164] ;
 wire \ConfigBits_N[165] ;
 wire \ConfigBits_N[166] ;
 wire \ConfigBits_N[167] ;
 wire \ConfigBits_N[168] ;
 wire \ConfigBits_N[169] ;
 wire \ConfigBits_N[16] ;
 wire \ConfigBits_N[170] ;
 wire \ConfigBits_N[171] ;
 wire \ConfigBits_N[172] ;
 wire \ConfigBits_N[173] ;
 wire \ConfigBits_N[174] ;
 wire \ConfigBits_N[175] ;
 wire \ConfigBits_N[176] ;
 wire \ConfigBits_N[177] ;
 wire \ConfigBits_N[178] ;
 wire \ConfigBits_N[179] ;
 wire \ConfigBits_N[17] ;
 wire \ConfigBits_N[180] ;
 wire \ConfigBits_N[181] ;
 wire \ConfigBits_N[182] ;
 wire \ConfigBits_N[183] ;
 wire \ConfigBits_N[184] ;
 wire \ConfigBits_N[185] ;
 wire \ConfigBits_N[186] ;
 wire \ConfigBits_N[187] ;
 wire \ConfigBits_N[188] ;
 wire \ConfigBits_N[189] ;
 wire \ConfigBits_N[18] ;
 wire \ConfigBits_N[190] ;
 wire \ConfigBits_N[191] ;
 wire \ConfigBits_N[192] ;
 wire \ConfigBits_N[193] ;
 wire \ConfigBits_N[194] ;
 wire \ConfigBits_N[195] ;
 wire \ConfigBits_N[196] ;
 wire \ConfigBits_N[197] ;
 wire \ConfigBits_N[198] ;
 wire \ConfigBits_N[199] ;
 wire \ConfigBits_N[19] ;
 wire \ConfigBits_N[1] ;
 wire \ConfigBits_N[200] ;
 wire \ConfigBits_N[201] ;
 wire \ConfigBits_N[202] ;
 wire \ConfigBits_N[203] ;
 wire \ConfigBits_N[204] ;
 wire \ConfigBits_N[205] ;
 wire \ConfigBits_N[206] ;
 wire \ConfigBits_N[207] ;
 wire \ConfigBits_N[208] ;
 wire \ConfigBits_N[209] ;
 wire \ConfigBits_N[20] ;
 wire \ConfigBits_N[210] ;
 wire \ConfigBits_N[211] ;
 wire \ConfigBits_N[212] ;
 wire \ConfigBits_N[213] ;
 wire \ConfigBits_N[214] ;
 wire \ConfigBits_N[215] ;
 wire \ConfigBits_N[216] ;
 wire \ConfigBits_N[217] ;
 wire \ConfigBits_N[218] ;
 wire \ConfigBits_N[219] ;
 wire \ConfigBits_N[21] ;
 wire \ConfigBits_N[220] ;
 wire \ConfigBits_N[221] ;
 wire \ConfigBits_N[222] ;
 wire \ConfigBits_N[223] ;
 wire \ConfigBits_N[224] ;
 wire \ConfigBits_N[225] ;
 wire \ConfigBits_N[226] ;
 wire \ConfigBits_N[227] ;
 wire \ConfigBits_N[228] ;
 wire \ConfigBits_N[229] ;
 wire \ConfigBits_N[22] ;
 wire \ConfigBits_N[230] ;
 wire \ConfigBits_N[231] ;
 wire \ConfigBits_N[232] ;
 wire \ConfigBits_N[233] ;
 wire \ConfigBits_N[234] ;
 wire \ConfigBits_N[235] ;
 wire \ConfigBits_N[236] ;
 wire \ConfigBits_N[237] ;
 wire \ConfigBits_N[238] ;
 wire \ConfigBits_N[239] ;
 wire \ConfigBits_N[23] ;
 wire \ConfigBits_N[240] ;
 wire \ConfigBits_N[241] ;
 wire \ConfigBits_N[242] ;
 wire \ConfigBits_N[243] ;
 wire \ConfigBits_N[244] ;
 wire \ConfigBits_N[245] ;
 wire \ConfigBits_N[246] ;
 wire \ConfigBits_N[247] ;
 wire \ConfigBits_N[248] ;
 wire \ConfigBits_N[249] ;
 wire \ConfigBits_N[24] ;
 wire \ConfigBits_N[250] ;
 wire \ConfigBits_N[251] ;
 wire \ConfigBits_N[252] ;
 wire \ConfigBits_N[253] ;
 wire \ConfigBits_N[254] ;
 wire \ConfigBits_N[255] ;
 wire \ConfigBits_N[256] ;
 wire \ConfigBits_N[257] ;
 wire \ConfigBits_N[258] ;
 wire \ConfigBits_N[259] ;
 wire \ConfigBits_N[25] ;
 wire \ConfigBits_N[260] ;
 wire \ConfigBits_N[261] ;
 wire \ConfigBits_N[262] ;
 wire \ConfigBits_N[263] ;
 wire \ConfigBits_N[264] ;
 wire \ConfigBits_N[265] ;
 wire \ConfigBits_N[266] ;
 wire \ConfigBits_N[267] ;
 wire \ConfigBits_N[268] ;
 wire \ConfigBits_N[269] ;
 wire \ConfigBits_N[26] ;
 wire \ConfigBits_N[270] ;
 wire \ConfigBits_N[271] ;
 wire \ConfigBits_N[272] ;
 wire \ConfigBits_N[273] ;
 wire \ConfigBits_N[274] ;
 wire \ConfigBits_N[275] ;
 wire \ConfigBits_N[276] ;
 wire \ConfigBits_N[277] ;
 wire \ConfigBits_N[278] ;
 wire \ConfigBits_N[279] ;
 wire \ConfigBits_N[27] ;
 wire \ConfigBits_N[280] ;
 wire \ConfigBits_N[281] ;
 wire \ConfigBits_N[282] ;
 wire \ConfigBits_N[283] ;
 wire \ConfigBits_N[284] ;
 wire \ConfigBits_N[285] ;
 wire \ConfigBits_N[286] ;
 wire \ConfigBits_N[287] ;
 wire \ConfigBits_N[288] ;
 wire \ConfigBits_N[289] ;
 wire \ConfigBits_N[28] ;
 wire \ConfigBits_N[290] ;
 wire \ConfigBits_N[291] ;
 wire \ConfigBits_N[292] ;
 wire \ConfigBits_N[293] ;
 wire \ConfigBits_N[294] ;
 wire \ConfigBits_N[295] ;
 wire \ConfigBits_N[296] ;
 wire \ConfigBits_N[297] ;
 wire \ConfigBits_N[298] ;
 wire \ConfigBits_N[299] ;
 wire \ConfigBits_N[29] ;
 wire \ConfigBits_N[2] ;
 wire \ConfigBits_N[300] ;
 wire \ConfigBits_N[301] ;
 wire \ConfigBits_N[302] ;
 wire \ConfigBits_N[303] ;
 wire \ConfigBits_N[304] ;
 wire \ConfigBits_N[305] ;
 wire \ConfigBits_N[306] ;
 wire \ConfigBits_N[307] ;
 wire \ConfigBits_N[308] ;
 wire \ConfigBits_N[309] ;
 wire \ConfigBits_N[30] ;
 wire \ConfigBits_N[310] ;
 wire \ConfigBits_N[311] ;
 wire \ConfigBits_N[312] ;
 wire \ConfigBits_N[313] ;
 wire \ConfigBits_N[314] ;
 wire \ConfigBits_N[315] ;
 wire \ConfigBits_N[316] ;
 wire \ConfigBits_N[317] ;
 wire \ConfigBits_N[318] ;
 wire \ConfigBits_N[319] ;
 wire \ConfigBits_N[31] ;
 wire \ConfigBits_N[320] ;
 wire \ConfigBits_N[321] ;
 wire \ConfigBits_N[322] ;
 wire \ConfigBits_N[323] ;
 wire \ConfigBits_N[324] ;
 wire \ConfigBits_N[325] ;
 wire \ConfigBits_N[326] ;
 wire \ConfigBits_N[327] ;
 wire \ConfigBits_N[32] ;
 wire \ConfigBits_N[33] ;
 wire \ConfigBits_N[34] ;
 wire \ConfigBits_N[35] ;
 wire \ConfigBits_N[36] ;
 wire \ConfigBits_N[37] ;
 wire \ConfigBits_N[38] ;
 wire \ConfigBits_N[39] ;
 wire \ConfigBits_N[3] ;
 wire \ConfigBits_N[40] ;
 wire \ConfigBits_N[41] ;
 wire \ConfigBits_N[42] ;
 wire \ConfigBits_N[43] ;
 wire \ConfigBits_N[44] ;
 wire \ConfigBits_N[45] ;
 wire \ConfigBits_N[46] ;
 wire \ConfigBits_N[47] ;
 wire \ConfigBits_N[48] ;
 wire \ConfigBits_N[49] ;
 wire \ConfigBits_N[4] ;
 wire \ConfigBits_N[50] ;
 wire \ConfigBits_N[51] ;
 wire \ConfigBits_N[52] ;
 wire \ConfigBits_N[53] ;
 wire \ConfigBits_N[54] ;
 wire \ConfigBits_N[55] ;
 wire \ConfigBits_N[56] ;
 wire \ConfigBits_N[57] ;
 wire \ConfigBits_N[58] ;
 wire \ConfigBits_N[59] ;
 wire \ConfigBits_N[5] ;
 wire \ConfigBits_N[60] ;
 wire \ConfigBits_N[61] ;
 wire \ConfigBits_N[62] ;
 wire \ConfigBits_N[63] ;
 wire \ConfigBits_N[64] ;
 wire \ConfigBits_N[65] ;
 wire \ConfigBits_N[66] ;
 wire \ConfigBits_N[67] ;
 wire \ConfigBits_N[68] ;
 wire \ConfigBits_N[69] ;
 wire \ConfigBits_N[6] ;
 wire \ConfigBits_N[70] ;
 wire \ConfigBits_N[71] ;
 wire \ConfigBits_N[72] ;
 wire \ConfigBits_N[73] ;
 wire \ConfigBits_N[74] ;
 wire \ConfigBits_N[75] ;
 wire \ConfigBits_N[76] ;
 wire \ConfigBits_N[77] ;
 wire \ConfigBits_N[78] ;
 wire \ConfigBits_N[79] ;
 wire \ConfigBits_N[7] ;
 wire \ConfigBits_N[80] ;
 wire \ConfigBits_N[81] ;
 wire \ConfigBits_N[82] ;
 wire \ConfigBits_N[83] ;
 wire \ConfigBits_N[84] ;
 wire \ConfigBits_N[85] ;
 wire \ConfigBits_N[86] ;
 wire \ConfigBits_N[87] ;
 wire \ConfigBits_N[88] ;
 wire \ConfigBits_N[89] ;
 wire \ConfigBits_N[8] ;
 wire \ConfigBits_N[90] ;
 wire \ConfigBits_N[91] ;
 wire \ConfigBits_N[92] ;
 wire \ConfigBits_N[93] ;
 wire \ConfigBits_N[94] ;
 wire \ConfigBits_N[95] ;
 wire \ConfigBits_N[96] ;
 wire \ConfigBits_N[97] ;
 wire \ConfigBits_N[98] ;
 wire \ConfigBits_N[99] ;
 wire \ConfigBits_N[9] ;
 wire FAB2RAM_A0_I0;
 wire FAB2RAM_A0_I1;
 wire FAB2RAM_A0_I2;
 wire FAB2RAM_A0_I3;
 wire FAB2RAM_A1_I0;
 wire FAB2RAM_A1_I1;
 wire FAB2RAM_A1_I2;
 wire FAB2RAM_A1_I3;
 wire FAB2RAM_C_I0;
 wire FAB2RAM_C_I1;
 wire FAB2RAM_C_I2;
 wire FAB2RAM_C_I3;
 wire FAB2RAM_D0_I0;
 wire FAB2RAM_D0_I1;
 wire FAB2RAM_D0_I2;
 wire FAB2RAM_D0_I3;
 wire FAB2RAM_D1_I0;
 wire FAB2RAM_D1_I1;
 wire FAB2RAM_D1_I2;
 wire FAB2RAM_D1_I3;
 wire FAB2RAM_D2_I0;
 wire FAB2RAM_D2_I1;
 wire FAB2RAM_D2_I2;
 wire FAB2RAM_D2_I3;
 wire FAB2RAM_D3_I0;
 wire FAB2RAM_D3_I1;
 wire FAB2RAM_D3_I2;
 wire FAB2RAM_D3_I3;
 wire \FrameData_O_i[0] ;
 wire \FrameData_O_i[10] ;
 wire \FrameData_O_i[11] ;
 wire \FrameData_O_i[12] ;
 wire \FrameData_O_i[13] ;
 wire \FrameData_O_i[14] ;
 wire \FrameData_O_i[15] ;
 wire \FrameData_O_i[16] ;
 wire \FrameData_O_i[17] ;
 wire \FrameData_O_i[18] ;
 wire \FrameData_O_i[19] ;
 wire \FrameData_O_i[1] ;
 wire \FrameData_O_i[20] ;
 wire \FrameData_O_i[21] ;
 wire \FrameData_O_i[22] ;
 wire \FrameData_O_i[23] ;
 wire \FrameData_O_i[24] ;
 wire \FrameData_O_i[25] ;
 wire \FrameData_O_i[26] ;
 wire \FrameData_O_i[27] ;
 wire \FrameData_O_i[28] ;
 wire \FrameData_O_i[29] ;
 wire \FrameData_O_i[2] ;
 wire \FrameData_O_i[30] ;
 wire \FrameData_O_i[31] ;
 wire \FrameData_O_i[3] ;
 wire \FrameData_O_i[4] ;
 wire \FrameData_O_i[5] ;
 wire \FrameData_O_i[6] ;
 wire \FrameData_O_i[7] ;
 wire \FrameData_O_i[8] ;
 wire \FrameData_O_i[9] ;
 wire \FrameStrobe_O_i[0] ;
 wire \FrameStrobe_O_i[10] ;
 wire \FrameStrobe_O_i[11] ;
 wire \FrameStrobe_O_i[12] ;
 wire \FrameStrobe_O_i[13] ;
 wire \FrameStrobe_O_i[14] ;
 wire \FrameStrobe_O_i[15] ;
 wire \FrameStrobe_O_i[16] ;
 wire \FrameStrobe_O_i[17] ;
 wire \FrameStrobe_O_i[18] ;
 wire \FrameStrobe_O_i[19] ;
 wire \FrameStrobe_O_i[1] ;
 wire \FrameStrobe_O_i[2] ;
 wire \FrameStrobe_O_i[3] ;
 wire \FrameStrobe_O_i[4] ;
 wire \FrameStrobe_O_i[5] ;
 wire \FrameStrobe_O_i[6] ;
 wire \FrameStrobe_O_i[7] ;
 wire \FrameStrobe_O_i[8] ;
 wire \FrameStrobe_O_i[9] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[2] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[3] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[2] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[3] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[2] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[3] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[2] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[3] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[2] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[3] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[2] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[3] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[2] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[3] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[2] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[3] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[2] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[3] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[2] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[3] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[2] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[3] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ;
 wire \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_0_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_0_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_0_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_0_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_out1 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_0_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_out0 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_out1 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_0_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_out0 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_out1 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_0_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_out0 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_out1 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/AIN[0] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/AIN[1] ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_0_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_1_ ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_out0 ;
 wire \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_out1 ;
 wire \J_NS1_BEG[0] ;
 wire \J_NS1_BEG[1] ;
 wire \J_NS1_BEG[2] ;
 wire \J_NS1_BEG[3] ;
 wire \J_NS2_BEG[0] ;
 wire \J_NS2_BEG[1] ;
 wire \J_NS2_BEG[2] ;
 wire \J_NS2_BEG[3] ;
 wire \J_NS2_BEG[4] ;
 wire \J_NS2_BEG[5] ;
 wire \J_NS2_BEG[6] ;
 wire \J_NS2_BEG[7] ;
 wire \J_NS4_BEG[0] ;
 wire \J_NS4_BEG[10] ;
 wire \J_NS4_BEG[11] ;
 wire \J_NS4_BEG[12] ;
 wire \J_NS4_BEG[13] ;
 wire \J_NS4_BEG[14] ;
 wire \J_NS4_BEG[15] ;
 wire \J_NS4_BEG[1] ;
 wire \J_NS4_BEG[2] ;
 wire \J_NS4_BEG[3] ;
 wire \J_NS4_BEG[4] ;
 wire \J_NS4_BEG[5] ;
 wire \J_NS4_BEG[6] ;
 wire \J_NS4_BEG[7] ;
 wire \J_NS4_BEG[8] ;
 wire \J_NS4_BEG[9] ;
 wire \N4BEG_i[0] ;
 wire \N4BEG_i[10] ;
 wire \N4BEG_i[11] ;
 wire \N4BEG_i[1] ;
 wire \N4BEG_i[2] ;
 wire \N4BEG_i[3] ;
 wire \N4BEG_i[4] ;
 wire \N4BEG_i[5] ;
 wire \N4BEG_i[6] ;
 wire \N4BEG_i[7] ;
 wire \N4BEG_i[8] ;
 wire \N4BEG_i[9] ;
 wire RAM2FAB_D0_O0;
 wire RAM2FAB_D0_O1;
 wire RAM2FAB_D0_O2;
 wire RAM2FAB_D0_O3;
 wire RAM2FAB_D1_O0;
 wire RAM2FAB_D1_O1;
 wire RAM2FAB_D1_O2;
 wire RAM2FAB_D1_O3;
 wire RAM2FAB_D2_O0;
 wire RAM2FAB_D2_O1;
 wire RAM2FAB_D2_O2;
 wire RAM2FAB_D2_O3;
 wire RAM2FAB_D3_O0;
 wire RAM2FAB_D3_O1;
 wire RAM2FAB_D3_O2;
 wire RAM2FAB_D3_O3;
 wire \S4BEG_i[0] ;
 wire \S4BEG_i[10] ;
 wire \S4BEG_i[11] ;
 wire \S4BEG_i[1] ;
 wire \S4BEG_i[2] ;
 wire \S4BEG_i[3] ;
 wire \S4BEG_i[4] ;
 wire \S4BEG_i[5] ;
 wire \S4BEG_i[6] ;
 wire \S4BEG_i[7] ;
 wire \S4BEG_i[8] ;
 wire \S4BEG_i[9] ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(\N4BEG_i[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(\S4BEG_i[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\N4BEG_i[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\S4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(RAM2FAB_D3_O2));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(RAM2FAB_D3_O2));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\S4BEG_i[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(net106));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_112 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_198 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_34 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_90 ();
 sky130_fd_sc_hd__clkbuf_1 \Inst_Config_accessConfig_access/_0_  (.A(\ConfigBits[44] ),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 \Inst_Config_accessConfig_access/_1_  (.A(\ConfigBits[45] ),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 \Inst_Config_accessConfig_access/_2_  (.A(\ConfigBits[46] ),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 \Inst_Config_accessConfig_access/_3_  (.A(\ConfigBits[47] ),
    .X(net192));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(FAB2RAM_A0_I0),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(FAB2RAM_A0_I1),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(FAB2RAM_A0_I2),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(FAB2RAM_A0_I3),
    .Q(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[32] ),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[32] ),
    .A2(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(net193));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(FAB2RAM_A0_I0),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[0] ),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[33] ),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[33] ),
    .A2(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(net194));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(FAB2RAM_A0_I1),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[1] ),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[34] ),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[34] ),
    .A2(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(net195));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(FAB2RAM_A0_I2),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[2] ),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[35] ),
    .Y(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[35] ),
    .A2(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(net196));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(FAB2RAM_A0_I3),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q[3] ),
    .X(\Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(FAB2RAM_A1_I0),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(FAB2RAM_A1_I1),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(FAB2RAM_A1_I2),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(FAB2RAM_A1_I3),
    .Q(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[36] ),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[36] ),
    .A2(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(net197));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(FAB2RAM_A1_I0),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[0] ),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[37] ),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[37] ),
    .A2(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(net198));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(FAB2RAM_A1_I1),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[1] ),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[38] ),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[38] ),
    .A2(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(net199));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(FAB2RAM_A1_I2),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[2] ),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[39] ),
    .Y(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[39] ),
    .A2(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(net200));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(FAB2RAM_A1_I3),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q[3] ),
    .X(\Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(FAB2RAM_C_I0),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(FAB2RAM_C_I1),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(FAB2RAM_C_I2),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(FAB2RAM_C_I3),
    .Q(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[40] ),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[40] ),
    .A2(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(net201));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(FAB2RAM_C_I0),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[0] ),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[41] ),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[41] ),
    .A2(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(net202));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(FAB2RAM_C_I1),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[1] ),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[42] ),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[42] ),
    .A2(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(net203));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(FAB2RAM_C_I2),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[2] ),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[43] ),
    .Y(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[43] ),
    .A2(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(net204));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(FAB2RAM_C_I3),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q[3] ),
    .X(\Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(FAB2RAM_D0_I0),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(FAB2RAM_D0_I1),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(FAB2RAM_D0_I2),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(FAB2RAM_D0_I3),
    .Q(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[16] ),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[16] ),
    .A2(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(net205));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D0_I0),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[0] ),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[17] ),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[17] ),
    .A2(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(net206));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D0_I1),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[1] ),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[18] ),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[18] ),
    .A2(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(net207));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D0_I2),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[2] ),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[19] ),
    .Y(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[19] ),
    .A2(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(net208));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D0_I3),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q[3] ),
    .X(\Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(FAB2RAM_D1_I0),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(FAB2RAM_D1_I1),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(FAB2RAM_D1_I2),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(FAB2RAM_D1_I3),
    .Q(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[20] ),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[20] ),
    .A2(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(net209));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D1_I0),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[0] ),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[21] ),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[21] ),
    .A2(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(net210));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D1_I1),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[1] ),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[22] ),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[22] ),
    .A2(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(net211));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D1_I2),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[2] ),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[23] ),
    .Y(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[23] ),
    .A2(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(net212));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D1_I3),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q[3] ),
    .X(\Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(FAB2RAM_D2_I0),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(FAB2RAM_D2_I1),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(FAB2RAM_D2_I2),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(FAB2RAM_D2_I3),
    .Q(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[24] ),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[24] ),
    .A2(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(net213));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D2_I0),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[0] ),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[25] ),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[25] ),
    .A2(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(net214));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D2_I1),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[1] ),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[26] ),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[26] ),
    .A2(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(net215));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D2_I2),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[2] ),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[27] ),
    .Y(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[27] ),
    .A2(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(net216));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D2_I3),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q[3] ),
    .X(\Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(FAB2RAM_D3_I0),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(FAB2RAM_D3_I1),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(FAB2RAM_D3_I2),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(FAB2RAM_D3_I3),
    .Q(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[28] ),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[28] ),
    .A2(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(net217));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D3_I0),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[0] ),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[29] ),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[29] ),
    .A2(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(net218));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D3_I1),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[1] ),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[30] ),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[30] ),
    .A2(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(net219));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D3_I2),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[2] ),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[31] ),
    .Y(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[31] ),
    .A2(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(net220));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(FAB2RAM_D3_I3),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q[3] ),
    .X(\Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(net137),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(net138),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(net139),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(net140),
    .Q(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[0] ),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[0] ),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(RAM2FAB_D0_O0));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(net137),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[0] ),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[1] ),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[1] ),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(RAM2FAB_D0_O1));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(net138),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[1] ),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[2] ),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[2] ),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(RAM2FAB_D0_O2));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(net139),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[2] ),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[3] ),
    .Y(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[3] ),
    .A2(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(RAM2FAB_D0_O3));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(net140),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q[3] ),
    .X(\Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(net141),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(net142),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(net143),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(net144),
    .Q(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[4] ),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[4] ),
    .A2(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(RAM2FAB_D1_O0));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(net141),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[0] ),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[5] ),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[5] ),
    .A2(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(RAM2FAB_D1_O1));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(net142),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[1] ),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[6] ),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[6] ),
    .A2(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(RAM2FAB_D1_O2));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(net143),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[2] ),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[7] ),
    .Y(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[7] ),
    .A2(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(RAM2FAB_D1_O3));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(net144),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q[3] ),
    .X(\Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(net145),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(net146),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(net147),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(net148),
    .Q(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[8] ),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[8] ),
    .A2(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(RAM2FAB_D2_O0));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(net145),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[0] ),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[9] ),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[9] ),
    .A2(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(RAM2FAB_D2_O1));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(net146),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[1] ),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[10] ),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[10] ),
    .A2(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(RAM2FAB_D2_O2));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(net147),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[2] ),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[11] ),
    .Y(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[11] ),
    .A2(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(RAM2FAB_D2_O3));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(net148),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q[3] ),
    .X(\Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/_0_  (.CLK(UserCLK),
    .D(net149),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[0] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/_1_  (.CLK(UserCLK),
    .D(net150),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[1] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/_2_  (.CLK(UserCLK),
    .D(net151),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[2] ));
 sky130_fd_sc_hd__dfxtp_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/_3_  (.CLK(UserCLK),
    .D(net152),
    .Q(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[3] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_2_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_3_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ),
    .B(\ConfigBits[12] ),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_4_  (.A1(\ConfigBits[12] ),
    .A2(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_0_ ),
    .B1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_1_ ),
    .Y(RAM2FAB_D3_O0));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst0/_0_  (.A(net149),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[0] ),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_2_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_3_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ),
    .B(\ConfigBits[13] ),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_4_  (.A1(\ConfigBits[13] ),
    .A2(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_0_ ),
    .B1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_1_ ),
    .Y(RAM2FAB_D3_O1));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst0/_0_  (.A(net150),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[1] ),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_2_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_3_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ),
    .B(\ConfigBits[14] ),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ));
 sky130_fd_sc_hd__o21ai_4 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_4_  (.A1(\ConfigBits[14] ),
    .A2(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_0_ ),
    .B1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_1_ ),
    .Y(RAM2FAB_D3_O2));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst0/_0_  (.A(net151),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[2] ),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/AIN[1] ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_2_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_3_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ),
    .B(\ConfigBits[15] ),
    .Y(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_4_  (.A1(\ConfigBits[15] ),
    .A2(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_0_ ),
    .B1(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_1_ ),
    .Y(RAM2FAB_D3_O3));
 sky130_fd_sc_hd__buf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst0/_0_  (.A(net152),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/break_comb_loop_inst1/_0_  (.A(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q[3] ),
    .X(\Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/AIN[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit0  (.D(net49),
    .GATE(net81),
    .Q(\ConfigBits[296] ),
    .Q_N(\ConfigBits_N[296] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit1  (.D(net60),
    .GATE(net81),
    .Q(\ConfigBits[297] ),
    .Q_N(\ConfigBits_N[297] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit10  (.D(net50),
    .GATE(net81),
    .Q(\ConfigBits[306] ),
    .Q_N(\ConfigBits_N[306] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit11  (.D(net51),
    .GATE(net81),
    .Q(\ConfigBits[307] ),
    .Q_N(\ConfigBits_N[307] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit12  (.D(net52),
    .GATE(net81),
    .Q(\ConfigBits[308] ),
    .Q_N(\ConfigBits_N[308] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit13  (.D(net53),
    .GATE(net81),
    .Q(\ConfigBits[309] ),
    .Q_N(\ConfigBits_N[309] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit14  (.D(net54),
    .GATE(net81),
    .Q(\ConfigBits[310] ),
    .Q_N(\ConfigBits_N[310] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit15  (.D(net55),
    .GATE(net81),
    .Q(\ConfigBits[311] ),
    .Q_N(\ConfigBits_N[311] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit16  (.D(net56),
    .GATE(net81),
    .Q(\ConfigBits[312] ),
    .Q_N(\ConfigBits_N[312] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit17  (.D(net57),
    .GATE(net81),
    .Q(\ConfigBits[313] ),
    .Q_N(\ConfigBits_N[313] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit18  (.D(net58),
    .GATE(net81),
    .Q(\ConfigBits[314] ),
    .Q_N(\ConfigBits_N[314] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit19  (.D(net59),
    .GATE(net81),
    .Q(\ConfigBits[315] ),
    .Q_N(\ConfigBits_N[315] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit2  (.D(net71),
    .GATE(net81),
    .Q(\ConfigBits[298] ),
    .Q_N(\ConfigBits_N[298] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit20  (.D(net61),
    .GATE(net81),
    .Q(\ConfigBits[316] ),
    .Q_N(\ConfigBits_N[316] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit21  (.D(net62),
    .GATE(net81),
    .Q(\ConfigBits[317] ),
    .Q_N(\ConfigBits_N[317] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit22  (.D(net63),
    .GATE(net81),
    .Q(\ConfigBits[318] ),
    .Q_N(\ConfigBits_N[318] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit23  (.D(net64),
    .GATE(net81),
    .Q(\ConfigBits[319] ),
    .Q_N(\ConfigBits_N[319] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit24  (.D(net65),
    .GATE(net81),
    .Q(\ConfigBits[320] ),
    .Q_N(\ConfigBits_N[320] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit25  (.D(net66),
    .GATE(net81),
    .Q(\ConfigBits[321] ),
    .Q_N(\ConfigBits_N[321] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit26  (.D(net67),
    .GATE(net81),
    .Q(\ConfigBits[322] ),
    .Q_N(\ConfigBits_N[322] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit27  (.D(net68),
    .GATE(net81),
    .Q(\ConfigBits[323] ),
    .Q_N(\ConfigBits_N[323] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit28  (.D(net69),
    .GATE(net81),
    .Q(\ConfigBits[324] ),
    .Q_N(\ConfigBits_N[324] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit29  (.D(net70),
    .GATE(net81),
    .Q(\ConfigBits[325] ),
    .Q_N(\ConfigBits_N[325] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit3  (.D(net74),
    .GATE(net81),
    .Q(\ConfigBits[299] ),
    .Q_N(\ConfigBits_N[299] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit30  (.D(net72),
    .GATE(net81),
    .Q(\ConfigBits[326] ),
    .Q_N(\ConfigBits_N[326] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit31  (.D(net73),
    .GATE(net81),
    .Q(\ConfigBits[327] ),
    .Q_N(\ConfigBits_N[327] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit4  (.D(net75),
    .GATE(net81),
    .Q(\ConfigBits[300] ),
    .Q_N(\ConfigBits_N[300] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit5  (.D(net76),
    .GATE(net81),
    .Q(\ConfigBits[301] ),
    .Q_N(\ConfigBits_N[301] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit6  (.D(net77),
    .GATE(net81),
    .Q(\ConfigBits[302] ),
    .Q_N(\ConfigBits_N[302] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit7  (.D(net78),
    .GATE(net81),
    .Q(\ConfigBits[303] ),
    .Q_N(\ConfigBits_N[303] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit8  (.D(net79),
    .GATE(net81),
    .Q(\ConfigBits[304] ),
    .Q_N(\ConfigBits_N[304] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame0_bit9  (.D(net80),
    .GATE(net81),
    .Q(\ConfigBits[305] ),
    .Q_N(\ConfigBits_N[305] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame10_bit24  (.D(net65),
    .GATE(net82),
    .Q(\ConfigBits[0] ),
    .Q_N(\ConfigBits_N[0] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame10_bit25  (.D(net66),
    .GATE(net82),
    .Q(\ConfigBits[1] ),
    .Q_N(\ConfigBits_N[1] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame10_bit26  (.D(net67),
    .GATE(net82),
    .Q(\ConfigBits[2] ),
    .Q_N(\ConfigBits_N[2] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame10_bit27  (.D(net68),
    .GATE(net82),
    .Q(\ConfigBits[3] ),
    .Q_N(\ConfigBits_N[3] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame10_bit28  (.D(net69),
    .GATE(net82),
    .Q(\ConfigBits[4] ),
    .Q_N(\ConfigBits_N[4] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame10_bit29  (.D(net70),
    .GATE(net82),
    .Q(\ConfigBits[5] ),
    .Q_N(\ConfigBits_N[5] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame10_bit30  (.D(net72),
    .GATE(net82),
    .Q(\ConfigBits[6] ),
    .Q_N(\ConfigBits_N[6] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame10_bit31  (.D(net73),
    .GATE(net82),
    .Q(\ConfigBits[7] ),
    .Q_N(\ConfigBits_N[7] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit0  (.D(net49),
    .GATE(net92),
    .Q(\ConfigBits[264] ),
    .Q_N(\ConfigBits_N[264] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit1  (.D(net60),
    .GATE(net92),
    .Q(\ConfigBits[265] ),
    .Q_N(\ConfigBits_N[265] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit10  (.D(net50),
    .GATE(net92),
    .Q(\ConfigBits[274] ),
    .Q_N(\ConfigBits_N[274] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit11  (.D(net51),
    .GATE(net92),
    .Q(\ConfigBits[275] ),
    .Q_N(\ConfigBits_N[275] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit12  (.D(net52),
    .GATE(net92),
    .Q(\ConfigBits[276] ),
    .Q_N(\ConfigBits_N[276] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit13  (.D(net53),
    .GATE(net92),
    .Q(\ConfigBits[277] ),
    .Q_N(\ConfigBits_N[277] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit14  (.D(net54),
    .GATE(net92),
    .Q(\ConfigBits[278] ),
    .Q_N(\ConfigBits_N[278] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit15  (.D(net55),
    .GATE(net92),
    .Q(\ConfigBits[279] ),
    .Q_N(\ConfigBits_N[279] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit16  (.D(net56),
    .GATE(net92),
    .Q(\ConfigBits[280] ),
    .Q_N(\ConfigBits_N[280] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit17  (.D(net57),
    .GATE(net92),
    .Q(\ConfigBits[281] ),
    .Q_N(\ConfigBits_N[281] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit18  (.D(net58),
    .GATE(net92),
    .Q(\ConfigBits[282] ),
    .Q_N(\ConfigBits_N[282] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit19  (.D(net59),
    .GATE(net92),
    .Q(\ConfigBits[283] ),
    .Q_N(\ConfigBits_N[283] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit2  (.D(net71),
    .GATE(net92),
    .Q(\ConfigBits[266] ),
    .Q_N(\ConfigBits_N[266] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit20  (.D(net61),
    .GATE(net92),
    .Q(\ConfigBits[284] ),
    .Q_N(\ConfigBits_N[284] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit21  (.D(net62),
    .GATE(net92),
    .Q(\ConfigBits[285] ),
    .Q_N(\ConfigBits_N[285] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit22  (.D(net63),
    .GATE(net92),
    .Q(\ConfigBits[286] ),
    .Q_N(\ConfigBits_N[286] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit23  (.D(net64),
    .GATE(net92),
    .Q(\ConfigBits[287] ),
    .Q_N(\ConfigBits_N[287] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit24  (.D(net65),
    .GATE(net92),
    .Q(\ConfigBits[288] ),
    .Q_N(\ConfigBits_N[288] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit25  (.D(net66),
    .GATE(net92),
    .Q(\ConfigBits[289] ),
    .Q_N(\ConfigBits_N[289] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit26  (.D(net67),
    .GATE(net92),
    .Q(\ConfigBits[290] ),
    .Q_N(\ConfigBits_N[290] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit27  (.D(net68),
    .GATE(net92),
    .Q(\ConfigBits[291] ),
    .Q_N(\ConfigBits_N[291] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit28  (.D(net69),
    .GATE(net92),
    .Q(\ConfigBits[292] ),
    .Q_N(\ConfigBits_N[292] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit29  (.D(net70),
    .GATE(net92),
    .Q(\ConfigBits[293] ),
    .Q_N(\ConfigBits_N[293] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit3  (.D(net74),
    .GATE(net92),
    .Q(\ConfigBits[267] ),
    .Q_N(\ConfigBits_N[267] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit30  (.D(net72),
    .GATE(net92),
    .Q(\ConfigBits[294] ),
    .Q_N(\ConfigBits_N[294] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit31  (.D(net73),
    .GATE(net92),
    .Q(\ConfigBits[295] ),
    .Q_N(\ConfigBits_N[295] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit4  (.D(net75),
    .GATE(net92),
    .Q(\ConfigBits[268] ),
    .Q_N(\ConfigBits_N[268] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit5  (.D(net76),
    .GATE(net92),
    .Q(\ConfigBits[269] ),
    .Q_N(\ConfigBits_N[269] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit6  (.D(net77),
    .GATE(net92),
    .Q(\ConfigBits[270] ),
    .Q_N(\ConfigBits_N[270] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit7  (.D(net78),
    .GATE(net92),
    .Q(\ConfigBits[271] ),
    .Q_N(\ConfigBits_N[271] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit8  (.D(net79),
    .GATE(net92),
    .Q(\ConfigBits[272] ),
    .Q_N(\ConfigBits_N[272] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame1_bit9  (.D(net80),
    .GATE(net92),
    .Q(\ConfigBits[273] ),
    .Q_N(\ConfigBits_N[273] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit0  (.D(net49),
    .GATE(net93),
    .Q(\ConfigBits[232] ),
    .Q_N(\ConfigBits_N[232] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit1  (.D(net60),
    .GATE(net93),
    .Q(\ConfigBits[233] ),
    .Q_N(\ConfigBits_N[233] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit10  (.D(net50),
    .GATE(net93),
    .Q(\ConfigBits[242] ),
    .Q_N(\ConfigBits_N[242] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit11  (.D(net51),
    .GATE(net93),
    .Q(\ConfigBits[243] ),
    .Q_N(\ConfigBits_N[243] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit12  (.D(net52),
    .GATE(net93),
    .Q(\ConfigBits[244] ),
    .Q_N(\ConfigBits_N[244] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit13  (.D(net53),
    .GATE(net93),
    .Q(\ConfigBits[245] ),
    .Q_N(\ConfigBits_N[245] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit14  (.D(net54),
    .GATE(net93),
    .Q(\ConfigBits[246] ),
    .Q_N(\ConfigBits_N[246] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit15  (.D(net55),
    .GATE(net93),
    .Q(\ConfigBits[247] ),
    .Q_N(\ConfigBits_N[247] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit16  (.D(net56),
    .GATE(net93),
    .Q(\ConfigBits[248] ),
    .Q_N(\ConfigBits_N[248] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit17  (.D(net57),
    .GATE(net93),
    .Q(\ConfigBits[249] ),
    .Q_N(\ConfigBits_N[249] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit18  (.D(net58),
    .GATE(net93),
    .Q(\ConfigBits[250] ),
    .Q_N(\ConfigBits_N[250] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit19  (.D(net59),
    .GATE(net93),
    .Q(\ConfigBits[251] ),
    .Q_N(\ConfigBits_N[251] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit2  (.D(net71),
    .GATE(net93),
    .Q(\ConfigBits[234] ),
    .Q_N(\ConfigBits_N[234] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit20  (.D(net61),
    .GATE(net93),
    .Q(\ConfigBits[252] ),
    .Q_N(\ConfigBits_N[252] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit21  (.D(net62),
    .GATE(net93),
    .Q(\ConfigBits[253] ),
    .Q_N(\ConfigBits_N[253] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit22  (.D(net63),
    .GATE(net93),
    .Q(\ConfigBits[254] ),
    .Q_N(\ConfigBits_N[254] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit23  (.D(net64),
    .GATE(net93),
    .Q(\ConfigBits[255] ),
    .Q_N(\ConfigBits_N[255] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit24  (.D(net65),
    .GATE(net93),
    .Q(\ConfigBits[256] ),
    .Q_N(\ConfigBits_N[256] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit25  (.D(net66),
    .GATE(net93),
    .Q(\ConfigBits[257] ),
    .Q_N(\ConfigBits_N[257] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit26  (.D(net67),
    .GATE(net93),
    .Q(\ConfigBits[258] ),
    .Q_N(\ConfigBits_N[258] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit27  (.D(net68),
    .GATE(net93),
    .Q(\ConfigBits[259] ),
    .Q_N(\ConfigBits_N[259] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit28  (.D(net69),
    .GATE(net93),
    .Q(\ConfigBits[260] ),
    .Q_N(\ConfigBits_N[260] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit29  (.D(net70),
    .GATE(net93),
    .Q(\ConfigBits[261] ),
    .Q_N(\ConfigBits_N[261] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit3  (.D(net74),
    .GATE(net93),
    .Q(\ConfigBits[235] ),
    .Q_N(\ConfigBits_N[235] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit30  (.D(net72),
    .GATE(net93),
    .Q(\ConfigBits[262] ),
    .Q_N(\ConfigBits_N[262] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit31  (.D(net73),
    .GATE(net93),
    .Q(\ConfigBits[263] ),
    .Q_N(\ConfigBits_N[263] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit4  (.D(net75),
    .GATE(net93),
    .Q(\ConfigBits[236] ),
    .Q_N(\ConfigBits_N[236] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit5  (.D(net76),
    .GATE(net93),
    .Q(\ConfigBits[237] ),
    .Q_N(\ConfigBits_N[237] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit6  (.D(net77),
    .GATE(net93),
    .Q(\ConfigBits[238] ),
    .Q_N(\ConfigBits_N[238] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit7  (.D(net78),
    .GATE(net93),
    .Q(\ConfigBits[239] ),
    .Q_N(\ConfigBits_N[239] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit8  (.D(net79),
    .GATE(net93),
    .Q(\ConfigBits[240] ),
    .Q_N(\ConfigBits_N[240] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame2_bit9  (.D(net80),
    .GATE(net93),
    .Q(\ConfigBits[241] ),
    .Q_N(\ConfigBits_N[241] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit0  (.D(net49),
    .GATE(net94),
    .Q(\ConfigBits[200] ),
    .Q_N(\ConfigBits_N[200] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit1  (.D(net60),
    .GATE(net94),
    .Q(\ConfigBits[201] ),
    .Q_N(\ConfigBits_N[201] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit10  (.D(net50),
    .GATE(net94),
    .Q(\ConfigBits[210] ),
    .Q_N(\ConfigBits_N[210] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit11  (.D(net51),
    .GATE(net94),
    .Q(\ConfigBits[211] ),
    .Q_N(\ConfigBits_N[211] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit12  (.D(net52),
    .GATE(net94),
    .Q(\ConfigBits[212] ),
    .Q_N(\ConfigBits_N[212] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit13  (.D(net53),
    .GATE(net94),
    .Q(\ConfigBits[213] ),
    .Q_N(\ConfigBits_N[213] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit14  (.D(net54),
    .GATE(net94),
    .Q(\ConfigBits[214] ),
    .Q_N(\ConfigBits_N[214] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit15  (.D(net55),
    .GATE(net94),
    .Q(\ConfigBits[215] ),
    .Q_N(\ConfigBits_N[215] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit16  (.D(net56),
    .GATE(net94),
    .Q(\ConfigBits[216] ),
    .Q_N(\ConfigBits_N[216] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit17  (.D(net57),
    .GATE(net94),
    .Q(\ConfigBits[217] ),
    .Q_N(\ConfigBits_N[217] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit18  (.D(net58),
    .GATE(net94),
    .Q(\ConfigBits[218] ),
    .Q_N(\ConfigBits_N[218] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit19  (.D(net59),
    .GATE(net94),
    .Q(\ConfigBits[219] ),
    .Q_N(\ConfigBits_N[219] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit2  (.D(net71),
    .GATE(net94),
    .Q(\ConfigBits[202] ),
    .Q_N(\ConfigBits_N[202] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit20  (.D(net61),
    .GATE(net94),
    .Q(\ConfigBits[220] ),
    .Q_N(\ConfigBits_N[220] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit21  (.D(net62),
    .GATE(net94),
    .Q(\ConfigBits[221] ),
    .Q_N(\ConfigBits_N[221] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit22  (.D(net63),
    .GATE(net94),
    .Q(\ConfigBits[222] ),
    .Q_N(\ConfigBits_N[222] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit23  (.D(net64),
    .GATE(net94),
    .Q(\ConfigBits[223] ),
    .Q_N(\ConfigBits_N[223] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit24  (.D(net65),
    .GATE(net94),
    .Q(\ConfigBits[224] ),
    .Q_N(\ConfigBits_N[224] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit25  (.D(net66),
    .GATE(net94),
    .Q(\ConfigBits[225] ),
    .Q_N(\ConfigBits_N[225] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit26  (.D(net67),
    .GATE(net94),
    .Q(\ConfigBits[226] ),
    .Q_N(\ConfigBits_N[226] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit27  (.D(net68),
    .GATE(net94),
    .Q(\ConfigBits[227] ),
    .Q_N(\ConfigBits_N[227] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit28  (.D(net69),
    .GATE(net94),
    .Q(\ConfigBits[228] ),
    .Q_N(\ConfigBits_N[228] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit29  (.D(net70),
    .GATE(net94),
    .Q(\ConfigBits[229] ),
    .Q_N(\ConfigBits_N[229] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit3  (.D(net74),
    .GATE(net94),
    .Q(\ConfigBits[203] ),
    .Q_N(\ConfigBits_N[203] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit30  (.D(net72),
    .GATE(net94),
    .Q(\ConfigBits[230] ),
    .Q_N(\ConfigBits_N[230] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit31  (.D(net73),
    .GATE(net94),
    .Q(\ConfigBits[231] ),
    .Q_N(\ConfigBits_N[231] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit4  (.D(net75),
    .GATE(net94),
    .Q(\ConfigBits[204] ),
    .Q_N(\ConfigBits_N[204] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit5  (.D(net76),
    .GATE(net94),
    .Q(\ConfigBits[205] ),
    .Q_N(\ConfigBits_N[205] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit6  (.D(net77),
    .GATE(net94),
    .Q(\ConfigBits[206] ),
    .Q_N(\ConfigBits_N[206] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit7  (.D(net78),
    .GATE(net94),
    .Q(\ConfigBits[207] ),
    .Q_N(\ConfigBits_N[207] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit8  (.D(net79),
    .GATE(net94),
    .Q(\ConfigBits[208] ),
    .Q_N(\ConfigBits_N[208] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame3_bit9  (.D(net80),
    .GATE(net94),
    .Q(\ConfigBits[209] ),
    .Q_N(\ConfigBits_N[209] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit0  (.D(net49),
    .GATE(net95),
    .Q(\ConfigBits[168] ),
    .Q_N(\ConfigBits_N[168] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit1  (.D(net60),
    .GATE(net95),
    .Q(\ConfigBits[169] ),
    .Q_N(\ConfigBits_N[169] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit10  (.D(net50),
    .GATE(net95),
    .Q(\ConfigBits[178] ),
    .Q_N(\ConfigBits_N[178] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit11  (.D(net51),
    .GATE(net95),
    .Q(\ConfigBits[179] ),
    .Q_N(\ConfigBits_N[179] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit12  (.D(net52),
    .GATE(net95),
    .Q(\ConfigBits[180] ),
    .Q_N(\ConfigBits_N[180] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit13  (.D(net53),
    .GATE(net95),
    .Q(\ConfigBits[181] ),
    .Q_N(\ConfigBits_N[181] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit14  (.D(net54),
    .GATE(net95),
    .Q(\ConfigBits[182] ),
    .Q_N(\ConfigBits_N[182] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit15  (.D(net55),
    .GATE(net95),
    .Q(\ConfigBits[183] ),
    .Q_N(\ConfigBits_N[183] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit16  (.D(net56),
    .GATE(net95),
    .Q(\ConfigBits[184] ),
    .Q_N(\ConfigBits_N[184] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit17  (.D(net57),
    .GATE(net95),
    .Q(\ConfigBits[185] ),
    .Q_N(\ConfigBits_N[185] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit18  (.D(net58),
    .GATE(net95),
    .Q(\ConfigBits[186] ),
    .Q_N(\ConfigBits_N[186] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit19  (.D(net59),
    .GATE(net95),
    .Q(\ConfigBits[187] ),
    .Q_N(\ConfigBits_N[187] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit2  (.D(net71),
    .GATE(net95),
    .Q(\ConfigBits[170] ),
    .Q_N(\ConfigBits_N[170] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit20  (.D(net61),
    .GATE(net95),
    .Q(\ConfigBits[188] ),
    .Q_N(\ConfigBits_N[188] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit21  (.D(net62),
    .GATE(net95),
    .Q(\ConfigBits[189] ),
    .Q_N(\ConfigBits_N[189] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit22  (.D(net63),
    .GATE(net95),
    .Q(\ConfigBits[190] ),
    .Q_N(\ConfigBits_N[190] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit23  (.D(net64),
    .GATE(net95),
    .Q(\ConfigBits[191] ),
    .Q_N(\ConfigBits_N[191] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit24  (.D(net65),
    .GATE(net95),
    .Q(\ConfigBits[192] ),
    .Q_N(\ConfigBits_N[192] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit25  (.D(net66),
    .GATE(net95),
    .Q(\ConfigBits[193] ),
    .Q_N(\ConfigBits_N[193] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit26  (.D(net67),
    .GATE(net95),
    .Q(\ConfigBits[194] ),
    .Q_N(\ConfigBits_N[194] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit27  (.D(net68),
    .GATE(net95),
    .Q(\ConfigBits[195] ),
    .Q_N(\ConfigBits_N[195] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit28  (.D(net69),
    .GATE(net95),
    .Q(\ConfigBits[196] ),
    .Q_N(\ConfigBits_N[196] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit29  (.D(net70),
    .GATE(net95),
    .Q(\ConfigBits[197] ),
    .Q_N(\ConfigBits_N[197] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit3  (.D(net74),
    .GATE(net95),
    .Q(\ConfigBits[171] ),
    .Q_N(\ConfigBits_N[171] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit30  (.D(net72),
    .GATE(net95),
    .Q(\ConfigBits[198] ),
    .Q_N(\ConfigBits_N[198] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit31  (.D(net73),
    .GATE(net95),
    .Q(\ConfigBits[199] ),
    .Q_N(\ConfigBits_N[199] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit4  (.D(net75),
    .GATE(net95),
    .Q(\ConfigBits[172] ),
    .Q_N(\ConfigBits_N[172] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit5  (.D(net76),
    .GATE(net95),
    .Q(\ConfigBits[173] ),
    .Q_N(\ConfigBits_N[173] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit6  (.D(net77),
    .GATE(net95),
    .Q(\ConfigBits[174] ),
    .Q_N(\ConfigBits_N[174] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit7  (.D(net78),
    .GATE(net95),
    .Q(\ConfigBits[175] ),
    .Q_N(\ConfigBits_N[175] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit8  (.D(net79),
    .GATE(net95),
    .Q(\ConfigBits[176] ),
    .Q_N(\ConfigBits_N[176] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame4_bit9  (.D(net80),
    .GATE(net95),
    .Q(\ConfigBits[177] ),
    .Q_N(\ConfigBits_N[177] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit0  (.D(net49),
    .GATE(net96),
    .Q(\ConfigBits[136] ),
    .Q_N(\ConfigBits_N[136] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit1  (.D(net60),
    .GATE(net96),
    .Q(\ConfigBits[137] ),
    .Q_N(\ConfigBits_N[137] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit10  (.D(net50),
    .GATE(net96),
    .Q(\ConfigBits[146] ),
    .Q_N(\ConfigBits_N[146] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit11  (.D(net51),
    .GATE(net96),
    .Q(\ConfigBits[147] ),
    .Q_N(\ConfigBits_N[147] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit12  (.D(net52),
    .GATE(net96),
    .Q(\ConfigBits[148] ),
    .Q_N(\ConfigBits_N[148] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit13  (.D(net53),
    .GATE(net96),
    .Q(\ConfigBits[149] ),
    .Q_N(\ConfigBits_N[149] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit14  (.D(net54),
    .GATE(net96),
    .Q(\ConfigBits[150] ),
    .Q_N(\ConfigBits_N[150] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit15  (.D(net55),
    .GATE(net96),
    .Q(\ConfigBits[151] ),
    .Q_N(\ConfigBits_N[151] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit16  (.D(net56),
    .GATE(net96),
    .Q(\ConfigBits[152] ),
    .Q_N(\ConfigBits_N[152] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit17  (.D(net57),
    .GATE(net96),
    .Q(\ConfigBits[153] ),
    .Q_N(\ConfigBits_N[153] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit18  (.D(net58),
    .GATE(net96),
    .Q(\ConfigBits[154] ),
    .Q_N(\ConfigBits_N[154] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit19  (.D(net59),
    .GATE(net96),
    .Q(\ConfigBits[155] ),
    .Q_N(\ConfigBits_N[155] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit2  (.D(net71),
    .GATE(net96),
    .Q(\ConfigBits[138] ),
    .Q_N(\ConfigBits_N[138] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit20  (.D(net61),
    .GATE(net96),
    .Q(\ConfigBits[156] ),
    .Q_N(\ConfigBits_N[156] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit21  (.D(net62),
    .GATE(net96),
    .Q(\ConfigBits[157] ),
    .Q_N(\ConfigBits_N[157] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit22  (.D(net63),
    .GATE(net96),
    .Q(\ConfigBits[158] ),
    .Q_N(\ConfigBits_N[158] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit23  (.D(net64),
    .GATE(net96),
    .Q(\ConfigBits[159] ),
    .Q_N(\ConfigBits_N[159] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit24  (.D(net65),
    .GATE(net96),
    .Q(\ConfigBits[160] ),
    .Q_N(\ConfigBits_N[160] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit25  (.D(net66),
    .GATE(net96),
    .Q(\ConfigBits[161] ),
    .Q_N(\ConfigBits_N[161] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit26  (.D(net67),
    .GATE(net96),
    .Q(\ConfigBits[162] ),
    .Q_N(\ConfigBits_N[162] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit27  (.D(net68),
    .GATE(net96),
    .Q(\ConfigBits[163] ),
    .Q_N(\ConfigBits_N[163] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit28  (.D(net69),
    .GATE(net96),
    .Q(\ConfigBits[164] ),
    .Q_N(\ConfigBits_N[164] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit29  (.D(net70),
    .GATE(net96),
    .Q(\ConfigBits[165] ),
    .Q_N(\ConfigBits_N[165] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit3  (.D(net74),
    .GATE(net96),
    .Q(\ConfigBits[139] ),
    .Q_N(\ConfigBits_N[139] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit30  (.D(net72),
    .GATE(net96),
    .Q(\ConfigBits[166] ),
    .Q_N(\ConfigBits_N[166] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit31  (.D(net73),
    .GATE(net96),
    .Q(\ConfigBits[167] ),
    .Q_N(\ConfigBits_N[167] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit4  (.D(net75),
    .GATE(net96),
    .Q(\ConfigBits[140] ),
    .Q_N(\ConfigBits_N[140] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit5  (.D(net76),
    .GATE(net96),
    .Q(\ConfigBits[141] ),
    .Q_N(\ConfigBits_N[141] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit6  (.D(net77),
    .GATE(net96),
    .Q(\ConfigBits[142] ),
    .Q_N(\ConfigBits_N[142] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit7  (.D(net78),
    .GATE(net96),
    .Q(\ConfigBits[143] ),
    .Q_N(\ConfigBits_N[143] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit8  (.D(net79),
    .GATE(net96),
    .Q(\ConfigBits[144] ),
    .Q_N(\ConfigBits_N[144] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame5_bit9  (.D(net80),
    .GATE(net96),
    .Q(\ConfigBits[145] ),
    .Q_N(\ConfigBits_N[145] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit0  (.D(net49),
    .GATE(net97),
    .Q(\ConfigBits[104] ),
    .Q_N(\ConfigBits_N[104] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit1  (.D(net60),
    .GATE(net97),
    .Q(\ConfigBits[105] ),
    .Q_N(\ConfigBits_N[105] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit10  (.D(net50),
    .GATE(net97),
    .Q(\ConfigBits[114] ),
    .Q_N(\ConfigBits_N[114] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit11  (.D(net51),
    .GATE(net97),
    .Q(\ConfigBits[115] ),
    .Q_N(\ConfigBits_N[115] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit12  (.D(net52),
    .GATE(net97),
    .Q(\ConfigBits[116] ),
    .Q_N(\ConfigBits_N[116] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit13  (.D(net53),
    .GATE(net97),
    .Q(\ConfigBits[117] ),
    .Q_N(\ConfigBits_N[117] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit14  (.D(net54),
    .GATE(net97),
    .Q(\ConfigBits[118] ),
    .Q_N(\ConfigBits_N[118] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit15  (.D(net55),
    .GATE(net97),
    .Q(\ConfigBits[119] ),
    .Q_N(\ConfigBits_N[119] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit16  (.D(net56),
    .GATE(net97),
    .Q(\ConfigBits[120] ),
    .Q_N(\ConfigBits_N[120] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit17  (.D(net57),
    .GATE(net97),
    .Q(\ConfigBits[121] ),
    .Q_N(\ConfigBits_N[121] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit18  (.D(net58),
    .GATE(net97),
    .Q(\ConfigBits[122] ),
    .Q_N(\ConfigBits_N[122] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit19  (.D(net59),
    .GATE(net97),
    .Q(\ConfigBits[123] ),
    .Q_N(\ConfigBits_N[123] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit2  (.D(net71),
    .GATE(net97),
    .Q(\ConfigBits[106] ),
    .Q_N(\ConfigBits_N[106] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit20  (.D(net61),
    .GATE(net97),
    .Q(\ConfigBits[124] ),
    .Q_N(\ConfigBits_N[124] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit21  (.D(net62),
    .GATE(net97),
    .Q(\ConfigBits[125] ),
    .Q_N(\ConfigBits_N[125] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit22  (.D(net63),
    .GATE(net97),
    .Q(\ConfigBits[126] ),
    .Q_N(\ConfigBits_N[126] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit23  (.D(net64),
    .GATE(net97),
    .Q(\ConfigBits[127] ),
    .Q_N(\ConfigBits_N[127] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit24  (.D(net65),
    .GATE(net97),
    .Q(\ConfigBits[128] ),
    .Q_N(\ConfigBits_N[128] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit25  (.D(net66),
    .GATE(net97),
    .Q(\ConfigBits[129] ),
    .Q_N(\ConfigBits_N[129] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit26  (.D(net67),
    .GATE(net97),
    .Q(\ConfigBits[130] ),
    .Q_N(\ConfigBits_N[130] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit27  (.D(net68),
    .GATE(net97),
    .Q(\ConfigBits[131] ),
    .Q_N(\ConfigBits_N[131] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit28  (.D(net69),
    .GATE(net97),
    .Q(\ConfigBits[132] ),
    .Q_N(\ConfigBits_N[132] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit29  (.D(net70),
    .GATE(net97),
    .Q(\ConfigBits[133] ),
    .Q_N(\ConfigBits_N[133] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit3  (.D(net74),
    .GATE(net97),
    .Q(\ConfigBits[107] ),
    .Q_N(\ConfigBits_N[107] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit30  (.D(net72),
    .GATE(net97),
    .Q(\ConfigBits[134] ),
    .Q_N(\ConfigBits_N[134] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit31  (.D(net73),
    .GATE(net97),
    .Q(\ConfigBits[135] ),
    .Q_N(\ConfigBits_N[135] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit4  (.D(net75),
    .GATE(net97),
    .Q(\ConfigBits[108] ),
    .Q_N(\ConfigBits_N[108] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit5  (.D(net76),
    .GATE(net97),
    .Q(\ConfigBits[109] ),
    .Q_N(\ConfigBits_N[109] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit6  (.D(net77),
    .GATE(net97),
    .Q(\ConfigBits[110] ),
    .Q_N(\ConfigBits_N[110] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit7  (.D(net78),
    .GATE(net97),
    .Q(\ConfigBits[111] ),
    .Q_N(\ConfigBits_N[111] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit8  (.D(net79),
    .GATE(net97),
    .Q(\ConfigBits[112] ),
    .Q_N(\ConfigBits_N[112] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame6_bit9  (.D(net80),
    .GATE(net97),
    .Q(\ConfigBits[113] ),
    .Q_N(\ConfigBits_N[113] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit0  (.D(net49),
    .GATE(net98),
    .Q(\ConfigBits[72] ),
    .Q_N(\ConfigBits_N[72] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit1  (.D(net60),
    .GATE(net98),
    .Q(\ConfigBits[73] ),
    .Q_N(\ConfigBits_N[73] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit10  (.D(net50),
    .GATE(net98),
    .Q(\ConfigBits[82] ),
    .Q_N(\ConfigBits_N[82] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit11  (.D(net51),
    .GATE(net98),
    .Q(\ConfigBits[83] ),
    .Q_N(\ConfigBits_N[83] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit12  (.D(net52),
    .GATE(net98),
    .Q(\ConfigBits[84] ),
    .Q_N(\ConfigBits_N[84] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit13  (.D(net53),
    .GATE(net98),
    .Q(\ConfigBits[85] ),
    .Q_N(\ConfigBits_N[85] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit14  (.D(net54),
    .GATE(net98),
    .Q(\ConfigBits[86] ),
    .Q_N(\ConfigBits_N[86] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit15  (.D(net55),
    .GATE(net98),
    .Q(\ConfigBits[87] ),
    .Q_N(\ConfigBits_N[87] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit16  (.D(net56),
    .GATE(net98),
    .Q(\ConfigBits[88] ),
    .Q_N(\ConfigBits_N[88] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit17  (.D(net57),
    .GATE(net98),
    .Q(\ConfigBits[89] ),
    .Q_N(\ConfigBits_N[89] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit18  (.D(net58),
    .GATE(net98),
    .Q(\ConfigBits[90] ),
    .Q_N(\ConfigBits_N[90] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit19  (.D(net59),
    .GATE(net98),
    .Q(\ConfigBits[91] ),
    .Q_N(\ConfigBits_N[91] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit2  (.D(net71),
    .GATE(net98),
    .Q(\ConfigBits[74] ),
    .Q_N(\ConfigBits_N[74] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit20  (.D(net61),
    .GATE(net98),
    .Q(\ConfigBits[92] ),
    .Q_N(\ConfigBits_N[92] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit21  (.D(net62),
    .GATE(net98),
    .Q(\ConfigBits[93] ),
    .Q_N(\ConfigBits_N[93] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit22  (.D(net63),
    .GATE(net98),
    .Q(\ConfigBits[94] ),
    .Q_N(\ConfigBits_N[94] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit23  (.D(net64),
    .GATE(net98),
    .Q(\ConfigBits[95] ),
    .Q_N(\ConfigBits_N[95] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit24  (.D(net65),
    .GATE(net98),
    .Q(\ConfigBits[96] ),
    .Q_N(\ConfigBits_N[96] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit25  (.D(net66),
    .GATE(net98),
    .Q(\ConfigBits[97] ),
    .Q_N(\ConfigBits_N[97] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit26  (.D(net67),
    .GATE(net98),
    .Q(\ConfigBits[98] ),
    .Q_N(\ConfigBits_N[98] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit27  (.D(net68),
    .GATE(net98),
    .Q(\ConfigBits[99] ),
    .Q_N(\ConfigBits_N[99] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit28  (.D(net69),
    .GATE(net98),
    .Q(\ConfigBits[100] ),
    .Q_N(\ConfigBits_N[100] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit29  (.D(net70),
    .GATE(net98),
    .Q(\ConfigBits[101] ),
    .Q_N(\ConfigBits_N[101] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit3  (.D(net74),
    .GATE(net98),
    .Q(\ConfigBits[75] ),
    .Q_N(\ConfigBits_N[75] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit30  (.D(net72),
    .GATE(net98),
    .Q(\ConfigBits[102] ),
    .Q_N(\ConfigBits_N[102] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit31  (.D(net73),
    .GATE(net98),
    .Q(\ConfigBits[103] ),
    .Q_N(\ConfigBits_N[103] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit4  (.D(net75),
    .GATE(net98),
    .Q(\ConfigBits[76] ),
    .Q_N(\ConfigBits_N[76] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit5  (.D(net76),
    .GATE(net98),
    .Q(\ConfigBits[77] ),
    .Q_N(\ConfigBits_N[77] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit6  (.D(net77),
    .GATE(net98),
    .Q(\ConfigBits[78] ),
    .Q_N(\ConfigBits_N[78] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit7  (.D(net78),
    .GATE(net98),
    .Q(\ConfigBits[79] ),
    .Q_N(\ConfigBits_N[79] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit8  (.D(net79),
    .GATE(net98),
    .Q(\ConfigBits[80] ),
    .Q_N(\ConfigBits_N[80] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame7_bit9  (.D(net80),
    .GATE(net98),
    .Q(\ConfigBits[81] ),
    .Q_N(\ConfigBits_N[81] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit0  (.D(net49),
    .GATE(net99),
    .Q(\ConfigBits[40] ),
    .Q_N(\ConfigBits_N[40] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit1  (.D(net60),
    .GATE(net99),
    .Q(\ConfigBits[41] ),
    .Q_N(\ConfigBits_N[41] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit10  (.D(net50),
    .GATE(net99),
    .Q(\ConfigBits[50] ),
    .Q_N(\ConfigBits_N[50] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit11  (.D(net51),
    .GATE(net99),
    .Q(\ConfigBits[51] ),
    .Q_N(\ConfigBits_N[51] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit12  (.D(net52),
    .GATE(net99),
    .Q(\ConfigBits[52] ),
    .Q_N(\ConfigBits_N[52] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit13  (.D(net53),
    .GATE(net99),
    .Q(\ConfigBits[53] ),
    .Q_N(\ConfigBits_N[53] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit14  (.D(net54),
    .GATE(net99),
    .Q(\ConfigBits[54] ),
    .Q_N(\ConfigBits_N[54] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit15  (.D(net55),
    .GATE(net99),
    .Q(\ConfigBits[55] ),
    .Q_N(\ConfigBits_N[55] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit16  (.D(net56),
    .GATE(net99),
    .Q(\ConfigBits[56] ),
    .Q_N(\ConfigBits_N[56] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit17  (.D(net57),
    .GATE(net99),
    .Q(\ConfigBits[57] ),
    .Q_N(\ConfigBits_N[57] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit18  (.D(net58),
    .GATE(net99),
    .Q(\ConfigBits[58] ),
    .Q_N(\ConfigBits_N[58] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit19  (.D(net59),
    .GATE(net99),
    .Q(\ConfigBits[59] ),
    .Q_N(\ConfigBits_N[59] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit2  (.D(net71),
    .GATE(net99),
    .Q(\ConfigBits[42] ),
    .Q_N(\ConfigBits_N[42] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit20  (.D(net61),
    .GATE(net99),
    .Q(\ConfigBits[60] ),
    .Q_N(\ConfigBits_N[60] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit21  (.D(net62),
    .GATE(net99),
    .Q(\ConfigBits[61] ),
    .Q_N(\ConfigBits_N[61] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit22  (.D(net63),
    .GATE(net99),
    .Q(\ConfigBits[62] ),
    .Q_N(\ConfigBits_N[62] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit23  (.D(net64),
    .GATE(net99),
    .Q(\ConfigBits[63] ),
    .Q_N(\ConfigBits_N[63] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit24  (.D(net65),
    .GATE(net99),
    .Q(\ConfigBits[64] ),
    .Q_N(\ConfigBits_N[64] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit25  (.D(net66),
    .GATE(net99),
    .Q(\ConfigBits[65] ),
    .Q_N(\ConfigBits_N[65] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit26  (.D(net67),
    .GATE(net99),
    .Q(\ConfigBits[66] ),
    .Q_N(\ConfigBits_N[66] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit27  (.D(net68),
    .GATE(net99),
    .Q(\ConfigBits[67] ),
    .Q_N(\ConfigBits_N[67] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit28  (.D(net69),
    .GATE(net99),
    .Q(\ConfigBits[68] ),
    .Q_N(\ConfigBits_N[68] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit29  (.D(net70),
    .GATE(net99),
    .Q(\ConfigBits[69] ),
    .Q_N(\ConfigBits_N[69] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit3  (.D(net74),
    .GATE(net99),
    .Q(\ConfigBits[43] ),
    .Q_N(\ConfigBits_N[43] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit30  (.D(net72),
    .GATE(net99),
    .Q(\ConfigBits[70] ),
    .Q_N(\ConfigBits_N[70] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit31  (.D(net73),
    .GATE(net99),
    .Q(\ConfigBits[71] ),
    .Q_N(\ConfigBits_N[71] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit4  (.D(net75),
    .GATE(net99),
    .Q(\ConfigBits[44] ),
    .Q_N(\ConfigBits_N[44] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit5  (.D(net76),
    .GATE(net99),
    .Q(\ConfigBits[45] ),
    .Q_N(\ConfigBits_N[45] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit6  (.D(net77),
    .GATE(net99),
    .Q(\ConfigBits[46] ),
    .Q_N(\ConfigBits_N[46] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit7  (.D(net78),
    .GATE(net99),
    .Q(\ConfigBits[47] ),
    .Q_N(\ConfigBits_N[47] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit8  (.D(net79),
    .GATE(net99),
    .Q(\ConfigBits[48] ),
    .Q_N(\ConfigBits_N[48] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame8_bit9  (.D(net80),
    .GATE(net99),
    .Q(\ConfigBits[49] ),
    .Q_N(\ConfigBits_N[49] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit0  (.D(net49),
    .GATE(net100),
    .Q(\ConfigBits[8] ),
    .Q_N(\ConfigBits_N[8] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit1  (.D(net60),
    .GATE(net100),
    .Q(\ConfigBits[9] ),
    .Q_N(\ConfigBits_N[9] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit10  (.D(net50),
    .GATE(net100),
    .Q(\ConfigBits[18] ),
    .Q_N(\ConfigBits_N[18] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit11  (.D(net51),
    .GATE(net100),
    .Q(\ConfigBits[19] ),
    .Q_N(\ConfigBits_N[19] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit12  (.D(net52),
    .GATE(net100),
    .Q(\ConfigBits[20] ),
    .Q_N(\ConfigBits_N[20] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit13  (.D(net53),
    .GATE(net100),
    .Q(\ConfigBits[21] ),
    .Q_N(\ConfigBits_N[21] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit14  (.D(net54),
    .GATE(net100),
    .Q(\ConfigBits[22] ),
    .Q_N(\ConfigBits_N[22] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit15  (.D(net55),
    .GATE(net100),
    .Q(\ConfigBits[23] ),
    .Q_N(\ConfigBits_N[23] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit16  (.D(net56),
    .GATE(net100),
    .Q(\ConfigBits[24] ),
    .Q_N(\ConfigBits_N[24] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit17  (.D(net57),
    .GATE(net100),
    .Q(\ConfigBits[25] ),
    .Q_N(\ConfigBits_N[25] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit18  (.D(net58),
    .GATE(net100),
    .Q(\ConfigBits[26] ),
    .Q_N(\ConfigBits_N[26] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit19  (.D(net59),
    .GATE(net100),
    .Q(\ConfigBits[27] ),
    .Q_N(\ConfigBits_N[27] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit2  (.D(net71),
    .GATE(net100),
    .Q(\ConfigBits[10] ),
    .Q_N(\ConfigBits_N[10] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit20  (.D(net61),
    .GATE(net100),
    .Q(\ConfigBits[28] ),
    .Q_N(\ConfigBits_N[28] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit21  (.D(net62),
    .GATE(net100),
    .Q(\ConfigBits[29] ),
    .Q_N(\ConfigBits_N[29] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit22  (.D(net63),
    .GATE(net100),
    .Q(\ConfigBits[30] ),
    .Q_N(\ConfigBits_N[30] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit23  (.D(net64),
    .GATE(net100),
    .Q(\ConfigBits[31] ),
    .Q_N(\ConfigBits_N[31] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit24  (.D(net65),
    .GATE(net100),
    .Q(\ConfigBits[32] ),
    .Q_N(\ConfigBits_N[32] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit25  (.D(net66),
    .GATE(net100),
    .Q(\ConfigBits[33] ),
    .Q_N(\ConfigBits_N[33] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit26  (.D(net67),
    .GATE(net100),
    .Q(\ConfigBits[34] ),
    .Q_N(\ConfigBits_N[34] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit27  (.D(net68),
    .GATE(net100),
    .Q(\ConfigBits[35] ),
    .Q_N(\ConfigBits_N[35] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit28  (.D(net69),
    .GATE(net100),
    .Q(\ConfigBits[36] ),
    .Q_N(\ConfigBits_N[36] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit29  (.D(net70),
    .GATE(net100),
    .Q(\ConfigBits[37] ),
    .Q_N(\ConfigBits_N[37] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit3  (.D(net74),
    .GATE(net100),
    .Q(\ConfigBits[11] ),
    .Q_N(\ConfigBits_N[11] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit30  (.D(net72),
    .GATE(net100),
    .Q(\ConfigBits[38] ),
    .Q_N(\ConfigBits_N[38] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit31  (.D(net73),
    .GATE(net100),
    .Q(\ConfigBits[39] ),
    .Q_N(\ConfigBits_N[39] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit4  (.D(net75),
    .GATE(net100),
    .Q(\ConfigBits[12] ),
    .Q_N(\ConfigBits_N[12] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit5  (.D(net76),
    .GATE(net100),
    .Q(\ConfigBits[13] ),
    .Q_N(\ConfigBits_N[13] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit6  (.D(net77),
    .GATE(net100),
    .Q(\ConfigBits[14] ),
    .Q_N(\ConfigBits_N[14] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit7  (.D(net78),
    .GATE(net100),
    .Q(\ConfigBits[15] ),
    .Q_N(\ConfigBits_N[15] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit8  (.D(net79),
    .GATE(net100),
    .Q(\ConfigBits[16] ),
    .Q_N(\ConfigBits_N[16] ));
 sky130_fd_sc_hd__dlxbp_1 \Inst_RAM_IO_ConfigMem/Inst_frame9_bit9  (.D(net80),
    .GATE(net100),
    .Q(\ConfigBits[17] ),
    .Q_N(\ConfigBits_N[17] ));
 sky130_fd_sc_hd__buf_2 \Inst_RAM_IO_switch_matrix/_32_  (.A(net113),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/_33_  (.A(net114),
    .X(net286));
 sky130_fd_sc_hd__buf_1 \Inst_RAM_IO_switch_matrix/_34_  (.A(net115),
    .X(net287));
 sky130_fd_sc_hd__buf_1 \Inst_RAM_IO_switch_matrix/_35_  (.A(net116),
    .X(net288));
 sky130_fd_sc_hd__buf_2 \Inst_RAM_IO_switch_matrix/_36_  (.A(net117),
    .X(net289));
 sky130_fd_sc_hd__dlymetal6s2s_1 \Inst_RAM_IO_switch_matrix/_37_  (.A(net118),
    .X(net290));
 sky130_fd_sc_hd__buf_1 \Inst_RAM_IO_switch_matrix/_38_  (.A(net119),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix/_39_  (.A(net120),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/_40_  (.A(net165),
    .X(net321));
 sky130_fd_sc_hd__buf_2 \Inst_RAM_IO_switch_matrix/_41_  (.A(net166),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix/_42_  (.A(net167),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix/_43_  (.A(net168),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/_44_  (.A(net169),
    .X(net325));
 sky130_fd_sc_hd__buf_1 \Inst_RAM_IO_switch_matrix/_45_  (.A(net170),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 \Inst_RAM_IO_switch_matrix/_46_  (.A(net171),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/_47_  (.A(net172),
    .X(net328));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A0_I0  (.A0(net13),
    .A1(net5),
    .A2(\J_NS2_BEG[0] ),
    .A3(net395),
    .S0(\ConfigBits[248] ),
    .S1(\ConfigBits[249] ),
    .X(FAB2RAM_A0_I0));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A0_I0_395  (.LO(net395));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A0_I1  (.A0(net14),
    .A1(net6),
    .A2(\J_NS2_BEG[1] ),
    .A3(net396),
    .S0(\ConfigBits[250] ),
    .S1(\ConfigBits[251] ),
    .X(FAB2RAM_A0_I1));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A0_I1_396  (.LO(net396));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A0_I2  (.A0(net15),
    .A1(net7),
    .A2(\J_NS2_BEG[2] ),
    .A3(net397),
    .S0(\ConfigBits[252] ),
    .S1(\ConfigBits[253] ),
    .X(FAB2RAM_A0_I2));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A0_I2_397  (.LO(net397));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A0_I3  (.A0(net16),
    .A1(net8),
    .A2(\J_NS2_BEG[3] ),
    .A3(net398),
    .S0(\ConfigBits[254] ),
    .S1(\ConfigBits[255] ),
    .X(FAB2RAM_A0_I3));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A0_I3_398  (.LO(net398));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A1_I0  (.A0(net17),
    .A1(net9),
    .A2(\J_NS2_BEG[4] ),
    .A3(net399),
    .S0(\ConfigBits[256] ),
    .S1(\ConfigBits[257] ),
    .X(FAB2RAM_A1_I0));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A1_I0_399  (.LO(net399));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A1_I1  (.A0(net18),
    .A1(net10),
    .A2(\J_NS2_BEG[5] ),
    .A3(net400),
    .S0(\ConfigBits[258] ),
    .S1(\ConfigBits[259] ),
    .X(FAB2RAM_A1_I1));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A1_I1_400  (.LO(net400));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A1_I2  (.A0(net19),
    .A1(net11),
    .A2(\J_NS2_BEG[6] ),
    .A3(net401),
    .S0(\ConfigBits[260] ),
    .S1(\ConfigBits[261] ),
    .X(FAB2RAM_A1_I2));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A1_I2_401  (.LO(net401));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A1_I3  (.A0(net20),
    .A1(net12),
    .A2(\J_NS2_BEG[7] ),
    .A3(net402),
    .S0(\ConfigBits[262] ),
    .S1(\ConfigBits[263] ),
    .X(FAB2RAM_A1_I3));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_A1_I3_402  (.LO(net402));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_C_I0  (.A0(net1),
    .A1(net21),
    .A2(\J_NS1_BEG[0] ),
    .A3(net403),
    .S0(\ConfigBits[264] ),
    .S1(\ConfigBits[265] ),
    .X(FAB2RAM_C_I0));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_C_I0_403  (.LO(net403));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_C_I1  (.A0(net2),
    .A1(net24),
    .A2(\J_NS1_BEG[1] ),
    .A3(net404),
    .S0(\ConfigBits[266] ),
    .S1(\ConfigBits[267] ),
    .X(FAB2RAM_C_I1));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_C_I1_404  (.LO(net404));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_C_I2  (.A0(net3),
    .A1(net25),
    .A2(\J_NS1_BEG[2] ),
    .A3(net405),
    .S0(\ConfigBits[268] ),
    .S1(\ConfigBits[269] ),
    .X(FAB2RAM_C_I2));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_C_I2_405  (.LO(net405));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_C_I3  (.A0(net4),
    .A1(net26),
    .A2(\J_NS1_BEG[3] ),
    .A3(net409),
    .S0(\ConfigBits[270] ),
    .S1(\ConfigBits[271] ),
    .X(FAB2RAM_C_I3));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_C_I3_409  (.LO(net409));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D0_I0  (.A0(net33),
    .A1(net47),
    .A2(net21),
    .A3(\J_NS4_BEG[0] ),
    .S0(\ConfigBits[216] ),
    .S1(\ConfigBits[217] ),
    .X(FAB2RAM_D0_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D0_I1  (.A0(net40),
    .A1(net48),
    .A2(net24),
    .A3(\J_NS4_BEG[1] ),
    .S0(\ConfigBits[218] ),
    .S1(\ConfigBits[219] ),
    .X(FAB2RAM_D0_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D0_I2  (.A0(net41),
    .A1(net34),
    .A2(net25),
    .A3(\J_NS4_BEG[2] ),
    .S0(\ConfigBits[220] ),
    .S1(\ConfigBits[221] ),
    .X(FAB2RAM_D0_I2));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D0_I3  (.A0(net42),
    .A1(net35),
    .A2(net26),
    .A3(\J_NS4_BEG[3] ),
    .S0(\ConfigBits[222] ),
    .S1(\ConfigBits[223] ),
    .X(FAB2RAM_D0_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D1_I0  (.A0(net43),
    .A1(net36),
    .A2(net27),
    .A3(\J_NS4_BEG[4] ),
    .S0(\ConfigBits[224] ),
    .S1(\ConfigBits[225] ),
    .X(FAB2RAM_D1_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D1_I1  (.A0(net44),
    .A1(net37),
    .A2(net28),
    .A3(\J_NS4_BEG[5] ),
    .S0(\ConfigBits[226] ),
    .S1(\ConfigBits[227] ),
    .X(FAB2RAM_D1_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D1_I2  (.A0(net45),
    .A1(net38),
    .A2(net29),
    .A3(\J_NS4_BEG[6] ),
    .S0(\ConfigBits[228] ),
    .S1(\ConfigBits[229] ),
    .X(FAB2RAM_D1_I2));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D1_I3  (.A0(net46),
    .A1(net39),
    .A2(net30),
    .A3(\J_NS4_BEG[7] ),
    .S0(\ConfigBits[230] ),
    .S1(\ConfigBits[231] ),
    .X(FAB2RAM_D1_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D2_I0  (.A0(net33),
    .A1(net47),
    .A2(net31),
    .A3(\J_NS4_BEG[8] ),
    .S0(\ConfigBits[232] ),
    .S1(\ConfigBits[233] ),
    .X(FAB2RAM_D2_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D2_I1  (.A0(net40),
    .A1(net48),
    .A2(net32),
    .A3(\J_NS4_BEG[9] ),
    .S0(\ConfigBits[234] ),
    .S1(\ConfigBits[235] ),
    .X(FAB2RAM_D2_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D2_I2  (.A0(net41),
    .A1(net34),
    .A2(net22),
    .A3(\J_NS4_BEG[10] ),
    .S0(\ConfigBits[236] ),
    .S1(\ConfigBits[237] ),
    .X(FAB2RAM_D2_I2));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D2_I3  (.A0(net42),
    .A1(net35),
    .A2(net23),
    .A3(\J_NS4_BEG[11] ),
    .S0(\ConfigBits[238] ),
    .S1(\ConfigBits[239] ),
    .X(FAB2RAM_D2_I3));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D3_I0  (.A0(net1),
    .A1(net43),
    .A2(net36),
    .A3(\J_NS4_BEG[12] ),
    .S0(\ConfigBits[240] ),
    .S1(\ConfigBits[241] ),
    .X(FAB2RAM_D3_I0));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D3_I1  (.A0(net2),
    .A1(net44),
    .A2(net37),
    .A3(\J_NS4_BEG[13] ),
    .S0(\ConfigBits[242] ),
    .S1(\ConfigBits[243] ),
    .X(FAB2RAM_D3_I1));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D3_I2  (.A0(net3),
    .A1(net45),
    .A2(net38),
    .A3(\J_NS4_BEG[14] ),
    .S0(\ConfigBits[244] ),
    .S1(\ConfigBits[245] ),
    .X(FAB2RAM_D3_I2));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_FAB2RAM_D3_I3  (.A0(net4),
    .A1(net46),
    .A2(net39),
    .A3(\J_NS4_BEG[15] ),
    .S0(\ConfigBits[246] ),
    .S1(\ConfigBits[247] ),
    .X(FAB2RAM_D3_I3));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS1_BEG0  (.A0(net101),
    .A1(net21),
    .A2(net153),
    .A3(net406),
    .S0(\ConfigBits[320] ),
    .S1(\ConfigBits[321] ),
    .X(\J_NS1_BEG[0] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS1_BEG0_406  (.LO(net406));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS1_BEG1  (.A0(net102),
    .A1(net24),
    .A2(net154),
    .A3(net407),
    .S0(\ConfigBits[322] ),
    .S1(\ConfigBits[323] ),
    .X(\J_NS1_BEG[1] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS1_BEG1_407  (.LO(net407));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS1_BEG2  (.A0(net103),
    .A1(net25),
    .A2(net155),
    .A3(net408),
    .S0(\ConfigBits[324] ),
    .S1(\ConfigBits[325] ),
    .X(\J_NS1_BEG[2] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS1_BEG2_408  (.LO(net408));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS1_BEG3  (.A0(net104),
    .A1(net26),
    .A2(net156),
    .A3(net394),
    .S0(\ConfigBits[326] ),
    .S1(\ConfigBits[327] ),
    .X(\J_NS1_BEG[3] ));
 sky130_fd_sc_hd__conb_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS1_BEG3_394  (.LO(net394));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS2_BEG0  (.A0(net113),
    .A1(net105),
    .A2(net165),
    .A3(net157),
    .S0(\ConfigBits[304] ),
    .S1(\ConfigBits[305] ),
    .X(\J_NS2_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS2_BEG1  (.A0(net114),
    .A1(net106),
    .A2(net166),
    .A3(net158),
    .S0(\ConfigBits[306] ),
    .S1(\ConfigBits[307] ),
    .X(\J_NS2_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS2_BEG2  (.A0(net115),
    .A1(net107),
    .A2(net167),
    .A3(net159),
    .S0(\ConfigBits[308] ),
    .S1(\ConfigBits[309] ),
    .X(\J_NS2_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS2_BEG3  (.A0(net116),
    .A1(net108),
    .A2(net168),
    .A3(net160),
    .S0(\ConfigBits[310] ),
    .S1(\ConfigBits[311] ),
    .X(\J_NS2_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS2_BEG4  (.A0(net117),
    .A1(net109),
    .A2(net169),
    .A3(net161),
    .S0(\ConfigBits[312] ),
    .S1(\ConfigBits[313] ),
    .X(\J_NS2_BEG[4] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS2_BEG5  (.A0(net118),
    .A1(net110),
    .A2(net170),
    .A3(net162),
    .S0(\ConfigBits[314] ),
    .S1(\ConfigBits[315] ),
    .X(\J_NS2_BEG[5] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS2_BEG6  (.A0(net119),
    .A1(net111),
    .A2(net171),
    .A3(net163),
    .S0(\ConfigBits[316] ),
    .S1(\ConfigBits[317] ),
    .X(\J_NS2_BEG[6] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS2_BEG7  (.A0(net120),
    .A1(net112),
    .A2(net172),
    .A3(net164),
    .S0(\ConfigBits[318] ),
    .S1(\ConfigBits[319] ),
    .X(\J_NS2_BEG[7] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG0  (.A0(net101),
    .A1(net121),
    .A2(net153),
    .A3(net173),
    .S0(\ConfigBits[272] ),
    .S1(\ConfigBits[273] ),
    .X(\J_NS4_BEG[0] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG1  (.A0(net102),
    .A1(net128),
    .A2(net154),
    .A3(net180),
    .S0(\ConfigBits[274] ),
    .S1(\ConfigBits[275] ),
    .X(\J_NS4_BEG[1] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG10  (.A0(net103),
    .A1(net129),
    .A2(net155),
    .A3(net181),
    .S0(\ConfigBits[292] ),
    .S1(\ConfigBits[293] ),
    .X(\J_NS4_BEG[10] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG11  (.A0(net104),
    .A1(net130),
    .A2(net156),
    .A3(net182),
    .S0(\ConfigBits[294] ),
    .S1(\ConfigBits[295] ),
    .X(\J_NS4_BEG[11] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG12  (.A0(net101),
    .A1(net121),
    .A2(net153),
    .A3(net173),
    .S0(\ConfigBits[296] ),
    .S1(\ConfigBits[297] ),
    .X(\J_NS4_BEG[12] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG13  (.A0(net102),
    .A1(net128),
    .A2(net154),
    .A3(net180),
    .S0(\ConfigBits[298] ),
    .S1(\ConfigBits[299] ),
    .X(\J_NS4_BEG[13] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG14  (.A0(net103),
    .A1(net129),
    .A2(net155),
    .A3(net181),
    .S0(\ConfigBits[300] ),
    .S1(\ConfigBits[301] ),
    .X(\J_NS4_BEG[14] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG15  (.A0(net104),
    .A1(net130),
    .A2(net156),
    .A3(net182),
    .S0(\ConfigBits[302] ),
    .S1(\ConfigBits[303] ),
    .X(\J_NS4_BEG[15] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG2  (.A0(net103),
    .A1(net129),
    .A2(net155),
    .A3(net181),
    .S0(\ConfigBits[276] ),
    .S1(\ConfigBits[277] ),
    .X(\J_NS4_BEG[2] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG3  (.A0(net104),
    .A1(net130),
    .A2(net156),
    .A3(net182),
    .S0(\ConfigBits[278] ),
    .S1(\ConfigBits[279] ),
    .X(\J_NS4_BEG[3] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG4  (.A0(net101),
    .A1(net121),
    .A2(net153),
    .A3(net173),
    .S0(\ConfigBits[280] ),
    .S1(\ConfigBits[281] ),
    .X(\J_NS4_BEG[4] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG5  (.A0(net102),
    .A1(net128),
    .A2(net154),
    .A3(net180),
    .S0(\ConfigBits[282] ),
    .S1(\ConfigBits[283] ),
    .X(\J_NS4_BEG[5] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG6  (.A0(net103),
    .A1(net129),
    .A2(net155),
    .A3(net181),
    .S0(\ConfigBits[284] ),
    .S1(\ConfigBits[285] ),
    .X(\J_NS4_BEG[6] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG7  (.A0(net104),
    .A1(net130),
    .A2(net156),
    .A3(net182),
    .S0(\ConfigBits[286] ),
    .S1(\ConfigBits[287] ),
    .X(\J_NS4_BEG[7] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG8  (.A0(net101),
    .A1(net121),
    .A2(net153),
    .A3(net173),
    .S0(\ConfigBits[288] ),
    .S1(\ConfigBits[289] ),
    .X(\J_NS4_BEG[8] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_J_NS4_BEG9  (.A0(net102),
    .A1(net128),
    .A2(net154),
    .A3(net180),
    .S0(\ConfigBits[290] ),
    .S1(\ConfigBits[291] ),
    .X(\J_NS4_BEG[9] ));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N1BEG0  (.A0(net1),
    .A1(net27),
    .A2(\J_NS4_BEG[12] ),
    .A3(\J_NS1_BEG[0] ),
    .S0(\ConfigBits[48] ),
    .S1(\ConfigBits[49] ),
    .X(net273));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N1BEG1  (.A0(net2),
    .A1(net28),
    .A2(\J_NS4_BEG[13] ),
    .A3(\J_NS1_BEG[1] ),
    .S0(\ConfigBits[50] ),
    .S1(\ConfigBits[51] ),
    .X(net274));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N1BEG2  (.A0(net3),
    .A1(net29),
    .A2(\J_NS4_BEG[14] ),
    .A3(\J_NS1_BEG[2] ),
    .S0(\ConfigBits[52] ),
    .S1(\ConfigBits[53] ),
    .X(net275));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N1BEG3  (.A0(net4),
    .A1(net30),
    .A2(\J_NS4_BEG[15] ),
    .A3(\J_NS1_BEG[3] ),
    .S0(\ConfigBits[54] ),
    .S1(\ConfigBits[55] ),
    .X(net276));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N2BEG0  (.A0(net20),
    .A1(net12),
    .A2(net30),
    .A3(\J_NS2_BEG[0] ),
    .S0(\ConfigBits[56] ),
    .S1(\ConfigBits[57] ),
    .X(net277));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N2BEG1  (.A0(net19),
    .A1(net11),
    .A2(net29),
    .A3(\J_NS2_BEG[1] ),
    .S0(\ConfigBits[58] ),
    .S1(\ConfigBits[59] ),
    .X(net278));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N2BEG2  (.A0(net18),
    .A1(net10),
    .A2(net28),
    .A3(\J_NS2_BEG[2] ),
    .S0(\ConfigBits[60] ),
    .S1(\ConfigBits[61] ),
    .X(net279));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N2BEG3  (.A0(net17),
    .A1(net9),
    .A2(net27),
    .A3(\J_NS2_BEG[3] ),
    .S0(\ConfigBits[62] ),
    .S1(\ConfigBits[63] ),
    .X(net280));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N2BEG4  (.A0(net16),
    .A1(net8),
    .A2(net26),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[64] ),
    .S1(\ConfigBits[65] ),
    .X(net281));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N2BEG5  (.A0(net15),
    .A1(net7),
    .A2(net25),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[66] ),
    .S1(\ConfigBits[67] ),
    .X(net282));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N2BEG6  (.A0(net14),
    .A1(net6),
    .A2(net24),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[68] ),
    .S1(\ConfigBits[69] ),
    .X(net283));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_N2BEG7  (.A0(net13),
    .A1(net5),
    .A2(net21),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[70] ),
    .S1(\ConfigBits[71] ),
    .X(net284));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S1BEG0  (.A0(net1),
    .A1(net31),
    .A2(\J_NS4_BEG[12] ),
    .A3(\J_NS1_BEG[0] ),
    .S0(\ConfigBits[84] ),
    .S1(\ConfigBits[85] ),
    .X(net309));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S1BEG1  (.A0(net2),
    .A1(net32),
    .A2(\J_NS4_BEG[13] ),
    .A3(\J_NS1_BEG[1] ),
    .S0(\ConfigBits[86] ),
    .S1(\ConfigBits[87] ),
    .X(net310));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S1BEG2  (.A0(net3),
    .A1(net22),
    .A2(\J_NS4_BEG[14] ),
    .A3(\J_NS1_BEG[2] ),
    .S0(\ConfigBits[88] ),
    .S1(\ConfigBits[89] ),
    .X(net311));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S1BEG3  (.A0(net4),
    .A1(net23),
    .A2(\J_NS4_BEG[15] ),
    .A3(\J_NS1_BEG[3] ),
    .S0(\ConfigBits[90] ),
    .S1(\ConfigBits[91] ),
    .X(net312));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S2BEG0  (.A0(net20),
    .A1(net12),
    .A2(net31),
    .A3(\J_NS2_BEG[0] ),
    .S0(\ConfigBits[92] ),
    .S1(\ConfigBits[93] ),
    .X(net313));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S2BEG1  (.A0(net19),
    .A1(net11),
    .A2(net32),
    .A3(\J_NS2_BEG[1] ),
    .S0(\ConfigBits[94] ),
    .S1(\ConfigBits[95] ),
    .X(net314));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S2BEG2  (.A0(net18),
    .A1(net10),
    .A2(net22),
    .A3(\J_NS2_BEG[2] ),
    .S0(\ConfigBits[96] ),
    .S1(\ConfigBits[97] ),
    .X(net315));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S2BEG3  (.A0(net17),
    .A1(net9),
    .A2(net23),
    .A3(\J_NS2_BEG[3] ),
    .S0(\ConfigBits[98] ),
    .S1(\ConfigBits[99] ),
    .X(net316));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S2BEG4  (.A0(net1),
    .A1(net16),
    .A2(net8),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[100] ),
    .S1(\ConfigBits[101] ),
    .X(net317));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S2BEG5  (.A0(net2),
    .A1(net15),
    .A2(net7),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[102] ),
    .S1(\ConfigBits[103] ),
    .X(net318));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S2BEG6  (.A0(net3),
    .A1(net14),
    .A2(net6),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[104] ),
    .S1(\ConfigBits[105] ),
    .X(net319));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_S2BEG7  (.A0(net4),
    .A1(net13),
    .A2(net5),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[106] ),
    .S1(\ConfigBits[107] ),
    .X(net320));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W1BEG0  (.A0(net101),
    .A1(net153),
    .A2(RAM2FAB_D0_O2),
    .A3(RAM2FAB_D1_O3),
    .S0(\ConfigBits[120] ),
    .S1(\ConfigBits[121] ),
    .X(net346));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W1BEG1  (.A0(net102),
    .A1(net154),
    .A2(RAM2FAB_D0_O3),
    .A3(RAM2FAB_D1_O2),
    .S0(\ConfigBits[122] ),
    .S1(\ConfigBits[123] ),
    .X(net347));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W1BEG2  (.A0(net103),
    .A1(net155),
    .A2(RAM2FAB_D0_O0),
    .A3(RAM2FAB_D1_O1),
    .S0(\ConfigBits[124] ),
    .S1(\ConfigBits[125] ),
    .X(net348));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W1BEG3  (.A0(net104),
    .A1(net156),
    .A2(RAM2FAB_D0_O1),
    .A3(RAM2FAB_D1_O0),
    .S0(\ConfigBits[126] ),
    .S1(\ConfigBits[127] ),
    .X(net349));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEG0  (.A0(RAM2FAB_D0_O0),
    .A1(RAM2FAB_D2_O0),
    .A2(\J_NS2_BEG[0] ),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[128] ),
    .S1(\ConfigBits[129] ),
    .X(net350));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEG1  (.A0(RAM2FAB_D0_O1),
    .A1(RAM2FAB_D2_O1),
    .A2(\J_NS2_BEG[1] ),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[130] ),
    .S1(\ConfigBits[131] ),
    .X(net351));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEG2  (.A0(RAM2FAB_D0_O2),
    .A1(RAM2FAB_D2_O2),
    .A2(\J_NS2_BEG[2] ),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[132] ),
    .S1(\ConfigBits[133] ),
    .X(net352));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEG3  (.A0(RAM2FAB_D0_O3),
    .A1(RAM2FAB_D2_O3),
    .A2(\J_NS2_BEG[3] ),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[134] ),
    .S1(\ConfigBits[135] ),
    .X(net353));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEG4  (.A0(RAM2FAB_D1_O0),
    .A1(RAM2FAB_D3_O0),
    .A2(\J_NS2_BEG[3] ),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[136] ),
    .S1(\ConfigBits[137] ),
    .X(net354));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEG5  (.A0(RAM2FAB_D1_O1),
    .A1(RAM2FAB_D3_O1),
    .A2(\J_NS2_BEG[2] ),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[138] ),
    .S1(\ConfigBits[139] ),
    .X(net355));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEG6  (.A0(RAM2FAB_D1_O2),
    .A1(RAM2FAB_D3_O2),
    .A2(\J_NS2_BEG[1] ),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[140] ),
    .S1(\ConfigBits[141] ),
    .X(net356));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEG7  (.A0(RAM2FAB_D1_O3),
    .A1(RAM2FAB_D3_O3),
    .A2(\J_NS2_BEG[0] ),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[142] ),
    .S1(\ConfigBits[143] ),
    .X(net357));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEGb0  (.A0(RAM2FAB_D0_O0),
    .A1(RAM2FAB_D2_O0),
    .A2(\J_NS2_BEG[0] ),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[144] ),
    .S1(\ConfigBits[145] ),
    .X(net358));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEGb1  (.A0(RAM2FAB_D0_O1),
    .A1(RAM2FAB_D2_O1),
    .A2(\J_NS2_BEG[1] ),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[146] ),
    .S1(\ConfigBits[147] ),
    .X(net359));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEGb2  (.A0(RAM2FAB_D0_O2),
    .A1(RAM2FAB_D2_O2),
    .A2(\J_NS2_BEG[2] ),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[148] ),
    .S1(\ConfigBits[149] ),
    .X(net360));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEGb3  (.A0(RAM2FAB_D0_O3),
    .A1(RAM2FAB_D2_O3),
    .A2(\J_NS2_BEG[3] ),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[150] ),
    .S1(\ConfigBits[151] ),
    .X(net361));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEGb4  (.A0(RAM2FAB_D1_O0),
    .A1(RAM2FAB_D3_O0),
    .A2(\J_NS2_BEG[3] ),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[152] ),
    .S1(\ConfigBits[153] ),
    .X(net362));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEGb5  (.A0(RAM2FAB_D1_O1),
    .A1(RAM2FAB_D3_O1),
    .A2(\J_NS2_BEG[2] ),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[154] ),
    .S1(\ConfigBits[155] ),
    .X(net363));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEGb6  (.A0(RAM2FAB_D1_O2),
    .A1(RAM2FAB_D3_O2),
    .A2(\J_NS2_BEG[1] ),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[156] ),
    .S1(\ConfigBits[157] ),
    .X(net364));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W2BEGb7  (.A0(RAM2FAB_D1_O3),
    .A1(RAM2FAB_D3_O3),
    .A2(\J_NS2_BEG[0] ),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[158] ),
    .S1(\ConfigBits[159] ),
    .X(net365));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG0  (.A0(net121),
    .A1(net173),
    .A2(\J_NS4_BEG[11] ),
    .A3(\J_NS4_BEG[15] ),
    .S0(\ConfigBits[192] ),
    .S1(\ConfigBits[193] ),
    .X(net366));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG1  (.A0(net128),
    .A1(net180),
    .A2(\J_NS4_BEG[10] ),
    .A3(\J_NS4_BEG[14] ),
    .S0(\ConfigBits[194] ),
    .S1(\ConfigBits[195] ),
    .X(net369));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG10  (.A0(RAM2FAB_D0_O2),
    .A1(\J_NS4_BEG[1] ),
    .A2(\J_NS4_BEG[5] ),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[212] ),
    .S1(\ConfigBits[213] ),
    .X(net367));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG11  (.A0(RAM2FAB_D0_O3),
    .A1(\J_NS4_BEG[0] ),
    .A2(\J_NS4_BEG[4] ),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[214] ),
    .S1(\ConfigBits[215] ),
    .X(net368));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG2  (.A0(net129),
    .A1(net181),
    .A2(\J_NS4_BEG[9] ),
    .A3(\J_NS4_BEG[13] ),
    .S0(\ConfigBits[196] ),
    .S1(\ConfigBits[197] ),
    .X(net370));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG3  (.A0(net130),
    .A1(net182),
    .A2(\J_NS4_BEG[8] ),
    .A3(\J_NS4_BEG[12] ),
    .S0(\ConfigBits[198] ),
    .S1(\ConfigBits[199] ),
    .X(net371));
 sky130_fd_sc_hd__mux4_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG4  (.A0(RAM2FAB_D1_O0),
    .A1(\J_NS4_BEG[7] ),
    .A2(\J_NS4_BEG[11] ),
    .A3(\J_NS2_BEG[0] ),
    .S0(\ConfigBits[200] ),
    .S1(\ConfigBits[201] ),
    .X(net372));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG5  (.A0(RAM2FAB_D1_O1),
    .A1(\J_NS4_BEG[6] ),
    .A2(\J_NS4_BEG[10] ),
    .A3(\J_NS2_BEG[1] ),
    .S0(\ConfigBits[202] ),
    .S1(\ConfigBits[203] ),
    .X(net373));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG6  (.A0(RAM2FAB_D1_O2),
    .A1(\J_NS4_BEG[5] ),
    .A2(\J_NS4_BEG[9] ),
    .A3(\J_NS2_BEG[2] ),
    .S0(\ConfigBits[204] ),
    .S1(\ConfigBits[205] ),
    .X(net374));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG7  (.A0(RAM2FAB_D1_O3),
    .A1(\J_NS4_BEG[4] ),
    .A2(\J_NS4_BEG[8] ),
    .A3(\J_NS2_BEG[3] ),
    .S0(\ConfigBits[206] ),
    .S1(\ConfigBits[207] ),
    .X(net375));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG8  (.A0(RAM2FAB_D0_O0),
    .A1(\J_NS4_BEG[3] ),
    .A2(\J_NS4_BEG[7] ),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[208] ),
    .S1(\ConfigBits[209] ),
    .X(net376));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_W6BEG9  (.A0(RAM2FAB_D0_O1),
    .A1(\J_NS4_BEG[2] ),
    .A2(\J_NS4_BEG[6] ),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[210] ),
    .S1(\ConfigBits[211] ),
    .X(net377));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG0  (.A0(RAM2FAB_D0_O0),
    .A1(RAM2FAB_D3_O0),
    .A2(\J_NS4_BEG[15] ),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[160] ),
    .S1(\ConfigBits[161] ),
    .X(net378));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG1  (.A0(RAM2FAB_D0_O1),
    .A1(RAM2FAB_D3_O1),
    .A2(\J_NS4_BEG[14] ),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[162] ),
    .S1(\ConfigBits[163] ),
    .X(net385));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG10  (.A0(RAM2FAB_D1_O2),
    .A1(RAM2FAB_D2_O2),
    .A2(\J_NS4_BEG[5] ),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[180] ),
    .S1(\ConfigBits[181] ),
    .X(net379));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG11  (.A0(RAM2FAB_D1_O3),
    .A1(RAM2FAB_D2_O3),
    .A2(\J_NS4_BEG[4] ),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[182] ),
    .S1(\ConfigBits[183] ),
    .X(net380));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG12  (.A0(RAM2FAB_D0_O0),
    .A1(RAM2FAB_D3_O0),
    .A2(\J_NS4_BEG[3] ),
    .A3(\J_NS2_BEG[3] ),
    .S0(\ConfigBits[184] ),
    .S1(\ConfigBits[185] ),
    .X(net381));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG13  (.A0(RAM2FAB_D0_O1),
    .A1(RAM2FAB_D3_O1),
    .A2(\J_NS4_BEG[2] ),
    .A3(\J_NS2_BEG[2] ),
    .S0(\ConfigBits[186] ),
    .S1(\ConfigBits[187] ),
    .X(net382));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG14  (.A0(RAM2FAB_D0_O2),
    .A1(RAM2FAB_D3_O2),
    .A2(\J_NS4_BEG[1] ),
    .A3(\J_NS2_BEG[1] ),
    .S0(\ConfigBits[188] ),
    .S1(\ConfigBits[189] ),
    .X(net383));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG15  (.A0(RAM2FAB_D0_O3),
    .A1(RAM2FAB_D3_O3),
    .A2(\J_NS4_BEG[0] ),
    .A3(\J_NS2_BEG[0] ),
    .S0(\ConfigBits[190] ),
    .S1(\ConfigBits[191] ),
    .X(net384));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG2  (.A0(RAM2FAB_D0_O2),
    .A1(RAM2FAB_D3_O2),
    .A2(\J_NS4_BEG[13] ),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[164] ),
    .S1(\ConfigBits[165] ),
    .X(net386));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG3  (.A0(RAM2FAB_D0_O3),
    .A1(RAM2FAB_D3_O3),
    .A2(\J_NS4_BEG[12] ),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[166] ),
    .S1(\ConfigBits[167] ),
    .X(net387));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG4  (.A0(RAM2FAB_D1_O0),
    .A1(RAM2FAB_D2_O0),
    .A2(\J_NS4_BEG[11] ),
    .A3(\J_NS2_BEG[3] ),
    .S0(\ConfigBits[168] ),
    .S1(\ConfigBits[169] ),
    .X(net388));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG5  (.A0(RAM2FAB_D1_O1),
    .A1(RAM2FAB_D2_O1),
    .A2(\J_NS4_BEG[10] ),
    .A3(\J_NS2_BEG[2] ),
    .S0(\ConfigBits[170] ),
    .S1(\ConfigBits[171] ),
    .X(net389));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG6  (.A0(RAM2FAB_D1_O2),
    .A1(RAM2FAB_D2_O2),
    .A2(\J_NS4_BEG[9] ),
    .A3(\J_NS2_BEG[1] ),
    .S0(\ConfigBits[172] ),
    .S1(\ConfigBits[173] ),
    .X(net390));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG7  (.A0(RAM2FAB_D1_O3),
    .A1(RAM2FAB_D2_O3),
    .A2(\J_NS4_BEG[8] ),
    .A3(\J_NS2_BEG[0] ),
    .S0(\ConfigBits[174] ),
    .S1(\ConfigBits[175] ),
    .X(net391));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG8  (.A0(RAM2FAB_D1_O0),
    .A1(RAM2FAB_D2_O0),
    .A2(\J_NS4_BEG[7] ),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[176] ),
    .S1(\ConfigBits[177] ),
    .X(net392));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux41_buf_WW4BEG9  (.A0(RAM2FAB_D1_O1),
    .A1(RAM2FAB_D2_O1),
    .A2(\J_NS4_BEG[6] ),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[178] ),
    .S1(\ConfigBits[179] ),
    .X(net393));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_2_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_3_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[74] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_4_  (.A1(\ConfigBits[74] ),
    .A2(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_0_ ),
    .B1(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_1_ ),
    .Y(net296));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_out0 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_out1 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_inst0  (.A0(net1),
    .A1(net33),
    .A2(net31),
    .A3(\J_NS4_BEG[0] ),
    .S0(\ConfigBits[72] ),
    .S1(\ConfigBits[73] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_inst1  (.A0(\J_NS4_BEG[4] ),
    .A1(\J_NS4_BEG[8] ),
    .A2(\J_NS4_BEG[12] ),
    .A3(\J_NS2_BEG[0] ),
    .S0(\ConfigBits[72] ),
    .S1(\ConfigBits[73] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_2_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_3_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[77] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_4_  (.A1(\ConfigBits[77] ),
    .A2(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_0_ ),
    .B1(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_1_ ),
    .Y(net297));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_out0 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_out1 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_inst0  (.A0(net2),
    .A1(net40),
    .A2(net32),
    .A3(\J_NS4_BEG[1] ),
    .S0(\ConfigBits[75] ),
    .S1(\ConfigBits[76] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_inst1  (.A0(\J_NS4_BEG[5] ),
    .A1(\J_NS4_BEG[9] ),
    .A2(\J_NS4_BEG[13] ),
    .A3(\J_NS2_BEG[1] ),
    .S0(\ConfigBits[75] ),
    .S1(\ConfigBits[76] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_2_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_3_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[80] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_4_  (.A1(\ConfigBits[80] ),
    .A2(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_0_ ),
    .B1(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_1_ ),
    .Y(net298));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_out0 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_out1 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_inst0  (.A0(net3),
    .A1(net41),
    .A2(net22),
    .A3(\J_NS4_BEG[2] ),
    .S0(\ConfigBits[78] ),
    .S1(\ConfigBits[79] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_inst1  (.A0(\J_NS4_BEG[6] ),
    .A1(\J_NS4_BEG[10] ),
    .A2(\J_NS4_BEG[14] ),
    .A3(\J_NS2_BEG[2] ),
    .S0(\ConfigBits[78] ),
    .S1(\ConfigBits[79] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_2_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_3_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[83] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_4_  (.A1(\ConfigBits[83] ),
    .A2(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_0_ ),
    .B1(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_1_ ),
    .Y(net299));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_out0 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_out1 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_inst0  (.A0(net4),
    .A1(net42),
    .A2(net23),
    .A3(\J_NS4_BEG[3] ),
    .S0(\ConfigBits[81] ),
    .S1(\ConfigBits[82] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_inst1  (.A0(\J_NS4_BEG[7] ),
    .A1(\J_NS4_BEG[11] ),
    .A2(\J_NS4_BEG[15] ),
    .A3(\J_NS2_BEG[3] ),
    .S0(\ConfigBits[81] ),
    .S1(\ConfigBits[82] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_2_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_3_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[110] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_4_  (.A1(\ConfigBits[110] ),
    .A2(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_0_ ),
    .B1(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_1_ ),
    .Y(net332));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_out0 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_out1 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_inst0  (.A0(net1),
    .A1(net36),
    .A2(net27),
    .A3(\J_NS4_BEG[0] ),
    .S0(\ConfigBits[108] ),
    .S1(\ConfigBits[109] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_inst1  (.A0(\J_NS4_BEG[4] ),
    .A1(\J_NS4_BEG[8] ),
    .A2(\J_NS4_BEG[12] ),
    .A3(\J_NS2_BEG[4] ),
    .S0(\ConfigBits[108] ),
    .S1(\ConfigBits[109] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_2_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_3_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[113] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_4_  (.A1(\ConfigBits[113] ),
    .A2(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_0_ ),
    .B1(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_1_ ),
    .Y(net333));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_out0 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_out1 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_inst0  (.A0(net2),
    .A1(net37),
    .A2(net28),
    .A3(\J_NS4_BEG[1] ),
    .S0(\ConfigBits[111] ),
    .S1(\ConfigBits[112] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_inst1  (.A0(\J_NS4_BEG[5] ),
    .A1(\J_NS4_BEG[9] ),
    .A2(\J_NS4_BEG[13] ),
    .A3(\J_NS2_BEG[5] ),
    .S0(\ConfigBits[111] ),
    .S1(\ConfigBits[112] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_2_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_3_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[116] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_4_  (.A1(\ConfigBits[116] ),
    .A2(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_0_ ),
    .B1(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_1_ ),
    .Y(net334));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_out0 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_out1 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_inst0  (.A0(net3),
    .A1(net38),
    .A2(net29),
    .A3(\J_NS4_BEG[2] ),
    .S0(\ConfigBits[114] ),
    .S1(\ConfigBits[115] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_inst1  (.A0(\J_NS4_BEG[6] ),
    .A1(\J_NS4_BEG[10] ),
    .A2(\J_NS4_BEG[14] ),
    .A3(\J_NS2_BEG[6] ),
    .S0(\ConfigBits[114] ),
    .S1(\ConfigBits[115] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__inv_2 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_2_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/AIN[0] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_0_ ));
 sky130_fd_sc_hd__nand2_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_3_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/AIN[1] ),
    .B(\ConfigBits[119] ),
    .Y(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_1_ ));
 sky130_fd_sc_hd__o21ai_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_4_  (.A1(\ConfigBits[119] ),
    .A2(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_0_ ),
    .B1(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_1_ ),
    .Y(net335));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/break_comb_loop_inst0/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_out0 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/AIN[0] ));
 sky130_fd_sc_hd__clkbuf_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/break_comb_loop_inst1/_0_  (.A(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_out1 ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/AIN[1] ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_inst0  (.A0(net4),
    .A1(net39),
    .A2(net30),
    .A3(\J_NS4_BEG[3] ),
    .S0(\ConfigBits[117] ),
    .S1(\ConfigBits[118] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_out0 ));
 sky130_fd_sc_hd__mux4_1 \Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_inst1  (.A0(\J_NS4_BEG[7] ),
    .A1(\J_NS4_BEG[11] ),
    .A2(\J_NS4_BEG[15] ),
    .A3(\J_NS2_BEG[7] ),
    .S0(\ConfigBits[117] ),
    .S1(\ConfigBits[118] ),
    .X(\Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_out1 ));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_0/_0_  (.A(\N4BEG_i[0] ),
    .X(net293));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_1/_0_  (.A(\N4BEG_i[1] ),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_10/_0_  (.A(\N4BEG_i[10] ),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_11/_0_  (.A(\N4BEG_i[11] ),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_2/_0_  (.A(\N4BEG_i[2] ),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_3/_0_  (.A(\N4BEG_i[3] ),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_4/_0_  (.A(\N4BEG_i[4] ),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_5/_0_  (.A(\N4BEG_i[5] ),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_6/_0_  (.A(\N4BEG_i[6] ),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_7/_0_  (.A(\N4BEG_i[7] ),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_8/_0_  (.A(\N4BEG_i[8] ),
    .X(net307));
 sky130_fd_sc_hd__clkbuf_1 \N4BEG_outbuf_9/_0_  (.A(\N4BEG_i[9] ),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_0/_0_  (.A(net131),
    .X(\N4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_1/_0_  (.A(net132),
    .X(\N4BEG_i[1] ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_10/_0_  (.A(net126),
    .X(\N4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_11/_0_  (.A(net127),
    .X(\N4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_2/_0_  (.A(net133),
    .X(\N4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_3/_0_  (.A(net134),
    .X(\N4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_4/_0_  (.A(net135),
    .X(\N4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_5/_0_  (.A(net136),
    .X(\N4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_6/_0_  (.A(net122),
    .X(\N4BEG_i[6] ));
 sky130_fd_sc_hd__buf_2 \N4END_inbuf_7/_0_  (.A(net123),
    .X(\N4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_8/_0_  (.A(net124),
    .X(\N4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \N4END_inbuf_9/_0_  (.A(net125),
    .X(\N4BEG_i[9] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_0/_0_  (.A(\S4BEG_i[0] ),
    .X(net329));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_1/_0_  (.A(\S4BEG_i[1] ),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_10/_0_  (.A(\S4BEG_i[10] ),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_11/_0_  (.A(\S4BEG_i[11] ),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_2/_0_  (.A(\S4BEG_i[2] ),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_3/_0_  (.A(\S4BEG_i[3] ),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_4/_0_  (.A(\S4BEG_i[4] ),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_5/_0_  (.A(\S4BEG_i[5] ),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_6/_0_  (.A(\S4BEG_i[6] ),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_7/_0_  (.A(\S4BEG_i[7] ),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_8/_0_  (.A(\S4BEG_i[8] ),
    .X(net343));
 sky130_fd_sc_hd__clkbuf_1 \S4BEG_outbuf_9/_0_  (.A(\S4BEG_i[9] ),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_0/_0_  (.A(net183),
    .X(\S4BEG_i[0] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_1/_0_  (.A(net184),
    .X(\S4BEG_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_10/_0_  (.A(net178),
    .X(\S4BEG_i[10] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_11/_0_  (.A(net179),
    .X(\S4BEG_i[11] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_2/_0_  (.A(net185),
    .X(\S4BEG_i[2] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_3/_0_  (.A(net186),
    .X(\S4BEG_i[3] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_4/_0_  (.A(net187),
    .X(\S4BEG_i[4] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_5/_0_  (.A(net188),
    .X(\S4BEG_i[5] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_6/_0_  (.A(net174),
    .X(\S4BEG_i[6] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_7/_0_  (.A(net175),
    .X(\S4BEG_i[7] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_8/_0_  (.A(net176),
    .X(\S4BEG_i[8] ));
 sky130_fd_sc_hd__clkbuf_2 \S4END_inbuf_9/_0_  (.A(net177),
    .X(\S4BEG_i[9] ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_0/_0_  (.A(net49),
    .X(\FrameData_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_1/_0_  (.A(net60),
    .X(\FrameData_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_10/_0_  (.A(net50),
    .X(\FrameData_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_11/_0_  (.A(net51),
    .X(\FrameData_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_12/_0_  (.A(net52),
    .X(\FrameData_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_13/_0_  (.A(net53),
    .X(\FrameData_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_14/_0_  (.A(net54),
    .X(\FrameData_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_15/_0_  (.A(net55),
    .X(\FrameData_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_16/_0_  (.A(net56),
    .X(\FrameData_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_17/_0_  (.A(net57),
    .X(\FrameData_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_18/_0_  (.A(net58),
    .X(\FrameData_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_19/_0_  (.A(net59),
    .X(\FrameData_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_2/_0_  (.A(net71),
    .X(\FrameData_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_20/_0_  (.A(net61),
    .X(\FrameData_O_i[20] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_21/_0_  (.A(net62),
    .X(\FrameData_O_i[21] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_22/_0_  (.A(net63),
    .X(\FrameData_O_i[22] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_23/_0_  (.A(net64),
    .X(\FrameData_O_i[23] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_24/_0_  (.A(net65),
    .X(\FrameData_O_i[24] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_25/_0_  (.A(net66),
    .X(\FrameData_O_i[25] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_26/_0_  (.A(net67),
    .X(\FrameData_O_i[26] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_27/_0_  (.A(net68),
    .X(\FrameData_O_i[27] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_28/_0_  (.A(net69),
    .X(\FrameData_O_i[28] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_29/_0_  (.A(net70),
    .X(\FrameData_O_i[29] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_3/_0_  (.A(net74),
    .X(\FrameData_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_30/_0_  (.A(net72),
    .X(\FrameData_O_i[30] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_31/_0_  (.A(net73),
    .X(\FrameData_O_i[31] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_4/_0_  (.A(net75),
    .X(\FrameData_O_i[4] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_5/_0_  (.A(net76),
    .X(\FrameData_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_6/_0_  (.A(net77),
    .X(\FrameData_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_7/_0_  (.A(net78),
    .X(\FrameData_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_8/_0_  (.A(net79),
    .X(\FrameData_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \data_inbuf_9/_0_  (.A(net80),
    .X(\FrameData_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_0/_0_  (.A(\FrameData_O_i[0] ),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_1/_0_  (.A(\FrameData_O_i[1] ),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_10/_0_  (.A(\FrameData_O_i[10] ),
    .X(net222));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_11/_0_  (.A(\FrameData_O_i[11] ),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_12/_0_  (.A(\FrameData_O_i[12] ),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_13/_0_  (.A(\FrameData_O_i[13] ),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_14/_0_  (.A(\FrameData_O_i[14] ),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_15/_0_  (.A(\FrameData_O_i[15] ),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_16/_0_  (.A(\FrameData_O_i[16] ),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_17/_0_  (.A(\FrameData_O_i[17] ),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_18/_0_  (.A(\FrameData_O_i[18] ),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_19/_0_  (.A(\FrameData_O_i[19] ),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_2/_0_  (.A(\FrameData_O_i[2] ),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_20/_0_  (.A(\FrameData_O_i[20] ),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_21/_0_  (.A(\FrameData_O_i[21] ),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_22/_0_  (.A(\FrameData_O_i[22] ),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_23/_0_  (.A(\FrameData_O_i[23] ),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_24/_0_  (.A(\FrameData_O_i[24] ),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_25/_0_  (.A(\FrameData_O_i[25] ),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_26/_0_  (.A(\FrameData_O_i[26] ),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_27/_0_  (.A(\FrameData_O_i[27] ),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_28/_0_  (.A(\FrameData_O_i[28] ),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_29/_0_  (.A(\FrameData_O_i[29] ),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_3/_0_  (.A(\FrameData_O_i[3] ),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_30/_0_  (.A(\FrameData_O_i[30] ),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_31/_0_  (.A(\FrameData_O_i[31] ),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_4/_0_  (.A(\FrameData_O_i[4] ),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_5/_0_  (.A(\FrameData_O_i[5] ),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_6/_0_  (.A(\FrameData_O_i[6] ),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_7/_0_  (.A(\FrameData_O_i[7] ),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_8/_0_  (.A(\FrameData_O_i[8] ),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 \data_outbuf_9/_0_  (.A(\FrameData_O_i[9] ),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(E1END[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(E2END[5]),
    .X(net10));
 sky130_fd_sc_hd__buf_8 input100 (.A(FrameStrobe[9]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_2 input101 (.A(N1END[0]),
    .X(net101));
 sky130_fd_sc_hd__buf_2 input102 (.A(N1END[1]),
    .X(net102));
 sky130_fd_sc_hd__buf_2 input103 (.A(N1END[2]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 input104 (.A(N1END[3]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(N2END[0]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(N2END[1]),
    .X(net106));
 sky130_fd_sc_hd__dlymetal6s2s_1 input107 (.A(N2END[2]),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 input108 (.A(N2END[3]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_1 input109 (.A(N2END[4]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(E2END[6]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input110 (.A(N2END[5]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 input111 (.A(N2END[6]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(N2END[7]),
    .X(net112));
 sky130_fd_sc_hd__buf_1 input113 (.A(N2MID[0]),
    .X(net113));
 sky130_fd_sc_hd__buf_2 input114 (.A(N2MID[1]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(N2MID[2]),
    .X(net115));
 sky130_fd_sc_hd__clkbuf_2 input116 (.A(N2MID[3]),
    .X(net116));
 sky130_fd_sc_hd__buf_1 input117 (.A(N2MID[4]),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(N2MID[5]),
    .X(net118));
 sky130_fd_sc_hd__buf_2 input119 (.A(N2MID[6]),
    .X(net119));
 sky130_fd_sc_hd__buf_1 input12 (.A(E2END[7]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input120 (.A(N2MID[7]),
    .X(net120));
 sky130_fd_sc_hd__dlymetal6s2s_1 input121 (.A(N4END[0]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(N4END[10]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(N4END[11]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(N4END[12]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(N4END[13]),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 input126 (.A(N4END[14]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 input127 (.A(N4END[15]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(N4END[1]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_2 input129 (.A(N4END[2]),
    .X(net129));
 sky130_fd_sc_hd__buf_1 input13 (.A(E2MID[0]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input130 (.A(N4END[3]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 input131 (.A(N4END[4]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 input132 (.A(N4END[5]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 input133 (.A(N4END[6]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 input134 (.A(N4END[7]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(N4END[8]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(N4END[9]),
    .X(net136));
 sky130_fd_sc_hd__buf_1 input137 (.A(RAM2FAB_D0_I0),
    .X(net137));
 sky130_fd_sc_hd__buf_1 input138 (.A(RAM2FAB_D0_I1),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 input139 (.A(RAM2FAB_D0_I2),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(E2MID[1]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input140 (.A(RAM2FAB_D0_I3),
    .X(net140));
 sky130_fd_sc_hd__buf_1 input141 (.A(RAM2FAB_D1_I0),
    .X(net141));
 sky130_fd_sc_hd__buf_1 input142 (.A(RAM2FAB_D1_I1),
    .X(net142));
 sky130_fd_sc_hd__buf_1 input143 (.A(RAM2FAB_D1_I2),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(RAM2FAB_D1_I3),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(RAM2FAB_D2_I0),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(RAM2FAB_D2_I1),
    .X(net146));
 sky130_fd_sc_hd__buf_1 input147 (.A(RAM2FAB_D2_I2),
    .X(net147));
 sky130_fd_sc_hd__buf_1 input148 (.A(RAM2FAB_D2_I3),
    .X(net148));
 sky130_fd_sc_hd__buf_1 input149 (.A(RAM2FAB_D3_I0),
    .X(net149));
 sky130_fd_sc_hd__buf_1 input15 (.A(E2MID[2]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input150 (.A(RAM2FAB_D3_I1),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(RAM2FAB_D3_I2),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 input152 (.A(RAM2FAB_D3_I3),
    .X(net152));
 sky130_fd_sc_hd__buf_2 input153 (.A(S1END[0]),
    .X(net153));
 sky130_fd_sc_hd__buf_2 input154 (.A(S1END[1]),
    .X(net154));
 sky130_fd_sc_hd__buf_2 input155 (.A(S1END[2]),
    .X(net155));
 sky130_fd_sc_hd__buf_2 input156 (.A(S1END[3]),
    .X(net156));
 sky130_fd_sc_hd__buf_2 input157 (.A(S2END[0]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 input158 (.A(S2END[1]),
    .X(net158));
 sky130_fd_sc_hd__buf_1 input159 (.A(S2END[2]),
    .X(net159));
 sky130_fd_sc_hd__buf_1 input16 (.A(E2MID[3]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input160 (.A(S2END[3]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 input161 (.A(S2END[4]),
    .X(net161));
 sky130_fd_sc_hd__buf_1 input162 (.A(S2END[5]),
    .X(net162));
 sky130_fd_sc_hd__buf_1 input163 (.A(S2END[6]),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_2 input164 (.A(S2END[7]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 input165 (.A(S2MID[0]),
    .X(net165));
 sky130_fd_sc_hd__buf_1 input166 (.A(S2MID[1]),
    .X(net166));
 sky130_fd_sc_hd__buf_1 input167 (.A(S2MID[2]),
    .X(net167));
 sky130_fd_sc_hd__buf_1 input168 (.A(S2MID[3]),
    .X(net168));
 sky130_fd_sc_hd__buf_2 input169 (.A(S2MID[4]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(E2MID[4]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input170 (.A(S2MID[5]),
    .X(net170));
 sky130_fd_sc_hd__buf_1 input171 (.A(S2MID[6]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_2 input172 (.A(S2MID[7]),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(S4END[0]),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 input174 (.A(S4END[10]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(S4END[11]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(S4END[12]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(S4END[13]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 input178 (.A(S4END[14]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 input179 (.A(S4END[15]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(E2MID[5]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input180 (.A(S4END[1]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(S4END[2]),
    .X(net181));
 sky130_fd_sc_hd__buf_2 input182 (.A(S4END[3]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 input183 (.A(S4END[4]),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 input184 (.A(S4END[5]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 input185 (.A(S4END[6]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 input186 (.A(S4END[7]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 input187 (.A(S4END[8]),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 input188 (.A(S4END[9]),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(E2MID[6]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input2 (.A(E1END[1]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(E2MID[7]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(E6END[0]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(E6END[10]),
    .X(net22));
 sky130_fd_sc_hd__buf_1 input23 (.A(E6END[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(E6END[1]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(E6END[2]),
    .X(net25));
 sky130_fd_sc_hd__dlymetal6s2s_1 input26 (.A(E6END[3]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(E6END[4]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(E6END[5]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(E6END[6]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(E1END[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(E6END[7]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(E6END[8]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(E6END[9]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(EE4END[0]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(EE4END[10]),
    .X(net34));
 sky130_fd_sc_hd__buf_1 input35 (.A(EE4END[11]),
    .X(net35));
 sky130_fd_sc_hd__buf_1 input36 (.A(EE4END[12]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(EE4END[13]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(EE4END[14]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(EE4END[15]),
    .X(net39));
 sky130_fd_sc_hd__buf_2 input4 (.A(E1END[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(EE4END[1]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(EE4END[2]),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(EE4END[3]),
    .X(net42));
 sky130_fd_sc_hd__buf_1 input43 (.A(EE4END[4]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(EE4END[5]),
    .X(net44));
 sky130_fd_sc_hd__buf_1 input45 (.A(EE4END[6]),
    .X(net45));
 sky130_fd_sc_hd__buf_1 input46 (.A(EE4END[7]),
    .X(net46));
 sky130_fd_sc_hd__buf_1 input47 (.A(EE4END[8]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(EE4END[9]),
    .X(net48));
 sky130_fd_sc_hd__buf_4 input49 (.A(FrameData[0]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(E2END[0]),
    .X(net5));
 sky130_fd_sc_hd__buf_4 input50 (.A(FrameData[10]),
    .X(net50));
 sky130_fd_sc_hd__buf_4 input51 (.A(FrameData[11]),
    .X(net51));
 sky130_fd_sc_hd__buf_4 input52 (.A(FrameData[12]),
    .X(net52));
 sky130_fd_sc_hd__buf_4 input53 (.A(FrameData[13]),
    .X(net53));
 sky130_fd_sc_hd__buf_4 input54 (.A(FrameData[14]),
    .X(net54));
 sky130_fd_sc_hd__buf_4 input55 (.A(FrameData[15]),
    .X(net55));
 sky130_fd_sc_hd__buf_4 input56 (.A(FrameData[16]),
    .X(net56));
 sky130_fd_sc_hd__buf_4 input57 (.A(FrameData[17]),
    .X(net57));
 sky130_fd_sc_hd__buf_4 input58 (.A(FrameData[18]),
    .X(net58));
 sky130_fd_sc_hd__buf_4 input59 (.A(FrameData[19]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(E2END[1]),
    .X(net6));
 sky130_fd_sc_hd__buf_4 input60 (.A(FrameData[1]),
    .X(net60));
 sky130_fd_sc_hd__buf_4 input61 (.A(FrameData[20]),
    .X(net61));
 sky130_fd_sc_hd__buf_4 input62 (.A(FrameData[21]),
    .X(net62));
 sky130_fd_sc_hd__buf_4 input63 (.A(FrameData[22]),
    .X(net63));
 sky130_fd_sc_hd__buf_4 input64 (.A(FrameData[23]),
    .X(net64));
 sky130_fd_sc_hd__buf_4 input65 (.A(FrameData[24]),
    .X(net65));
 sky130_fd_sc_hd__buf_4 input66 (.A(FrameData[25]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_8 input67 (.A(FrameData[26]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_8 input68 (.A(FrameData[27]),
    .X(net68));
 sky130_fd_sc_hd__buf_4 input69 (.A(FrameData[28]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input7 (.A(E2END[2]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input70 (.A(FrameData[29]),
    .X(net70));
 sky130_fd_sc_hd__buf_4 input71 (.A(FrameData[2]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_8 input72 (.A(FrameData[30]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_8 input73 (.A(FrameData[31]),
    .X(net73));
 sky130_fd_sc_hd__buf_4 input74 (.A(FrameData[3]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_8 input75 (.A(FrameData[4]),
    .X(net75));
 sky130_fd_sc_hd__buf_4 input76 (.A(FrameData[5]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_8 input77 (.A(FrameData[6]),
    .X(net77));
 sky130_fd_sc_hd__buf_4 input78 (.A(FrameData[7]),
    .X(net78));
 sky130_fd_sc_hd__buf_4 input79 (.A(FrameData[8]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input8 (.A(E2END[3]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input80 (.A(FrameData[9]),
    .X(net80));
 sky130_fd_sc_hd__buf_8 input81 (.A(FrameStrobe[0]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input82 (.A(FrameStrobe[10]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(FrameStrobe[11]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_2 input84 (.A(FrameStrobe[12]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(FrameStrobe[13]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(FrameStrobe[14]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(FrameStrobe[15]),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(FrameStrobe[16]),
    .X(net88));
 sky130_fd_sc_hd__dlymetal6s2s_1 input89 (.A(FrameStrobe[17]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(E2END[4]),
    .X(net9));
 sky130_fd_sc_hd__dlymetal6s2s_1 input90 (.A(FrameStrobe[18]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 input91 (.A(FrameStrobe[19]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_16 input92 (.A(FrameStrobe[1]),
    .X(net92));
 sky130_fd_sc_hd__buf_8 input93 (.A(FrameStrobe[2]),
    .X(net93));
 sky130_fd_sc_hd__buf_8 input94 (.A(FrameStrobe[3]),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_16 input95 (.A(FrameStrobe[4]),
    .X(net95));
 sky130_fd_sc_hd__buf_8 input96 (.A(FrameStrobe[5]),
    .X(net96));
 sky130_fd_sc_hd__buf_8 input97 (.A(FrameStrobe[6]),
    .X(net97));
 sky130_fd_sc_hd__buf_8 input98 (.A(FrameStrobe[7]),
    .X(net98));
 sky130_fd_sc_hd__buf_8 input99 (.A(FrameStrobe[8]),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_16 inst_clk_buf (.A(UserCLK),
    .X(net345));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(Config_accessC_bit0));
 sky130_fd_sc_hd__clkbuf_4 output190 (.A(net190),
    .X(Config_accessC_bit1));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(Config_accessC_bit2));
 sky130_fd_sc_hd__clkbuf_4 output192 (.A(net192),
    .X(Config_accessC_bit3));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(FAB2RAM_A0_O0));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(FAB2RAM_A0_O1));
 sky130_fd_sc_hd__clkbuf_4 output195 (.A(net195),
    .X(FAB2RAM_A0_O2));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(FAB2RAM_A0_O3));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(FAB2RAM_A1_O0));
 sky130_fd_sc_hd__clkbuf_4 output198 (.A(net198),
    .X(FAB2RAM_A1_O1));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(FAB2RAM_A1_O2));
 sky130_fd_sc_hd__clkbuf_4 output200 (.A(net200),
    .X(FAB2RAM_A1_O3));
 sky130_fd_sc_hd__clkbuf_4 output201 (.A(net201),
    .X(FAB2RAM_C_O0));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(FAB2RAM_C_O1));
 sky130_fd_sc_hd__clkbuf_4 output203 (.A(net203),
    .X(FAB2RAM_C_O2));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(FAB2RAM_C_O3));
 sky130_fd_sc_hd__clkbuf_4 output205 (.A(net205),
    .X(FAB2RAM_D0_O0));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(FAB2RAM_D0_O1));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(FAB2RAM_D0_O2));
 sky130_fd_sc_hd__clkbuf_4 output208 (.A(net208),
    .X(FAB2RAM_D0_O3));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(FAB2RAM_D1_O0));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(FAB2RAM_D1_O1));
 sky130_fd_sc_hd__clkbuf_4 output211 (.A(net211),
    .X(FAB2RAM_D1_O2));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(FAB2RAM_D1_O3));
 sky130_fd_sc_hd__clkbuf_4 output213 (.A(net213),
    .X(FAB2RAM_D2_O0));
 sky130_fd_sc_hd__clkbuf_4 output214 (.A(net214),
    .X(FAB2RAM_D2_O1));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(FAB2RAM_D2_O2));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(FAB2RAM_D2_O3));
 sky130_fd_sc_hd__clkbuf_4 output217 (.A(net217),
    .X(FAB2RAM_D3_O0));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(FAB2RAM_D3_O1));
 sky130_fd_sc_hd__clkbuf_4 output219 (.A(net219),
    .X(FAB2RAM_D3_O2));
 sky130_fd_sc_hd__clkbuf_4 output220 (.A(net220),
    .X(FAB2RAM_D3_O3));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(FrameData_O[0]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(FrameData_O[10]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(FrameData_O[11]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(FrameData_O[12]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(FrameData_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output226 (.A(net226),
    .X(FrameData_O[14]));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(FrameData_O[15]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(FrameData_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output229 (.A(net229),
    .X(FrameData_O[17]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(FrameData_O[18]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(FrameData_O[19]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(FrameData_O[1]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(FrameData_O[20]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(FrameData_O[21]));
 sky130_fd_sc_hd__clkbuf_4 output235 (.A(net235),
    .X(FrameData_O[22]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(FrameData_O[23]));
 sky130_fd_sc_hd__clkbuf_4 output237 (.A(net237),
    .X(FrameData_O[24]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(FrameData_O[25]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(FrameData_O[26]));
 sky130_fd_sc_hd__clkbuf_4 output240 (.A(net240),
    .X(FrameData_O[27]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(FrameData_O[28]));
 sky130_fd_sc_hd__clkbuf_4 output242 (.A(net242),
    .X(FrameData_O[29]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(FrameData_O[2]));
 sky130_fd_sc_hd__clkbuf_4 output244 (.A(net244),
    .X(FrameData_O[30]));
 sky130_fd_sc_hd__clkbuf_4 output245 (.A(net245),
    .X(FrameData_O[31]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(FrameData_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output247 (.A(net247),
    .X(FrameData_O[4]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(FrameData_O[5]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(FrameData_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output250 (.A(net250),
    .X(FrameData_O[7]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(FrameData_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output252 (.A(net252),
    .X(FrameData_O[9]));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(FrameStrobe_O[0]));
 sky130_fd_sc_hd__clkbuf_4 output254 (.A(net254),
    .X(FrameStrobe_O[10]));
 sky130_fd_sc_hd__clkbuf_4 output255 (.A(net255),
    .X(FrameStrobe_O[11]));
 sky130_fd_sc_hd__clkbuf_4 output256 (.A(net256),
    .X(FrameStrobe_O[12]));
 sky130_fd_sc_hd__clkbuf_4 output257 (.A(net257),
    .X(FrameStrobe_O[13]));
 sky130_fd_sc_hd__clkbuf_4 output258 (.A(net258),
    .X(FrameStrobe_O[14]));
 sky130_fd_sc_hd__clkbuf_4 output259 (.A(net259),
    .X(FrameStrobe_O[15]));
 sky130_fd_sc_hd__clkbuf_4 output260 (.A(net260),
    .X(FrameStrobe_O[16]));
 sky130_fd_sc_hd__clkbuf_4 output261 (.A(net261),
    .X(FrameStrobe_O[17]));
 sky130_fd_sc_hd__clkbuf_4 output262 (.A(net262),
    .X(FrameStrobe_O[18]));
 sky130_fd_sc_hd__clkbuf_4 output263 (.A(net263),
    .X(FrameStrobe_O[19]));
 sky130_fd_sc_hd__clkbuf_4 output264 (.A(net264),
    .X(FrameStrobe_O[1]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net265),
    .X(FrameStrobe_O[2]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net266),
    .X(FrameStrobe_O[3]));
 sky130_fd_sc_hd__clkbuf_4 output267 (.A(net267),
    .X(FrameStrobe_O[4]));
 sky130_fd_sc_hd__clkbuf_4 output268 (.A(net268),
    .X(FrameStrobe_O[5]));
 sky130_fd_sc_hd__clkbuf_4 output269 (.A(net269),
    .X(FrameStrobe_O[6]));
 sky130_fd_sc_hd__clkbuf_4 output270 (.A(net270),
    .X(FrameStrobe_O[7]));
 sky130_fd_sc_hd__clkbuf_4 output271 (.A(net271),
    .X(FrameStrobe_O[8]));
 sky130_fd_sc_hd__clkbuf_4 output272 (.A(net272),
    .X(FrameStrobe_O[9]));
 sky130_fd_sc_hd__clkbuf_4 output273 (.A(net273),
    .X(N1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output274 (.A(net274),
    .X(N1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output275 (.A(net275),
    .X(N1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output276 (.A(net276),
    .X(N1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output277 (.A(net277),
    .X(N2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output278 (.A(net278),
    .X(N2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output279 (.A(net279),
    .X(N2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output280 (.A(net280),
    .X(N2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output281 (.A(net281),
    .X(N2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output282 (.A(net282),
    .X(N2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output283 (.A(net283),
    .X(N2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output284 (.A(net284),
    .X(N2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output285 (.A(net285),
    .X(N2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output286 (.A(net286),
    .X(N2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output287 (.A(net287),
    .X(N2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output288 (.A(net288),
    .X(N2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output289 (.A(net289),
    .X(N2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output290 (.A(net290),
    .X(N2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(N2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(N2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output293 (.A(net293),
    .X(N4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output294 (.A(net294),
    .X(N4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output295 (.A(net295),
    .X(N4BEG[11]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net296),
    .X(N4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output297 (.A(net297),
    .X(N4BEG[13]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net298),
    .X(N4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output299 (.A(net299),
    .X(N4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output300 (.A(net300),
    .X(N4BEG[1]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net301),
    .X(N4BEG[2]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(N4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output303 (.A(net303),
    .X(N4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output304 (.A(net304),
    .X(N4BEG[5]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(N4BEG[6]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(N4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output307 (.A(net307),
    .X(N4BEG[8]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(N4BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output309 (.A(net309),
    .X(S1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output310 (.A(net310),
    .X(S1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output311 (.A(net311),
    .X(S1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output312 (.A(net312),
    .X(S1BEG[3]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(S2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output314 (.A(net314),
    .X(S2BEG[1]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net315),
    .X(S2BEG[2]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net316),
    .X(S2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output317 (.A(net317),
    .X(S2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output318 (.A(net318),
    .X(S2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output319 (.A(net319),
    .X(S2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output320 (.A(net320),
    .X(S2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output321 (.A(net321),
    .X(S2BEGb[0]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(S2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output323 (.A(net323),
    .X(S2BEGb[2]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(S2BEGb[3]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(S2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output326 (.A(net326),
    .X(S2BEGb[5]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(S2BEGb[6]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(S2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output329 (.A(net329),
    .X(S4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output330 (.A(net330),
    .X(S4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output331 (.A(net331),
    .X(S4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output332 (.A(net332),
    .X(S4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output333 (.A(net333),
    .X(S4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output334 (.A(net334),
    .X(S4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output335 (.A(net335),
    .X(S4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output336 (.A(net336),
    .X(S4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output337 (.A(net337),
    .X(S4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output338 (.A(net338),
    .X(S4BEG[3]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(S4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output340 (.A(net340),
    .X(S4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output341 (.A(net341),
    .X(S4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output342 (.A(net342),
    .X(S4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output343 (.A(net343),
    .X(S4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output344 (.A(net344),
    .X(S4BEG[9]));
 sky130_fd_sc_hd__buf_1 output345 (.A(net345),
    .X(UserCLKo));
 sky130_fd_sc_hd__clkbuf_4 output346 (.A(net346),
    .X(W1BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output347 (.A(net347),
    .X(W1BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output348 (.A(net348),
    .X(W1BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output349 (.A(net349),
    .X(W1BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output350 (.A(net350),
    .X(W2BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output351 (.A(net351),
    .X(W2BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output352 (.A(net352),
    .X(W2BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output353 (.A(net353),
    .X(W2BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output354 (.A(net354),
    .X(W2BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output355 (.A(net355),
    .X(W2BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output356 (.A(net356),
    .X(W2BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output357 (.A(net357),
    .X(W2BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output358 (.A(net358),
    .X(W2BEGb[0]));
 sky130_fd_sc_hd__clkbuf_4 output359 (.A(net359),
    .X(W2BEGb[1]));
 sky130_fd_sc_hd__clkbuf_4 output360 (.A(net360),
    .X(W2BEGb[2]));
 sky130_fd_sc_hd__clkbuf_4 output361 (.A(net361),
    .X(W2BEGb[3]));
 sky130_fd_sc_hd__clkbuf_4 output362 (.A(net362),
    .X(W2BEGb[4]));
 sky130_fd_sc_hd__clkbuf_4 output363 (.A(net363),
    .X(W2BEGb[5]));
 sky130_fd_sc_hd__clkbuf_4 output364 (.A(net364),
    .X(W2BEGb[6]));
 sky130_fd_sc_hd__clkbuf_4 output365 (.A(net365),
    .X(W2BEGb[7]));
 sky130_fd_sc_hd__clkbuf_4 output366 (.A(net366),
    .X(W6BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output367 (.A(net367),
    .X(W6BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output368 (.A(net368),
    .X(W6BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output369 (.A(net369),
    .X(W6BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output370 (.A(net370),
    .X(W6BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output371 (.A(net371),
    .X(W6BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output372 (.A(net372),
    .X(W6BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output373 (.A(net373),
    .X(W6BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output374 (.A(net374),
    .X(W6BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output375 (.A(net375),
    .X(W6BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output376 (.A(net376),
    .X(W6BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output377 (.A(net377),
    .X(W6BEG[9]));
 sky130_fd_sc_hd__clkbuf_4 output378 (.A(net378),
    .X(WW4BEG[0]));
 sky130_fd_sc_hd__clkbuf_4 output379 (.A(net379),
    .X(WW4BEG[10]));
 sky130_fd_sc_hd__clkbuf_4 output380 (.A(net380),
    .X(WW4BEG[11]));
 sky130_fd_sc_hd__clkbuf_4 output381 (.A(net381),
    .X(WW4BEG[12]));
 sky130_fd_sc_hd__clkbuf_4 output382 (.A(net382),
    .X(WW4BEG[13]));
 sky130_fd_sc_hd__clkbuf_4 output383 (.A(net383),
    .X(WW4BEG[14]));
 sky130_fd_sc_hd__clkbuf_4 output384 (.A(net384),
    .X(WW4BEG[15]));
 sky130_fd_sc_hd__clkbuf_4 output385 (.A(net385),
    .X(WW4BEG[1]));
 sky130_fd_sc_hd__clkbuf_4 output386 (.A(net386),
    .X(WW4BEG[2]));
 sky130_fd_sc_hd__clkbuf_4 output387 (.A(net387),
    .X(WW4BEG[3]));
 sky130_fd_sc_hd__clkbuf_4 output388 (.A(net388),
    .X(WW4BEG[4]));
 sky130_fd_sc_hd__clkbuf_4 output389 (.A(net389),
    .X(WW4BEG[5]));
 sky130_fd_sc_hd__clkbuf_4 output390 (.A(net390),
    .X(WW4BEG[6]));
 sky130_fd_sc_hd__clkbuf_4 output391 (.A(net391),
    .X(WW4BEG[7]));
 sky130_fd_sc_hd__clkbuf_4 output392 (.A(net392),
    .X(WW4BEG[8]));
 sky130_fd_sc_hd__clkbuf_4 output393 (.A(net393),
    .X(WW4BEG[9]));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_0/_0_  (.A(net81),
    .X(\FrameStrobe_O_i[0] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_1/_0_  (.A(net92),
    .X(\FrameStrobe_O_i[1] ));
 sky130_fd_sc_hd__clkbuf_2 \strobe_inbuf_10/_0_  (.A(net82),
    .X(\FrameStrobe_O_i[10] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_11/_0_  (.A(net83),
    .X(\FrameStrobe_O_i[11] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_12/_0_  (.A(net84),
    .X(\FrameStrobe_O_i[12] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_13/_0_  (.A(net85),
    .X(\FrameStrobe_O_i[13] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_14/_0_  (.A(net86),
    .X(\FrameStrobe_O_i[14] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_15/_0_  (.A(net87),
    .X(\FrameStrobe_O_i[15] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_16/_0_  (.A(net88),
    .X(\FrameStrobe_O_i[16] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_17/_0_  (.A(net89),
    .X(\FrameStrobe_O_i[17] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_18/_0_  (.A(net90),
    .X(\FrameStrobe_O_i[18] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_19/_0_  (.A(net91),
    .X(\FrameStrobe_O_i[19] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_2/_0_  (.A(net93),
    .X(\FrameStrobe_O_i[2] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_3/_0_  (.A(net94),
    .X(\FrameStrobe_O_i[3] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_4/_0_  (.A(net95),
    .X(\FrameStrobe_O_i[4] ));
 sky130_fd_sc_hd__buf_1 \strobe_inbuf_5/_0_  (.A(net96),
    .X(\FrameStrobe_O_i[5] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_6/_0_  (.A(net97),
    .X(\FrameStrobe_O_i[6] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_7/_0_  (.A(net98),
    .X(\FrameStrobe_O_i[7] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_8/_0_  (.A(net99),
    .X(\FrameStrobe_O_i[8] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_inbuf_9/_0_  (.A(net100),
    .X(\FrameStrobe_O_i[9] ));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_0/_0_  (.A(\FrameStrobe_O_i[0] ),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_1/_0_  (.A(\FrameStrobe_O_i[1] ),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_10/_0_  (.A(\FrameStrobe_O_i[10] ),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_11/_0_  (.A(\FrameStrobe_O_i[11] ),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_12/_0_  (.A(\FrameStrobe_O_i[12] ),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_13/_0_  (.A(\FrameStrobe_O_i[13] ),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_14/_0_  (.A(\FrameStrobe_O_i[14] ),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_15/_0_  (.A(\FrameStrobe_O_i[15] ),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_16/_0_  (.A(\FrameStrobe_O_i[16] ),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_17/_0_  (.A(\FrameStrobe_O_i[17] ),
    .X(net261));
 sky130_fd_sc_hd__buf_1 \strobe_outbuf_18/_0_  (.A(\FrameStrobe_O_i[18] ),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_19/_0_  (.A(\FrameStrobe_O_i[19] ),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_2/_0_  (.A(\FrameStrobe_O_i[2] ),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_3/_0_  (.A(\FrameStrobe_O_i[3] ),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_4/_0_  (.A(\FrameStrobe_O_i[4] ),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_5/_0_  (.A(\FrameStrobe_O_i[5] ),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_6/_0_  (.A(\FrameStrobe_O_i[6] ),
    .X(net269));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_7/_0_  (.A(\FrameStrobe_O_i[7] ),
    .X(net270));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_8/_0_  (.A(\FrameStrobe_O_i[8] ),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_1 \strobe_outbuf_9/_0_  (.A(\FrameStrobe_O_i[9] ),
    .X(net272));
endmodule

