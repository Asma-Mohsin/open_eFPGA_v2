* NGSPICE file created from W_IO.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxbp_1 abstract view
.subckt sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt W_IO A_I_top A_O_top A_T_top A_config_C_bit0 A_config_C_bit1 A_config_C_bit2
+ A_config_C_bit3 B_I_top B_O_top B_T_top B_config_C_bit0 B_config_C_bit1 B_config_C_bit2
+ B_config_C_bit3 E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3]
+ E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7] E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4]
+ E2BEGb[5] E2BEGb[6] E2BEGb[7] E6BEG[0] E6BEG[10] E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3]
+ E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8] E6BEG[9] EE4BEG[0] EE4BEG[10] EE4BEG[11]
+ EE4BEG[12] EE4BEG[13] EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4]
+ EE4BEG[5] EE4BEG[6] EE4BEG[7] EE4BEG[8] EE4BEG[9] FrameData[0] FrameData[10] FrameData[11]
+ FrameData[12] FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17]
+ FrameData[18] FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22]
+ FrameData[23] FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28]
+ FrameData[29] FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4]
+ FrameData[5] FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0]
+ FrameData_O[10] FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14]
+ FrameData_O[15] FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19]
+ FrameData_O[1] FrameData_O[20] FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24]
+ FrameData_O[25] FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29]
+ FrameData_O[2] FrameData_O[30] FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5]
+ FrameData_O[6] FrameData_O[7] FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10]
+ FrameStrobe[11] FrameStrobe[12] FrameStrobe[13] FrameStrobe[14] FrameStrobe[15]
+ FrameStrobe[16] FrameStrobe[17] FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2]
+ FrameStrobe[3] FrameStrobe[4] FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8]
+ FrameStrobe[9] FrameStrobe_O[0] FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12]
+ FrameStrobe_O[13] FrameStrobe_O[14] FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17]
+ FrameStrobe_O[18] FrameStrobe_O[19] FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3]
+ FrameStrobe_O[4] FrameStrobe_O[5] FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8]
+ FrameStrobe_O[9] UserCLK UserCLKo VGND VPWR W1END[0] W1END[1] W1END[2] W1END[3]
+ W2END[0] W2END[1] W2END[2] W2END[3] W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0]
+ W2MID[1] W2MID[2] W2MID[3] W2MID[4] W2MID[5] W2MID[6] W2MID[7] W6END[0] W6END[10]
+ W6END[11] W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8]
+ W6END[9] WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15]
+ WW4END[1] WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8]
+ WW4END[9]
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst_break_comb_loop_inst0__0_
+ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst0/X VGND VGND VPWR
+ VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__2_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1_217 VGND VGND
+ VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1_217/HI
+ net217 sky130_fd_sc_hd__conb_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_B_config_Config_access__0_ ConfigBits\[4\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_20__0_ net15 VGND VGND VPWR VPWR FrameData_O_i\[20\] sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG6 net67 net69 net71 net73 ConfigBits\[56\]
+ ConfigBits\[57\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__mux4_1
XFILLER_0_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_inbuf_11__0_ net5 VGND VGND VPWR VPWR FrameData_O_i\[11\] sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_ConfigMem_Inst_frame1_bit0 net3 net46 VGND VGND VPWR VPWR ConfigBits\[50\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__2_ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__2_/A
+ VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__2_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_14__0_ FrameStrobe_O_i\[14\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_9__0_ FrameData_O_i\[9\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput210 net210 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__buf_2
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_11__0_ net37 VGND VGND VPWR VPWR FrameStrobe_O_i\[11\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_9__0_ FrameStrobe_O_i\[9\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG7 net68 net70 net72 net74 ConfigBits\[58\]
+ ConfigBits\[59\] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__mux4_1
XFILLER_0_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_A_IO_1_bidirectional_frame_config_pass__3_ net1 VGND VGND VPWR VPWR A_O sky130_fd_sc_hd__clkbuf_2
XInst_W_IO_ConfigMem_Inst_frame1_bit1 net14 net46 VGND VGND VPWR VPWR ConfigBits\[51\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_inbuf_3__0_ net28 VGND VGND VPWR VPWR FrameData_O_i\[3\] sky130_fd_sc_hd__clkbuf_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1_219 VGND VGND
+ VPWR VPWR net219 Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1_219/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput200 net200 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__buf_2
Xoutput211 net211 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__buf_2
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_30__0_ FrameData_O_i\[30\] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_21__0_ FrameData_O_i\[21\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_12__0_ FrameData_O_i\[12\] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst0 net74 net59 net60
+ net61 ConfigBits\[104\] ConfigBits\[105\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG8 net81 net83 net85 net76 ConfigBits\[60\]
+ ConfigBits\[61\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__mux4_1
XInst_A_IO_1_bidirectional_frame_config_pass__2_ A_I VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_ConfigMem_Inst_frame1_bit2 net25 net46 VGND VGND VPWR VPWR ConfigBits\[52\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput100 WW4END[7] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_37_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput201 net201 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput212 net212 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__buf_2
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_23__0_ net18 VGND VGND VPWR VPWR FrameData_O_i\[23\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xstrobe_inbuf_2__0_ net47 VGND VGND VPWR VPWR FrameStrobe_O_i\[2\] sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_14__0_ net8 VGND VGND VPWR VPWR FrameData_O_i\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1 net62 net63 net216
+ net218 ConfigBits\[104\] ConfigBits\[105\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG9 net78 net80 net82 net84 ConfigBits\[62\]
+ ConfigBits\[63\] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__mux4_1
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame1_bit3 net28 net46 VGND VGND VPWR VPWR ConfigBits\[53\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_A_IO_1_bidirectional_frame_config_pass__1_ UserCLK net1 VGND VGND VPWR VPWR
+ A_Q sky130_fd_sc_hd__dfxtp_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_17__0_ FrameStrobe_O_i\[17\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput101 WW4END[8] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_14__0_ net40 VGND VGND VPWR VPWR FrameStrobe_O_i\[14\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput202 net202 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__buf_2
Xoutput213 net213 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__buf_2
XFILLER_0_71_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_W_IO_ConfigMem_Inst_frame3_bit30 net26 net48 VGND VGND VPWR VPWR ConfigBits\[16\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_6__0_ net31 VGND VGND VPWR VPWR FrameData_O_i\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_A_IO_1_bidirectional_frame_config_pass__0_ A_T VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__inv_2
XInst_W_IO_ConfigMem_Inst_frame1_bit4 net29 net46 VGND VGND VPWR VPWR ConfigBits\[54\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput102 WW4END[9] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput214 net214 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__buf_2
Xoutput203 net203 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_24__0_ FrameData_O_i\[24\] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_15__0_ FrameData_O_i\[15\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_ConfigMem_Inst_frame3_bit20 net15 net48 VGND VGND VPWR VPWR ConfigBits\[6\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame3_bit31 net27 net48 VGND VGND VPWR VPWR ConfigBits\[17\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame1_bit5 net30 net46 VGND VGND VPWR VPWR ConfigBits\[55\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit30 net26 net47 VGND VGND VPWR VPWR ConfigBits\[48\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1_break_comb_loop_inst1__0_ A_Q VGND
+ VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__3_/A sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_2__0_ FrameData_O_i\[2\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
Xoutput215 net215 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_1
Xoutput204 net204 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_inbuf_26__0_ net21 VGND VGND VPWR VPWR FrameData_O_i\[26\] sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_5__0_ net50 VGND VGND VPWR VPWR FrameStrobe_O_i\[5\] sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_17__0_ net11 VGND VGND VPWR VPWR FrameData_O_i\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame3_bit21 net16 net48 VGND VGND VPWR VPWR ConfigBits\[7\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2_break_comb_loop_inst0__0_ net56 VGND
+ VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__2_/A sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_ConfigMem_Inst_frame1_bit6 net31 net46 VGND VGND VPWR VPWR ConfigBits\[56\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit20 net15 net47 VGND VGND VPWR VPWR ConfigBits\[38\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit31 net27 net47 VGND VGND VPWR VPWR ConfigBits\[49\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_2__0_ FrameStrobe_O_i\[2\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__buf_1
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_17__0_ net43 VGND VGND VPWR VPWR FrameStrobe_O_i\[17\] sky130_fd_sc_hd__clkbuf_2
XInst_W_IO_ConfigMem_Inst_frame1_bit30 net26 net46 VGND VGND VPWR VPWR ConfigBits\[80\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput205 net205 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_9__0_ net34 VGND VGND VPWR VPWR FrameData_O_i\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_ConfigMem_Inst_frame3_bit22 net17 net48 VGND VGND VPWR VPWR ConfigBits\[8\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_ConfigMem_Inst_frame1_bit7 net32 net46 VGND VGND VPWR VPWR ConfigBits\[57\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit21 net16 net47 VGND VGND VPWR VPWR ConfigBits\[39\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit10 net4 net47 VGND VGND VPWR VPWR ConfigBits\[28\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_ConfigMem_Inst_frame1_bit31 net27 net46 VGND VGND VPWR VPWR ConfigBits\[81\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame1_bit20 net15 net46 VGND VGND VPWR VPWR ConfigBits\[70\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_49_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_A_config_Config_access__3_ ConfigBits\[3\] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_27__0_ FrameData_O_i\[27\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput206 net206 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__buf_2
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_18__0_ FrameData_O_i\[18\] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_ConfigMem_Inst_frame0_bit30 net26 net35 VGND VGND VPWR VPWR ConfigBits\[112\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit30/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_ConfigMem_Inst_frame3_bit23 net18 net48 VGND VGND VPWR VPWR ConfigBits\[9\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_W_IO_ConfigMem_Inst_frame1_bit8 net33 net46 VGND VGND VPWR VPWR ConfigBits\[58\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit22 net17 net47 VGND VGND VPWR VPWR ConfigBits\[40\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit11 net5 net47 VGND VGND VPWR VPWR ConfigBits\[29\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_10__0_ FrameStrobe_O_i\[10\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_outbuf_5__0_ FrameData_O_i\[5\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_ConfigMem_Inst_frame1_bit10 net4 net46 VGND VGND VPWR VPWR ConfigBits\[60\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame1_bit21 net16 net46 VGND VGND VPWR VPWR ConfigBits\[71\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_inbuf_29__0_ net24 VGND VGND VPWR VPWR FrameData_O_i\[29\] sky130_fd_sc_hd__clkbuf_1
XInst_A_config_Config_access__2_ ConfigBits\[2\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_8__0_ net53 VGND VGND VPWR VPWR FrameStrobe_O_i\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput207 net207 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_ConfigMem_Inst_frame0_bit20 net15 net35 VGND VGND VPWR VPWR ConfigBits\[102\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit20/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit31 net27 net35 VGND VGND VPWR VPWR ConfigBits\[113\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit31/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame3_bit24 net19 net48 VGND VGND VPWR VPWR ConfigBits\[10\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame1_bit9 net34 net46 VGND VGND VPWR VPWR ConfigBits\[59\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_5__0_ FrameStrobe_O_i\[5\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__4_ ConfigBits\[10\] Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__2_/Y
+ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__3_/Y VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__o21ai_1
XInst_W_IO_ConfigMem_Inst_frame2_bit12 net6 net47 VGND VGND VPWR VPWR ConfigBits\[30\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit23 net18 net47 VGND VGND VPWR VPWR ConfigBits\[41\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1_216 VGND VGND
+ VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1_216/HI
+ net216 sky130_fd_sc_hd__conb_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG10 net75 net79 net81 A_O ConfigBits\[64\]
+ ConfigBits\[65\] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__mux4_1
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_ConfigMem_Inst_frame1_bit22 net17 net46 VGND VGND VPWR VPWR ConfigBits\[72\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame1_bit11 net5 net46 VGND VGND VPWR VPWR ConfigBits\[61\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_A_config_Config_access__1_ ConfigBits\[1\] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput208 net208 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__buf_2
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_ConfigMem_Inst_frame0_bit21 net16 net35 VGND VGND VPWR VPWR ConfigBits\[103\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit21/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit10 net4 net35 VGND VGND VPWR VPWR ConfigBits\[92\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit10/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame3_bit14 net8 net48 VGND VGND VPWR VPWR ConfigBits\[0\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame3_bit25 net20 net48 VGND VGND VPWR VPWR ConfigBits\[11\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit24 net19 net47 VGND VGND VPWR VPWR ConfigBits\[42\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__3_ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__3_/A
+ ConfigBits\[10\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__3_/Y
+ sky130_fd_sc_hd__nand2_1
XInst_W_IO_ConfigMem_Inst_frame2_bit13 net7 net47 VGND VGND VPWR VPWR ConfigBits\[31\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG11 net83 net85 net76 B_O ConfigBits\[66\]
+ ConfigBits\[67\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__mux4_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput90 WW4END[12] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_1
XInst_W_IO_ConfigMem_Inst_frame1_bit23 net18 net46 VGND VGND VPWR VPWR ConfigBits\[73\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_ConfigMem_Inst_frame1_bit12 net6 net46 VGND VGND VPWR VPWR ConfigBits\[62\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_A_config_Config_access__0_ ConfigBits\[0\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput209 net209 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_ConfigMem_Inst_frame0_bit11 net5 net35 VGND VGND VPWR VPWR ConfigBits\[93\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit11/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit22 net17 net35 VGND VGND VPWR VPWR ConfigBits\[104\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit22/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_ConfigMem_Inst_frame3_bit15 net9 net48 VGND VGND VPWR VPWR ConfigBits\[1\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame3_bit26 net21 net48 VGND VGND VPWR VPWR ConfigBits\[12\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__4_ ConfigBits\[106\]
+ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__2_/Y Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__3_/Y
+ VGND VGND VPWR VPWR A_T sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_inbuf_10__0_ net4 VGND VGND VPWR VPWR FrameData_O_i\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame0_bit0 net3 net35 VGND VGND VPWR VPWR ConfigBits\[82\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__2_ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__2_/A
+ VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__2_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_57_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit25 net20 net47 VGND VGND VPWR VPWR ConfigBits\[43\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit14 net8 net47 VGND VGND VPWR VPWR ConfigBits\[32\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1_218 VGND VGND
+ VPWR VPWR net218 Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1_218/LO
+ sky130_fd_sc_hd__conb_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG12 net78 net80 net82 A_Q ConfigBits\[68\]
+ ConfigBits\[69\] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__mux4_1
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_13__0_ FrameStrobe_O_i\[13\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_8__0_ FrameData_O_i\[8\] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
Xinput91 WW4END[13] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_1
Xinput80 W6END[3] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_2
XInst_W_IO_ConfigMem_Inst_frame1_bit24 net19 net46 VGND VGND VPWR VPWR ConfigBits\[74\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame1_bit13 net7 net46 VGND VGND VPWR VPWR ConfigBits\[63\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_ConfigMem_Inst_frame0_bit23 net18 net35 VGND VGND VPWR VPWR ConfigBits\[105\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit23/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit12 net6 net35 VGND VGND VPWR VPWR ConfigBits\[94\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit12/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_10__0_ net36 VGND VGND VPWR VPWR FrameStrobe_O_i\[10\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_ConfigMem_Inst_frame3_bit16 net10 net48 VGND VGND VPWR VPWR ConfigBits\[2\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame3_bit27 net22 net48 VGND VGND VPWR VPWR ConfigBits\[13\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__3_ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__3_/A
+ ConfigBits\[106\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_8__0_ FrameStrobe_O_i\[8\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
Xinput1 A_O_top VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XFILLER_0_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_2__0_ net25 VGND VGND VPWR VPWR FrameData_O_i\[2\] sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_ConfigMem_Inst_frame0_bit1 net14 net35 VGND VGND VPWR VPWR ConfigBits\[83\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_W_IO_ConfigMem_Inst_frame2_bit15 net9 net47 VGND VGND VPWR VPWR ConfigBits\[33\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit26 net21 net47 VGND VGND VPWR VPWR ConfigBits\[44\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG13 net84 net86 net77 B_Q ConfigBits\[70\]
+ ConfigBits\[71\] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__mux4_1
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput190 net190 VGND VGND VPWR VPWR FrameData_O[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput70 W2MID[3] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
Xinput92 WW4END[14] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_1
Xinput81 W6END[4] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlymetal6s2s_1
XInst_W_IO_ConfigMem_Inst_frame1_bit25 net20 net46 VGND VGND VPWR VPWR ConfigBits\[75\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame1_bit14 net8 net46 VGND VGND VPWR VPWR ConfigBits\[64\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_ConfigMem_Inst_frame0_bit24 net19 net35 VGND VGND VPWR VPWR ConfigBits\[106\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit24/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit13 net7 net35 VGND VGND VPWR VPWR ConfigBits\[95\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit13/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame3_bit28 net23 net48 VGND VGND VPWR VPWR ConfigBits\[14\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame3_bit17 net11 net48 VGND VGND VPWR VPWR ConfigBits\[3\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_outbuf_20__0_ FrameData_O_i\[20\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_11__0_ FrameData_O_i\[11\] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__2_ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__2_/A
+ VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XFILLER_0_46_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput2 B_O_top VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_1
XFILLER_0_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_W_IO_ConfigMem_Inst_frame0_bit2 net25 net35 VGND VGND VPWR VPWR ConfigBits\[84\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit16 net10 net47 VGND VGND VPWR VPWR ConfigBits\[34\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit27 net22 net47 VGND VGND VPWR VPWR ConfigBits\[45\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG14 net67 net69 net71 net73 ConfigBits\[72\]
+ ConfigBits\[73\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__mux4_2
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput180 net180 VGND VGND VPWR VPWR FrameData_O[25] sky130_fd_sc_hd__buf_2
Xoutput191 net191 VGND VGND VPWR VPWR FrameData_O[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput60 W2END[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput71 W2MID[4] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput93 WW4END[15] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__buf_1
Xinput82 W6END[5] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_66_103 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame1_bit26 net21 net46 VGND VGND VPWR VPWR ConfigBits\[76\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame1_bit15 net9 net46 VGND VGND VPWR VPWR ConfigBits\[65\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame0_bit25 net20 net35 VGND VGND VPWR VPWR ConfigBits\[107\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit25/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit14 net8 net35 VGND VGND VPWR VPWR ConfigBits\[96\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit14/Q_N sky130_fd_sc_hd__dlxbp_1
Xdata_inbuf_31__0_ net27 VGND VGND VPWR VPWR FrameData_O_i\[31\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_inbuf_22__0_ net17 VGND VGND VPWR VPWR FrameData_O_i\[22\] sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_ConfigMem_Inst_frame3_bit18 net12 net48 VGND VGND VPWR VPWR ConfigBits\[4\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame3_bit29 net24 net48 VGND VGND VPWR VPWR ConfigBits\[15\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_1__0_ net46 VGND VGND VPWR VPWR FrameStrobe_O_i\[1\] sky130_fd_sc_hd__buf_1
Xdata_inbuf_13__0_ net7 VGND VGND VPWR VPWR FrameData_O_i\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput3 FrameData[0] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame0_bit3 net28 net35 VGND VGND VPWR VPWR ConfigBits\[85\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_16__0_ FrameStrobe_O_i\[16\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_ConfigMem_Inst_frame2_bit17 net11 net47 VGND VGND VPWR VPWR ConfigBits\[35\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame2_bit28 net23 net47 VGND VGND VPWR VPWR ConfigBits\[46\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG15 net68 net70 net72 net74 ConfigBits\[74\]
+ ConfigBits\[75\] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__mux4_2
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinst_clk_buf UserCLK VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_16
Xoutput181 net181 VGND VGND VPWR VPWR FrameData_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput192 net192 VGND VGND VPWR VPWR FrameData_O[7] sky130_fd_sc_hd__clkbuf_4
Xoutput170 net170 VGND VGND VPWR VPWR FrameData_O[16] sky130_fd_sc_hd__clkbuf_4
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput61 W2END[2] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_1
Xinput72 W2MID[5] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_2
Xinput50 FrameStrobe[5] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_2
Xinput94 WW4END[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput83 W6END[6] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_W_IO_ConfigMem_Inst_frame1_bit27 net22 net46 VGND VGND VPWR VPWR ConfigBits\[77\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame1_bit16 net10 net46 VGND VGND VPWR VPWR ConfigBits\[66\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_13__0_ net39 VGND VGND VPWR VPWR FrameStrobe_O_i\[13\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame0_bit26 net21 net35 VGND VGND VPWR VPWR ConfigBits\[108\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit26/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit15 net9 net35 VGND VGND VPWR VPWR ConfigBits\[97\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit15/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame3_bit19 net13 net48 VGND VGND VPWR VPWR ConfigBits\[5\]
+ Inst_W_IO_ConfigMem_Inst_frame3_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_5_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_5__0_ net30 VGND VGND VPWR VPWR FrameData_O_i\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput4 FrameData[10] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame0_bit4 net29 net35 VGND VGND VPWR VPWR ConfigBits\[86\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit18 net12 net47 VGND VGND VPWR VPWR ConfigBits\[36\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit29 net24 net47 VGND VGND VPWR VPWR ConfigBits\[47\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput182 net182 VGND VGND VPWR VPWR FrameData_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput160 net160 VGND VGND VPWR VPWR EE4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput193 net193 VGND VGND VPWR VPWR FrameData_O[8] sky130_fd_sc_hd__clkbuf_4
Xoutput171 net171 VGND VGND VPWR VPWR FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput62 W2END[3] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput95 WW4END[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 W2MID[6] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_2
Xinput51 FrameStrobe[6] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput40 FrameStrobe[14] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput84 W6END[7] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame1_bit17 net11 net46 VGND VGND VPWR VPWR ConfigBits\[67\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame1_bit28 net23 net46 VGND VGND VPWR VPWR ConfigBits\[78\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_ConfigMem_Inst_frame0_bit16 net10 net35 VGND VGND VPWR VPWR ConfigBits\[98\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit16/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit27 net22 net35 VGND VGND VPWR VPWR ConfigBits\[109\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit27/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_23__0_ FrameData_O_i\[23\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_14__0_ FrameData_O_i\[14\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst_break_comb_loop_inst1__0_
+ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst1/X VGND VGND VPWR
+ VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__3_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput5 FrameData[11] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame0_bit5 net30 net35 VGND VGND VPWR VPWR ConfigBits\[87\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame2_bit19 net13 net47 VGND VGND VPWR VPWR ConfigBits\[37\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0_break_comb_loop_inst1__0_ A_O VGND
+ VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__3_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput150 net150 VGND VGND VPWR VPWR EE4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput161 net161 VGND VGND VPWR VPWR EE4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput183 net183 VGND VGND VPWR VPWR FrameData_O[28] sky130_fd_sc_hd__clkbuf_4
Xoutput194 net194 VGND VGND VPWR VPWR FrameData_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput172 net172 VGND VGND VPWR VPWR FrameData_O[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput63 W2END[4] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_2
Xinput74 W2MID[7] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput52 FrameStrobe[7] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput41 FrameStrobe[15] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput96 WW4END[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_1
Xinput85 W6END[8] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
Xinput30 FrameData[5] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame1_bit18 net12 net46 VGND VGND VPWR VPWR ConfigBits\[68\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame1_bit29 net24 net46 VGND VGND VPWR VPWR ConfigBits\[79\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1_break_comb_loop_inst0__0_ net57 VGND
+ VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__2_/A sky130_fd_sc_hd__clkbuf_1
Xdata_outbuf_1__0_ FrameData_O_i\[1\] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_inbuf_25__0_ net20 VGND VGND VPWR VPWR FrameData_O_i\[25\] sky130_fd_sc_hd__clkbuf_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_ConfigMem_Inst_frame0_bit28 net23 net35 VGND VGND VPWR VPWR ConfigBits\[110\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit28/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame0_bit17 net11 net35 VGND VGND VPWR VPWR ConfigBits\[99\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit17/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_4__0_ net49 VGND VGND VPWR VPWR FrameStrobe_O_i\[4\] sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_16__0_ net10 VGND VGND VPWR VPWR FrameData_O_i\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_19__0_ FrameStrobe_O_i\[19\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
Xinput6 FrameData[12] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_ConfigMem_Inst_frame0_bit6 net31 net35 VGND VGND VPWR VPWR ConfigBits\[88\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput195 net195 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput184 net184 VGND VGND VPWR VPWR FrameData_O[29] sky130_fd_sc_hd__buf_2
Xoutput151 net151 VGND VGND VPWR VPWR EE4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput162 net162 VGND VGND VPWR VPWR EE4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput140 net140 VGND VGND VPWR VPWR E6BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput173 net173 VGND VGND VPWR VPWR FrameData_O[19] sky130_fd_sc_hd__buf_2
XFILLER_0_68_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_1__0_ FrameStrobe_O_i\[1\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput31 FrameData[6] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput20 FrameData[25] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput64 W2END[5] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_2
Xinput53 FrameStrobe[8] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
Xinput42 FrameStrobe[16] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xinput97 WW4END[4] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__buf_1
Xinput75 W6END[0] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__clkbuf_2
Xinput86 W6END[9] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame1_bit19 net13 net46 VGND VGND VPWR VPWR ConfigBits\[69\]
+ Inst_W_IO_ConfigMem_Inst_frame1_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_16__0_ net42 VGND VGND VPWR VPWR FrameStrobe_O_i\[16\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame0_bit18 net12 net35 VGND VGND VPWR VPWR ConfigBits\[100\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit18/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_ConfigMem_Inst_frame0_bit29 net24 net35 VGND VGND VPWR VPWR ConfigBits\[111\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit29/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG0 net57 net89 net77 A_O ConfigBits\[76\]
+ ConfigBits\[77\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__mux4_1
XFILLER_0_25_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_8__0_ net33 VGND VGND VPWR VPWR FrameData_O_i\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 FrameData[13] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_ConfigMem_Inst_frame0_bit7 net32 net35 VGND VGND VPWR VPWR ConfigBits\[89\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput196 net196 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__buf_2
Xoutput130 net130 VGND VGND VPWR VPWR E2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput141 net141 VGND VGND VPWR VPWR E6BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput163 net163 VGND VGND VPWR VPWR FrameData_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput152 net152 VGND VGND VPWR VPWR EE4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput185 net185 VGND VGND VPWR VPWR FrameData_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput174 net174 VGND VGND VPWR VPWR FrameData_O[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput54 FrameStrobe[9] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xinput43 FrameStrobe[17] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput32 FrameData[7] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_2
Xinput10 FrameData[16] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__buf_2
Xinput21 FrameData[26] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_2
Xinput65 W2END[6] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_2
Xinput87 WW4END[0] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput98 WW4END[5] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 W6END[10] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_1
XFILLER_0_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_26__0_ FrameData_O_i\[26\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xdata_outbuf_17__0_ FrameData_O_i\[17\] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame0_bit19 net13 net35 VGND VGND VPWR VPWR ConfigBits\[101\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit19/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG1 net58 net88 net76 B_O ConfigBits\[78\]
+ ConfigBits\[79\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__mux4_1
XFILLER_0_25_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput8 FrameData[14] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XInst_W_IO_ConfigMem_Inst_frame0_bit8 net33 net35 VGND VGND VPWR VPWR ConfigBits\[90\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput197 net197 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__buf_2
Xoutput186 net186 VGND VGND VPWR VPWR FrameData_O[30] sky130_fd_sc_hd__clkbuf_4
Xoutput175 net175 VGND VGND VPWR VPWR FrameData_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput120 net120 VGND VGND VPWR VPWR E2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput131 net131 VGND VGND VPWR VPWR E2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput142 net142 VGND VGND VPWR VPWR E6BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput153 net153 VGND VGND VPWR VPWR EE4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput164 net164 VGND VGND VPWR VPWR FrameData_O[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput55 W1END[0] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput44 FrameStrobe[18] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput66 W2END[7] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_1
Xinput88 WW4END[10] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput77 W6END[11] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
Xinput33 FrameData[8] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
Xinput11 FrameData[17] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
Xinput22 FrameData[27] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__buf_2
Xinput99 WW4END[6] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__buf_1
XFILLER_0_58_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xdata_outbuf_4__0_ FrameData_O_i\[4\] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xdata_inbuf_28__0_ net23 VGND VGND VPWR VPWR FrameData_O_i\[28\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_7__0_ net52 VGND VGND VPWR VPWR FrameStrobe_O_i\[7\] sky130_fd_sc_hd__clkbuf_2
Xdata_inbuf_19__0_ net13 VGND VGND VPWR VPWR FrameData_O_i\[19\] sky130_fd_sc_hd__clkbuf_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG2 net100 net93 net84 A_O ConfigBits\[80\]
+ ConfigBits\[81\] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__mux4_1
XFILLER_0_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput9 FrameData[15] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_0_52_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame0_bit9 net34 net35 VGND VGND VPWR VPWR ConfigBits\[91\]
+ Inst_W_IO_ConfigMem_Inst_frame0_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__4_ ConfigBits\[9\] Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__2_/Y
+ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__3_/Y VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_4__0_ FrameStrobe_O_i\[4\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
Xoutput110 net110 VGND VGND VPWR VPWR B_T_top sky130_fd_sc_hd__clkbuf_4
Xoutput121 net121 VGND VGND VPWR VPWR E2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput132 net132 VGND VGND VPWR VPWR E2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput143 net143 VGND VGND VPWR VPWR E6BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput198 net198 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__buf_2
Xoutput187 net187 VGND VGND VPWR VPWR FrameData_O[31] sky130_fd_sc_hd__clkbuf_4
Xoutput176 net176 VGND VGND VPWR VPWR FrameData_O[21] sky130_fd_sc_hd__clkbuf_4
Xoutput154 net154 VGND VGND VPWR VPWR EE4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput165 net165 VGND VGND VPWR VPWR FrameData_O[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xstrobe_inbuf_19__0_ net45 VGND VGND VPWR VPWR FrameStrobe_O_i\[19\] sky130_fd_sc_hd__clkbuf_2
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3_break_comb_loop_inst1__0_ B_Q VGND
+ VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__3_/A sky130_fd_sc_hd__clkbuf_1
Xinput23 FrameData[28] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_2
Xinput67 W2MID[0] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_2
Xinput56 W1END[1] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput45 FrameStrobe[19] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput89 WW4END[11] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_1
Xinput78 W6END[1] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_2
Xinput34 FrameData[9] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
Xinput12 FrameData[18] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XFILLER_0_58_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG3 net99 net92 net83 B_O ConfigBits\[82\]
+ ConfigBits\[83\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__mux4_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb0 net66 net100 net93 net84 ConfigBits\[28\]
+ ConfigBits\[29\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__mux4_1
XFILLER_0_36_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__3_ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__3_/A
+ ConfigBits\[9\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__3_/Y
+ sky130_fd_sc_hd__nand2_1
Xoutput177 net177 VGND VGND VPWR VPWR FrameData_O[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput111 net111 VGND VGND VPWR VPWR B_config_C_bit0 sky130_fd_sc_hd__clkbuf_4
Xoutput122 net122 VGND VGND VPWR VPWR E2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput133 net133 VGND VGND VPWR VPWR E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput155 net155 VGND VGND VPWR VPWR EE4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput144 net144 VGND VGND VPWR VPWR E6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput166 net166 VGND VGND VPWR VPWR FrameData_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput199 net199 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput188 net188 VGND VGND VPWR VPWR FrameData_O[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 FrameData[19] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
Xinput24 FrameData[29] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_4
Xinput68 W2MID[1] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_2
Xinput57 W1END[2] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput35 FrameStrobe[0] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_8
Xinput46 FrameStrobe[1] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_8
Xinput79 W6END[2] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_29__0_ FrameData_O_i\[29\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG4 net57 net96 net80 A_O ConfigBits\[84\]
+ ConfigBits\[85\] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst0 net67 net68 net69
+ net70 ConfigBits\[107\] ConfigBits\[108\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb1 net65 net99 net92 net83 ConfigBits\[30\]
+ ConfigBits\[31\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__mux4_1
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__2_ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__2_/A
+ VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG1__2_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput178 net178 VGND VGND VPWR VPWR FrameData_O[23] sky130_fd_sc_hd__buf_2
Xoutput112 net112 VGND VGND VPWR VPWR B_config_C_bit1 sky130_fd_sc_hd__clkbuf_4
Xoutput123 net123 VGND VGND VPWR VPWR E2BEG[4] sky130_fd_sc_hd__buf_2
Xoutput156 net156 VGND VGND VPWR VPWR EE4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput134 net134 VGND VGND VPWR VPWR E2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput145 net145 VGND VGND VPWR VPWR E6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput189 net189 VGND VGND VPWR VPWR FrameData_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput167 net167 VGND VGND VPWR VPWR FrameData_O[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_12__0_ FrameStrobe_O_i\[12\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
Xinput36 FrameStrobe[10] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput14 FrameData[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 FrameData[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_2
Xinput58 W1END[3] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_2
Xinput69 W2MID[2] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput47 FrameStrobe[2] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_8
Xdata_outbuf_7__0_ FrameData_O_i\[7\] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_B_IO_1_bidirectional_frame_config_pass__3_ net2 VGND VGND VPWR VPWR B_O sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG5 net58 net95 net79 B_O ConfigBits\[86\]
+ ConfigBits\[87\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__mux4_1
XFILLER_0_31_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst1 net71 net72 net73
+ net74 ConfigBits\[107\] ConfigBits\[108\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb2 net64 net98 net91 net82 ConfigBits\[32\]
+ ConfigBits\[33\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__mux4_1
XFILLER_0_36_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_7__0_ FrameStrobe_O_i\[7\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xdata_inbuf_1__0_ net14 VGND VGND VPWR VPWR FrameData_O_i\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput179 net179 VGND VGND VPWR VPWR FrameData_O[24] sky130_fd_sc_hd__clkbuf_4
Xoutput113 net113 VGND VGND VPWR VPWR B_config_C_bit2 sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 VGND VGND VPWR VPWR E2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput157 net157 VGND VGND VPWR VPWR EE4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput135 net135 VGND VGND VPWR VPWR E6BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput146 net146 VGND VGND VPWR VPWR E6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput168 net168 VGND VGND VPWR VPWR FrameData_O[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput26 FrameData[30] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_2
Xinput59 W2END[0] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput48 FrameStrobe[3] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_4
Xinput37 FrameStrobe[11] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput15 FrameData[20] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_B_IO_1_bidirectional_frame_config_pass__2_ B_I VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG6 net56 net102 net86 A_Q ConfigBits\[88\]
+ ConfigBits\[89\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__mux4_1
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb3 net63 net97 net90 net81 ConfigBits\[34\]
+ ConfigBits\[35\] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst2 net59 net60 net61
+ net62 ConfigBits\[107\] ConfigBits\[108\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
Xdata_outbuf_10__0_ FrameData_O_i\[10\] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput114 net114 VGND VGND VPWR VPWR B_config_C_bit3 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput103 net103 VGND VGND VPWR VPWR A_I_top sky130_fd_sc_hd__clkbuf_4
Xoutput125 net125 VGND VGND VPWR VPWR E2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput158 net158 VGND VGND VPWR VPWR EE4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput147 net147 VGND VGND VPWR VPWR EE4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput136 net136 VGND VGND VPWR VPWR E6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput169 net169 VGND VGND VPWR VPWR FrameData_O[15] sky130_fd_sc_hd__buf_2
XFILLER_0_53_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst_break_comb_loop_inst1__0_
+ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1/X VGND VGND VPWR
+ VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__3_/A sky130_fd_sc_hd__clkbuf_1
Xinput27 FrameData[31] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_2
Xinput49 FrameStrobe[4] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_2
Xinput38 FrameStrobe[12] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput16 FrameData[21] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_B_IO_1_bidirectional_frame_config_pass__1_ UserCLK net2 VGND VGND VPWR VPWR
+ B_Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG7 net55 net101 net85 B_Q ConfigBits\[90\]
+ ConfigBits\[91\] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__mux4_1
Xdata_inbuf_30__0_ net26 VGND VGND VPWR VPWR FrameData_O_i\[30\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_21__0_ net16 VGND VGND VPWR VPWR FrameData_O_i\[21\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit0 net3 net47 VGND VGND VPWR VPWR ConfigBits\[18\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit0/Q_N sky130_fd_sc_hd__dlxbp_1
Xstrobe_inbuf_0__0_ net35 VGND VGND VPWR VPWR FrameStrobe_O_i\[0\] sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb4 net62 net96 net89 net80 ConfigBits\[36\]
+ ConfigBits\[37\] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__mux4_1
Xdata_inbuf_12__0_ net6 VGND VGND VPWR VPWR FrameData_O_i\[12\] sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst3 net63 net64 net65
+ net66 ConfigBits\[107\] ConfigBits\[108\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_15__0_ FrameStrobe_O_i\[15\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput104 net104 VGND VGND VPWR VPWR A_T_top sky130_fd_sc_hd__clkbuf_4
Xoutput115 net115 VGND VGND VPWR VPWR E1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput126 net126 VGND VGND VPWR VPWR E2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput159 net159 VGND VGND VPWR VPWR EE4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput148 net148 VGND VGND VPWR VPWR EE4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput137 net137 VGND VGND VPWR VPWR E6BEG[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput39 FrameStrobe[13] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
Xinput28 FrameData[3] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput17 FrameData[22] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_2
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG10 net56 net94 net78 A_Q ConfigBits\[96\]
+ ConfigBits\[97\] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__mux4_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_B_IO_1_bidirectional_frame_config_pass__0_ B_T VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__inv_2
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xstrobe_inbuf_12__0_ net38 VGND VGND VPWR VPWR FrameStrobe_O_i\[12\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG8 net98 net91 net82 A_Q ConfigBits\[92\]
+ ConfigBits\[93\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__mux4_2
XFILLER_0_41_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit1 net14 net47 VGND VGND VPWR VPWR ConfigBits\[19\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit1/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst4 Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst0/X
+ Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst1/X Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst2/X
+ Inst_W_IO_switch_matrix_inst_cus_mux161_buf_B_I_cus_mux41_buf_inst3/X ConfigBits\[109\]
+ ConfigBits\[110\] VGND VGND VPWR VPWR B_I sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb5 net61 net95 net88 net79 ConfigBits\[38\]
+ ConfigBits\[39\] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__mux4_1
XFILLER_0_31_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG0 net74 net100 net93 net84 ConfigBits\[12\]
+ ConfigBits\[13\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__mux4_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_4__0_ net29 VGND VGND VPWR VPWR FrameData_O_i\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput105 net105 VGND VGND VPWR VPWR A_config_C_bit0 sky130_fd_sc_hd__clkbuf_4
Xoutput116 net116 VGND VGND VPWR VPWR E1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput127 net127 VGND VGND VPWR VPWR E2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput149 net149 VGND VGND VPWR VPWR EE4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput138 net138 VGND VGND VPWR VPWR E6BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 FrameData[23] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__buf_2
Xinput29 FrameData[4] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG11 net55 net87 net75 B_Q ConfigBits\[98\]
+ ConfigBits\[99\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__mux4_1
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_31__0_ FrameData_O_i\[31\] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E6BEG9 net97 net90 net81 B_Q ConfigBits\[94\]
+ ConfigBits\[95\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__mux4_1
Xdata_outbuf_22__0_ FrameData_O_i\[22\] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_13__0_ FrameData_O_i\[13\] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_W_IO_ConfigMem_Inst_frame2_bit2 net25 net47 VGND VGND VPWR VPWR ConfigBits\[20\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit2/Q_N sky130_fd_sc_hd__dlxbp_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst_break_comb_loop_inst0__0_
+ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux41_buf_inst0/X VGND VGND VPWR
+ VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_A_T_cus_mux21_inst__2_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb6 net60 net94 net102 net78 ConfigBits\[40\]
+ ConfigBits\[41\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG1 net73 net99 net92 net83 ConfigBits\[14\]
+ ConfigBits\[15\] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__mux4_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput106 net106 VGND VGND VPWR VPWR A_config_C_bit1 sky130_fd_sc_hd__clkbuf_4
Xoutput117 net117 VGND VGND VPWR VPWR E1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput128 net128 VGND VGND VPWR VPWR E2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput139 net139 VGND VGND VPWR VPWR E6BEG[2] sky130_fd_sc_hd__clkbuf_4
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0_break_comb_loop_inst0__0_ net58 VGND
+ VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__2_/A sky130_fd_sc_hd__clkbuf_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 FrameData[24] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_0__0_ FrameData_O_i\[0\] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_inbuf_24__0_ net19 VGND VGND VPWR VPWR FrameData_O_i\[24\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_3__0_ net48 VGND VGND VPWR VPWR FrameStrobe_O_i\[3\] sky130_fd_sc_hd__buf_1
Xdata_inbuf_15__0_ net9 VGND VGND VPWR VPWR FrameData_O_i\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_ConfigMem_Inst_frame2_bit3 net28 net47 VGND VGND VPWR VPWR ConfigBits\[21\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit3/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEGb7 net59 net87 net101 net75 ConfigBits\[42\]
+ ConfigBits\[43\] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG2 net72 net98 net91 net82 ConfigBits\[16\]
+ ConfigBits\[17\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__mux4_1
XFILLER_0_22_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xstrobe_outbuf_18__0_ FrameStrobe_O_i\[18\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput107 net107 VGND VGND VPWR VPWR A_config_C_bit2 sky130_fd_sc_hd__clkbuf_4
Xoutput118 net118 VGND VGND VPWR VPWR E1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput129 net129 VGND VGND VPWR VPWR E2BEGb[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_0__0_ FrameStrobe_O_i\[0\] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_15__0_ net41 VGND VGND VPWR VPWR FrameStrobe_O_i\[15\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_34_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_10 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_7__0_ net32 VGND VGND VPWR VPWR FrameData_O_i\[7\] sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst0 net67 net68 net69
+ net70 ConfigBits\[100\] ConfigBits\[101\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_ConfigMem_Inst_frame2_bit4 net29 net47 VGND VGND VPWR VPWR ConfigBits\[22\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit4/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG3 net71 net97 net90 net81 ConfigBits\[18\]
+ ConfigBits\[19\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__4_ ConfigBits\[113\]
+ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__2_/Y Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__3_/Y
+ VGND VGND VPWR VPWR B_T sky130_fd_sc_hd__o21ai_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput108 net108 VGND VGND VPWR VPWR A_config_C_bit3 sky130_fd_sc_hd__clkbuf_4
Xoutput119 net119 VGND VGND VPWR VPWR E2BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_25__0_ FrameData_O_i\[25\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_22 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_16__0_ FrameData_O_i\[16\] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst1 net71 net72 net73
+ net74 ConfigBits\[100\] ConfigBits\[101\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XInst_W_IO_ConfigMem_Inst_frame2_bit5 net30 net47 VGND VGND VPWR VPWR ConfigBits\[23\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit5/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG4 net70 net96 net89 net80 ConfigBits\[20\]
+ ConfigBits\[21\] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG0 net75 net79 net81 A_O ConfigBits\[44\]
+ ConfigBits\[45\] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__3_ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__3_/A
+ ConfigBits\[113\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__3_/Y
+ sky130_fd_sc_hd__nand2_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput109 net109 VGND VGND VPWR VPWR B_I_top sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_outbuf_3__0_ FrameData_O_i\[3\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xdata_inbuf_27__0_ net22 VGND VGND VPWR VPWR FrameData_O_i\[27\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_6__0_ net51 VGND VGND VPWR VPWR FrameStrobe_O_i\[6\] sky130_fd_sc_hd__clkbuf_1
Xdata_inbuf_18__0_ net12 VGND VGND VPWR VPWR FrameData_O_i\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst2 net59 net60 net61
+ net62 ConfigBits\[100\] ConfigBits\[101\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst2/X
+ sky130_fd_sc_hd__mux4_1
XInst_W_IO_ConfigMem_Inst_frame2_bit6 net31 net47 VGND VGND VPWR VPWR ConfigBits\[24\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit6/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2_break_comb_loop_inst1__0_ B_O VGND
+ VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG2__3_/A sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG5 net69 net95 net88 net79 ConfigBits\[22\]
+ ConfigBits\[23\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG1 net83 net85 net76 B_O ConfigBits\[46\]
+ ConfigBits\[47\] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst0 net73 net74 net59
+ net63 ConfigBits\[111\] ConfigBits\[112\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst0/X
+ sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__2_ Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__2_/A
+ VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux21_inst__2_/Y
+ sky130_fd_sc_hd__inv_2
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xstrobe_outbuf_3__0_ FrameStrobe_O_i\[3\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__4_ ConfigBits\[8\] Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__2_/Y
+ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__3_/Y VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3_break_comb_loop_inst0__0_ net55 VGND
+ VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__2_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_inbuf_18__0_ net44 VGND VGND VPWR VPWR FrameStrobe_O_i\[18\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst3 net63 net64 net65
+ net66 ConfigBits\[100\] ConfigBits\[101\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst3/X
+ sky130_fd_sc_hd__mux4_1
XInst_W_IO_ConfigMem_Inst_frame2_bit7 net32 net47 VGND VGND VPWR VPWR ConfigBits\[25\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit7/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG6 net68 net94 net102 net78 ConfigBits\[24\]
+ ConfigBits\[25\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG2 net78 net80 net82 A_Q ConfigBits\[48\]
+ ConfigBits\[49\] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1 net64 net65 net217
+ net219 ConfigBits\[111\] ConfigBits\[112\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux81_buf_B_T_cus_mux41_buf_inst1/X
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 FrameStrobe_O_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__3_ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__3_/A
+ ConfigBits\[8\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xdata_outbuf_28__0_ FrameData_O_i\[28\] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_19__0_ FrameData_O_i\[19\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_B_config_Config_access__3_ ConfigBits\[7\] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst4 Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst0/X
+ Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst1/X Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst2/X
+ Inst_W_IO_switch_matrix_inst_cus_mux161_buf_A_I_cus_mux41_buf_inst3/X ConfigBits\[102\]
+ ConfigBits\[103\] VGND VGND VPWR VPWR A_I sky130_fd_sc_hd__mux4_1
XInst_W_IO_ConfigMem_Inst_frame2_bit8 net33 net47 VGND VGND VPWR VPWR ConfigBits\[26\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit8/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_E2BEG7 net67 net87 net101 net75 ConfigBits\[26\]
+ ConfigBits\[27\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__mux4_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG3 net84 net86 net77 B_Q ConfigBits\[50\]
+ ConfigBits\[51\] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__mux4_1
XFILLER_0_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_2 FrameStrobe_O_i\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__2_ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__2_/A
+ VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG0__2_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_11__0_ FrameStrobe_O_i\[11\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xdata_outbuf_6__0_ FrameData_O_i\[6\] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_9__0_ net54 VGND VGND VPWR VPWR FrameStrobe_O_i\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_B_config_Config_access__2_ ConfigBits\[6\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
XInst_W_IO_ConfigMem_Inst_frame2_bit9 net34 net47 VGND VGND VPWR VPWR ConfigBits\[27\]
+ Inst_W_IO_ConfigMem_Inst_frame2_bit9/Q_N sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG4 net59 net61 net63 net65 ConfigBits\[52\]
+ ConfigBits\[53\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__mux4_2
XFILLER_0_1_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 FrameStrobe_O_i\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__4_ ConfigBits\[11\] Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__2_/Y
+ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__3_/Y VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__o21ai_1
Xstrobe_outbuf_6__0_ FrameStrobe_O_i\[6\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xdata_inbuf_0__0_ net3 VGND VGND VPWR VPWR FrameData_O_i\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_B_config_Config_access__1_ ConfigBits\[5\] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_W_IO_switch_matrix_inst_cus_mux41_buf_EE4BEG5 net60 net62 net64 net66 ConfigBits\[54\]
+ ConfigBits\[55\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__mux4_1
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__3_ Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__3_/A
+ ConfigBits\[11\] VGND VGND VPWR VPWR Inst_W_IO_switch_matrix_inst_cus_mux21_E1BEG3__3_/Y
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

