magic
tech sky130A
magscale 1 2
timestamp 1734836625
<< viali >>
rect 1685 43401 1719 43435
rect 3157 43401 3191 43435
rect 4169 43401 4203 43435
rect 4537 43401 4571 43435
rect 5917 43401 5951 43435
rect 7021 43401 7055 43435
rect 8309 43401 8343 43435
rect 9321 43401 9355 43435
rect 11345 43401 11379 43435
rect 11897 43401 11931 43435
rect 15853 43401 15887 43435
rect 16865 43401 16899 43435
rect 17417 43401 17451 43435
rect 18337 43401 18371 43435
rect 19441 43401 19475 43435
rect 19809 43401 19843 43435
rect 2881 43333 2915 43367
rect 7849 43333 7883 43367
rect 9965 43333 9999 43367
rect 10333 43333 10367 43367
rect 11805 43333 11839 43367
rect 13461 43333 13495 43367
rect 1501 43265 1535 43299
rect 1961 43265 1995 43299
rect 2513 43265 2547 43299
rect 3065 43265 3099 43299
rect 3985 43265 4019 43299
rect 4445 43265 4479 43299
rect 5089 43265 5123 43299
rect 5273 43265 5307 43299
rect 5825 43265 5859 43299
rect 6561 43265 6595 43299
rect 6745 43265 6779 43299
rect 7481 43265 7515 43299
rect 8033 43265 8067 43299
rect 8493 43265 8527 43299
rect 9137 43265 9171 43299
rect 9505 43265 9539 43299
rect 10793 43265 10827 43299
rect 11069 43265 11103 43299
rect 11161 43265 11195 43299
rect 12265 43265 12299 43299
rect 12633 43265 12667 43299
rect 13001 43265 13035 43299
rect 13921 43265 13955 43299
rect 14105 43265 14139 43299
rect 14657 43265 14691 43299
rect 14933 43265 14967 43299
rect 15209 43265 15243 43299
rect 15485 43265 15519 43299
rect 15669 43265 15703 43299
rect 16129 43265 16163 43299
rect 16773 43265 16807 43299
rect 17325 43265 17359 43299
rect 17785 43265 17819 43299
rect 18245 43265 18279 43299
rect 18705 43265 18739 43299
rect 19349 43265 19383 43299
rect 19993 43265 20027 43299
rect 20177 43265 20211 43299
rect 2237 43197 2271 43231
rect 16405 43197 16439 43231
rect 5549 43129 5583 43163
rect 6377 43129 6411 43163
rect 10517 43129 10551 43163
rect 14749 43129 14783 43163
rect 15025 43129 15059 43163
rect 18889 43129 18923 43163
rect 4905 43061 4939 43095
rect 8677 43061 8711 43095
rect 9689 43061 9723 43095
rect 10057 43061 10091 43095
rect 10609 43061 10643 43095
rect 10885 43061 10919 43095
rect 12449 43061 12483 43095
rect 12817 43061 12851 43095
rect 13185 43061 13219 43095
rect 13553 43061 13587 43095
rect 13737 43061 13771 43095
rect 14289 43061 14323 43095
rect 14473 43061 14507 43095
rect 15301 43061 15335 43095
rect 17969 43061 18003 43095
rect 20453 43061 20487 43095
rect 7297 42857 7331 42891
rect 10425 42857 10459 42891
rect 10885 42857 10919 42891
rect 11161 42857 11195 42891
rect 16497 42857 16531 42891
rect 19257 42857 19291 42891
rect 19901 42857 19935 42891
rect 1777 42789 1811 42823
rect 13369 42789 13403 42823
rect 3525 42721 3559 42755
rect 4169 42721 4203 42755
rect 4721 42721 4755 42755
rect 5273 42721 5307 42755
rect 5825 42721 5859 42755
rect 6377 42721 6411 42755
rect 8033 42721 8067 42755
rect 8585 42721 8619 42755
rect 17233 42721 17267 42755
rect 17785 42721 17819 42755
rect 18889 42721 18923 42755
rect 1685 42653 1719 42687
rect 1961 42653 1995 42687
rect 2513 42653 2547 42687
rect 3065 42653 3099 42687
rect 6653 42653 6687 42687
rect 7205 42653 7239 42687
rect 9045 42653 9079 42687
rect 9493 42653 9527 42687
rect 10057 42653 10091 42687
rect 10333 42653 10367 42687
rect 10609 42653 10643 42687
rect 10701 42653 10735 42687
rect 11069 42653 11103 42687
rect 11345 42653 11379 42687
rect 11621 42653 11655 42687
rect 12081 42653 12115 42687
rect 12541 42653 12575 42687
rect 12817 42653 12851 42687
rect 12909 42653 12943 42687
rect 13185 42653 13219 42687
rect 13737 42653 13771 42687
rect 14841 42653 14875 42687
rect 15117 42653 15151 42687
rect 15393 42653 15427 42687
rect 15669 42653 15703 42687
rect 15945 42653 15979 42687
rect 16221 42653 16255 42687
rect 19441 42653 19475 42687
rect 20177 42653 20211 42687
rect 2145 42585 2179 42619
rect 2697 42585 2731 42619
rect 3249 42585 3283 42619
rect 3893 42585 3927 42619
rect 4445 42585 4479 42619
rect 4997 42585 5031 42619
rect 5549 42585 5583 42619
rect 6101 42585 6135 42619
rect 7021 42585 7055 42619
rect 7757 42585 7791 42619
rect 8309 42585 8343 42619
rect 14381 42585 14415 42619
rect 16405 42585 16439 42619
rect 16957 42585 16991 42619
rect 17509 42585 17543 42619
rect 18061 42585 18095 42619
rect 18613 42585 18647 42619
rect 19625 42585 19659 42619
rect 1501 42517 1535 42551
rect 9137 42517 9171 42551
rect 9689 42517 9723 42551
rect 9873 42517 9907 42551
rect 10149 42517 10183 42551
rect 11529 42517 11563 42551
rect 11805 42517 11839 42551
rect 11897 42517 11931 42551
rect 12357 42517 12391 42551
rect 12633 42517 12667 42551
rect 13093 42517 13127 42551
rect 13553 42517 13587 42551
rect 14473 42517 14507 42551
rect 14657 42517 14691 42551
rect 14933 42517 14967 42551
rect 15209 42517 15243 42551
rect 15485 42517 15519 42551
rect 15761 42517 15795 42551
rect 16037 42517 16071 42551
rect 18337 42517 18371 42551
rect 20269 42517 20303 42551
rect 1961 42313 1995 42347
rect 2605 42313 2639 42347
rect 3157 42313 3191 42347
rect 3525 42313 3559 42347
rect 4169 42313 4203 42347
rect 5089 42313 5123 42347
rect 5641 42313 5675 42347
rect 6009 42313 6043 42347
rect 6745 42313 6779 42347
rect 7849 42313 7883 42347
rect 8401 42313 8435 42347
rect 8953 42313 8987 42347
rect 9229 42313 9263 42347
rect 10885 42313 10919 42347
rect 12725 42313 12759 42347
rect 15945 42313 15979 42347
rect 16681 42313 16715 42347
rect 20269 42313 20303 42347
rect 2329 42245 2363 42279
rect 7757 42245 7791 42279
rect 15669 42245 15703 42279
rect 18061 42245 18095 42279
rect 18245 42245 18279 42279
rect 18613 42245 18647 42279
rect 2145 42177 2179 42211
rect 2973 42177 3007 42211
rect 3341 42177 3375 42211
rect 3893 42177 3927 42211
rect 3985 42177 4019 42211
rect 4445 42177 4479 42211
rect 4905 42177 4939 42211
rect 5549 42177 5583 42211
rect 6193 42177 6227 42211
rect 6653 42177 6687 42211
rect 7113 42177 7147 42211
rect 8217 42177 8251 42211
rect 8861 42177 8895 42211
rect 9137 42177 9171 42211
rect 9413 42177 9447 42211
rect 9689 42177 9723 42211
rect 10057 42177 10091 42211
rect 10609 42177 10643 42211
rect 10701 42177 10735 42211
rect 11345 42177 11379 42211
rect 12357 42177 12391 42211
rect 12633 42177 12667 42211
rect 12909 42177 12943 42211
rect 13001 42177 13035 42211
rect 13369 42177 13403 42211
rect 13737 42177 13771 42211
rect 14197 42177 14231 42211
rect 14473 42177 14507 42211
rect 14841 42177 14875 42211
rect 15209 42177 15243 42211
rect 16129 42177 16163 42211
rect 16405 42177 16439 42211
rect 16865 42177 16899 42211
rect 17141 42177 17175 42211
rect 17693 42177 17727 42211
rect 18889 42177 18923 42211
rect 19073 42177 19107 42211
rect 19809 42177 19843 42211
rect 19993 42177 20027 42211
rect 4721 42109 4755 42143
rect 3709 42041 3743 42075
rect 7297 42041 7331 42075
rect 8677 42041 8711 42075
rect 12449 42041 12483 42075
rect 16221 42041 16255 42075
rect 18705 42041 18739 42075
rect 9505 41973 9539 42007
rect 10241 41973 10275 42007
rect 10425 41973 10459 42007
rect 11161 41973 11195 42007
rect 12173 41973 12207 42007
rect 13185 41973 13219 42007
rect 13553 41973 13587 42007
rect 13921 41973 13955 42007
rect 14289 41973 14323 42007
rect 14657 41973 14691 42007
rect 15025 41973 15059 42007
rect 15393 41973 15427 42007
rect 15761 41973 15795 42007
rect 17417 41973 17451 42007
rect 19349 41973 19383 42007
rect 19625 41973 19659 42007
rect 2329 41769 2363 41803
rect 2881 41769 2915 41803
rect 3157 41769 3191 41803
rect 3433 41769 3467 41803
rect 4169 41769 4203 41803
rect 4721 41769 4755 41803
rect 6009 41769 6043 41803
rect 7941 41769 7975 41803
rect 8309 41769 8343 41803
rect 13185 41769 13219 41803
rect 17693 41769 17727 41803
rect 18429 41769 18463 41803
rect 18981 41769 19015 41803
rect 2605 41701 2639 41735
rect 3893 41701 3927 41735
rect 5273 41701 5307 41735
rect 6745 41701 6779 41735
rect 7297 41701 7331 41735
rect 8585 41701 8619 41735
rect 8953 41701 8987 41735
rect 13461 41701 13495 41735
rect 13737 41701 13771 41735
rect 15669 41701 15703 41735
rect 17141 41701 17175 41735
rect 19717 41633 19751 41667
rect 2513 41565 2547 41599
rect 2789 41565 2823 41599
rect 3065 41565 3099 41599
rect 3341 41565 3375 41599
rect 3617 41565 3651 41599
rect 4077 41565 4111 41599
rect 4353 41565 4387 41599
rect 4629 41565 4663 41599
rect 4905 41565 4939 41599
rect 5181 41565 5215 41599
rect 5457 41565 5491 41599
rect 5733 41565 5767 41599
rect 5825 41565 5859 41599
rect 6929 41565 6963 41599
rect 7205 41565 7239 41599
rect 7481 41565 7515 41599
rect 7757 41565 7791 41599
rect 8125 41565 8159 41599
rect 8493 41565 8527 41599
rect 8769 41565 8803 41599
rect 9137 41565 9171 41599
rect 13369 41565 13403 41599
rect 13645 41565 13679 41599
rect 13921 41565 13955 41599
rect 14197 41565 14231 41599
rect 14657 41565 14691 41599
rect 15117 41565 15151 41599
rect 15301 41565 15335 41599
rect 15577 41565 15611 41599
rect 15853 41565 15887 41599
rect 16137 41565 16171 41599
rect 16405 41565 16439 41599
rect 16773 41565 16807 41599
rect 17049 41565 17083 41599
rect 17325 41565 17359 41599
rect 17601 41565 17635 41599
rect 17877 41565 17911 41599
rect 18153 41497 18187 41531
rect 18705 41497 18739 41531
rect 19441 41497 19475 41531
rect 20177 41497 20211 41531
rect 20545 41497 20579 41531
rect 4445 41429 4479 41463
rect 4997 41429 5031 41463
rect 5549 41429 5583 41463
rect 6377 41429 6411 41463
rect 7021 41429 7055 41463
rect 14289 41429 14323 41463
rect 14841 41429 14875 41463
rect 15393 41429 15427 41463
rect 15945 41429 15979 41463
rect 16221 41429 16255 41463
rect 16589 41429 16623 41463
rect 16865 41429 16899 41463
rect 17417 41429 17451 41463
rect 3433 41225 3467 41259
rect 3709 41225 3743 41259
rect 3985 41225 4019 41259
rect 4261 41225 4295 41259
rect 5089 41225 5123 41259
rect 5825 41225 5859 41259
rect 6561 41225 6595 41259
rect 6837 41225 6871 41259
rect 7205 41225 7239 41259
rect 14381 41225 14415 41259
rect 14657 41225 14691 41259
rect 14933 41225 14967 41259
rect 15209 41225 15243 41259
rect 15853 41225 15887 41259
rect 16129 41225 16163 41259
rect 16681 41225 16715 41259
rect 17049 41225 17083 41259
rect 17601 41225 17635 41259
rect 18889 41225 18923 41259
rect 20269 41225 20303 41259
rect 20177 41157 20211 41191
rect 1409 41089 1443 41123
rect 3617 41089 3651 41123
rect 3893 41089 3927 41123
rect 4169 41089 4203 41123
rect 4445 41089 4479 41123
rect 4997 41089 5031 41123
rect 5273 41089 5307 41123
rect 5733 41089 5767 41123
rect 6009 41089 6043 41123
rect 6745 41089 6779 41123
rect 7021 41089 7055 41123
rect 7389 41089 7423 41123
rect 7665 41089 7699 41123
rect 7941 41089 7975 41123
rect 14289 41089 14323 41123
rect 14565 41089 14599 41123
rect 14841 41089 14875 41123
rect 15117 41089 15151 41123
rect 15393 41089 15427 41123
rect 15761 41089 15795 41123
rect 16037 41089 16071 41123
rect 16313 41089 16347 41123
rect 16865 41089 16899 41123
rect 17233 41089 17267 41123
rect 17509 41089 17543 41123
rect 17785 41089 17819 41123
rect 18245 41089 18279 41123
rect 18521 41089 18555 41123
rect 18797 41089 18831 41123
rect 19073 41089 19107 41123
rect 19533 41089 19567 41123
rect 19993 41089 20027 41123
rect 2145 41021 2179 41055
rect 4813 40953 4847 40987
rect 5549 40953 5583 40987
rect 7481 40953 7515 40987
rect 15577 40953 15611 40987
rect 18337 40953 18371 40987
rect 18613 40953 18647 40987
rect 7757 40885 7791 40919
rect 14105 40885 14139 40919
rect 17325 40885 17359 40919
rect 18061 40885 18095 40919
rect 19809 40885 19843 40919
rect 15209 40681 15243 40715
rect 15485 40681 15519 40715
rect 15761 40681 15795 40715
rect 16221 40681 16255 40715
rect 16405 40681 16439 40715
rect 16865 40681 16899 40715
rect 18613 40681 18647 40715
rect 19533 40681 19567 40715
rect 17325 40613 17359 40647
rect 18153 40613 18187 40647
rect 19257 40613 19291 40647
rect 1409 40477 1443 40511
rect 1685 40477 1719 40511
rect 15117 40477 15151 40511
rect 15393 40477 15427 40511
rect 15669 40477 15703 40511
rect 15945 40477 15979 40511
rect 16037 40477 16071 40511
rect 16589 40477 16623 40511
rect 17049 40477 17083 40511
rect 17509 40477 17543 40511
rect 17785 40477 17819 40511
rect 18061 40477 18095 40511
rect 18337 40477 18371 40511
rect 18797 40477 18831 40511
rect 19073 40477 19107 40511
rect 19441 40477 19475 40511
rect 19717 40477 19751 40511
rect 19993 40477 20027 40511
rect 1961 40409 1995 40443
rect 2697 40409 2731 40443
rect 20177 40409 20211 40443
rect 20545 40409 20579 40443
rect 14933 40341 14967 40375
rect 17601 40341 17635 40375
rect 17877 40341 17911 40375
rect 18889 40341 18923 40375
rect 19809 40341 19843 40375
rect 16129 40137 16163 40171
rect 16865 40137 16899 40171
rect 17141 40137 17175 40171
rect 17417 40137 17451 40171
rect 17969 40137 18003 40171
rect 1409 40069 1443 40103
rect 2789 40069 2823 40103
rect 20177 40069 20211 40103
rect 2513 40001 2547 40035
rect 3065 40001 3099 40035
rect 3341 40001 3375 40035
rect 4811 40001 4845 40035
rect 7907 40001 7941 40035
rect 14657 40001 14691 40035
rect 17049 40001 17083 40035
rect 17325 40001 17359 40035
rect 17601 40001 17635 40035
rect 17877 40001 17911 40035
rect 18153 40001 18187 40035
rect 18613 40001 18647 40035
rect 19073 40001 19107 40035
rect 19441 40001 19475 40035
rect 19717 40001 19751 40035
rect 19993 40001 20027 40035
rect 2145 39933 2179 39967
rect 4537 39933 4571 39967
rect 7665 39933 7699 39967
rect 17693 39865 17727 39899
rect 19257 39865 19291 39899
rect 5549 39797 5583 39831
rect 8677 39797 8711 39831
rect 18429 39797 18463 39831
rect 18889 39797 18923 39831
rect 19533 39797 19567 39831
rect 19809 39797 19843 39831
rect 20453 39797 20487 39831
rect 15301 39593 15335 39627
rect 16957 39593 16991 39627
rect 17233 39593 17267 39627
rect 17785 39593 17819 39627
rect 18337 39593 18371 39627
rect 18889 39593 18923 39627
rect 19625 39593 19659 39627
rect 7389 39525 7423 39559
rect 16221 39525 16255 39559
rect 16405 39525 16439 39559
rect 16681 39525 16715 39559
rect 18061 39525 18095 39559
rect 18613 39525 18647 39559
rect 6377 39457 6411 39491
rect 1409 39389 1443 39423
rect 1961 39389 1995 39423
rect 2235 39389 2269 39423
rect 3801 39389 3835 39423
rect 4075 39389 4109 39423
rect 6651 39389 6685 39423
rect 15485 39389 15519 39423
rect 16589 39389 16623 39423
rect 16865 39389 16899 39423
rect 17141 39389 17175 39423
rect 17417 39389 17451 39423
rect 17693 39389 17727 39423
rect 17969 39389 18003 39423
rect 18245 39389 18279 39423
rect 18521 39389 18555 39423
rect 18797 39389 18831 39423
rect 19073 39389 19107 39423
rect 19533 39389 19567 39423
rect 19809 39389 19843 39423
rect 1685 39321 1719 39355
rect 20177 39321 20211 39355
rect 20545 39321 20579 39355
rect 2973 39253 3007 39287
rect 4813 39253 4847 39287
rect 17509 39253 17543 39287
rect 19349 39253 19383 39287
rect 16497 39049 16531 39083
rect 17049 39049 17083 39083
rect 17693 39049 17727 39083
rect 18521 39049 18555 39083
rect 18797 39049 18831 39083
rect 19073 39049 19107 39083
rect 19441 39049 19475 39083
rect 2237 38981 2271 39015
rect 4537 38981 4571 39015
rect 4813 38981 4847 39015
rect 4905 38981 4939 39015
rect 20177 38981 20211 39015
rect 1409 38913 1443 38947
rect 1961 38913 1995 38947
rect 2955 38943 2989 38977
rect 5273 38913 5307 38947
rect 5655 38913 5689 38947
rect 7941 38913 7975 38947
rect 15373 38913 15407 38947
rect 17233 38913 17267 38947
rect 17509 38913 17543 38947
rect 17877 38913 17911 38947
rect 18153 38913 18187 38947
rect 18437 38913 18471 38947
rect 18705 38913 18739 38947
rect 18981 38913 19015 38947
rect 19257 38913 19291 38947
rect 19625 38913 19659 38947
rect 19993 38913 20027 38947
rect 1685 38845 1719 38879
rect 2697 38845 2731 38879
rect 4261 38845 4295 38879
rect 6745 38845 6779 38879
rect 6929 38845 6963 38879
rect 7389 38845 7423 38879
rect 7665 38845 7699 38879
rect 7803 38845 7837 38879
rect 15117 38845 15151 38879
rect 17325 38777 17359 38811
rect 18245 38777 18279 38811
rect 3709 38709 3743 38743
rect 5825 38709 5859 38743
rect 8585 38709 8619 38743
rect 17969 38709 18003 38743
rect 19809 38709 19843 38743
rect 20453 38709 20487 38743
rect 18521 38505 18555 38539
rect 15485 38437 15519 38471
rect 18245 38437 18279 38471
rect 18889 38437 18923 38471
rect 2329 38369 2363 38403
rect 16865 38369 16899 38403
rect 1409 38301 1443 38335
rect 2603 38301 2637 38335
rect 4353 38301 4387 38335
rect 10517 38301 10551 38335
rect 10791 38301 10825 38335
rect 13921 38301 13955 38335
rect 14105 38301 14139 38335
rect 15761 38301 15795 38335
rect 16221 38301 16255 38335
rect 16773 38301 16807 38335
rect 17509 38301 17543 38335
rect 17693 38301 17727 38335
rect 17969 38301 18003 38335
rect 18153 38301 18187 38335
rect 18429 38301 18463 38335
rect 18705 38301 18739 38335
rect 19073 38301 19107 38335
rect 19441 38301 19475 38335
rect 19533 38301 19567 38335
rect 19809 38301 19843 38335
rect 19993 38301 20027 38335
rect 20177 38301 20211 38335
rect 1685 38233 1719 38267
rect 4261 38233 4295 38267
rect 4721 38233 4755 38267
rect 11989 38233 12023 38267
rect 12173 38233 12207 38267
rect 14350 38233 14384 38267
rect 17785 38233 17819 38267
rect 17877 38233 17911 38267
rect 18061 38233 18095 38267
rect 20545 38233 20579 38267
rect 3341 38165 3375 38199
rect 3985 38165 4019 38199
rect 5089 38165 5123 38199
rect 5273 38165 5307 38199
rect 11529 38165 11563 38199
rect 13737 38165 13771 38199
rect 15577 38165 15611 38199
rect 16037 38165 16071 38199
rect 19257 38165 19291 38199
rect 19625 38165 19659 38199
rect 19993 38165 20027 38199
rect 2881 37961 2915 37995
rect 3985 37961 4019 37995
rect 5365 37961 5399 37995
rect 9965 37961 9999 37995
rect 12541 37961 12575 37995
rect 17693 37961 17727 37995
rect 18705 37961 18739 37995
rect 19257 37961 19291 37995
rect 1685 37893 1719 37927
rect 3249 37893 3283 37927
rect 10241 37893 10275 37927
rect 11069 37893 11103 37927
rect 1409 37825 1443 37859
rect 1961 37825 1995 37859
rect 3157 37825 3191 37859
rect 3617 37825 3651 37859
rect 5549 37825 5583 37859
rect 7295 37825 7329 37859
rect 10333 37825 10367 37859
rect 10701 37825 10735 37859
rect 11803 37825 11837 37859
rect 14473 37825 14507 37859
rect 14565 37825 14599 37859
rect 15025 37825 15059 37859
rect 15209 37825 15243 37859
rect 15301 37825 15335 37859
rect 15393 37825 15427 37859
rect 15485 37825 15519 37859
rect 15669 37825 15703 37859
rect 16955 37825 16989 37859
rect 18889 37825 18923 37859
rect 19165 37825 19199 37859
rect 19441 37825 19475 37859
rect 19717 37825 19751 37859
rect 19993 37825 20027 37859
rect 20177 37825 20211 37859
rect 2237 37757 2271 37791
rect 7021 37757 7055 37791
rect 11529 37757 11563 37791
rect 15577 37757 15611 37791
rect 16681 37757 16715 37791
rect 18981 37689 19015 37723
rect 19533 37689 19567 37723
rect 4169 37621 4203 37655
rect 8033 37621 8067 37655
rect 8953 37621 8987 37655
rect 11253 37621 11287 37655
rect 19809 37621 19843 37655
rect 20453 37621 20487 37655
rect 2697 37417 2731 37451
rect 15117 37417 15151 37451
rect 18797 37417 18831 37451
rect 18245 37349 18279 37383
rect 18521 37349 18555 37383
rect 1685 37281 1719 37315
rect 5917 37281 5951 37315
rect 7481 37281 7515 37315
rect 14105 37281 14139 37315
rect 20269 37281 20303 37315
rect 1959 37213 1993 37247
rect 3065 37213 3099 37247
rect 3801 37213 3835 37247
rect 6191 37213 6225 37247
rect 7739 37183 7773 37217
rect 8953 37213 8987 37247
rect 9227 37213 9261 37247
rect 11069 37213 11103 37247
rect 11343 37213 11377 37247
rect 14379 37213 14413 37247
rect 18153 37213 18187 37247
rect 18429 37213 18463 37247
rect 18705 37213 18739 37247
rect 18981 37213 19015 37247
rect 19993 37213 20027 37247
rect 3341 37145 3375 37179
rect 4077 37145 4111 37179
rect 19441 37145 19475 37179
rect 19809 37145 19843 37179
rect 6929 37077 6963 37111
rect 8493 37077 8527 37111
rect 9965 37077 9999 37111
rect 12081 37077 12115 37111
rect 17969 37077 18003 37111
rect 9689 36873 9723 36907
rect 17969 36873 18003 36907
rect 19901 36873 19935 36907
rect 3341 36805 3375 36839
rect 18788 36805 18822 36839
rect 1501 36737 1535 36771
rect 1961 36737 1995 36771
rect 3065 36737 3099 36771
rect 3617 36737 3651 36771
rect 4261 36737 4295 36771
rect 8769 36737 8803 36771
rect 9045 36737 9079 36771
rect 10055 36737 10089 36771
rect 11803 36737 11837 36771
rect 13995 36767 14029 36801
rect 15117 36737 15151 36771
rect 15301 36737 15335 36771
rect 15761 36737 15795 36771
rect 18153 36737 18187 36771
rect 18429 36737 18463 36771
rect 20177 36737 20211 36771
rect 2789 36669 2823 36703
rect 3801 36669 3835 36703
rect 7849 36669 7883 36703
rect 8033 36669 8067 36703
rect 8493 36669 8527 36703
rect 8886 36669 8920 36703
rect 9781 36669 9815 36703
rect 11529 36669 11563 36703
rect 13737 36669 13771 36703
rect 18521 36669 18555 36703
rect 1777 36533 1811 36567
rect 4537 36533 4571 36567
rect 10793 36533 10827 36567
rect 12541 36533 12575 36567
rect 14749 36533 14783 36567
rect 15209 36533 15243 36567
rect 15577 36533 15611 36567
rect 18245 36533 18279 36567
rect 20453 36533 20487 36567
rect 3433 36329 3467 36363
rect 8401 36329 8435 36363
rect 18061 36329 18095 36363
rect 18613 36329 18647 36363
rect 5549 36261 5583 36295
rect 7205 36261 7239 36295
rect 17141 36261 17175 36295
rect 18889 36261 18923 36295
rect 20269 36261 20303 36295
rect 2237 36193 2271 36227
rect 2513 36193 2547 36227
rect 7598 36193 7632 36227
rect 7757 36193 7791 36227
rect 9505 36193 9539 36227
rect 11253 36193 11287 36227
rect 14105 36193 14139 36227
rect 19257 36193 19291 36227
rect 1593 36125 1627 36159
rect 1777 36125 1811 36159
rect 2630 36125 2664 36159
rect 2789 36125 2823 36159
rect 4537 36125 4571 36159
rect 6561 36125 6595 36159
rect 6745 36125 6779 36159
rect 7481 36125 7515 36159
rect 9747 36125 9781 36159
rect 11527 36125 11561 36159
rect 13921 36125 13955 36159
rect 15669 36125 15703 36159
rect 17325 36125 17359 36159
rect 17417 36125 17451 36159
rect 17877 36125 17911 36159
rect 18245 36101 18279 36135
rect 18521 36125 18555 36159
rect 18797 36125 18831 36159
rect 19073 36125 19107 36159
rect 19499 36125 19533 36159
rect 4629 36057 4663 36091
rect 4997 36057 5031 36091
rect 14350 36057 14384 36091
rect 15914 36057 15948 36091
rect 4261 35989 4295 36023
rect 5365 35989 5399 36023
rect 10517 35989 10551 36023
rect 12265 35989 12299 36023
rect 13737 35989 13771 36023
rect 15485 35989 15519 36023
rect 17049 35989 17083 36023
rect 17509 35989 17543 36023
rect 17693 35989 17727 36023
rect 18337 35989 18371 36023
rect 2513 35785 2547 35819
rect 3893 35785 3927 35819
rect 5365 35785 5399 35819
rect 10701 35785 10735 35819
rect 13369 35785 13403 35819
rect 15393 35785 15427 35819
rect 16129 35785 16163 35819
rect 18429 35785 18463 35819
rect 9413 35717 9447 35751
rect 9689 35717 9723 35751
rect 9781 35717 9815 35751
rect 10517 35717 10551 35751
rect 15301 35717 15335 35751
rect 20269 35717 20303 35751
rect 1775 35649 1809 35683
rect 2881 35649 2915 35683
rect 3155 35649 3189 35683
rect 4627 35649 4661 35683
rect 10149 35649 10183 35683
rect 10977 35649 11011 35683
rect 12725 35649 12759 35683
rect 14473 35649 14507 35683
rect 14565 35649 14599 35683
rect 14933 35649 14967 35683
rect 15577 35649 15611 35683
rect 16313 35649 16347 35683
rect 17049 35649 17083 35683
rect 17417 35649 17451 35683
rect 17601 35649 17635 35683
rect 17877 35649 17911 35683
rect 18153 35649 18187 35683
rect 18613 35649 18647 35683
rect 18889 35649 18923 35683
rect 19349 35649 19383 35683
rect 19625 35649 19659 35683
rect 19901 35649 19935 35683
rect 20085 35649 20119 35683
rect 20545 35649 20579 35683
rect 1501 35581 1535 35615
rect 4353 35581 4387 35615
rect 11529 35581 11563 35615
rect 11713 35581 11747 35615
rect 12173 35581 12207 35615
rect 12449 35581 12483 35615
rect 12587 35581 12621 35615
rect 14749 35581 14783 35615
rect 17141 35581 17175 35615
rect 17325 35581 17359 35615
rect 17509 35581 17543 35615
rect 11161 35513 11195 35547
rect 15117 35513 15151 35547
rect 17969 35513 18003 35547
rect 20177 35513 20211 35547
rect 17233 35445 17267 35479
rect 17693 35445 17727 35479
rect 18705 35445 18739 35479
rect 19165 35445 19199 35479
rect 19441 35445 19475 35479
rect 20361 35445 20395 35479
rect 2421 35241 2455 35275
rect 4813 35241 4847 35275
rect 13369 35241 13403 35275
rect 17141 35241 17175 35275
rect 18889 35241 18923 35275
rect 20269 35241 20303 35275
rect 12173 35173 12207 35207
rect 15853 35173 15887 35207
rect 1409 35105 1443 35139
rect 3065 35105 3099 35139
rect 11713 35105 11747 35139
rect 13645 35105 13679 35139
rect 1683 35037 1717 35071
rect 2789 35037 2823 35071
rect 3801 35037 3835 35071
rect 4997 35037 5031 35071
rect 5089 35037 5123 35071
rect 5363 35037 5397 35071
rect 6469 35037 6503 35071
rect 6743 35037 6777 35071
rect 8585 35037 8619 35071
rect 9505 35037 9539 35071
rect 9763 35007 9797 35041
rect 11529 35037 11563 35071
rect 12449 35037 12483 35071
rect 12587 35037 12621 35071
rect 12725 35037 12759 35071
rect 14381 35037 14415 35071
rect 14655 35037 14689 35071
rect 16037 35037 16071 35071
rect 16129 35037 16163 35071
rect 16371 35037 16405 35071
rect 17509 35037 17543 35071
rect 17783 35037 17817 35071
rect 19073 35037 19107 35071
rect 19993 35037 20027 35071
rect 4077 34969 4111 35003
rect 19441 34969 19475 35003
rect 19809 34969 19843 35003
rect 6101 34901 6135 34935
rect 7481 34901 7515 34935
rect 8401 34901 8435 34935
rect 10517 34901 10551 34935
rect 15393 34901 15427 34935
rect 18521 34901 18555 34935
rect 5457 34697 5491 34731
rect 8217 34697 8251 34731
rect 8861 34697 8895 34731
rect 10425 34697 10459 34731
rect 12817 34697 12851 34731
rect 18429 34697 18463 34731
rect 19441 34697 19475 34731
rect 4169 34629 4203 34663
rect 7113 34629 7147 34663
rect 7389 34629 7423 34663
rect 7481 34629 7515 34663
rect 9321 34629 9355 34663
rect 9597 34629 9631 34663
rect 9689 34629 9723 34663
rect 10885 34629 10919 34663
rect 20177 34629 20211 34663
rect 1409 34561 1443 34595
rect 1961 34561 1995 34595
rect 2513 34561 2547 34595
rect 2787 34561 2821 34595
rect 3893 34561 3927 34595
rect 4445 34561 4479 34595
rect 4719 34561 4753 34595
rect 7849 34561 7883 34595
rect 8585 34561 8619 34595
rect 10057 34561 10091 34595
rect 11793 34561 11827 34595
rect 12079 34561 12113 34595
rect 13921 34561 13955 34595
rect 14195 34561 14229 34595
rect 16681 34561 16715 34595
rect 16948 34561 16982 34595
rect 18153 34561 18187 34595
rect 18705 34561 18739 34595
rect 18797 34561 18831 34595
rect 18981 34561 19015 34595
rect 19349 34561 19383 34595
rect 19625 34561 19659 34595
rect 19901 34561 19935 34595
rect 1685 34493 1719 34527
rect 2237 34493 2271 34527
rect 8861 34493 8895 34527
rect 11069 34493 11103 34527
rect 18429 34493 18463 34527
rect 18889 34493 18923 34527
rect 18061 34425 18095 34459
rect 18521 34425 18555 34459
rect 3525 34357 3559 34391
rect 8401 34357 8435 34391
rect 8677 34357 8711 34391
rect 10609 34357 10643 34391
rect 14933 34357 14967 34391
rect 18245 34357 18279 34391
rect 19165 34357 19199 34391
rect 19717 34357 19751 34391
rect 20453 34357 20487 34391
rect 4629 34153 4663 34187
rect 8677 34153 8711 34187
rect 10057 34153 10091 34187
rect 13737 34153 13771 34187
rect 17601 34153 17635 34187
rect 17785 34153 17819 34187
rect 18613 34153 18647 34187
rect 19533 34153 19567 34187
rect 7205 34085 7239 34119
rect 8401 34085 8435 34119
rect 10517 34085 10551 34119
rect 13829 34085 13863 34119
rect 18061 34085 18095 34119
rect 1685 34017 1719 34051
rect 2329 34017 2363 34051
rect 4997 34017 5031 34051
rect 7481 34017 7515 34051
rect 7619 34017 7653 34051
rect 13921 34017 13955 34051
rect 1409 33949 1443 33983
rect 2587 33919 2621 33953
rect 3801 33949 3835 33983
rect 4813 33949 4847 33983
rect 5271 33949 5305 33983
rect 6561 33949 6595 33983
rect 6745 33949 6779 33983
rect 7757 33949 7791 33983
rect 8585 33949 8619 33983
rect 8769 33949 8803 33983
rect 9045 33949 9079 33983
rect 9319 33939 9353 33973
rect 10425 33949 10459 33983
rect 10793 33949 10827 33983
rect 11067 33949 11101 33983
rect 13645 33949 13679 33983
rect 14105 33949 14139 33983
rect 14379 33949 14413 33983
rect 15485 33949 15519 33983
rect 15759 33949 15793 33983
rect 17049 33949 17083 33983
rect 17509 33949 17543 33983
rect 17969 33949 18003 33983
rect 18245 33949 18279 33983
rect 18521 33949 18555 33983
rect 18797 33949 18831 33983
rect 19073 33949 19107 33983
rect 19441 33949 19475 33983
rect 19625 33949 19659 33983
rect 19993 33949 20027 33983
rect 20269 33949 20303 33983
rect 4077 33881 4111 33915
rect 3341 33813 3375 33847
rect 6009 33813 6043 33847
rect 11805 33813 11839 33847
rect 15117 33813 15151 33847
rect 16497 33813 16531 33847
rect 16865 33813 16899 33847
rect 18337 33813 18371 33847
rect 18889 33813 18923 33847
rect 19809 33813 19843 33847
rect 20453 33813 20487 33847
rect 9965 33609 9999 33643
rect 15853 33609 15887 33643
rect 18613 33609 18647 33643
rect 19165 33609 19199 33643
rect 3709 33541 3743 33575
rect 3985 33541 4019 33575
rect 4077 33541 4111 33575
rect 4813 33541 4847 33575
rect 8493 33541 8527 33575
rect 20177 33541 20211 33575
rect 1667 33503 1701 33537
rect 2789 33473 2823 33507
rect 3065 33473 3099 33507
rect 4445 33473 4479 33507
rect 6653 33473 6687 33507
rect 7573 33473 7607 33507
rect 7690 33473 7724 33507
rect 8585 33473 8619 33507
rect 8859 33473 8893 33507
rect 10149 33473 10183 33507
rect 11529 33473 11563 33507
rect 11803 33473 11837 33507
rect 15209 33473 15243 33507
rect 15945 33473 15979 33507
rect 16129 33473 16163 33507
rect 18797 33473 18831 33507
rect 19073 33473 19107 33507
rect 19349 33473 19383 33507
rect 19809 33473 19843 33507
rect 1409 33405 1443 33439
rect 6837 33405 6871 33439
rect 7849 33405 7883 33439
rect 14013 33405 14047 33439
rect 14197 33405 14231 33439
rect 14657 33405 14691 33439
rect 14933 33405 14967 33439
rect 15050 33405 15084 33439
rect 4997 33337 5031 33371
rect 7297 33337 7331 33371
rect 9597 33337 9631 33371
rect 19625 33337 19659 33371
rect 2421 33269 2455 33303
rect 12541 33269 12575 33303
rect 16037 33269 16071 33303
rect 18889 33269 18923 33303
rect 20453 33269 20487 33303
rect 4721 33065 4755 33099
rect 8309 33065 8343 33099
rect 13001 33065 13035 33099
rect 15485 33065 15519 33099
rect 18797 33065 18831 33099
rect 11805 32997 11839 33031
rect 15853 32997 15887 33031
rect 19901 32997 19935 33031
rect 1961 32929 1995 32963
rect 8953 32929 8987 32963
rect 12081 32929 12115 32963
rect 12357 32929 12391 32963
rect 14105 32929 14139 32963
rect 19533 32929 19567 32963
rect 1409 32861 1443 32895
rect 2235 32861 2269 32895
rect 3801 32861 3835 32895
rect 4077 32861 4111 32895
rect 4905 32861 4939 32895
rect 5549 32861 5583 32895
rect 7297 32861 7331 32895
rect 7539 32861 7573 32895
rect 9195 32861 9229 32895
rect 11161 32861 11195 32895
rect 11345 32861 11379 32895
rect 12198 32861 12232 32895
rect 14347 32861 14381 32895
rect 15669 32861 15703 32895
rect 15761 32861 15795 32895
rect 17785 32861 17819 32895
rect 18027 32861 18061 32895
rect 19257 32861 19291 32895
rect 19349 32861 19383 32895
rect 19717 32861 19751 32895
rect 20177 32861 20211 32895
rect 1685 32793 1719 32827
rect 5457 32793 5491 32827
rect 5917 32793 5951 32827
rect 20545 32793 20579 32827
rect 2973 32725 3007 32759
rect 5181 32725 5215 32759
rect 6285 32725 6319 32759
rect 6469 32725 6503 32759
rect 9965 32725 9999 32759
rect 15117 32725 15151 32759
rect 19533 32725 19567 32759
rect 8125 32521 8159 32555
rect 13829 32521 13863 32555
rect 16037 32521 16071 32555
rect 17141 32521 17175 32555
rect 18797 32521 18831 32555
rect 20361 32521 20395 32555
rect 2237 32453 2271 32487
rect 2513 32453 2547 32487
rect 2605 32453 2639 32487
rect 3341 32453 3375 32487
rect 1409 32385 1443 32419
rect 2973 32385 3007 32419
rect 3709 32385 3743 32419
rect 3985 32385 4019 32419
rect 4719 32385 4753 32419
rect 7113 32385 7147 32419
rect 7387 32385 7421 32419
rect 9229 32385 9263 32419
rect 9779 32385 9813 32419
rect 12631 32385 12665 32419
rect 14013 32385 14047 32419
rect 15301 32385 15335 32419
rect 16221 32385 16255 32419
rect 16313 32385 16347 32419
rect 17325 32385 17359 32419
rect 17417 32385 17451 32419
rect 17673 32385 17707 32419
rect 18889 32385 18923 32419
rect 19145 32385 19179 32419
rect 20545 32385 20579 32419
rect 1685 32317 1719 32351
rect 4445 32317 4479 32351
rect 9505 32317 9539 32351
rect 12357 32317 12391 32351
rect 14105 32317 14139 32351
rect 14289 32317 14323 32351
rect 15025 32317 15059 32351
rect 15142 32317 15176 32351
rect 3525 32249 3559 32283
rect 14749 32249 14783 32283
rect 20269 32249 20303 32283
rect 5457 32181 5491 32215
rect 9321 32181 9355 32215
rect 10517 32181 10551 32215
rect 13369 32181 13403 32215
rect 15945 32181 15979 32215
rect 16405 32181 16439 32215
rect 6469 31977 6503 32011
rect 15945 31977 15979 32011
rect 18337 31977 18371 32011
rect 3249 31909 3283 31943
rect 10793 31909 10827 31943
rect 14749 31909 14783 31943
rect 17601 31909 17635 31943
rect 1501 31841 1535 31875
rect 9781 31841 9815 31875
rect 14289 31841 14323 31875
rect 15025 31841 15059 31875
rect 15142 31841 15176 31875
rect 15301 31841 15335 31875
rect 16037 31841 16071 31875
rect 19257 31841 19291 31875
rect 1759 31743 1793 31777
rect 3065 31773 3099 31807
rect 4629 31773 4663 31807
rect 5549 31773 5583 31807
rect 5917 31773 5951 31807
rect 6929 31773 6963 31807
rect 7203 31773 7237 31807
rect 10023 31773 10057 31807
rect 11621 31773 11655 31807
rect 11713 31773 11747 31807
rect 14105 31773 14139 31807
rect 16295 31743 16329 31777
rect 17785 31773 17819 31807
rect 18245 31773 18279 31807
rect 18521 31773 18555 31807
rect 18705 31773 18739 31807
rect 19531 31773 19565 31807
rect 3433 31705 3467 31739
rect 3617 31705 3651 31739
rect 3801 31705 3835 31739
rect 5181 31705 5215 31739
rect 5457 31705 5491 31739
rect 6285 31705 6319 31739
rect 12081 31705 12115 31739
rect 2513 31637 2547 31671
rect 7941 31637 7975 31671
rect 11345 31637 11379 31671
rect 12449 31637 12483 31671
rect 12633 31637 12667 31671
rect 17049 31637 17083 31671
rect 18061 31637 18095 31671
rect 18981 31637 19015 31671
rect 20269 31637 20303 31671
rect 5917 31433 5951 31467
rect 10977 31433 11011 31467
rect 12541 31433 12575 31467
rect 14749 31433 14783 31467
rect 15853 31433 15887 31467
rect 16221 31433 16255 31467
rect 18153 31433 18187 31467
rect 18613 31433 18647 31467
rect 20177 31365 20211 31399
rect 1685 31297 1719 31331
rect 2755 31297 2789 31331
rect 3893 31297 3927 31331
rect 5179 31297 5213 31331
rect 7297 31297 7331 31331
rect 7555 31327 7589 31361
rect 10057 31297 10091 31331
rect 10333 31297 10367 31331
rect 11529 31297 11563 31331
rect 11803 31297 11837 31331
rect 13093 31297 13127 31331
rect 15083 31297 15117 31331
rect 16405 31297 16439 31331
rect 16681 31297 16715 31331
rect 16865 31297 16899 31331
rect 18061 31297 18095 31331
rect 18337 31297 18371 31331
rect 18429 31297 18463 31331
rect 18613 31297 18647 31331
rect 18705 31297 18739 31331
rect 19165 31303 19199 31337
rect 19625 31297 19659 31331
rect 19717 31297 19751 31331
rect 1409 31229 1443 31263
rect 2513 31229 2547 31263
rect 4169 31229 4203 31263
rect 4905 31229 4939 31263
rect 9137 31229 9171 31263
rect 9321 31229 9355 31263
rect 10195 31229 10229 31263
rect 12909 31229 12943 31263
rect 13553 31229 13587 31263
rect 13829 31229 13863 31263
rect 13967 31229 14001 31263
rect 14105 31229 14139 31263
rect 14841 31229 14875 31263
rect 19993 31229 20027 31263
rect 9781 31161 9815 31195
rect 19257 31161 19291 31195
rect 19809 31161 19843 31195
rect 3525 31093 3559 31127
rect 8309 31093 8343 31127
rect 16773 31093 16807 31127
rect 17877 31093 17911 31127
rect 18797 31093 18831 31127
rect 19441 31093 19475 31127
rect 19901 31093 19935 31127
rect 20453 31093 20487 31127
rect 3433 30889 3467 30923
rect 15945 30889 15979 30923
rect 19257 30889 19291 30923
rect 8309 30821 8343 30855
rect 14749 30821 14783 30855
rect 17969 30821 18003 30855
rect 18613 30821 18647 30855
rect 18889 30821 18923 30855
rect 2237 30753 2271 30787
rect 2630 30753 2664 30787
rect 9413 30753 9447 30787
rect 10793 30753 10827 30787
rect 15301 30753 15335 30787
rect 16221 30753 16255 30787
rect 1593 30685 1627 30719
rect 1777 30685 1811 30719
rect 2513 30685 2547 30719
rect 2789 30685 2823 30719
rect 3801 30685 3835 30719
rect 4077 30685 4111 30719
rect 4351 30685 4385 30719
rect 7297 30685 7331 30719
rect 7389 30685 7423 30719
rect 8493 30685 8527 30719
rect 8677 30685 8711 30719
rect 9687 30685 9721 30719
rect 11035 30685 11069 30719
rect 14105 30685 14139 30719
rect 14289 30685 14323 30719
rect 15025 30685 15059 30719
rect 15142 30685 15176 30719
rect 16405 30685 16439 30719
rect 16865 30685 16899 30719
rect 17233 30685 17267 30719
rect 17785 30685 17819 30719
rect 18153 30685 18187 30719
rect 18797 30685 18831 30719
rect 19073 30685 19107 30719
rect 19441 30685 19475 30719
rect 19717 30685 19751 30719
rect 19993 30685 20027 30719
rect 7021 30617 7055 30651
rect 7757 30617 7791 30651
rect 17141 30617 17175 30651
rect 20177 30617 20211 30651
rect 20545 30617 20579 30651
rect 3985 30549 4019 30583
rect 5089 30549 5123 30583
rect 8125 30549 8159 30583
rect 8585 30549 8619 30583
rect 10425 30549 10459 30583
rect 11805 30549 11839 30583
rect 17325 30549 17359 30583
rect 17601 30549 17635 30583
rect 19533 30549 19567 30583
rect 19809 30549 19843 30583
rect 16313 30345 16347 30379
rect 18061 30345 18095 30379
rect 19073 30345 19107 30379
rect 19441 30345 19475 30379
rect 1501 30277 1535 30311
rect 5825 30277 5859 30311
rect 8585 30277 8619 30311
rect 14841 30277 14875 30311
rect 16926 30277 16960 30311
rect 2991 30209 3025 30243
rect 3985 30209 4019 30243
rect 5181 30209 5215 30243
rect 7171 30209 7205 30243
rect 8309 30209 8343 30243
rect 8677 30209 8711 30243
rect 8951 30209 8985 30243
rect 14038 30209 14072 30243
rect 14933 30209 14967 30243
rect 15207 30209 15241 30243
rect 16497 30209 16531 30243
rect 16681 30209 16715 30243
rect 18153 30209 18187 30243
rect 18521 30209 18555 30243
rect 18705 30209 18739 30243
rect 18981 30209 19015 30243
rect 19257 30209 19291 30243
rect 19625 30209 19659 30243
rect 19717 30209 19751 30243
rect 19901 30209 19935 30243
rect 20177 30209 20211 30243
rect 2053 30141 2087 30175
rect 2237 30141 2271 30175
rect 3090 30141 3124 30175
rect 3235 30141 3269 30175
rect 4169 30141 4203 30175
rect 4905 30141 4939 30175
rect 5043 30141 5077 30175
rect 6929 30141 6963 30175
rect 8585 30141 8619 30175
rect 13001 30141 13035 30175
rect 13185 30141 13219 30175
rect 13921 30141 13955 30175
rect 14197 30141 14231 30175
rect 18245 30141 18279 30175
rect 18429 30141 18463 30175
rect 18613 30141 18647 30175
rect 2697 30073 2731 30107
rect 3893 30073 3927 30107
rect 4629 30073 4663 30107
rect 7941 30073 7975 30107
rect 8401 30073 8435 30107
rect 13645 30073 13679 30107
rect 18797 30073 18831 30107
rect 1777 30005 1811 30039
rect 9689 30005 9723 30039
rect 15945 30005 15979 30039
rect 18337 30005 18371 30039
rect 19809 30005 19843 30039
rect 20453 30005 20487 30039
rect 2881 29801 2915 29835
rect 4813 29801 4847 29835
rect 8309 29801 8343 29835
rect 13461 29801 13495 29835
rect 17785 29801 17819 29835
rect 18613 29801 18647 29835
rect 19809 29801 19843 29835
rect 6009 29733 6043 29767
rect 19257 29733 19291 29767
rect 1869 29665 1903 29699
rect 3801 29665 3835 29699
rect 6402 29665 6436 29699
rect 6561 29665 6595 29699
rect 7297 29665 7331 29699
rect 9045 29665 9079 29699
rect 12449 29665 12483 29699
rect 16773 29665 16807 29699
rect 2143 29597 2177 29631
rect 3341 29597 3375 29631
rect 4075 29597 4109 29631
rect 5365 29597 5399 29631
rect 5549 29597 5583 29631
rect 6285 29597 6319 29631
rect 7539 29597 7573 29631
rect 9319 29597 9353 29631
rect 10885 29597 10919 29631
rect 10977 29597 11011 29631
rect 12691 29597 12725 29631
rect 14289 29597 14323 29631
rect 14563 29597 14597 29631
rect 17047 29597 17081 29631
rect 18797 29597 18831 29631
rect 19073 29597 19107 29631
rect 19441 29597 19475 29631
rect 1501 29529 1535 29563
rect 1685 29529 1719 29563
rect 3525 29529 3559 29563
rect 11345 29529 11379 29563
rect 20177 29529 20211 29563
rect 20545 29529 20579 29563
rect 7205 29461 7239 29495
rect 10057 29461 10091 29495
rect 10609 29461 10643 29495
rect 11713 29461 11747 29495
rect 11897 29461 11931 29495
rect 15301 29461 15335 29495
rect 18889 29461 18923 29495
rect 2421 29257 2455 29291
rect 4445 29257 4479 29291
rect 4721 29257 4755 29291
rect 9781 29257 9815 29291
rect 18429 29257 18463 29291
rect 18705 29257 18739 29291
rect 18981 29257 19015 29291
rect 8677 29189 8711 29223
rect 8953 29189 8987 29223
rect 9045 29189 9079 29223
rect 9413 29189 9447 29223
rect 10241 29189 10275 29223
rect 20177 29189 20211 29223
rect 1409 29121 1443 29155
rect 1683 29131 1717 29165
rect 2881 29121 2915 29155
rect 3123 29121 3157 29155
rect 4261 29121 4295 29155
rect 4537 29121 4571 29155
rect 4905 29121 4939 29155
rect 5179 29121 5213 29155
rect 7021 29121 7055 29155
rect 7371 29151 7405 29185
rect 11803 29121 11837 29155
rect 13427 29121 13461 29155
rect 14807 29121 14841 29155
rect 18613 29121 18647 29155
rect 18889 29121 18923 29155
rect 19165 29121 19199 29155
rect 19441 29121 19475 29155
rect 19533 29121 19567 29155
rect 19993 29121 20027 29155
rect 7113 29053 7147 29087
rect 11529 29053 11563 29087
rect 13185 29053 13219 29087
rect 14565 29053 14599 29087
rect 3893 28985 3927 29019
rect 6837 28985 6871 29019
rect 8125 28985 8159 29019
rect 10425 28985 10459 29019
rect 12541 28985 12575 29019
rect 20453 28985 20487 29019
rect 5917 28917 5951 28951
rect 9965 28917 9999 28951
rect 14197 28917 14231 28951
rect 15577 28917 15611 28951
rect 19257 28917 19291 28951
rect 19625 28917 19659 28951
rect 19809 28917 19843 28951
rect 8125 28713 8159 28747
rect 15945 28713 15979 28747
rect 19073 28713 19107 28747
rect 19257 28713 19291 28747
rect 19993 28713 20027 28747
rect 6193 28645 6227 28679
rect 7757 28645 7791 28679
rect 14749 28645 14783 28679
rect 2329 28577 2363 28611
rect 2605 28577 2639 28611
rect 3985 28577 4019 28611
rect 14289 28577 14323 28611
rect 15025 28577 15059 28611
rect 15301 28577 15335 28611
rect 20177 28577 20211 28611
rect 1501 28509 1535 28543
rect 3249 28509 3283 28543
rect 4259 28509 4293 28543
rect 5549 28509 5583 28543
rect 5733 28509 5767 28543
rect 6469 28509 6503 28543
rect 6586 28509 6620 28543
rect 6745 28509 6779 28543
rect 7389 28509 7423 28543
rect 7941 28509 7975 28543
rect 8033 28509 8067 28543
rect 9689 28509 9723 28543
rect 10149 28509 10183 28543
rect 11529 28509 11563 28543
rect 11803 28509 11837 28543
rect 14105 28509 14139 28543
rect 15163 28509 15197 28543
rect 16037 28509 16071 28543
rect 17693 28509 17727 28543
rect 17949 28509 17983 28543
rect 19441 28509 19475 28543
rect 19809 28509 19843 28543
rect 19901 28509 19935 28543
rect 20269 28509 20303 28543
rect 1685 28441 1719 28475
rect 9781 28441 9815 28475
rect 16293 28441 16327 28475
rect 3433 28373 3467 28407
rect 4997 28373 5031 28407
rect 9413 28373 9447 28407
rect 10517 28373 10551 28407
rect 10701 28373 10735 28407
rect 12541 28373 12575 28407
rect 17417 28373 17451 28407
rect 19625 28373 19659 28407
rect 20177 28373 20211 28407
rect 20453 28373 20487 28407
rect 9965 28169 9999 28203
rect 16313 28169 16347 28203
rect 19533 28169 19567 28203
rect 2881 28101 2915 28135
rect 20177 28101 20211 28135
rect 1651 28033 1685 28067
rect 3431 28033 3465 28067
rect 4811 28033 4845 28067
rect 9227 28033 9261 28067
rect 12725 28033 12759 28067
rect 14289 28033 14323 28067
rect 15326 28033 15360 28067
rect 16129 28033 16163 28067
rect 16497 28033 16531 28067
rect 16955 28033 16989 28067
rect 18061 28033 18095 28067
rect 18779 28063 18813 28097
rect 1409 27965 1443 27999
rect 3157 27965 3191 27999
rect 4537 27965 4571 27999
rect 8953 27965 8987 27999
rect 11529 27965 11563 27999
rect 11713 27965 11747 27999
rect 12173 27965 12207 27999
rect 12449 27965 12483 27999
rect 12587 27965 12621 27999
rect 14473 27965 14507 27999
rect 14933 27965 14967 27999
rect 15209 27965 15243 27999
rect 15485 27965 15519 27999
rect 16681 27965 16715 27999
rect 18521 27965 18555 27999
rect 3065 27897 3099 27931
rect 5549 27897 5583 27931
rect 13369 27897 13403 27931
rect 2421 27829 2455 27863
rect 4169 27829 4203 27863
rect 17693 27829 17727 27863
rect 18153 27829 18187 27863
rect 20453 27829 20487 27863
rect 3157 27625 3191 27659
rect 7849 27625 7883 27659
rect 16497 27625 16531 27659
rect 13921 27557 13955 27591
rect 17325 27557 17359 27591
rect 18153 27557 18187 27591
rect 18613 27557 18647 27591
rect 19257 27557 19291 27591
rect 14105 27489 14139 27523
rect 15485 27489 15519 27523
rect 17509 27489 17543 27523
rect 17693 27489 17727 27523
rect 19901 27489 19935 27523
rect 1409 27421 1443 27455
rect 3801 27421 3835 27455
rect 4077 27421 4111 27455
rect 4905 27421 4939 27455
rect 6837 27421 6871 27455
rect 7111 27421 7145 27455
rect 8401 27421 8435 27455
rect 8953 27421 8987 27455
rect 9227 27421 9261 27455
rect 14347 27421 14381 27455
rect 15727 27421 15761 27455
rect 16957 27421 16991 27455
rect 17233 27421 17267 27455
rect 17601 27421 17635 27455
rect 17785 27421 17819 27455
rect 18061 27421 18095 27455
rect 18337 27421 18371 27455
rect 18797 27421 18831 27455
rect 19073 27421 19107 27455
rect 19441 27421 19475 27455
rect 20177 27421 20211 27455
rect 2145 27353 2179 27387
rect 2237 27353 2271 27387
rect 2605 27353 2639 27387
rect 4813 27353 4847 27387
rect 5273 27353 5307 27387
rect 19625 27353 19659 27387
rect 20545 27353 20579 27387
rect 1593 27285 1627 27319
rect 1869 27285 1903 27319
rect 2973 27285 3007 27319
rect 3985 27285 4019 27319
rect 4261 27285 4295 27319
rect 4537 27285 4571 27319
rect 5641 27285 5675 27319
rect 5825 27285 5859 27319
rect 9965 27285 9999 27319
rect 15117 27285 15151 27319
rect 17049 27285 17083 27319
rect 17509 27285 17543 27319
rect 17877 27285 17911 27319
rect 18889 27285 18923 27319
rect 2605 27081 2639 27115
rect 3433 27081 3467 27115
rect 16681 27081 16715 27115
rect 18889 27081 18923 27115
rect 19165 27081 19199 27115
rect 4077 27013 4111 27047
rect 4445 27013 4479 27047
rect 7205 27013 7239 27047
rect 8309 27013 8343 27047
rect 14841 27013 14875 27047
rect 20177 27013 20211 27047
rect 1867 26945 1901 26979
rect 2973 26945 3007 26979
rect 3249 26945 3283 26979
rect 3525 26945 3559 26979
rect 4353 26945 4387 26979
rect 4813 26945 4847 26979
rect 5195 26945 5229 26979
rect 7481 26945 7515 26979
rect 7573 26945 7607 26979
rect 7941 26945 7975 26979
rect 10331 26945 10365 26979
rect 11529 26945 11563 26979
rect 11787 26975 11821 27009
rect 13001 26945 13035 26979
rect 13185 26945 13219 26979
rect 13921 26945 13955 26979
rect 14197 26945 14231 26979
rect 15117 26945 15151 26979
rect 15384 26945 15418 26979
rect 16865 26945 16899 26979
rect 17199 26945 17233 26979
rect 18337 26945 18371 26979
rect 18429 26945 18463 26979
rect 19073 26945 19107 26979
rect 19349 26945 19383 26979
rect 19625 26945 19659 26979
rect 1593 26877 1627 26911
rect 10057 26877 10091 26911
rect 14059 26877 14093 26911
rect 16957 26877 16991 26911
rect 18613 26877 18647 26911
rect 3157 26809 3191 26843
rect 5365 26809 5399 26843
rect 13645 26809 13679 26843
rect 3709 26741 3743 26775
rect 8493 26741 8527 26775
rect 11069 26741 11103 26775
rect 12541 26741 12575 26775
rect 16497 26741 16531 26775
rect 17969 26741 18003 26775
rect 18521 26741 18555 26775
rect 19901 26741 19935 26775
rect 20453 26741 20487 26775
rect 3433 26537 3467 26571
rect 5549 26537 5583 26571
rect 8217 26537 8251 26571
rect 13645 26537 13679 26571
rect 18705 26537 18739 26571
rect 3065 26469 3099 26503
rect 3341 26469 3375 26503
rect 11989 26469 12023 26503
rect 18337 26469 18371 26503
rect 18889 26469 18923 26503
rect 7205 26401 7239 26435
rect 19533 26401 19567 26435
rect 20361 26401 20395 26435
rect 20545 26401 20579 26435
rect 1501 26333 1535 26367
rect 1775 26333 1809 26367
rect 2881 26333 2915 26367
rect 3157 26333 3191 26367
rect 3617 26333 3651 26367
rect 4537 26333 4571 26367
rect 4811 26333 4845 26367
rect 7479 26333 7513 26367
rect 9137 26333 9171 26367
rect 9379 26333 9413 26367
rect 10977 26333 11011 26367
rect 12633 26333 12667 26367
rect 12907 26333 12941 26367
rect 15117 26333 15151 26367
rect 16773 26333 16807 26367
rect 16957 26333 16991 26367
rect 17509 26333 17543 26367
rect 17693 26333 17727 26367
rect 17877 26333 17911 26367
rect 18521 26333 18555 26367
rect 18613 26333 18647 26367
rect 18797 26333 18831 26367
rect 19073 26333 19107 26367
rect 19441 26333 19475 26367
rect 19791 26333 19825 26367
rect 20269 26333 20303 26367
rect 10701 26265 10735 26299
rect 11069 26265 11103 26299
rect 11437 26265 11471 26299
rect 15362 26265 15396 26299
rect 16865 26265 16899 26299
rect 20177 26265 20211 26299
rect 2513 26197 2547 26231
rect 10149 26197 10183 26231
rect 11805 26197 11839 26231
rect 16497 26197 16531 26231
rect 17325 26197 17359 26231
rect 17877 26197 17911 26231
rect 20545 26197 20579 26231
rect 1593 25993 1627 26027
rect 1869 25993 1903 26027
rect 8493 25993 8527 26027
rect 9413 25993 9447 26027
rect 15669 25993 15703 26027
rect 16497 25993 16531 26027
rect 17693 25993 17727 26027
rect 18153 25993 18187 26027
rect 19809 25993 19843 26027
rect 2145 25925 2179 25959
rect 2237 25925 2271 25959
rect 2973 25925 3007 25959
rect 9781 25925 9815 25959
rect 10149 25925 10183 25959
rect 13553 25925 13587 25959
rect 1409 25857 1443 25891
rect 2605 25857 2639 25891
rect 3525 25857 3559 25891
rect 3799 25857 3833 25891
rect 5179 25857 5213 25891
rect 6837 25857 6871 25891
rect 6929 25857 6963 25891
rect 7205 25857 7239 25891
rect 7389 25857 7423 25891
rect 7723 25857 7757 25891
rect 9689 25857 9723 25891
rect 10531 25857 10565 25891
rect 11955 25857 11989 25891
rect 13277 25857 13311 25891
rect 13645 25857 13679 25891
rect 13995 25887 14029 25921
rect 15853 25857 15887 25891
rect 15945 25857 15979 25891
rect 16221 25857 16255 25891
rect 16923 25867 16957 25901
rect 18337 25857 18371 25891
rect 18696 25857 18730 25891
rect 20177 25857 20211 25891
rect 4905 25789 4939 25823
rect 7481 25789 7515 25823
rect 11713 25789 11747 25823
rect 13093 25789 13127 25823
rect 13737 25789 13771 25823
rect 16497 25789 16531 25823
rect 16681 25789 16715 25823
rect 18429 25789 18463 25823
rect 6653 25721 6687 25755
rect 12725 25721 12759 25755
rect 3157 25653 3191 25687
rect 4537 25653 4571 25687
rect 5917 25653 5951 25687
rect 7021 25653 7055 25687
rect 7297 25653 7331 25687
rect 10701 25653 10735 25687
rect 14749 25653 14783 25687
rect 16037 25653 16071 25687
rect 16313 25653 16347 25687
rect 20453 25653 20487 25687
rect 2789 25449 2823 25483
rect 12173 25449 12207 25483
rect 12449 25449 12483 25483
rect 16865 25449 16899 25483
rect 20269 25449 20303 25483
rect 6285 25313 6319 25347
rect 6561 25313 6595 25347
rect 7757 25313 7791 25347
rect 15485 25313 15519 25347
rect 1409 25245 1443 25279
rect 1777 25245 1811 25279
rect 2051 25245 2085 25279
rect 3341 25245 3375 25279
rect 4721 25245 4755 25279
rect 5641 25245 5675 25279
rect 5825 25245 5859 25279
rect 6699 25245 6733 25279
rect 6837 25245 6871 25279
rect 8033 25245 8067 25279
rect 8493 25245 8527 25279
rect 8953 25245 8987 25279
rect 9211 25215 9245 25249
rect 12081 25245 12115 25279
rect 12265 25245 12299 25279
rect 12357 25245 12391 25279
rect 12633 25245 12667 25279
rect 12907 25245 12941 25279
rect 14105 25245 14139 25279
rect 14347 25235 14381 25269
rect 15743 25215 15777 25249
rect 17049 25245 17083 25279
rect 18981 25245 19015 25279
rect 19257 25245 19291 25279
rect 19531 25245 19565 25279
rect 4261 25177 4295 25211
rect 4353 25177 4387 25211
rect 8769 25177 8803 25211
rect 1593 25109 1627 25143
rect 3157 25109 3191 25143
rect 3985 25109 4019 25143
rect 5089 25109 5123 25143
rect 5273 25109 5307 25143
rect 7481 25109 7515 25143
rect 9965 25109 9999 25143
rect 13645 25109 13679 25143
rect 15117 25109 15151 25143
rect 16497 25109 16531 25143
rect 18797 25109 18831 25143
rect 3985 24905 4019 24939
rect 4537 24905 4571 24939
rect 5641 24905 5675 24939
rect 7389 24905 7423 24939
rect 7941 24905 7975 24939
rect 9229 24905 9263 24939
rect 13461 24905 13495 24939
rect 18490 24837 18524 24871
rect 2329 24769 2363 24803
rect 2605 24769 2639 24803
rect 3215 24769 3249 24803
rect 4813 24769 4847 24803
rect 4905 24769 4939 24803
rect 5273 24769 5307 24803
rect 6651 24769 6685 24803
rect 8125 24769 8159 24803
rect 8217 24769 8251 24803
rect 8491 24769 8525 24803
rect 9839 24769 9873 24803
rect 12047 24769 12081 24803
rect 13369 24769 13403 24803
rect 13645 24769 13679 24803
rect 13737 24769 13771 24803
rect 14795 24769 14829 24803
rect 17107 24769 17141 24803
rect 19993 24769 20027 24803
rect 1409 24701 1443 24735
rect 2973 24701 3007 24735
rect 6377 24701 6411 24735
rect 9597 24701 9631 24735
rect 11805 24701 11839 24735
rect 13921 24701 13955 24735
rect 14657 24701 14691 24735
rect 14933 24701 14967 24735
rect 16865 24701 16899 24735
rect 18245 24701 18279 24735
rect 2513 24633 2547 24667
rect 13185 24633 13219 24667
rect 14381 24633 14415 24667
rect 1639 24565 1673 24599
rect 2789 24565 2823 24599
rect 5825 24565 5859 24599
rect 10609 24565 10643 24599
rect 12817 24565 12851 24599
rect 15577 24565 15611 24599
rect 17877 24565 17911 24599
rect 19625 24565 19659 24599
rect 20269 24565 20303 24599
rect 4813 24361 4847 24395
rect 7113 24361 7147 24395
rect 10793 24361 10827 24395
rect 13277 24361 13311 24395
rect 18061 24361 18095 24395
rect 18889 24361 18923 24395
rect 5917 24293 5951 24327
rect 17969 24293 18003 24327
rect 18337 24293 18371 24327
rect 18521 24293 18555 24327
rect 1501 24225 1535 24259
rect 3801 24225 3835 24259
rect 5273 24225 5307 24259
rect 6310 24225 6344 24259
rect 6469 24225 6503 24259
rect 11437 24225 11471 24259
rect 12081 24225 12115 24259
rect 12474 24225 12508 24259
rect 12633 24225 12667 24259
rect 16405 24225 16439 24259
rect 18153 24225 18187 24259
rect 19257 24225 19291 24259
rect 1775 24157 1809 24191
rect 2881 24157 2915 24191
rect 4075 24157 4109 24191
rect 5457 24157 5491 24191
rect 6193 24157 6227 24191
rect 7205 24157 7239 24191
rect 7479 24157 7513 24191
rect 9781 24157 9815 24191
rect 9873 24157 9907 24191
rect 11621 24157 11655 24191
rect 12357 24157 12391 24191
rect 14565 24157 14599 24191
rect 14657 24157 14691 24191
rect 16313 24157 16347 24191
rect 16661 24157 16695 24191
rect 17877 24157 17911 24191
rect 18245 24157 18279 24191
rect 18705 24157 18739 24191
rect 18797 24157 18831 24191
rect 18981 24157 19015 24191
rect 19515 24127 19549 24161
rect 10241 24089 10275 24123
rect 10609 24089 10643 24123
rect 15025 24089 15059 24123
rect 2513 24021 2547 24055
rect 3065 24021 3099 24055
rect 8217 24021 8251 24055
rect 9505 24021 9539 24055
rect 14289 24021 14323 24055
rect 15393 24021 15427 24055
rect 15577 24021 15611 24055
rect 16129 24021 16163 24055
rect 17785 24021 17819 24055
rect 20269 24021 20303 24055
rect 1593 23817 1627 23851
rect 3249 23817 3283 23851
rect 9505 23817 9539 23851
rect 13369 23817 13403 23851
rect 2145 23749 2179 23783
rect 2421 23749 2455 23783
rect 9777 23749 9811 23783
rect 9873 23749 9907 23783
rect 10241 23749 10275 23783
rect 10609 23749 10643 23783
rect 19993 23749 20027 23783
rect 20177 23749 20211 23783
rect 1409 23681 1443 23715
rect 1685 23681 1719 23715
rect 2513 23681 2547 23715
rect 2881 23681 2915 23715
rect 4905 23681 4939 23715
rect 5179 23681 5213 23715
rect 6377 23681 6411 23715
rect 7573 23681 7607 23715
rect 11529 23681 11563 23715
rect 14197 23681 14231 23715
rect 14471 23681 14505 23715
rect 16681 23681 16715 23715
rect 16955 23691 16989 23725
rect 19257 23681 19291 23715
rect 19349 23681 19383 23715
rect 19717 23681 19751 23715
rect 6561 23613 6595 23647
rect 7297 23613 7331 23647
rect 7435 23613 7469 23647
rect 11713 23613 11747 23647
rect 12449 23613 12483 23647
rect 12566 23613 12600 23647
rect 12735 23613 12769 23647
rect 19993 23613 20027 23647
rect 1869 23545 1903 23579
rect 3433 23545 3467 23579
rect 5917 23545 5951 23579
rect 7021 23545 7055 23579
rect 12173 23545 12207 23579
rect 8217 23477 8251 23511
rect 10793 23477 10827 23511
rect 15209 23477 15243 23511
rect 17693 23477 17727 23511
rect 19073 23477 19107 23511
rect 19441 23477 19475 23511
rect 19809 23477 19843 23511
rect 20453 23477 20487 23511
rect 1869 23273 1903 23307
rect 2973 23273 3007 23307
rect 10609 23273 10643 23307
rect 12265 23273 12299 23307
rect 18613 23273 18647 23307
rect 1593 23205 1627 23239
rect 7113 23205 7147 23239
rect 15123 23205 15157 23239
rect 3801 23137 3835 23171
rect 6469 23137 6503 23171
rect 7389 23137 7423 23171
rect 7506 23137 7540 23171
rect 7665 23137 7699 23171
rect 14657 23137 14691 23171
rect 15393 23137 15427 23171
rect 19441 23137 19475 23171
rect 19809 23137 19843 23171
rect 19993 23137 20027 23171
rect 1409 23069 1443 23103
rect 1685 23069 1719 23103
rect 1961 23069 1995 23103
rect 2219 23039 2253 23073
rect 4075 23069 4109 23103
rect 6653 23069 6687 23103
rect 8585 23069 8619 23103
rect 9137 23085 9171 23119
rect 9597 23069 9631 23103
rect 9855 23039 9889 23073
rect 11253 23069 11287 23103
rect 11527 23069 11561 23103
rect 14473 23069 14507 23103
rect 15510 23069 15544 23103
rect 15669 23069 15703 23103
rect 18521 23069 18555 23103
rect 18705 23069 18739 23103
rect 18981 23069 19015 23103
rect 19349 23069 19383 23103
rect 19717 23069 19751 23103
rect 8309 23001 8343 23035
rect 16313 23001 16347 23035
rect 20177 23001 20211 23035
rect 20545 23001 20579 23035
rect 4813 22933 4847 22967
rect 8401 22933 8435 22967
rect 8953 22933 8987 22967
rect 18797 22933 18831 22967
rect 19993 22933 20027 22967
rect 2053 22729 2087 22763
rect 3341 22729 3375 22763
rect 3709 22729 3743 22763
rect 4997 22729 5031 22763
rect 2329 22661 2363 22695
rect 3157 22661 3191 22695
rect 4445 22661 4479 22695
rect 4813 22661 4847 22695
rect 18245 22661 18279 22695
rect 18696 22661 18730 22695
rect 20177 22661 20211 22695
rect 1409 22593 1443 22627
rect 2421 22593 2455 22627
rect 2789 22593 2823 22627
rect 3985 22593 4019 22627
rect 4077 22593 4111 22627
rect 8307 22593 8341 22627
rect 9597 22593 9631 22627
rect 9965 22593 9999 22627
rect 10331 22593 10365 22627
rect 11787 22623 11821 22657
rect 14473 22593 14507 22627
rect 16313 22593 16347 22627
rect 16681 22593 16715 22627
rect 16955 22593 16989 22627
rect 18153 22593 18187 22627
rect 18337 22593 18371 22627
rect 5181 22525 5215 22559
rect 5457 22525 5491 22559
rect 8033 22525 8067 22559
rect 9413 22525 9447 22559
rect 10057 22525 10091 22559
rect 11529 22525 11563 22559
rect 14657 22525 14691 22559
rect 15393 22525 15427 22559
rect 15531 22525 15565 22559
rect 15669 22525 15703 22559
rect 18429 22525 18463 22559
rect 9045 22457 9079 22491
rect 12541 22457 12575 22491
rect 15117 22457 15151 22491
rect 1593 22389 1627 22423
rect 6561 22389 6595 22423
rect 9873 22389 9907 22423
rect 11069 22389 11103 22423
rect 17693 22389 17727 22423
rect 19809 22389 19843 22423
rect 20453 22389 20487 22423
rect 1869 22185 1903 22219
rect 4445 22185 4479 22219
rect 9045 22185 9079 22219
rect 15393 22185 15427 22219
rect 18889 22185 18923 22219
rect 20269 22185 20303 22219
rect 6009 22117 6043 22151
rect 11621 22117 11655 22151
rect 13369 22117 13403 22151
rect 18153 22117 18187 22151
rect 6745 22049 6779 22083
rect 19257 22049 19291 22083
rect 1685 21981 1719 22015
rect 2053 21981 2087 22015
rect 2327 21981 2361 22015
rect 3433 21981 3467 22015
rect 4997 21981 5031 22015
rect 5089 21981 5123 22015
rect 6377 21981 6411 22015
rect 7019 21981 7053 22015
rect 8953 21981 8987 22015
rect 9229 21981 9263 22015
rect 9413 21981 9447 22015
rect 10609 21981 10643 22015
rect 10701 21981 10735 22015
rect 11451 21981 11485 22015
rect 12357 21981 12391 22015
rect 12631 21981 12665 22015
rect 14381 21981 14415 22015
rect 14655 21981 14689 22015
rect 16681 21981 16715 22015
rect 16773 21981 16807 22015
rect 18245 21981 18279 22015
rect 18705 21981 18739 22015
rect 19073 21981 19107 22015
rect 19531 21981 19565 22015
rect 5457 21913 5491 21947
rect 9321 21913 9355 21947
rect 10333 21913 10367 21947
rect 11069 21913 11103 21947
rect 17018 21913 17052 21947
rect 3065 21845 3099 21879
rect 3617 21845 3651 21879
rect 4721 21845 4755 21879
rect 5825 21845 5859 21879
rect 7757 21845 7791 21879
rect 16497 21845 16531 21879
rect 18337 21845 18371 21879
rect 18521 21845 18555 21879
rect 2513 21641 2547 21675
rect 4077 21641 4111 21675
rect 5641 21641 5675 21675
rect 8033 21641 8067 21675
rect 9137 21641 9171 21675
rect 20453 21641 20487 21675
rect 8309 21573 8343 21607
rect 8401 21573 8435 21607
rect 20177 21573 20211 21607
rect 1501 21505 1535 21539
rect 1775 21505 1809 21539
rect 3065 21505 3099 21539
rect 3339 21505 3373 21539
rect 4629 21505 4663 21539
rect 4903 21505 4937 21539
rect 6635 21535 6669 21569
rect 8769 21505 8803 21539
rect 10299 21505 10333 21539
rect 12081 21505 12115 21539
rect 13118 21505 13152 21539
rect 13277 21505 13311 21539
rect 14013 21505 14047 21539
rect 14197 21505 14231 21539
rect 15050 21505 15084 21539
rect 15853 21505 15887 21539
rect 16129 21505 16163 21539
rect 17567 21505 17601 21539
rect 18705 21505 18739 21539
rect 18797 21505 18831 21539
rect 19073 21505 19107 21539
rect 19257 21505 19291 21539
rect 19533 21505 19567 21539
rect 19717 21505 19751 21539
rect 6377 21437 6411 21471
rect 10057 21437 10091 21471
rect 12265 21437 12299 21471
rect 13001 21437 13035 21471
rect 14933 21437 14967 21471
rect 15209 21437 15243 21471
rect 17325 21437 17359 21471
rect 18981 21437 19015 21471
rect 19165 21437 19199 21471
rect 9321 21369 9355 21403
rect 11069 21369 11103 21403
rect 12725 21369 12759 21403
rect 14657 21369 14691 21403
rect 18337 21369 18371 21403
rect 7389 21301 7423 21335
rect 11989 21301 12023 21335
rect 13921 21301 13955 21335
rect 15945 21301 15979 21335
rect 18889 21301 18923 21335
rect 19349 21301 19383 21335
rect 19901 21301 19935 21335
rect 8493 21097 8527 21131
rect 9965 21097 9999 21131
rect 13185 21097 13219 21131
rect 3157 21029 3191 21063
rect 4813 21029 4847 21063
rect 10885 20961 10919 20995
rect 11529 20961 11563 20995
rect 11922 20961 11956 20995
rect 14289 20961 14323 20995
rect 14749 20961 14783 20995
rect 15142 20961 15176 20995
rect 1593 20893 1627 20927
rect 2145 20893 2179 20927
rect 3341 20893 3375 20927
rect 3801 20893 3835 20927
rect 4043 20893 4077 20927
rect 6009 20893 6043 20927
rect 6101 20893 6135 20927
rect 7481 20893 7515 20927
rect 7755 20893 7789 20927
rect 8953 20893 8987 20927
rect 9227 20893 9261 20927
rect 11069 20893 11103 20927
rect 11823 20893 11857 20927
rect 12081 20893 12115 20927
rect 12725 20893 12759 20927
rect 14105 20893 14139 20927
rect 15025 20893 15059 20927
rect 15301 20893 15335 20927
rect 16221 20893 16255 20927
rect 16405 20893 16439 20927
rect 16681 20893 16715 20927
rect 18613 20893 18647 20927
rect 18889 20893 18923 20927
rect 19073 20893 19107 20927
rect 19441 20893 19475 20927
rect 19993 20893 20027 20927
rect 1869 20825 1903 20859
rect 2237 20825 2271 20859
rect 2605 20825 2639 20859
rect 2973 20825 3007 20859
rect 6469 20825 6503 20859
rect 16497 20825 16531 20859
rect 16589 20825 16623 20859
rect 18705 20825 18739 20859
rect 19809 20825 19843 20859
rect 3525 20757 3559 20791
rect 5733 20757 5767 20791
rect 6837 20757 6871 20791
rect 7021 20757 7055 20791
rect 15945 20757 15979 20791
rect 16773 20757 16807 20791
rect 19073 20757 19107 20791
rect 20269 20757 20303 20791
rect 2605 20553 2639 20587
rect 12725 20553 12759 20587
rect 14289 20553 14323 20587
rect 15669 20553 15703 20587
rect 16497 20553 16531 20587
rect 18061 20553 18095 20587
rect 18880 20485 18914 20519
rect 1593 20417 1627 20451
rect 1867 20417 1901 20451
rect 3431 20417 3465 20451
rect 4537 20417 4571 20451
rect 4905 20417 4939 20451
rect 5179 20417 5213 20451
rect 7113 20417 7147 20451
rect 7387 20417 7421 20451
rect 9227 20417 9261 20451
rect 11971 20447 12005 20481
rect 13535 20447 13569 20481
rect 14931 20417 14965 20451
rect 16221 20417 16255 20451
rect 16313 20417 16347 20451
rect 16497 20417 16531 20451
rect 16937 20417 16971 20451
rect 20085 20417 20119 20451
rect 20177 20417 20211 20451
rect 3157 20349 3191 20383
rect 8953 20349 8987 20383
rect 11713 20349 11747 20383
rect 13277 20349 13311 20383
rect 14657 20349 14691 20383
rect 16681 20349 16715 20383
rect 18613 20349 18647 20383
rect 20361 20349 20395 20383
rect 5917 20281 5951 20315
rect 16037 20281 16071 20315
rect 4169 20213 4203 20247
rect 4721 20213 4755 20247
rect 8125 20213 8159 20247
rect 8861 20213 8895 20247
rect 9965 20213 9999 20247
rect 19993 20213 20027 20247
rect 20269 20213 20303 20247
rect 11621 20009 11655 20043
rect 16497 20009 16531 20043
rect 18889 20009 18923 20043
rect 20269 20009 20303 20043
rect 1409 19873 1443 19907
rect 1685 19873 1719 19907
rect 2329 19873 2363 19907
rect 5549 19873 5583 19907
rect 7481 19873 7515 19907
rect 9229 19873 9263 19907
rect 11989 19873 12023 19907
rect 15485 19873 15519 19907
rect 2603 19805 2637 19839
rect 4353 19805 4387 19839
rect 4445 19805 4479 19839
rect 5823 19805 5857 19839
rect 7723 19805 7757 19839
rect 9137 19805 9171 19839
rect 9503 19805 9537 19839
rect 10609 19805 10643 19839
rect 10883 19805 10917 19839
rect 12231 19805 12265 19839
rect 13553 19805 13587 19839
rect 13921 19805 13955 19839
rect 14105 19805 14139 19839
rect 14379 19805 14413 19839
rect 15727 19805 15761 19839
rect 17141 19805 17175 19839
rect 17509 19805 17543 19839
rect 18061 19805 18095 19839
rect 19073 19805 19107 19839
rect 19257 19805 19291 19839
rect 19499 19805 19533 19839
rect 4077 19737 4111 19771
rect 4813 19737 4847 19771
rect 3341 19669 3375 19703
rect 5181 19669 5215 19703
rect 5365 19669 5399 19703
rect 6561 19669 6595 19703
rect 8493 19669 8527 19703
rect 10241 19669 10275 19703
rect 13001 19669 13035 19703
rect 15117 19669 15151 19703
rect 16957 19669 16991 19703
rect 17601 19669 17635 19703
rect 17877 19669 17911 19703
rect 12173 19465 12207 19499
rect 17969 19465 18003 19499
rect 1501 19397 1535 19431
rect 3525 19397 3559 19431
rect 3801 19397 3835 19431
rect 4629 19397 4663 19431
rect 9781 19397 9815 19431
rect 10057 19397 10091 19431
rect 10149 19397 10183 19431
rect 10885 19397 10919 19431
rect 12449 19397 12483 19431
rect 13277 19397 13311 19431
rect 19809 19397 19843 19431
rect 20545 19397 20579 19431
rect 2235 19329 2269 19363
rect 3893 19329 3927 19363
rect 4261 19329 4295 19363
rect 7665 19329 7699 19363
rect 7849 19329 7883 19363
rect 8585 19329 8619 19363
rect 8702 19329 8736 19363
rect 8861 19329 8895 19363
rect 10517 19329 10551 19363
rect 12541 19329 12575 19363
rect 12909 19329 12943 19363
rect 13921 19329 13955 19363
rect 14105 19329 14139 19363
rect 14841 19329 14875 19363
rect 17231 19329 17265 19363
rect 18337 19329 18371 19363
rect 18705 19329 18739 19363
rect 18889 19329 18923 19363
rect 19625 19329 19659 19363
rect 20269 19329 20303 19363
rect 1961 19261 1995 19295
rect 8309 19261 8343 19295
rect 14565 19261 14599 19295
rect 14979 19261 15013 19295
rect 15117 19261 15151 19295
rect 16957 19261 16991 19295
rect 18429 19261 18463 19295
rect 18613 19261 18647 19295
rect 18797 19261 18831 19295
rect 20545 19261 20579 19295
rect 2973 19193 3007 19227
rect 4813 19193 4847 19227
rect 11069 19193 11103 19227
rect 15761 19193 15795 19227
rect 1593 19125 1627 19159
rect 9505 19125 9539 19159
rect 13461 19125 13495 19159
rect 16037 19125 16071 19159
rect 18521 19125 18555 19159
rect 19441 19125 19475 19159
rect 20085 19125 20119 19159
rect 20361 19125 20395 19159
rect 3157 18921 3191 18955
rect 3433 18921 3467 18955
rect 13277 18921 13311 18955
rect 17877 18921 17911 18955
rect 19349 18921 19383 18955
rect 5089 18853 5123 18887
rect 6101 18853 6135 18887
rect 20453 18853 20487 18887
rect 4077 18785 4111 18819
rect 5641 18785 5675 18819
rect 6377 18785 6411 18819
rect 12265 18785 12299 18819
rect 14933 18785 14967 18819
rect 15577 18785 15611 18819
rect 15970 18785 16004 18819
rect 16129 18785 16163 18819
rect 19901 18785 19935 18819
rect 1409 18717 1443 18751
rect 2329 18717 2363 18751
rect 2697 18717 2731 18751
rect 2973 18717 3007 18751
rect 3249 18717 3283 18751
rect 4319 18717 4353 18751
rect 5457 18717 5491 18751
rect 6515 18717 6549 18751
rect 6653 18717 6687 18751
rect 7481 18717 7515 18751
rect 7755 18717 7789 18751
rect 12539 18717 12573 18751
rect 15117 18717 15151 18751
rect 15853 18717 15887 18751
rect 16865 18717 16899 18751
rect 17107 18707 17141 18741
rect 19073 18717 19107 18751
rect 19257 18717 19291 18751
rect 19625 18717 19659 18751
rect 20177 18717 20211 18751
rect 1869 18649 1903 18683
rect 2053 18649 2087 18683
rect 10057 18649 10091 18683
rect 10333 18649 10367 18683
rect 10425 18649 10459 18683
rect 10793 18649 10827 18683
rect 1593 18581 1627 18615
rect 2513 18581 2547 18615
rect 2881 18581 2915 18615
rect 7297 18581 7331 18615
rect 8493 18581 8527 18615
rect 11161 18581 11195 18615
rect 11345 18581 11379 18615
rect 16773 18581 16807 18615
rect 18889 18581 18923 18615
rect 4813 18377 4847 18411
rect 9689 18377 9723 18411
rect 11069 18377 11103 18411
rect 15209 18377 15243 18411
rect 19809 18377 19843 18411
rect 1501 18309 1535 18343
rect 1685 18309 1719 18343
rect 3525 18309 3559 18343
rect 4629 18309 4663 18343
rect 18674 18309 18708 18343
rect 20177 18309 20211 18343
rect 2143 18241 2177 18275
rect 3801 18241 3835 18275
rect 3893 18241 3927 18275
rect 4261 18241 4295 18275
rect 7571 18241 7605 18275
rect 8677 18241 8711 18275
rect 8951 18241 8985 18275
rect 10299 18241 10333 18275
rect 11955 18241 11989 18275
rect 14439 18241 14473 18275
rect 18429 18241 18463 18275
rect 1869 18173 1903 18207
rect 7297 18173 7331 18207
rect 10057 18173 10091 18207
rect 11713 18173 11747 18207
rect 14197 18173 14231 18207
rect 2881 18105 2915 18139
rect 8309 18037 8343 18071
rect 12725 18037 12759 18071
rect 20453 18037 20487 18071
rect 1593 17833 1627 17867
rect 2697 17833 2731 17867
rect 3341 17833 3375 17867
rect 15761 17833 15795 17867
rect 20269 17833 20303 17867
rect 6193 17697 6227 17731
rect 6837 17697 6871 17731
rect 7230 17697 7264 17731
rect 12265 17697 12299 17731
rect 14749 17697 14783 17731
rect 1501 17629 1535 17663
rect 2053 17629 2087 17663
rect 3249 17629 3283 17663
rect 3525 17629 3559 17663
rect 4261 17629 4295 17663
rect 4721 17629 4755 17663
rect 6377 17629 6411 17663
rect 7113 17629 7147 17663
rect 7399 17629 7433 17663
rect 10425 17629 10459 17663
rect 12507 17629 12541 17663
rect 14991 17629 15025 17663
rect 16129 17629 16163 17663
rect 16403 17629 16437 17663
rect 18889 17629 18923 17663
rect 19073 17629 19107 17663
rect 19257 17629 19291 17663
rect 19499 17629 19533 17663
rect 2605 17561 2639 17595
rect 4353 17561 4387 17595
rect 5089 17561 5123 17595
rect 10149 17561 10183 17595
rect 10517 17561 10551 17595
rect 10885 17561 10919 17595
rect 18981 17561 19015 17595
rect 2145 17493 2179 17527
rect 3065 17493 3099 17527
rect 3985 17493 4019 17527
rect 5273 17493 5307 17527
rect 8033 17493 8067 17527
rect 11253 17493 11287 17527
rect 11437 17493 11471 17527
rect 13277 17493 13311 17527
rect 17141 17493 17175 17527
rect 1593 17289 1627 17323
rect 3065 17289 3099 17323
rect 4445 17289 4479 17323
rect 5917 17289 5951 17323
rect 7481 17289 7515 17323
rect 8861 17289 8895 17323
rect 9413 17289 9447 17323
rect 20453 17289 20487 17323
rect 10517 17221 10551 17255
rect 13737 17221 13771 17255
rect 20177 17221 20211 17255
rect 1501 17153 1535 17187
rect 2053 17153 2087 17187
rect 2311 17183 2345 17217
rect 3433 17153 3467 17187
rect 3707 17153 3741 17187
rect 5147 17153 5181 17187
rect 6711 17153 6745 17187
rect 8123 17153 8157 17187
rect 9689 17153 9723 17187
rect 9781 17153 9815 17187
rect 10149 17153 10183 17187
rect 11897 17153 11931 17187
rect 13093 17153 13127 17187
rect 14013 17153 14047 17187
rect 14866 17153 14900 17187
rect 16955 17153 16989 17187
rect 18501 17153 18535 17187
rect 19717 17153 19751 17187
rect 4905 17085 4939 17119
rect 6469 17085 6503 17119
rect 7849 17085 7883 17119
rect 12081 17085 12115 17119
rect 12817 17085 12851 17119
rect 12955 17085 12989 17119
rect 13829 17085 13863 17119
rect 14749 17085 14783 17119
rect 15025 17085 15059 17119
rect 16681 17085 16715 17119
rect 18245 17085 18279 17119
rect 12541 17017 12575 17051
rect 14473 17017 14507 17051
rect 10701 16949 10735 16983
rect 15669 16949 15703 16983
rect 17693 16949 17727 16983
rect 19625 16949 19659 16983
rect 19901 16949 19935 16983
rect 1777 16745 1811 16779
rect 3341 16745 3375 16779
rect 6745 16745 6779 16779
rect 3801 16677 3835 16711
rect 5365 16677 5399 16711
rect 8493 16677 8527 16711
rect 11253 16677 11287 16711
rect 13001 16677 13035 16711
rect 14841 16677 14875 16711
rect 16313 16677 16347 16711
rect 18797 16677 18831 16711
rect 2329 16609 2363 16643
rect 5733 16609 5767 16643
rect 14197 16609 14231 16643
rect 15234 16609 15268 16643
rect 16037 16609 16071 16643
rect 16405 16609 16439 16643
rect 19441 16609 19475 16643
rect 19809 16609 19843 16643
rect 19993 16609 20027 16643
rect 20453 16609 20487 16643
rect 2603 16541 2637 16575
rect 3985 16541 4019 16575
rect 4261 16541 4295 16575
rect 4353 16541 4387 16575
rect 4627 16541 4661 16575
rect 5975 16541 6009 16575
rect 7481 16541 7515 16575
rect 7755 16541 7789 16575
rect 10333 16541 10367 16575
rect 11989 16541 12023 16575
rect 12263 16531 12297 16565
rect 14381 16541 14415 16575
rect 15117 16541 15151 16575
rect 15403 16541 15437 16575
rect 16129 16541 16163 16575
rect 17877 16541 17911 16575
rect 18337 16541 18371 16575
rect 18429 16541 18463 16575
rect 18613 16541 18647 16575
rect 18981 16541 19015 16575
rect 19349 16541 19383 16575
rect 19717 16541 19751 16575
rect 1685 16473 1719 16507
rect 9965 16473 9999 16507
rect 10241 16473 10275 16507
rect 10701 16473 10735 16507
rect 16650 16473 16684 16507
rect 19993 16473 20027 16507
rect 20177 16473 20211 16507
rect 4077 16405 4111 16439
rect 11069 16405 11103 16439
rect 17785 16405 17819 16439
rect 17969 16405 18003 16439
rect 18153 16405 18187 16439
rect 18521 16405 18555 16439
rect 1593 16201 1627 16235
rect 2513 16201 2547 16235
rect 6101 16201 6135 16235
rect 13553 16201 13587 16235
rect 15945 16201 15979 16235
rect 19717 16201 19751 16235
rect 1501 16133 1535 16167
rect 2053 16065 2087 16099
rect 2697 16065 2731 16099
rect 3155 16075 3189 16109
rect 4261 16065 4295 16099
rect 5298 16065 5332 16099
rect 5457 16065 5491 16099
rect 7506 16065 7540 16099
rect 7665 16065 7699 16099
rect 8769 16065 8803 16099
rect 9806 16065 9840 16099
rect 12783 16065 12817 16099
rect 14105 16065 14139 16099
rect 15025 16065 15059 16099
rect 15301 16065 15335 16099
rect 17107 16065 17141 16099
rect 18245 16065 18279 16099
rect 18337 16065 18371 16099
rect 18947 16065 18981 16099
rect 20177 16065 20211 16099
rect 2881 15997 2915 16031
rect 4445 15997 4479 16031
rect 5181 15997 5215 16031
rect 6469 15997 6503 16031
rect 6653 15997 6687 16031
rect 7389 15997 7423 16031
rect 8953 15997 8987 16031
rect 9689 15997 9723 16031
rect 9965 15997 9999 16031
rect 10609 15997 10643 16031
rect 12541 15997 12575 16031
rect 14289 15997 14323 16031
rect 15142 15997 15176 16031
rect 16865 15997 16899 16031
rect 18521 15997 18555 16031
rect 18705 15997 18739 16031
rect 4905 15929 4939 15963
rect 7113 15929 7147 15963
rect 9413 15929 9447 15963
rect 14749 15929 14783 15963
rect 17877 15929 17911 15963
rect 2145 15861 2179 15895
rect 3893 15861 3927 15895
rect 8309 15861 8343 15895
rect 18429 15861 18463 15895
rect 20453 15861 20487 15895
rect 1501 15657 1535 15691
rect 3341 15657 3375 15691
rect 7113 15657 7147 15691
rect 8493 15657 8527 15691
rect 10057 15657 10091 15691
rect 11437 15657 11471 15691
rect 17049 15657 17083 15691
rect 19625 15657 19659 15691
rect 14749 15589 14783 15623
rect 18889 15589 18923 15623
rect 4721 15521 4755 15555
rect 9045 15521 9079 15555
rect 10425 15521 10459 15555
rect 14289 15521 14323 15555
rect 15025 15521 15059 15555
rect 15163 15521 15197 15555
rect 1685 15453 1719 15487
rect 1777 15453 1811 15487
rect 2051 15453 2085 15487
rect 3985 15453 4019 15487
rect 4261 15453 4295 15487
rect 4537 15453 4571 15487
rect 4995 15453 5029 15487
rect 6101 15453 6135 15487
rect 6375 15453 6409 15487
rect 7481 15453 7515 15487
rect 7755 15453 7789 15487
rect 9319 15453 9353 15487
rect 10699 15453 10733 15487
rect 11805 15453 11839 15487
rect 12079 15453 12113 15487
rect 14105 15453 14139 15487
rect 15301 15453 15335 15487
rect 16037 15453 16071 15487
rect 16311 15453 16345 15487
rect 18521 15453 18555 15487
rect 18705 15453 18739 15487
rect 19073 15453 19107 15487
rect 19257 15453 19291 15487
rect 19533 15453 19567 15487
rect 19717 15453 19751 15487
rect 19993 15453 20027 15487
rect 3249 15385 3283 15419
rect 15945 15385 15979 15419
rect 20177 15385 20211 15419
rect 20545 15385 20579 15419
rect 2789 15317 2823 15351
rect 3801 15317 3835 15351
rect 4077 15317 4111 15351
rect 4353 15317 4387 15351
rect 5733 15317 5767 15351
rect 12817 15317 12851 15351
rect 18705 15317 18739 15351
rect 19349 15317 19383 15351
rect 19809 15317 19843 15351
rect 1777 15113 1811 15147
rect 8217 15113 8251 15147
rect 15025 15113 15059 15147
rect 16405 15113 16439 15147
rect 16926 15045 16960 15079
rect 20177 15045 20211 15079
rect 1685 14977 1719 15011
rect 2145 14977 2179 15011
rect 2403 15007 2437 15041
rect 3799 14977 3833 15011
rect 4905 14977 4939 15011
rect 5179 14977 5213 15011
rect 7297 14977 7331 15011
rect 8919 14977 8953 15011
rect 10057 14977 10091 15011
rect 10331 14977 10365 15011
rect 12081 14977 12115 15011
rect 13001 14977 13035 15011
rect 14013 14977 14047 15011
rect 14287 14977 14321 15011
rect 16129 14977 16163 15011
rect 16313 14977 16347 15011
rect 16681 14977 16715 15011
rect 18153 14977 18187 15011
rect 18337 14977 18371 15011
rect 18685 14977 18719 15011
rect 3525 14909 3559 14943
rect 6377 14909 6411 14943
rect 6561 14909 6595 14943
rect 7021 14909 7055 14943
rect 7414 14909 7448 14943
rect 7573 14909 7607 14943
rect 8677 14909 8711 14943
rect 12265 14909 12299 14943
rect 13118 14909 13152 14943
rect 13277 14909 13311 14943
rect 18429 14909 18463 14943
rect 4537 14841 4571 14875
rect 11069 14841 11103 14875
rect 12725 14841 12759 14875
rect 3157 14773 3191 14807
rect 5917 14773 5951 14807
rect 9689 14773 9723 14807
rect 13921 14773 13955 14807
rect 15945 14773 15979 14807
rect 18061 14773 18095 14807
rect 18245 14773 18279 14807
rect 19809 14773 19843 14807
rect 20453 14773 20487 14807
rect 1593 14569 1627 14603
rect 3341 14569 3375 14603
rect 13093 14569 13127 14603
rect 15117 14569 15151 14603
rect 18889 14569 18923 14603
rect 4445 14501 4479 14535
rect 8493 14501 8527 14535
rect 2329 14433 2363 14467
rect 4721 14433 4755 14467
rect 4838 14433 4872 14467
rect 9965 14433 9999 14467
rect 10241 14433 10275 14467
rect 10358 14433 10392 14467
rect 14105 14433 14139 14467
rect 16865 14433 16899 14467
rect 18521 14433 18555 14467
rect 19257 14433 19291 14467
rect 2237 14365 2271 14399
rect 2603 14365 2637 14399
rect 3801 14365 3835 14399
rect 3985 14365 4019 14399
rect 4997 14365 5031 14399
rect 6101 14365 6135 14399
rect 6343 14365 6377 14399
rect 7481 14365 7515 14399
rect 7755 14365 7789 14399
rect 9321 14365 9355 14399
rect 9505 14365 9539 14399
rect 10517 14365 10551 14399
rect 12081 14365 12115 14399
rect 14379 14365 14413 14399
rect 15485 14365 15519 14399
rect 15759 14365 15793 14399
rect 17123 14335 17157 14369
rect 18245 14365 18279 14399
rect 18337 14365 18371 14399
rect 18613 14365 18647 14399
rect 19073 14365 19107 14399
rect 19515 14335 19549 14369
rect 1501 14297 1535 14331
rect 12173 14297 12207 14331
rect 12541 14297 12575 14331
rect 18705 14297 18739 14331
rect 2053 14229 2087 14263
rect 5641 14229 5675 14263
rect 7113 14229 7147 14263
rect 11161 14229 11195 14263
rect 11805 14229 11839 14263
rect 12909 14229 12943 14263
rect 16497 14229 16531 14263
rect 17877 14229 17911 14263
rect 18521 14229 18555 14263
rect 20269 14229 20303 14263
rect 1961 14025 1995 14059
rect 4261 14025 4295 14059
rect 13369 14025 13403 14059
rect 16313 14025 16347 14059
rect 20453 14025 20487 14059
rect 1685 13957 1719 13991
rect 19257 13957 19291 13991
rect 19993 13957 20027 13991
rect 3366 13889 3400 13923
rect 3525 13889 3559 13923
rect 4445 13889 4479 13923
rect 4721 13889 4755 13923
rect 5147 13889 5181 13923
rect 6561 13889 6595 13923
rect 7297 13889 7331 13923
rect 7414 13889 7448 13923
rect 10563 13889 10597 13923
rect 12631 13889 12665 13923
rect 14287 13889 14321 13923
rect 16221 13889 16255 13923
rect 16497 13889 16531 13923
rect 16681 13889 16715 13923
rect 16937 13889 16971 13923
rect 18337 13889 18371 13923
rect 18429 13889 18463 13923
rect 18613 13889 18647 13923
rect 18797 13889 18831 13923
rect 18981 13889 19015 13923
rect 19717 13889 19751 13923
rect 20177 13889 20211 13923
rect 2329 13821 2363 13855
rect 2513 13821 2547 13855
rect 2973 13821 3007 13855
rect 3249 13821 3283 13855
rect 4905 13821 4939 13855
rect 6377 13821 6411 13855
rect 7573 13821 7607 13855
rect 9505 13821 9539 13855
rect 9689 13821 9723 13855
rect 10425 13821 10459 13855
rect 10701 13821 10735 13855
rect 12357 13821 12391 13855
rect 14013 13821 14047 13855
rect 18889 13821 18923 13855
rect 19533 13821 19567 13855
rect 19993 13821 20027 13855
rect 5917 13753 5951 13787
rect 7021 13753 7055 13787
rect 10149 13753 10183 13787
rect 15025 13753 15059 13787
rect 16037 13753 16071 13787
rect 18061 13753 18095 13787
rect 19809 13753 19843 13787
rect 4169 13685 4203 13719
rect 4537 13685 4571 13719
rect 8217 13685 8251 13719
rect 11345 13685 11379 13719
rect 18153 13685 18187 13719
rect 18521 13685 18555 13719
rect 1593 13481 1627 13515
rect 3157 13481 3191 13515
rect 3985 13481 4019 13515
rect 13369 13481 13403 13515
rect 17049 13481 17083 13515
rect 18429 13481 18463 13515
rect 18889 13481 18923 13515
rect 5641 13413 5675 13447
rect 6653 13413 6687 13447
rect 14749 13413 14783 13447
rect 6009 13345 6043 13379
rect 7046 13345 7080 13379
rect 7205 13345 7239 13379
rect 9965 13345 9999 13379
rect 10425 13345 10459 13379
rect 14289 13345 14323 13379
rect 15142 13345 15176 13379
rect 15301 13345 15335 13379
rect 17417 13345 17451 13379
rect 19257 13345 19291 13379
rect 2145 13277 2179 13311
rect 2403 13247 2437 13281
rect 4537 13277 4571 13311
rect 4629 13277 4663 13311
rect 4903 13277 4937 13311
rect 6193 13277 6227 13311
rect 6929 13277 6963 13311
rect 9781 13277 9815 13311
rect 10701 13277 10735 13311
rect 10839 13277 10873 13311
rect 10977 13277 11011 13311
rect 12357 13277 12391 13311
rect 14105 13277 14139 13311
rect 15025 13277 15059 13311
rect 16037 13277 16071 13311
rect 16311 13277 16345 13311
rect 19073 13293 19107 13327
rect 17675 13247 17709 13281
rect 19499 13267 19533 13301
rect 1501 13209 1535 13243
rect 3893 13209 3927 13243
rect 12449 13209 12483 13243
rect 12817 13209 12851 13243
rect 15945 13209 15979 13243
rect 4353 13141 4387 13175
rect 7849 13141 7883 13175
rect 11621 13141 11655 13175
rect 12081 13141 12115 13175
rect 13185 13141 13219 13175
rect 20269 13141 20303 13175
rect 1593 12937 1627 12971
rect 6653 12937 6687 12971
rect 8309 12937 8343 12971
rect 9689 12937 9723 12971
rect 11069 12937 11103 12971
rect 16313 12937 16347 12971
rect 18889 12937 18923 12971
rect 20453 12937 20487 12971
rect 1961 12869 1995 12903
rect 2513 12869 2547 12903
rect 4629 12869 4663 12903
rect 12081 12869 12115 12903
rect 12357 12869 12391 12903
rect 12817 12869 12851 12903
rect 13185 12869 13219 12903
rect 1777 12801 1811 12835
rect 3247 12801 3281 12835
rect 5163 12831 5197 12865
rect 6561 12801 6595 12835
rect 6837 12801 6871 12835
rect 7571 12801 7605 12835
rect 8935 12831 8969 12865
rect 10299 12801 10333 12835
rect 12449 12801 12483 12835
rect 14473 12801 14507 12835
rect 15326 12801 15360 12835
rect 16497 12801 16531 12835
rect 16955 12801 16989 12835
rect 18061 12801 18095 12835
rect 18613 12801 18647 12835
rect 19073 12801 19107 12835
rect 19625 12801 19659 12835
rect 20177 12801 20211 12835
rect 2973 12733 3007 12767
rect 4905 12733 4939 12767
rect 7297 12733 7331 12767
rect 8677 12733 8711 12767
rect 10057 12733 10091 12767
rect 14289 12733 14323 12767
rect 15209 12733 15243 12767
rect 15485 12733 15519 12767
rect 16681 12733 16715 12767
rect 18337 12733 18371 12767
rect 18889 12733 18923 12767
rect 6377 12665 6411 12699
rect 13369 12665 13403 12699
rect 14933 12665 14967 12699
rect 16129 12665 16163 12699
rect 2053 12597 2087 12631
rect 2605 12597 2639 12631
rect 3985 12597 4019 12631
rect 5917 12597 5951 12631
rect 17693 12597 17727 12631
rect 18153 12597 18187 12631
rect 18245 12597 18279 12631
rect 18705 12597 18739 12631
rect 19349 12597 19383 12631
rect 19901 12597 19935 12631
rect 1777 12393 1811 12427
rect 4169 12393 4203 12427
rect 8493 12393 8527 12427
rect 13829 12393 13863 12427
rect 17141 12393 17175 12427
rect 18429 12393 18463 12427
rect 18981 12393 19015 12427
rect 3341 12325 3375 12359
rect 5273 12325 5307 12359
rect 13185 12325 13219 12359
rect 14841 12325 14875 12359
rect 2329 12257 2363 12291
rect 4629 12257 4663 12291
rect 5825 12257 5859 12291
rect 7481 12257 7515 12291
rect 9597 12257 9631 12291
rect 10057 12257 10091 12291
rect 10333 12257 10367 12291
rect 10450 12257 10484 12291
rect 15117 12257 15151 12291
rect 15255 12257 15289 12291
rect 15403 12257 15437 12291
rect 20361 12257 20395 12291
rect 1685 12189 1719 12223
rect 2587 12159 2621 12193
rect 4537 12189 4571 12223
rect 4813 12189 4847 12223
rect 5549 12189 5583 12223
rect 5687 12189 5721 12223
rect 6745 12189 6779 12223
rect 7021 12189 7055 12223
rect 7755 12189 7789 12223
rect 9413 12189 9447 12223
rect 10609 12189 10643 12223
rect 12173 12189 12207 12223
rect 13737 12189 13771 12223
rect 13921 12189 13955 12223
rect 14197 12189 14231 12223
rect 14381 12189 14415 12223
rect 16129 12189 16163 12223
rect 16403 12189 16437 12223
rect 17693 12189 17727 12223
rect 17877 12189 17911 12223
rect 18337 12189 18371 12223
rect 18705 12189 18739 12223
rect 19625 12189 19659 12223
rect 19809 12189 19843 12223
rect 20269 12189 20303 12223
rect 3893 12121 3927 12155
rect 12265 12121 12299 12155
rect 12633 12121 12667 12155
rect 4353 12053 4387 12087
rect 6469 12053 6503 12087
rect 6561 12053 6595 12087
rect 6837 12053 6871 12087
rect 11253 12053 11287 12087
rect 11897 12053 11931 12087
rect 13001 12053 13035 12087
rect 16037 12053 16071 12087
rect 17509 12053 17543 12087
rect 17969 12053 18003 12087
rect 1593 11849 1627 11883
rect 3065 11849 3099 11883
rect 5549 11849 5583 11883
rect 6101 11849 6135 11883
rect 9597 11849 9631 11883
rect 9781 11849 9815 11883
rect 10977 11849 11011 11883
rect 14749 11849 14783 11883
rect 16129 11849 16163 11883
rect 18521 11849 18555 11883
rect 19993 11849 20027 11883
rect 8493 11781 8527 11815
rect 8769 11781 8803 11815
rect 8861 11781 8895 11815
rect 18880 11781 18914 11815
rect 20177 11781 20211 11815
rect 1501 11713 1535 11747
rect 2295 11713 2329 11747
rect 3617 11713 3651 11747
rect 4491 11713 4525 11747
rect 4629 11713 4663 11747
rect 5457 11713 5491 11747
rect 6009 11713 6043 11747
rect 7414 11713 7448 11747
rect 9229 11713 9263 11747
rect 10239 11713 10273 11747
rect 12615 11713 12649 11747
rect 13737 11713 13771 11747
rect 14011 11713 14045 11747
rect 15359 11713 15393 11747
rect 16773 11713 16807 11747
rect 17029 11713 17063 11747
rect 18245 11713 18279 11747
rect 18337 11713 18371 11747
rect 18613 11713 18647 11747
rect 2053 11645 2087 11679
rect 3433 11645 3467 11679
rect 4353 11645 4387 11679
rect 6377 11645 6411 11679
rect 6561 11645 6595 11679
rect 7297 11645 7331 11679
rect 7573 11645 7607 11679
rect 9965 11645 9999 11679
rect 12357 11645 12391 11679
rect 15117 11645 15151 11679
rect 18521 11645 18555 11679
rect 4077 11577 4111 11611
rect 7021 11577 7055 11611
rect 5273 11509 5307 11543
rect 8217 11509 8251 11543
rect 13369 11509 13403 11543
rect 18153 11509 18187 11543
rect 20453 11509 20487 11543
rect 1685 11305 1719 11339
rect 3341 11305 3375 11339
rect 5641 11305 5675 11339
rect 6745 11305 6779 11339
rect 10793 11305 10827 11339
rect 13185 11305 13219 11339
rect 15117 11305 15151 11339
rect 17141 11305 17175 11339
rect 18337 11305 18371 11339
rect 18705 11305 18739 11339
rect 20269 11305 20303 11339
rect 2329 11169 2363 11203
rect 3985 11169 4019 11203
rect 4445 11169 4479 11203
rect 4721 11169 4755 11203
rect 4859 11169 4893 11203
rect 12173 11169 12207 11203
rect 19257 11169 19291 11203
rect 2237 11101 2271 11135
rect 2603 11101 2637 11135
rect 3801 11101 3835 11135
rect 4997 11101 5031 11135
rect 5733 11101 5767 11135
rect 6007 11101 6041 11135
rect 7481 11101 7515 11135
rect 7755 11101 7789 11135
rect 9689 11101 9723 11135
rect 9781 11101 9815 11135
rect 10055 11101 10089 11135
rect 12447 11101 12481 11135
rect 14105 11101 14139 11135
rect 14379 11101 14413 11135
rect 15485 11101 15519 11135
rect 15759 11101 15793 11135
rect 17325 11101 17359 11135
rect 17599 11101 17633 11135
rect 18889 11101 18923 11135
rect 19499 11101 19533 11135
rect 1593 11033 1627 11067
rect 17049 11033 17083 11067
rect 2053 10965 2087 10999
rect 8493 10965 8527 10999
rect 9505 10965 9539 10999
rect 16497 10965 16531 10999
rect 1593 10761 1627 10795
rect 3157 10761 3191 10795
rect 4537 10761 4571 10795
rect 5917 10761 5951 10795
rect 7757 10761 7791 10795
rect 9137 10761 9171 10795
rect 10517 10761 10551 10795
rect 12541 10761 12575 10795
rect 14841 10761 14875 10795
rect 1501 10625 1535 10659
rect 2145 10625 2179 10659
rect 2403 10655 2437 10689
rect 3767 10625 3801 10659
rect 5147 10625 5181 10659
rect 6987 10625 7021 10659
rect 8383 10655 8417 10689
rect 9747 10625 9781 10659
rect 11771 10625 11805 10659
rect 13001 10625 13035 10659
rect 13921 10625 13955 10659
rect 14038 10625 14072 10659
rect 14933 10625 14967 10659
rect 15207 10635 15241 10669
rect 16497 10625 16531 10659
rect 16939 10655 16973 10689
rect 18303 10625 18337 10659
rect 19809 10625 19843 10659
rect 20269 10625 20303 10659
rect 3525 10557 3559 10591
rect 4905 10557 4939 10591
rect 6745 10557 6779 10591
rect 8125 10557 8159 10591
rect 9505 10557 9539 10591
rect 11529 10557 11563 10591
rect 13185 10557 13219 10591
rect 13645 10557 13679 10591
rect 14197 10557 14231 10591
rect 16681 10557 16715 10591
rect 18061 10557 18095 10591
rect 19625 10557 19659 10591
rect 20269 10489 20303 10523
rect 15945 10421 15979 10455
rect 16313 10421 16347 10455
rect 17693 10421 17727 10455
rect 19073 10421 19107 10455
rect 1593 10217 1627 10251
rect 4169 10217 4203 10251
rect 7113 10217 7147 10251
rect 12541 10217 12575 10251
rect 17049 10217 17083 10251
rect 18797 10217 18831 10251
rect 20269 10217 20303 10251
rect 10241 10149 10275 10183
rect 14749 10149 14783 10183
rect 4721 10081 4755 10115
rect 6101 10081 6135 10115
rect 9597 10081 9631 10115
rect 10517 10081 10551 10115
rect 10634 10081 10668 10115
rect 11437 10081 11471 10115
rect 11529 10081 11563 10115
rect 14289 10081 14323 10115
rect 15025 10081 15059 10115
rect 15142 10081 15176 10115
rect 15301 10081 15335 10115
rect 17417 10081 17451 10115
rect 19257 10081 19291 10115
rect 1777 10013 1811 10047
rect 1869 10013 1903 10047
rect 2143 10013 2177 10047
rect 3617 10013 3651 10047
rect 4537 10013 4571 10047
rect 4963 10013 4997 10047
rect 6343 10013 6377 10047
rect 7481 10013 7515 10047
rect 7755 10013 7789 10047
rect 9781 10013 9815 10047
rect 10793 10013 10827 10047
rect 11803 10013 11837 10047
rect 14105 10013 14139 10047
rect 16037 10013 16071 10047
rect 16279 10013 16313 10047
rect 17659 10013 17693 10047
rect 18981 10013 19015 10047
rect 19499 10013 19533 10047
rect 3893 9945 3927 9979
rect 2881 9877 2915 9911
rect 3433 9877 3467 9911
rect 4353 9877 4387 9911
rect 5733 9877 5767 9911
rect 8493 9877 8527 9911
rect 15945 9877 15979 9911
rect 18429 9877 18463 9911
rect 1777 9673 1811 9707
rect 7757 9673 7791 9707
rect 15761 9673 15795 9707
rect 16405 9673 16439 9707
rect 19809 9673 19843 9707
rect 1501 9605 1535 9639
rect 20269 9605 20303 9639
rect 2329 9537 2363 9571
rect 2605 9537 2639 9571
rect 3479 9537 3513 9571
rect 4353 9537 4387 9571
rect 5291 9537 5325 9571
rect 6561 9537 6595 9571
rect 6745 9537 6779 9571
rect 6987 9537 7021 9571
rect 8125 9537 8159 9571
rect 8399 9537 8433 9571
rect 9505 9537 9539 9571
rect 10425 9537 10459 9571
rect 10563 9537 10597 9571
rect 11955 9537 11989 9571
rect 13829 9537 13863 9571
rect 14887 9537 14921 9571
rect 15945 9537 15979 9571
rect 16221 9537 16255 9571
rect 16313 9537 16347 9571
rect 16497 9537 16531 9571
rect 16937 9537 16971 9571
rect 18337 9537 18371 9571
rect 19039 9537 19073 9571
rect 20177 9537 20211 9571
rect 2421 9469 2455 9503
rect 3341 9469 3375 9503
rect 3617 9469 3651 9503
rect 4537 9469 4571 9503
rect 5411 9469 5445 9503
rect 5549 9469 5583 9503
rect 9689 9469 9723 9503
rect 10701 9469 10735 9503
rect 11713 9469 11747 9503
rect 14013 9469 14047 9503
rect 14749 9469 14783 9503
rect 15023 9469 15057 9503
rect 16681 9469 16715 9503
rect 18613 9469 18647 9503
rect 18797 9469 18831 9503
rect 3065 9401 3099 9435
rect 4997 9401 5031 9435
rect 10149 9401 10183 9435
rect 14473 9401 14507 9435
rect 2145 9333 2179 9367
rect 4261 9333 4295 9367
rect 6193 9333 6227 9367
rect 6377 9333 6411 9367
rect 9137 9333 9171 9367
rect 11345 9333 11379 9367
rect 12725 9333 12759 9367
rect 15669 9333 15703 9367
rect 16037 9333 16071 9367
rect 18061 9333 18095 9367
rect 1777 9129 1811 9163
rect 4169 9129 4203 9163
rect 4537 9129 4571 9163
rect 11897 9129 11931 9163
rect 15117 9129 15151 9163
rect 16497 9129 16531 9163
rect 16957 9129 16991 9163
rect 18981 9129 19015 9163
rect 5917 9061 5951 9095
rect 6929 9061 6963 9095
rect 12633 9061 12667 9095
rect 20269 9061 20303 9095
rect 4905 8993 4939 9027
rect 6469 8993 6503 9027
rect 7322 8993 7356 9027
rect 7481 8993 7515 9027
rect 10241 8993 10275 9027
rect 10701 8993 10735 9027
rect 11115 8993 11149 9027
rect 11989 8993 12023 9027
rect 12909 8993 12943 9027
rect 15485 8993 15519 9027
rect 19257 8993 19291 9027
rect 1685 8925 1719 8959
rect 2329 8925 2363 8959
rect 2603 8925 2637 8959
rect 3893 8925 3927 8959
rect 4445 8925 4479 8959
rect 5179 8925 5213 8959
rect 6285 8925 6319 8959
rect 7205 8925 7239 8959
rect 9965 8925 9999 8959
rect 10057 8925 10091 8959
rect 10977 8925 11011 8959
rect 11253 8925 11287 8959
rect 12173 8925 12207 8959
rect 13026 8925 13060 8959
rect 13185 8925 13219 8959
rect 14105 8925 14139 8959
rect 14379 8925 14413 8959
rect 15727 8925 15761 8959
rect 16865 8925 16899 8959
rect 17233 8925 17267 8959
rect 17507 8925 17541 8959
rect 19531 8925 19565 8959
rect 18705 8857 18739 8891
rect 3341 8789 3375 8823
rect 8125 8789 8159 8823
rect 9781 8789 9815 8823
rect 13829 8789 13863 8823
rect 18245 8789 18279 8823
rect 1777 8585 1811 8619
rect 5457 8585 5491 8619
rect 9229 8585 9263 8619
rect 10885 8585 10919 8619
rect 15209 8585 15243 8619
rect 16405 8585 16439 8619
rect 16865 8585 16899 8619
rect 17325 8585 17359 8619
rect 20545 8585 20579 8619
rect 2053 8517 2087 8551
rect 7941 8517 7975 8551
rect 8297 8517 8331 8551
rect 9045 8517 9079 8551
rect 19432 8517 19466 8551
rect 1501 8449 1535 8483
rect 2697 8449 2731 8483
rect 3433 8449 3467 8483
rect 3709 8449 3743 8483
rect 4445 8449 4479 8483
rect 4719 8449 4753 8483
rect 6009 8449 6043 8483
rect 6619 8449 6653 8483
rect 8217 8449 8251 8483
rect 8677 8449 8711 8483
rect 9781 8449 9815 8483
rect 10131 8479 10165 8513
rect 12507 8449 12541 8483
rect 13645 8449 13679 8483
rect 13919 8449 13953 8483
rect 15393 8449 15427 8483
rect 15669 8449 15703 8483
rect 15761 8449 15795 8483
rect 16221 8449 16255 8483
rect 16313 8449 16347 8483
rect 16681 8449 16715 8483
rect 16865 8449 16899 8483
rect 16957 8449 16991 8483
rect 17509 8449 17543 8483
rect 17785 8449 17819 8483
rect 18027 8449 18061 8483
rect 19165 8449 19199 8483
rect 2513 8381 2547 8415
rect 3157 8381 3191 8415
rect 3571 8381 3605 8415
rect 6377 8381 6411 8415
rect 9873 8381 9907 8415
rect 12265 8381 12299 8415
rect 17049 8381 17083 8415
rect 5825 8313 5859 8347
rect 7389 8313 7423 8347
rect 13277 8313 13311 8347
rect 18797 8313 18831 8347
rect 2145 8245 2179 8279
rect 4353 8245 4387 8279
rect 9597 8245 9631 8279
rect 14657 8245 14691 8279
rect 15485 8245 15519 8279
rect 15853 8245 15887 8279
rect 16037 8245 16071 8279
rect 1777 8041 1811 8075
rect 3341 8041 3375 8075
rect 5733 8041 5767 8075
rect 8493 8041 8527 8075
rect 11529 8041 11563 8075
rect 15117 8041 15151 8075
rect 15945 8041 15979 8075
rect 16221 8041 16255 8075
rect 12725 7973 12759 8007
rect 18889 7973 18923 8007
rect 20085 7973 20119 8007
rect 2329 7905 2363 7939
rect 4721 7905 4755 7939
rect 6101 7905 6135 7939
rect 7481 7905 7515 7939
rect 8953 7905 8987 7939
rect 10517 7905 10551 7939
rect 12081 7905 12115 7939
rect 13118 7905 13152 7939
rect 13277 7905 13311 7939
rect 14105 7905 14139 7939
rect 16497 7905 16531 7939
rect 19441 7905 19475 7939
rect 1501 7837 1535 7871
rect 2145 7837 2179 7871
rect 2603 7837 2637 7871
rect 4995 7837 5029 7871
rect 6375 7837 6409 7871
rect 7723 7837 7757 7871
rect 9227 7837 9261 7871
rect 10791 7827 10825 7861
rect 12265 7837 12299 7871
rect 13001 7837 13035 7871
rect 14379 7837 14413 7871
rect 15485 7837 15519 7871
rect 15669 7837 15703 7871
rect 16129 7837 16163 7871
rect 16405 7837 16439 7871
rect 16753 7837 16787 7871
rect 17969 7837 18003 7871
rect 18337 7837 18371 7871
rect 18797 7837 18831 7871
rect 19625 7837 19659 7871
rect 20085 7837 20119 7871
rect 3893 7769 3927 7803
rect 4261 7769 4295 7803
rect 1961 7701 1995 7735
rect 3985 7701 4019 7735
rect 4353 7701 4387 7735
rect 7113 7701 7147 7735
rect 9965 7701 9999 7735
rect 13921 7701 13955 7735
rect 15669 7701 15703 7735
rect 17877 7701 17911 7735
rect 1409 7497 1443 7531
rect 2697 7497 2731 7531
rect 3985 7497 4019 7531
rect 7665 7497 7699 7531
rect 10977 7497 11011 7531
rect 11529 7497 11563 7531
rect 16129 7497 16163 7531
rect 17693 7497 17727 7531
rect 19809 7497 19843 7531
rect 20453 7497 20487 7531
rect 3341 7429 3375 7463
rect 20177 7429 20211 7463
rect 1593 7361 1627 7395
rect 1959 7361 1993 7395
rect 3893 7361 3927 7395
rect 4353 7361 4387 7395
rect 5273 7361 5307 7395
rect 5549 7361 5583 7395
rect 6561 7361 6595 7395
rect 8033 7361 8067 7395
rect 9070 7361 9104 7395
rect 9229 7361 9263 7395
rect 10239 7361 10273 7395
rect 11713 7361 11747 7395
rect 11805 7361 11839 7395
rect 12725 7361 12759 7395
rect 12842 7361 12876 7395
rect 13001 7361 13035 7395
rect 13737 7361 13771 7395
rect 14363 7391 14397 7425
rect 15669 7361 15703 7395
rect 16037 7361 16071 7395
rect 16313 7361 16347 7395
rect 16955 7361 16989 7395
rect 18153 7361 18187 7395
rect 18409 7361 18443 7395
rect 19625 7361 19659 7395
rect 19809 7361 19843 7395
rect 1685 7293 1719 7327
rect 4537 7293 4571 7327
rect 5411 7293 5445 7327
rect 8217 7293 8251 7327
rect 8953 7293 8987 7327
rect 9965 7293 9999 7327
rect 11989 7293 12023 7327
rect 14105 7293 14139 7327
rect 15485 7293 15519 7327
rect 16681 7293 16715 7327
rect 4997 7225 5031 7259
rect 8677 7225 8711 7259
rect 12449 7225 12483 7259
rect 13921 7225 13955 7259
rect 15117 7225 15151 7259
rect 15669 7225 15703 7259
rect 3433 7157 3467 7191
rect 6193 7157 6227 7191
rect 6377 7157 6411 7191
rect 9873 7157 9907 7191
rect 13645 7157 13679 7191
rect 19533 7157 19567 7191
rect 1501 6953 1535 6987
rect 1961 6953 1995 6987
rect 3985 6953 4019 6987
rect 5641 6953 5675 6987
rect 11989 6953 12023 6987
rect 13093 6953 13127 6987
rect 13829 6953 13863 6987
rect 20085 6885 20119 6919
rect 2329 6817 2363 6851
rect 4629 6817 4663 6851
rect 6469 6817 6503 6851
rect 6929 6817 6963 6851
rect 7205 6817 7239 6851
rect 10333 6817 10367 6851
rect 10793 6817 10827 6851
rect 15669 6817 15703 6851
rect 17141 6817 17175 6851
rect 1685 6749 1719 6783
rect 1869 6749 1903 6783
rect 2571 6749 2605 6783
rect 4537 6749 4571 6783
rect 4903 6749 4937 6783
rect 6193 6749 6227 6783
rect 6285 6749 6319 6783
rect 7322 6749 7356 6783
rect 7481 6749 7515 6783
rect 9229 6749 9263 6783
rect 10149 6749 10183 6783
rect 11069 6749 11103 6783
rect 11186 6749 11220 6783
rect 11345 6749 11379 6783
rect 12081 6749 12115 6783
rect 12339 6749 12373 6783
rect 13461 6749 13495 6783
rect 13737 6749 13771 6783
rect 14289 6749 14323 6783
rect 14563 6749 14597 6783
rect 15925 6749 15959 6783
rect 17383 6749 17417 6783
rect 18521 6749 18555 6783
rect 18705 6749 18739 6783
rect 18797 6749 18831 6783
rect 18981 6749 19015 6783
rect 19349 6749 19383 6783
rect 19625 6749 19659 6783
rect 20085 6749 20119 6783
rect 3893 6681 3927 6715
rect 3341 6613 3375 6647
rect 4353 6613 4387 6647
rect 6009 6613 6043 6647
rect 8125 6613 8159 6647
rect 13645 6613 13679 6647
rect 15301 6613 15335 6647
rect 17049 6613 17083 6647
rect 18153 6613 18187 6647
rect 18613 6613 18647 6647
rect 18889 6613 18923 6647
rect 1593 6409 1627 6443
rect 2329 6409 2363 6443
rect 4445 6409 4479 6443
rect 5549 6409 5583 6443
rect 8217 6409 8251 6443
rect 9873 6409 9907 6443
rect 10057 6409 10091 6443
rect 12541 6409 12575 6443
rect 15853 6409 15887 6443
rect 15945 6409 15979 6443
rect 20269 6409 20303 6443
rect 1501 6341 1535 6375
rect 8769 6341 8803 6375
rect 9045 6341 9079 6375
rect 9505 6341 9539 6375
rect 18797 6341 18831 6375
rect 2053 6273 2087 6307
rect 2789 6273 2823 6307
rect 3801 6273 3835 6307
rect 4537 6273 4571 6307
rect 4811 6273 4845 6307
rect 6101 6273 6135 6307
rect 6561 6273 6595 6307
rect 7205 6273 7239 6307
rect 7479 6283 7513 6317
rect 9137 6273 9171 6307
rect 10241 6273 10275 6307
rect 11069 6273 11103 6307
rect 11161 6273 11195 6307
rect 11345 6273 11379 6307
rect 11529 6273 11563 6307
rect 11803 6273 11837 6307
rect 13335 6273 13369 6307
rect 14740 6273 14774 6307
rect 16129 6273 16163 6307
rect 16313 6273 16347 6307
rect 16497 6273 16531 6307
rect 16865 6273 16899 6307
rect 17139 6273 17173 6307
rect 18429 6273 18463 6307
rect 18613 6273 18647 6307
rect 19145 6273 19179 6307
rect 20361 6273 20395 6307
rect 2605 6205 2639 6239
rect 3525 6205 3559 6239
rect 3663 6205 3697 6239
rect 13093 6205 13127 6239
rect 14473 6205 14507 6239
rect 16405 6205 16439 6239
rect 18889 6205 18923 6239
rect 3249 6137 3283 6171
rect 14105 6137 14139 6171
rect 18429 6137 18463 6171
rect 5917 6069 5951 6103
rect 6377 6069 6411 6103
rect 10425 6069 10459 6103
rect 10885 6069 10919 6103
rect 11253 6069 11287 6103
rect 17877 6069 17911 6103
rect 20453 6069 20487 6103
rect 3065 5865 3099 5899
rect 3985 5865 4019 5899
rect 7021 5865 7055 5899
rect 9965 5865 9999 5899
rect 11345 5865 11379 5899
rect 12633 5865 12667 5899
rect 12909 5865 12943 5899
rect 18521 5865 18555 5899
rect 12449 5797 12483 5831
rect 13553 5797 13587 5831
rect 16313 5797 16347 5831
rect 16681 5797 16715 5831
rect 2053 5729 2087 5763
rect 6009 5729 6043 5763
rect 8953 5729 8987 5763
rect 13737 5729 13771 5763
rect 14105 5729 14139 5763
rect 19073 5729 19107 5763
rect 19257 5729 19291 5763
rect 1501 5661 1535 5695
rect 1869 5661 1903 5695
rect 2327 5661 2361 5695
rect 3617 5661 3651 5695
rect 4537 5661 4571 5695
rect 4629 5661 4663 5695
rect 4903 5661 4937 5695
rect 6283 5661 6317 5695
rect 9211 5631 9245 5665
rect 10333 5661 10367 5695
rect 10607 5661 10641 5695
rect 11989 5661 12023 5695
rect 12265 5661 12299 5695
rect 12541 5661 12575 5695
rect 12817 5661 12851 5695
rect 13093 5655 13127 5689
rect 13553 5661 13587 5695
rect 14379 5661 14413 5695
rect 15669 5661 15703 5695
rect 16037 5661 16071 5695
rect 16405 5661 16439 5695
rect 16865 5661 16899 5695
rect 17141 5661 17175 5695
rect 19531 5661 19565 5695
rect 3893 5593 3927 5627
rect 13921 5593 13955 5627
rect 17386 5593 17420 5627
rect 18889 5593 18923 5627
rect 3433 5525 3467 5559
rect 4353 5525 4387 5559
rect 5641 5525 5675 5559
rect 13185 5525 13219 5559
rect 15117 5525 15151 5559
rect 20269 5525 20303 5559
rect 1593 5321 1627 5355
rect 1961 5321 1995 5355
rect 6193 5321 6227 5355
rect 7849 5321 7883 5355
rect 9413 5321 9447 5355
rect 10793 5321 10827 5355
rect 11161 5321 11195 5355
rect 11805 5321 11839 5355
rect 12081 5321 12115 5355
rect 12541 5321 12575 5355
rect 15209 5321 15243 5355
rect 17509 5321 17543 5355
rect 6561 5253 6595 5287
rect 7665 5253 7699 5287
rect 13982 5253 14016 5287
rect 16033 5253 16067 5287
rect 1501 5185 1535 5219
rect 2145 5185 2179 5219
rect 2237 5185 2271 5219
rect 2421 5185 2455 5219
rect 3433 5185 3467 5219
rect 4537 5185 4571 5219
rect 5390 5185 5424 5219
rect 5549 5185 5583 5219
rect 6837 5185 6871 5219
rect 6929 5185 6963 5219
rect 7297 5185 7331 5219
rect 8401 5185 8435 5219
rect 8675 5185 8709 5219
rect 10023 5185 10057 5219
rect 11345 5185 11379 5219
rect 11713 5185 11747 5219
rect 11897 5185 11931 5219
rect 12265 5185 12299 5219
rect 12357 5185 12391 5219
rect 12817 5185 12851 5219
rect 13093 5185 13127 5219
rect 13553 5185 13587 5219
rect 13737 5185 13771 5219
rect 15393 5185 15427 5219
rect 15485 5185 15519 5219
rect 15669 5185 15703 5219
rect 16129 5185 16163 5219
rect 16865 5185 16899 5219
rect 17049 5185 17083 5219
rect 17417 5185 17451 5219
rect 17693 5185 17727 5219
rect 17967 5185 18001 5219
rect 19165 5185 19199 5219
rect 19432 5185 19466 5219
rect 3157 5117 3191 5151
rect 3295 5117 3329 5151
rect 4353 5117 4387 5151
rect 5273 5117 5307 5151
rect 9781 5117 9815 5151
rect 2881 5049 2915 5083
rect 4997 5049 5031 5083
rect 12633 5049 12667 5083
rect 13277 5049 13311 5083
rect 13369 5049 13403 5083
rect 15117 5049 15151 5083
rect 15669 5049 15703 5083
rect 17233 5049 17267 5083
rect 18705 5049 18739 5083
rect 4077 4981 4111 5015
rect 16221 4981 16255 5015
rect 16681 4981 16715 5015
rect 20545 4981 20579 5015
rect 1593 4777 1627 4811
rect 1961 4777 1995 4811
rect 3341 4777 3375 4811
rect 4537 4777 4571 4811
rect 5181 4777 5215 4811
rect 6377 4777 6411 4811
rect 7757 4777 7791 4811
rect 9873 4777 9907 4811
rect 10793 4777 10827 4811
rect 11161 4777 11195 4811
rect 12449 4777 12483 4811
rect 12633 4777 12667 4811
rect 13185 4777 13219 4811
rect 13829 4777 13863 4811
rect 14933 4777 14967 4811
rect 9413 4709 9447 4743
rect 10333 4709 10367 4743
rect 10977 4709 11011 4743
rect 11805 4709 11839 4743
rect 12909 4709 12943 4743
rect 14289 4709 14323 4743
rect 17601 4709 17635 4743
rect 20085 4709 20119 4743
rect 6745 4641 6779 4675
rect 12173 4641 12207 4675
rect 14473 4641 14507 4675
rect 15117 4641 15151 4675
rect 17417 4641 17451 4675
rect 1501 4573 1535 4607
rect 2145 4573 2179 4607
rect 2329 4573 2363 4607
rect 2603 4573 2637 4607
rect 3893 4573 3927 4607
rect 5365 4573 5399 4607
rect 5607 4573 5641 4607
rect 7003 4543 7037 4577
rect 10517 4573 10551 4607
rect 10609 4573 10643 4607
rect 10885 4573 10919 4607
rect 11345 4573 11379 4607
rect 11713 4573 11747 4607
rect 11989 4573 12023 4607
rect 12081 4573 12115 4607
rect 12357 4573 12391 4607
rect 12541 4573 12575 4607
rect 12817 4573 12851 4607
rect 13093 4573 13127 4607
rect 13369 4573 13403 4607
rect 13645 4573 13679 4607
rect 13737 4573 13771 4607
rect 13921 4573 13955 4607
rect 14289 4573 14323 4607
rect 14749 4573 14783 4607
rect 15025 4573 15059 4607
rect 15217 4573 15251 4607
rect 15393 4573 15427 4607
rect 17601 4573 17635 4607
rect 18061 4573 18095 4607
rect 18889 4573 18923 4607
rect 19257 4573 19291 4607
rect 19625 4573 19659 4607
rect 20085 4573 20119 4607
rect 4445 4505 4479 4539
rect 5089 4505 5123 4539
rect 14657 4505 14691 4539
rect 15638 4505 15672 4539
rect 16957 4505 16991 4539
rect 17969 4505 18003 4539
rect 3985 4437 4019 4471
rect 10149 4437 10183 4471
rect 11529 4437 11563 4471
rect 13461 4437 13495 4471
rect 16773 4437 16807 4471
rect 17049 4437 17083 4471
rect 5641 4233 5675 4267
rect 9597 4233 9631 4267
rect 10517 4233 10551 4267
rect 10885 4233 10919 4267
rect 12173 4233 12207 4267
rect 12449 4233 12483 4267
rect 13461 4233 13495 4267
rect 13921 4233 13955 4267
rect 19901 4233 19935 4267
rect 20453 4233 20487 4267
rect 1777 4165 1811 4199
rect 14372 4165 14406 4199
rect 16313 4165 16347 4199
rect 16865 4165 16899 4199
rect 1593 4097 1627 4131
rect 2513 4097 2547 4131
rect 3249 4097 3283 4131
rect 3387 4097 3421 4131
rect 4169 4097 4203 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 4903 4097 4937 4131
rect 10241 4097 10275 4131
rect 10333 4097 10367 4131
rect 10609 4097 10643 4131
rect 10793 4097 10827 4131
rect 11069 4097 11103 4131
rect 11345 4097 11379 4131
rect 11621 4097 11655 4131
rect 12081 4097 12115 4131
rect 12357 4097 12391 4131
rect 12633 4097 12667 4131
rect 12725 4097 12759 4131
rect 12909 4097 12943 4131
rect 13185 4097 13219 4131
rect 13645 4097 13679 4131
rect 13737 4097 13771 4131
rect 15761 4097 15795 4131
rect 16497 4097 16531 4131
rect 17141 4097 17175 4131
rect 17415 4097 17449 4131
rect 18521 4097 18555 4131
rect 18777 4097 18811 4131
rect 20085 4097 20119 4131
rect 20361 4097 20395 4131
rect 2329 4029 2363 4063
rect 3525 4029 3559 4063
rect 9965 4029 9999 4063
rect 14105 4029 14139 4063
rect 20269 4029 20303 4063
rect 1409 3961 1443 3995
rect 2973 3961 3007 3995
rect 12817 3961 12851 3995
rect 15485 3961 15519 3995
rect 1869 3893 1903 3927
rect 4261 3893 4295 3927
rect 8861 3893 8895 3927
rect 9229 3893 9263 3927
rect 10057 3893 10091 3927
rect 10701 3893 10735 3927
rect 11161 3893 11195 3927
rect 11713 3893 11747 3927
rect 11897 3893 11931 3927
rect 13369 3893 13403 3927
rect 15853 3893 15887 3927
rect 16957 3893 16991 3927
rect 18153 3893 18187 3927
rect 2605 3689 2639 3723
rect 3157 3689 3191 3723
rect 3985 3689 4019 3723
rect 4353 3689 4387 3723
rect 4629 3689 4663 3723
rect 7481 3689 7515 3723
rect 8309 3689 8343 3723
rect 8953 3689 8987 3723
rect 10793 3689 10827 3723
rect 11253 3689 11287 3723
rect 12081 3689 12115 3723
rect 6561 3621 6595 3655
rect 10333 3621 10367 3655
rect 11713 3621 11747 3655
rect 11805 3621 11839 3655
rect 12633 3621 12667 3655
rect 15485 3621 15519 3655
rect 17417 3621 17451 3655
rect 17877 3553 17911 3587
rect 19349 3553 19383 3587
rect 20177 3553 20211 3587
rect 1593 3485 1627 3519
rect 1867 3485 1901 3519
rect 4537 3485 4571 3519
rect 4813 3485 4847 3519
rect 6745 3485 6779 3519
rect 7021 3485 7055 3519
rect 7297 3485 7331 3519
rect 7665 3485 7699 3519
rect 7941 3485 7975 3519
rect 9137 3485 9171 3519
rect 9505 3485 9539 3519
rect 9873 3485 9907 3519
rect 10057 3485 10091 3519
rect 10149 3485 10183 3519
rect 10609 3485 10643 3519
rect 11161 3485 11195 3519
rect 11437 3485 11471 3519
rect 11529 3485 11563 3519
rect 11989 3485 12023 3519
rect 12265 3485 12299 3519
rect 12541 3485 12575 3519
rect 12817 3485 12851 3519
rect 13093 3485 13127 3519
rect 13461 3485 13495 3519
rect 13737 3485 13771 3519
rect 14105 3485 14139 3519
rect 14379 3485 14413 3519
rect 15669 3485 15703 3519
rect 15945 3485 15979 3519
rect 16405 3485 16439 3519
rect 16679 3485 16713 3519
rect 18153 3485 18187 3519
rect 18613 3485 18647 3519
rect 18889 3485 18923 3519
rect 19625 3485 19659 3519
rect 20085 3485 20119 3519
rect 3065 3417 3099 3451
rect 3893 3417 3927 3451
rect 8769 3417 8803 3451
rect 6837 3349 6871 3383
rect 7113 3349 7147 3383
rect 7757 3349 7791 3383
rect 9321 3349 9355 3383
rect 10057 3349 10091 3383
rect 10977 3349 11011 3383
rect 12357 3349 12391 3383
rect 12909 3349 12943 3383
rect 13277 3349 13311 3383
rect 13553 3349 13587 3383
rect 15117 3349 15151 3383
rect 16037 3349 16071 3383
rect 1593 3145 1627 3179
rect 2329 3145 2363 3179
rect 3709 3145 3743 3179
rect 4261 3145 4295 3179
rect 5825 3145 5859 3179
rect 12449 3145 12483 3179
rect 13461 3145 13495 3179
rect 18245 3145 18279 3179
rect 18521 3145 18555 3179
rect 20361 3145 20395 3179
rect 1501 3077 1535 3111
rect 15025 3077 15059 3111
rect 15761 3077 15795 3111
rect 16313 3077 16347 3111
rect 18950 3077 18984 3111
rect 20269 3077 20303 3111
rect 2053 3009 2087 3043
rect 2955 3009 2989 3043
rect 6009 3009 6043 3043
rect 6653 3009 6687 3043
rect 6929 3009 6963 3043
rect 7205 3009 7239 3043
rect 7481 3009 7515 3043
rect 7757 3009 7791 3043
rect 8033 3009 8067 3043
rect 8309 3009 8343 3043
rect 8585 3009 8619 3043
rect 8861 3009 8895 3043
rect 9137 3009 9171 3043
rect 9413 3009 9447 3043
rect 9689 3009 9723 3043
rect 9965 3009 9999 3043
rect 10057 3009 10091 3043
rect 10333 3009 10367 3043
rect 10793 3009 10827 3043
rect 11069 3009 11103 3043
rect 11161 3009 11195 3043
rect 11805 2993 11839 3027
rect 11923 3009 11957 3043
rect 12173 3009 12207 3043
rect 12625 3009 12659 3043
rect 12725 3009 12759 3043
rect 13185 3009 13219 3043
rect 13369 3009 13403 3043
rect 13645 3009 13679 3043
rect 13829 3009 13863 3043
rect 14105 3009 14139 3043
rect 14657 3009 14691 3043
rect 15209 3009 15243 3043
rect 16497 3009 16531 3043
rect 17121 3009 17155 3043
rect 18429 3009 18463 3043
rect 18705 3009 18739 3043
rect 2697 2941 2731 2975
rect 14473 2941 14507 2975
rect 14933 2941 14967 2975
rect 16865 2941 16899 2975
rect 7297 2873 7331 2907
rect 10241 2873 10275 2907
rect 11345 2873 11379 2907
rect 12081 2873 12115 2907
rect 12357 2873 12391 2907
rect 12909 2873 12943 2907
rect 13277 2873 13311 2907
rect 20085 2873 20119 2907
rect 6469 2805 6503 2839
rect 6745 2805 6779 2839
rect 7021 2805 7055 2839
rect 7573 2805 7607 2839
rect 7849 2805 7883 2839
rect 8125 2805 8159 2839
rect 8401 2805 8435 2839
rect 8677 2805 8711 2839
rect 8953 2805 8987 2839
rect 9229 2805 9263 2839
rect 9505 2805 9539 2839
rect 9781 2805 9815 2839
rect 10425 2805 10459 2839
rect 10609 2805 10643 2839
rect 10885 2805 10919 2839
rect 11621 2805 11655 2839
rect 13921 2805 13955 2839
rect 14289 2805 14323 2839
rect 15301 2805 15335 2839
rect 15853 2805 15887 2839
rect 1685 2601 1719 2635
rect 2881 2601 2915 2635
rect 3617 2601 3651 2635
rect 4353 2601 4387 2635
rect 4813 2601 4847 2635
rect 5365 2601 5399 2635
rect 6193 2601 6227 2635
rect 7021 2601 7055 2635
rect 7849 2601 7883 2635
rect 14105 2601 14139 2635
rect 16405 2601 16439 2635
rect 5733 2533 5767 2567
rect 7389 2533 7423 2567
rect 10517 2533 10551 2567
rect 11805 2533 11839 2567
rect 18889 2533 18923 2567
rect 1869 2465 1903 2499
rect 13829 2465 13863 2499
rect 17509 2465 17543 2499
rect 18521 2465 18555 2499
rect 1501 2397 1535 2431
rect 2143 2397 2177 2431
rect 3433 2397 3467 2431
rect 3801 2397 3835 2431
rect 4537 2397 4571 2431
rect 4629 2397 4663 2431
rect 5181 2397 5215 2431
rect 6837 2397 6871 2431
rect 7573 2397 7607 2431
rect 8401 2397 8435 2431
rect 8493 2397 8527 2431
rect 9229 2397 9263 2431
rect 9505 2397 9539 2431
rect 9597 2397 9631 2431
rect 10149 2397 10183 2431
rect 10425 2397 10459 2431
rect 10701 2397 10735 2431
rect 10977 2397 11011 2431
rect 11345 2397 11379 2431
rect 11437 2397 11471 2431
rect 11989 2397 12023 2431
rect 12265 2397 12299 2431
rect 12541 2397 12575 2431
rect 12817 2397 12851 2431
rect 13185 2397 13219 2431
rect 13553 2397 13587 2431
rect 14289 2397 14323 2431
rect 14749 2397 14783 2431
rect 15016 2397 15050 2431
rect 16313 2397 16347 2431
rect 16681 2397 16715 2431
rect 19073 2397 19107 2431
rect 20545 2397 20579 2431
rect 5549 2329 5583 2363
rect 6101 2329 6135 2363
rect 6561 2329 6595 2363
rect 17877 2329 17911 2363
rect 19349 2329 19383 2363
rect 3985 2261 4019 2295
rect 6653 2261 6687 2295
rect 8217 2261 8251 2295
rect 8677 2261 8711 2295
rect 9045 2261 9079 2295
rect 9321 2261 9355 2295
rect 9781 2261 9815 2295
rect 9965 2261 9999 2295
rect 10241 2261 10275 2295
rect 10793 2261 10827 2295
rect 11161 2261 11195 2295
rect 11621 2261 11655 2295
rect 12081 2261 12115 2295
rect 12357 2261 12391 2295
rect 12633 2261 12667 2295
rect 13001 2261 13035 2295
rect 14657 2261 14691 2295
rect 16129 2261 16163 2295
rect 17969 2261 18003 2295
rect 19441 2261 19475 2295
rect 19993 2261 20027 2295
rect 20361 2261 20395 2295
rect 1777 2057 1811 2091
rect 2697 2057 2731 2091
rect 3801 2057 3835 2091
rect 7021 2057 7055 2091
rect 15209 2057 15243 2091
rect 19809 2057 19843 2091
rect 2421 1989 2455 2023
rect 2605 1989 2639 2023
rect 6009 1989 6043 2023
rect 7665 1989 7699 2023
rect 8769 1989 8803 2023
rect 10977 1989 11011 2023
rect 12357 1989 12391 2023
rect 12909 1989 12943 2023
rect 13995 1989 14029 2023
rect 14565 1989 14599 2023
rect 1685 1921 1719 1955
rect 3249 1921 3283 1955
rect 3709 1921 3743 1955
rect 3985 1921 4019 1955
rect 4629 1921 4663 1955
rect 4997 1921 5031 1955
rect 5825 1921 5859 1955
rect 6469 1921 6503 1955
rect 6837 1921 6871 1955
rect 7205 1921 7239 1955
rect 7941 1921 7975 1955
rect 8309 1921 8343 1955
rect 9321 1921 9355 1955
rect 9873 1921 9907 1955
rect 10425 1921 10459 1955
rect 11805 1921 11839 1955
rect 13461 1921 13495 1955
rect 15025 1921 15059 1955
rect 15669 1921 15703 1955
rect 16681 1921 16715 1955
rect 18521 1921 18555 1955
rect 20545 1921 20579 1955
rect 4721 1853 4755 1887
rect 6193 1853 6227 1887
rect 16037 1853 16071 1887
rect 3433 1785 3467 1819
rect 4445 1785 4479 1819
rect 6653 1785 6687 1819
rect 14749 1785 14783 1819
rect 20361 1785 20395 1819
rect 4169 1717 4203 1751
rect 5641 1717 5675 1751
rect 7389 1717 7423 1751
rect 7757 1717 7791 1751
rect 8125 1717 8159 1751
rect 8493 1717 8527 1751
rect 9045 1717 9079 1751
rect 9597 1717 9631 1751
rect 10149 1717 10183 1751
rect 10517 1717 10551 1751
rect 11069 1717 11103 1751
rect 11897 1717 11931 1751
rect 12633 1717 12667 1751
rect 13001 1717 13035 1751
rect 13553 1717 13587 1751
rect 14105 1717 14139 1751
rect 17969 1717 18003 1751
rect 1869 1513 1903 1547
rect 2421 1513 2455 1547
rect 2789 1513 2823 1547
rect 4629 1513 4663 1547
rect 4997 1513 5031 1547
rect 5365 1513 5399 1547
rect 5733 1513 5767 1547
rect 6101 1513 6135 1547
rect 6653 1513 6687 1547
rect 7021 1513 7055 1547
rect 13185 1513 13219 1547
rect 20361 1513 20395 1547
rect 3249 1445 3283 1479
rect 3617 1445 3651 1479
rect 11713 1445 11747 1479
rect 14105 1445 14139 1479
rect 14749 1377 14783 1411
rect 17049 1377 17083 1411
rect 19625 1377 19659 1411
rect 3801 1309 3835 1343
rect 4077 1309 4111 1343
rect 6469 1309 6503 1343
rect 6929 1309 6963 1343
rect 7481 1309 7515 1343
rect 7849 1309 7883 1343
rect 8401 1309 8435 1343
rect 8953 1309 8987 1343
rect 10609 1309 10643 1343
rect 11069 1309 11103 1343
rect 11529 1309 11563 1343
rect 12541 1309 12575 1343
rect 13553 1309 13587 1343
rect 14289 1309 14323 1343
rect 14565 1309 14599 1343
rect 15669 1309 15703 1343
rect 16313 1309 16347 1343
rect 16681 1309 16715 1343
rect 17969 1309 18003 1343
rect 18061 1309 18095 1343
rect 18889 1309 18923 1343
rect 19349 1309 19383 1343
rect 20545 1309 20579 1343
rect 1777 1241 1811 1275
rect 2145 1241 2179 1275
rect 2697 1241 2731 1275
rect 3065 1241 3099 1275
rect 3433 1241 3467 1275
rect 4537 1241 4571 1275
rect 4905 1241 4939 1275
rect 5273 1241 5307 1275
rect 5641 1241 5675 1275
rect 6009 1241 6043 1275
rect 8217 1241 8251 1275
rect 8769 1241 8803 1275
rect 9413 1241 9447 1275
rect 9965 1241 9999 1275
rect 11989 1241 12023 1275
rect 12357 1241 12391 1275
rect 13093 1241 13127 1275
rect 3985 1173 4019 1207
rect 4261 1173 4295 1207
rect 7573 1173 7607 1207
rect 9137 1173 9171 1207
rect 9689 1173 9723 1207
rect 10057 1173 10091 1207
rect 10701 1173 10735 1207
rect 11253 1173 11287 1207
rect 12633 1173 12667 1207
rect 13737 1173 13771 1207
rect 17785 1173 17819 1207
<< metal1 >>
rect 11514 43976 11520 43988
rect 3252 43948 11520 43976
rect 1302 43800 1308 43852
rect 1360 43840 1366 43852
rect 3252 43840 3280 43948
rect 11514 43936 11520 43948
rect 11572 43936 11578 43988
rect 17770 43936 17776 43988
rect 17828 43976 17834 43988
rect 19426 43976 19432 43988
rect 17828 43948 19432 43976
rect 17828 43936 17834 43948
rect 19426 43936 19432 43948
rect 19484 43936 19490 43988
rect 12066 43908 12072 43920
rect 1360 43812 3280 43840
rect 7576 43880 12072 43908
rect 1360 43800 1366 43812
rect 2314 43732 2320 43784
rect 2372 43772 2378 43784
rect 7576 43772 7604 43880
rect 12066 43868 12072 43880
rect 12124 43868 12130 43920
rect 13538 43868 13544 43920
rect 13596 43908 13602 43920
rect 14918 43908 14924 43920
rect 13596 43880 14924 43908
rect 13596 43868 13602 43880
rect 14918 43868 14924 43880
rect 14976 43868 14982 43920
rect 18506 43868 18512 43920
rect 18564 43908 18570 43920
rect 19242 43908 19248 43920
rect 18564 43880 19248 43908
rect 18564 43868 18570 43880
rect 19242 43868 19248 43880
rect 19300 43868 19306 43920
rect 9858 43800 9864 43852
rect 9916 43840 9922 43852
rect 10134 43840 10140 43852
rect 9916 43812 10140 43840
rect 9916 43800 9922 43812
rect 10134 43800 10140 43812
rect 10192 43800 10198 43852
rect 19702 43840 19708 43852
rect 11716 43812 19708 43840
rect 2372 43744 7604 43772
rect 2372 43732 2378 43744
rect 5626 43664 5632 43716
rect 5684 43704 5690 43716
rect 9674 43704 9680 43716
rect 5684 43676 9680 43704
rect 5684 43664 5690 43676
rect 9674 43664 9680 43676
rect 9732 43664 9738 43716
rect 11716 43648 11744 43812
rect 19702 43800 19708 43812
rect 19760 43800 19766 43852
rect 12434 43732 12440 43784
rect 12492 43772 12498 43784
rect 12492 43744 19104 43772
rect 12492 43732 12498 43744
rect 19076 43716 19104 43744
rect 13814 43664 13820 43716
rect 13872 43704 13878 43716
rect 15194 43704 15200 43716
rect 13872 43676 15200 43704
rect 13872 43664 13878 43676
rect 15194 43664 15200 43676
rect 15252 43664 15258 43716
rect 19058 43664 19064 43716
rect 19116 43664 19122 43716
rect 1486 43596 1492 43648
rect 1544 43636 1550 43648
rect 10134 43636 10140 43648
rect 1544 43608 10140 43636
rect 1544 43596 1550 43608
rect 10134 43596 10140 43608
rect 10192 43596 10198 43648
rect 11698 43596 11704 43648
rect 11756 43596 11762 43648
rect 13630 43596 13636 43648
rect 13688 43636 13694 43648
rect 14182 43636 14188 43648
rect 13688 43608 14188 43636
rect 13688 43596 13694 43608
rect 14182 43596 14188 43608
rect 14240 43596 14246 43648
rect 14826 43596 14832 43648
rect 14884 43636 14890 43648
rect 19794 43636 19800 43648
rect 14884 43608 19800 43636
rect 14884 43596 14890 43608
rect 19794 43596 19800 43608
rect 19852 43596 19858 43648
rect 1104 43546 21043 43568
rect 1104 43494 5894 43546
rect 5946 43494 5958 43546
rect 6010 43494 6022 43546
rect 6074 43494 6086 43546
rect 6138 43494 6150 43546
rect 6202 43494 10839 43546
rect 10891 43494 10903 43546
rect 10955 43494 10967 43546
rect 11019 43494 11031 43546
rect 11083 43494 11095 43546
rect 11147 43494 15784 43546
rect 15836 43494 15848 43546
rect 15900 43494 15912 43546
rect 15964 43494 15976 43546
rect 16028 43494 16040 43546
rect 16092 43494 20729 43546
rect 20781 43494 20793 43546
rect 20845 43494 20857 43546
rect 20909 43494 20921 43546
rect 20973 43494 20985 43546
rect 21037 43494 21043 43546
rect 1104 43472 21043 43494
rect 1673 43435 1731 43441
rect 1673 43401 1685 43435
rect 1719 43432 1731 43435
rect 2406 43432 2412 43444
rect 1719 43404 2412 43432
rect 1719 43401 1731 43404
rect 1673 43395 1731 43401
rect 2406 43392 2412 43404
rect 2464 43392 2470 43444
rect 2774 43392 2780 43444
rect 2832 43432 2838 43444
rect 3145 43435 3203 43441
rect 3145 43432 3157 43435
rect 2832 43404 3157 43432
rect 2832 43392 2838 43404
rect 3145 43401 3157 43404
rect 3191 43401 3203 43435
rect 3145 43395 3203 43401
rect 3510 43392 3516 43444
rect 3568 43392 3574 43444
rect 4154 43392 4160 43444
rect 4212 43392 4218 43444
rect 4522 43392 4528 43444
rect 4580 43392 4586 43444
rect 5534 43392 5540 43444
rect 5592 43432 5598 43444
rect 5905 43435 5963 43441
rect 5905 43432 5917 43435
rect 5592 43404 5917 43432
rect 5592 43392 5598 43404
rect 5905 43401 5917 43404
rect 5951 43401 5963 43435
rect 5905 43395 5963 43401
rect 7009 43435 7067 43441
rect 7009 43401 7021 43435
rect 7055 43432 7067 43435
rect 7374 43432 7380 43444
rect 7055 43404 7380 43432
rect 7055 43401 7067 43404
rect 7009 43395 7067 43401
rect 7374 43392 7380 43404
rect 7432 43392 7438 43444
rect 8297 43435 8355 43441
rect 8297 43401 8309 43435
rect 8343 43432 8355 43435
rect 8662 43432 8668 43444
rect 8343 43404 8668 43432
rect 8343 43401 8355 43404
rect 8297 43395 8355 43401
rect 8662 43392 8668 43404
rect 8720 43392 8726 43444
rect 9309 43435 9367 43441
rect 9309 43401 9321 43435
rect 9355 43401 9367 43435
rect 10594 43432 10600 43444
rect 9309 43395 9367 43401
rect 9968 43404 10600 43432
rect 2869 43367 2927 43373
rect 2869 43333 2881 43367
rect 2915 43364 2927 43367
rect 3528 43364 3556 43392
rect 7190 43364 7196 43376
rect 2915 43336 3556 43364
rect 5092 43336 7196 43364
rect 2915 43333 2927 43336
rect 2869 43327 2927 43333
rect 1486 43256 1492 43308
rect 1544 43256 1550 43308
rect 1949 43299 2007 43305
rect 1949 43265 1961 43299
rect 1995 43296 2007 43299
rect 2130 43296 2136 43308
rect 1995 43268 2136 43296
rect 1995 43265 2007 43268
rect 1949 43259 2007 43265
rect 2130 43256 2136 43268
rect 2188 43256 2194 43308
rect 2498 43256 2504 43308
rect 2556 43256 2562 43308
rect 3050 43256 3056 43308
rect 3108 43256 3114 43308
rect 3973 43299 4031 43305
rect 3973 43265 3985 43299
rect 4019 43296 4031 43299
rect 4154 43296 4160 43308
rect 4019 43268 4160 43296
rect 4019 43265 4031 43268
rect 3973 43259 4031 43265
rect 4154 43256 4160 43268
rect 4212 43256 4218 43308
rect 4338 43256 4344 43308
rect 4396 43296 4402 43308
rect 5092 43305 5120 43336
rect 7190 43324 7196 43336
rect 7248 43324 7254 43376
rect 7837 43367 7895 43373
rect 7837 43333 7849 43367
rect 7883 43364 7895 43367
rect 8386 43364 8392 43376
rect 7883 43336 8392 43364
rect 7883 43333 7895 43336
rect 7837 43327 7895 43333
rect 8386 43324 8392 43336
rect 8444 43324 8450 43376
rect 8570 43324 8576 43376
rect 8628 43364 8634 43376
rect 9324 43364 9352 43395
rect 9968 43373 9996 43404
rect 10594 43392 10600 43404
rect 10652 43392 10658 43444
rect 11333 43435 11391 43441
rect 11333 43432 11345 43435
rect 10704 43404 11345 43432
rect 8628 43336 9352 43364
rect 9953 43367 10011 43373
rect 8628 43324 8634 43336
rect 9953 43333 9965 43367
rect 9999 43333 10011 43367
rect 10321 43367 10379 43373
rect 10321 43364 10333 43367
rect 9953 43327 10011 43333
rect 10060 43336 10333 43364
rect 4433 43299 4491 43305
rect 4433 43296 4445 43299
rect 4396 43268 4445 43296
rect 4396 43256 4402 43268
rect 4433 43265 4445 43268
rect 4479 43265 4491 43299
rect 4433 43259 4491 43265
rect 5077 43299 5135 43305
rect 5077 43265 5089 43299
rect 5123 43265 5135 43299
rect 5077 43259 5135 43265
rect 5258 43256 5264 43308
rect 5316 43256 5322 43308
rect 5442 43256 5448 43308
rect 5500 43296 5506 43308
rect 5813 43299 5871 43305
rect 5813 43296 5825 43299
rect 5500 43268 5825 43296
rect 5500 43256 5506 43268
rect 5813 43265 5825 43268
rect 5859 43265 5871 43299
rect 5813 43259 5871 43265
rect 6549 43299 6607 43305
rect 6549 43265 6561 43299
rect 6595 43265 6607 43299
rect 6549 43259 6607 43265
rect 2225 43231 2283 43237
rect 2225 43197 2237 43231
rect 2271 43228 2283 43231
rect 3142 43228 3148 43240
rect 2271 43200 3148 43228
rect 2271 43197 2283 43200
rect 2225 43191 2283 43197
rect 3142 43188 3148 43200
rect 3200 43188 3206 43240
rect 6564 43228 6592 43259
rect 6730 43256 6736 43308
rect 6788 43256 6794 43308
rect 7469 43299 7527 43305
rect 7469 43265 7481 43299
rect 7515 43265 7527 43299
rect 7469 43259 7527 43265
rect 8021 43299 8079 43305
rect 8021 43265 8033 43299
rect 8067 43265 8079 43299
rect 8021 43259 8079 43265
rect 8481 43299 8539 43305
rect 8481 43265 8493 43299
rect 8527 43296 8539 43299
rect 9030 43296 9036 43308
rect 8527 43268 9036 43296
rect 8527 43265 8539 43268
rect 8481 43259 8539 43265
rect 7374 43228 7380 43240
rect 6564 43200 7380 43228
rect 7374 43188 7380 43200
rect 7432 43188 7438 43240
rect 5537 43163 5595 43169
rect 5537 43129 5549 43163
rect 5583 43160 5595 43163
rect 5810 43160 5816 43172
rect 5583 43132 5816 43160
rect 5583 43129 5595 43132
rect 5537 43123 5595 43129
rect 5810 43120 5816 43132
rect 5868 43120 5874 43172
rect 6365 43163 6423 43169
rect 6365 43129 6377 43163
rect 6411 43160 6423 43163
rect 6914 43160 6920 43172
rect 6411 43132 6920 43160
rect 6411 43129 6423 43132
rect 6365 43123 6423 43129
rect 6914 43120 6920 43132
rect 6972 43120 6978 43172
rect 7484 43160 7512 43259
rect 8036 43228 8064 43259
rect 9030 43256 9036 43268
rect 9088 43256 9094 43308
rect 9125 43299 9183 43305
rect 9125 43265 9137 43299
rect 9171 43296 9183 43299
rect 9398 43296 9404 43308
rect 9171 43268 9404 43296
rect 9171 43265 9183 43268
rect 9125 43259 9183 43265
rect 9398 43256 9404 43268
rect 9456 43256 9462 43308
rect 9490 43256 9496 43308
rect 9548 43256 9554 43308
rect 9858 43256 9864 43308
rect 9916 43296 9922 43308
rect 10060 43296 10088 43336
rect 10321 43333 10333 43336
rect 10367 43333 10379 43367
rect 10321 43327 10379 43333
rect 10410 43324 10416 43376
rect 10468 43364 10474 43376
rect 10704 43364 10732 43404
rect 11333 43401 11345 43404
rect 11379 43401 11391 43435
rect 11333 43395 11391 43401
rect 11514 43392 11520 43444
rect 11572 43432 11578 43444
rect 11885 43435 11943 43441
rect 11885 43432 11897 43435
rect 11572 43404 11897 43432
rect 11572 43392 11578 43404
rect 11885 43401 11897 43404
rect 11931 43401 11943 43435
rect 11885 43395 11943 43401
rect 13262 43392 13268 43444
rect 13320 43432 13326 43444
rect 13320 43404 14044 43432
rect 13320 43392 13326 43404
rect 11698 43364 11704 43376
rect 10468 43336 10732 43364
rect 11072 43336 11704 43364
rect 10468 43324 10474 43336
rect 9916 43268 10088 43296
rect 9916 43256 9922 43268
rect 10778 43256 10784 43308
rect 10836 43256 10842 43308
rect 11072 43305 11100 43336
rect 11698 43324 11704 43336
rect 11756 43324 11762 43376
rect 11790 43324 11796 43376
rect 11848 43324 11854 43376
rect 12894 43324 12900 43376
rect 12952 43364 12958 43376
rect 13449 43367 13507 43373
rect 13449 43364 13461 43367
rect 12952 43336 13461 43364
rect 12952 43324 12958 43336
rect 13449 43333 13461 43336
rect 13495 43333 13507 43367
rect 13449 43327 13507 43333
rect 11057 43299 11115 43305
rect 11057 43265 11069 43299
rect 11103 43265 11115 43299
rect 11057 43259 11115 43265
rect 11149 43299 11207 43305
rect 11149 43265 11161 43299
rect 11195 43296 11207 43299
rect 11974 43296 11980 43308
rect 11195 43268 11980 43296
rect 11195 43265 11207 43268
rect 11149 43259 11207 43265
rect 11974 43256 11980 43268
rect 12032 43256 12038 43308
rect 12250 43256 12256 43308
rect 12308 43256 12314 43308
rect 12342 43256 12348 43308
rect 12400 43296 12406 43308
rect 12621 43299 12679 43305
rect 12621 43296 12633 43299
rect 12400 43268 12633 43296
rect 12400 43256 12406 43268
rect 12621 43265 12633 43268
rect 12667 43265 12679 43299
rect 12621 43259 12679 43265
rect 12710 43256 12716 43308
rect 12768 43296 12774 43308
rect 12989 43299 13047 43305
rect 12989 43296 13001 43299
rect 12768 43268 13001 43296
rect 12768 43256 12774 43268
rect 12989 43265 13001 43268
rect 13035 43265 13047 43299
rect 12989 43259 13047 43265
rect 13909 43299 13967 43305
rect 13909 43265 13921 43299
rect 13955 43265 13967 43299
rect 14016 43296 14044 43404
rect 14458 43392 14464 43444
rect 14516 43432 14522 43444
rect 15841 43435 15899 43441
rect 14516 43404 15332 43432
rect 14516 43392 14522 43404
rect 14182 43324 14188 43376
rect 14240 43364 14246 43376
rect 15304 43364 15332 43404
rect 15841 43401 15853 43435
rect 15887 43432 15899 43435
rect 16114 43432 16120 43444
rect 15887 43404 16120 43432
rect 15887 43401 15899 43404
rect 15841 43395 15899 43401
rect 16114 43392 16120 43404
rect 16172 43392 16178 43444
rect 16206 43392 16212 43444
rect 16264 43432 16270 43444
rect 16853 43435 16911 43441
rect 16853 43432 16865 43435
rect 16264 43404 16865 43432
rect 16264 43392 16270 43404
rect 16853 43401 16865 43404
rect 16899 43401 16911 43435
rect 16853 43395 16911 43401
rect 17405 43435 17463 43441
rect 17405 43401 17417 43435
rect 17451 43401 17463 43435
rect 17405 43395 17463 43401
rect 16298 43364 16304 43376
rect 14240 43336 15240 43364
rect 15304 43336 16304 43364
rect 14240 43324 14246 43336
rect 14093 43299 14151 43305
rect 14093 43296 14105 43299
rect 14016 43268 14105 43296
rect 13909 43259 13967 43265
rect 14093 43265 14105 43268
rect 14139 43265 14151 43299
rect 14093 43259 14151 43265
rect 14645 43299 14703 43305
rect 14645 43265 14657 43299
rect 14691 43296 14703 43299
rect 14826 43296 14832 43308
rect 14691 43268 14832 43296
rect 14691 43265 14703 43268
rect 14645 43259 14703 43265
rect 8754 43228 8760 43240
rect 8036 43200 8760 43228
rect 8754 43188 8760 43200
rect 8812 43188 8818 43240
rect 9674 43188 9680 43240
rect 9732 43228 9738 43240
rect 13924 43228 13952 43259
rect 14826 43256 14832 43268
rect 14884 43256 14890 43308
rect 14918 43256 14924 43308
rect 14976 43256 14982 43308
rect 15102 43256 15108 43308
rect 15160 43256 15166 43308
rect 15212 43305 15240 43336
rect 16298 43324 16304 43336
rect 16356 43324 16362 43376
rect 16390 43324 16396 43376
rect 16448 43364 16454 43376
rect 17420 43364 17448 43395
rect 17494 43392 17500 43444
rect 17552 43432 17558 43444
rect 18325 43435 18383 43441
rect 18325 43432 18337 43435
rect 17552 43404 18337 43432
rect 17552 43392 17558 43404
rect 18325 43401 18337 43404
rect 18371 43401 18383 43435
rect 18325 43395 18383 43401
rect 19426 43392 19432 43444
rect 19484 43392 19490 43444
rect 19794 43392 19800 43444
rect 19852 43392 19858 43444
rect 16448 43336 17448 43364
rect 16448 43324 16454 43336
rect 15197 43299 15255 43305
rect 15197 43265 15209 43299
rect 15243 43265 15255 43299
rect 15197 43259 15255 43265
rect 15470 43256 15476 43308
rect 15528 43256 15534 43308
rect 15654 43256 15660 43308
rect 15712 43256 15718 43308
rect 16114 43256 16120 43308
rect 16172 43256 16178 43308
rect 16761 43299 16819 43305
rect 16761 43265 16773 43299
rect 16807 43296 16819 43299
rect 17218 43296 17224 43308
rect 16807 43268 17224 43296
rect 16807 43265 16819 43268
rect 16761 43259 16819 43265
rect 17218 43256 17224 43268
rect 17276 43256 17282 43308
rect 17313 43299 17371 43305
rect 17313 43265 17325 43299
rect 17359 43296 17371 43299
rect 17494 43296 17500 43308
rect 17359 43268 17500 43296
rect 17359 43265 17371 43268
rect 17313 43259 17371 43265
rect 17494 43256 17500 43268
rect 17552 43256 17558 43308
rect 17773 43299 17831 43305
rect 17773 43265 17785 43299
rect 17819 43296 17831 43299
rect 17954 43296 17960 43308
rect 17819 43268 17960 43296
rect 17819 43265 17831 43268
rect 17773 43259 17831 43265
rect 17954 43256 17960 43268
rect 18012 43256 18018 43308
rect 18138 43256 18144 43308
rect 18196 43296 18202 43308
rect 18233 43299 18291 43305
rect 18233 43296 18245 43299
rect 18196 43268 18245 43296
rect 18196 43256 18202 43268
rect 18233 43265 18245 43268
rect 18279 43265 18291 43299
rect 18233 43259 18291 43265
rect 18598 43256 18604 43308
rect 18656 43256 18662 43308
rect 18690 43256 18696 43308
rect 18748 43256 18754 43308
rect 19058 43256 19064 43308
rect 19116 43296 19122 43308
rect 19337 43299 19395 43305
rect 19337 43296 19349 43299
rect 19116 43268 19349 43296
rect 19116 43256 19122 43268
rect 19337 43265 19349 43268
rect 19383 43265 19395 43299
rect 19337 43259 19395 43265
rect 19978 43256 19984 43308
rect 20036 43256 20042 43308
rect 20162 43256 20168 43308
rect 20220 43256 20226 43308
rect 15120 43228 15148 43256
rect 16393 43231 16451 43237
rect 9732 43200 10548 43228
rect 13924 43200 15056 43228
rect 15120 43200 15240 43228
rect 9732 43188 9738 43200
rect 8938 43160 8944 43172
rect 7484 43132 8944 43160
rect 8938 43120 8944 43132
rect 8996 43120 9002 43172
rect 10520 43169 10548 43200
rect 10505 43163 10563 43169
rect 10505 43129 10517 43163
rect 10551 43129 10563 43163
rect 11606 43160 11612 43172
rect 10505 43123 10563 43129
rect 10612 43132 11612 43160
rect 4893 43095 4951 43101
rect 4893 43061 4905 43095
rect 4939 43092 4951 43095
rect 5902 43092 5908 43104
rect 4939 43064 5908 43092
rect 4939 43061 4951 43064
rect 4893 43055 4951 43061
rect 5902 43052 5908 43064
rect 5960 43052 5966 43104
rect 5994 43052 6000 43104
rect 6052 43092 6058 43104
rect 8570 43092 8576 43104
rect 6052 43064 8576 43092
rect 6052 43052 6058 43064
rect 8570 43052 8576 43064
rect 8628 43052 8634 43104
rect 8665 43095 8723 43101
rect 8665 43061 8677 43095
rect 8711 43092 8723 43095
rect 9030 43092 9036 43104
rect 8711 43064 9036 43092
rect 8711 43061 8723 43064
rect 8665 43055 8723 43061
rect 9030 43052 9036 43064
rect 9088 43052 9094 43104
rect 9674 43052 9680 43104
rect 9732 43052 9738 43104
rect 9858 43052 9864 43104
rect 9916 43092 9922 43104
rect 10612 43101 10640 43132
rect 11606 43120 11612 43132
rect 11664 43120 11670 43172
rect 12710 43120 12716 43172
rect 12768 43160 12774 43172
rect 12768 43132 13216 43160
rect 12768 43120 12774 43132
rect 10045 43095 10103 43101
rect 10045 43092 10057 43095
rect 9916 43064 10057 43092
rect 9916 43052 9922 43064
rect 10045 43061 10057 43064
rect 10091 43061 10103 43095
rect 10045 43055 10103 43061
rect 10597 43095 10655 43101
rect 10597 43061 10609 43095
rect 10643 43061 10655 43095
rect 10597 43055 10655 43061
rect 10873 43095 10931 43101
rect 10873 43061 10885 43095
rect 10919 43092 10931 43095
rect 11146 43092 11152 43104
rect 10919 43064 11152 43092
rect 10919 43061 10931 43064
rect 10873 43055 10931 43061
rect 11146 43052 11152 43064
rect 11204 43052 11210 43104
rect 11974 43052 11980 43104
rect 12032 43092 12038 43104
rect 12437 43095 12495 43101
rect 12437 43092 12449 43095
rect 12032 43064 12449 43092
rect 12032 43052 12038 43064
rect 12437 43061 12449 43064
rect 12483 43061 12495 43095
rect 12437 43055 12495 43061
rect 12805 43095 12863 43101
rect 12805 43061 12817 43095
rect 12851 43092 12863 43095
rect 12986 43092 12992 43104
rect 12851 43064 12992 43092
rect 12851 43061 12863 43064
rect 12805 43055 12863 43061
rect 12986 43052 12992 43064
rect 13044 43052 13050 43104
rect 13188 43101 13216 43132
rect 13630 43120 13636 43172
rect 13688 43160 13694 43172
rect 15028 43169 15056 43200
rect 14737 43163 14795 43169
rect 14737 43160 14749 43163
rect 13688 43132 14749 43160
rect 13688 43120 13694 43132
rect 14737 43129 14749 43132
rect 14783 43129 14795 43163
rect 14737 43123 14795 43129
rect 15013 43163 15071 43169
rect 15013 43129 15025 43163
rect 15059 43129 15071 43163
rect 15212 43160 15240 43200
rect 16393 43197 16405 43231
rect 16439 43228 16451 43231
rect 18616 43228 18644 43256
rect 16439 43200 18644 43228
rect 16439 43197 16451 43200
rect 16393 43191 16451 43197
rect 15212 43132 16436 43160
rect 15013 43123 15071 43129
rect 16408 43104 16436 43132
rect 16942 43120 16948 43172
rect 17000 43160 17006 43172
rect 18877 43163 18935 43169
rect 18877 43160 18889 43163
rect 17000 43132 18889 43160
rect 17000 43120 17006 43132
rect 18877 43129 18889 43132
rect 18923 43129 18935 43163
rect 18877 43123 18935 43129
rect 13173 43095 13231 43101
rect 13173 43061 13185 43095
rect 13219 43061 13231 43095
rect 13173 43055 13231 43061
rect 13538 43052 13544 43104
rect 13596 43052 13602 43104
rect 13722 43052 13728 43104
rect 13780 43052 13786 43104
rect 14274 43052 14280 43104
rect 14332 43052 14338 43104
rect 14458 43052 14464 43104
rect 14516 43052 14522 43104
rect 14918 43052 14924 43104
rect 14976 43092 14982 43104
rect 15289 43095 15347 43101
rect 15289 43092 15301 43095
rect 14976 43064 15301 43092
rect 14976 43052 14982 43064
rect 15289 43061 15301 43064
rect 15335 43061 15347 43095
rect 15289 43055 15347 43061
rect 16390 43052 16396 43104
rect 16448 43052 16454 43104
rect 16574 43052 16580 43104
rect 16632 43092 16638 43104
rect 17957 43095 18015 43101
rect 17957 43092 17969 43095
rect 16632 43064 17969 43092
rect 16632 43052 16638 43064
rect 17957 43061 17969 43064
rect 18003 43061 18015 43095
rect 17957 43055 18015 43061
rect 18046 43052 18052 43104
rect 18104 43092 18110 43104
rect 18598 43092 18604 43104
rect 18104 43064 18604 43092
rect 18104 43052 18110 43064
rect 18598 43052 18604 43064
rect 18656 43052 18662 43104
rect 20441 43095 20499 43101
rect 20441 43061 20453 43095
rect 20487 43092 20499 43095
rect 21266 43092 21272 43104
rect 20487 43064 21272 43092
rect 20487 43061 20499 43064
rect 20441 43055 20499 43061
rect 21266 43052 21272 43064
rect 21324 43052 21330 43104
rect 1104 43002 20884 43024
rect 1104 42950 3422 43002
rect 3474 42950 3486 43002
rect 3538 42950 3550 43002
rect 3602 42950 3614 43002
rect 3666 42950 3678 43002
rect 3730 42950 8367 43002
rect 8419 42950 8431 43002
rect 8483 42950 8495 43002
rect 8547 42950 8559 43002
rect 8611 42950 8623 43002
rect 8675 42950 13312 43002
rect 13364 42950 13376 43002
rect 13428 42950 13440 43002
rect 13492 42950 13504 43002
rect 13556 42950 13568 43002
rect 13620 42950 18257 43002
rect 18309 42950 18321 43002
rect 18373 42950 18385 43002
rect 18437 42950 18449 43002
rect 18501 42950 18513 43002
rect 18565 42950 20884 43002
rect 1104 42928 20884 42950
rect 3694 42848 3700 42900
rect 3752 42888 3758 42900
rect 5258 42888 5264 42900
rect 3752 42860 5264 42888
rect 3752 42848 3758 42860
rect 5258 42848 5264 42860
rect 5316 42848 5322 42900
rect 6362 42848 6368 42900
rect 6420 42848 6426 42900
rect 7282 42848 7288 42900
rect 7340 42848 7346 42900
rect 7466 42848 7472 42900
rect 7524 42888 7530 42900
rect 7524 42860 9812 42888
rect 7524 42848 7530 42860
rect 1765 42823 1823 42829
rect 1765 42789 1777 42823
rect 1811 42789 1823 42823
rect 1765 42783 1823 42789
rect 1780 42752 1808 42783
rect 3602 42780 3608 42832
rect 3660 42820 3666 42832
rect 6380 42820 6408 42848
rect 9674 42820 9680 42832
rect 3660 42792 3924 42820
rect 6380 42792 9680 42820
rect 3660 42780 3666 42792
rect 3896 42764 3924 42792
rect 9674 42780 9680 42792
rect 9732 42780 9738 42832
rect 9784 42820 9812 42860
rect 10134 42848 10140 42900
rect 10192 42888 10198 42900
rect 10413 42891 10471 42897
rect 10413 42888 10425 42891
rect 10192 42860 10425 42888
rect 10192 42848 10198 42860
rect 10413 42857 10425 42860
rect 10459 42857 10471 42891
rect 10413 42851 10471 42857
rect 10870 42848 10876 42900
rect 10928 42848 10934 42900
rect 11149 42891 11207 42897
rect 11149 42857 11161 42891
rect 11195 42857 11207 42891
rect 11149 42851 11207 42857
rect 11164 42820 11192 42851
rect 12894 42848 12900 42900
rect 12952 42888 12958 42900
rect 14274 42888 14280 42900
rect 12952 42860 14280 42888
rect 12952 42848 12958 42860
rect 14274 42848 14280 42860
rect 14332 42848 14338 42900
rect 15120 42860 15976 42888
rect 15120 42832 15148 42860
rect 9784 42792 11192 42820
rect 11330 42780 11336 42832
rect 11388 42780 11394 42832
rect 12066 42780 12072 42832
rect 12124 42820 12130 42832
rect 13357 42823 13415 42829
rect 13357 42820 13369 42823
rect 12124 42792 13369 42820
rect 12124 42780 12130 42792
rect 13357 42789 13369 42792
rect 13403 42789 13415 42823
rect 13357 42783 13415 42789
rect 13446 42780 13452 42832
rect 13504 42820 13510 42832
rect 14642 42820 14648 42832
rect 13504 42792 14648 42820
rect 13504 42780 13510 42792
rect 14642 42780 14648 42792
rect 14700 42780 14706 42832
rect 15102 42780 15108 42832
rect 15160 42780 15166 42832
rect 3513 42755 3571 42761
rect 1780 42724 3464 42752
rect 1670 42644 1676 42696
rect 1728 42644 1734 42696
rect 1946 42644 1952 42696
rect 2004 42644 2010 42696
rect 2501 42687 2559 42693
rect 2501 42653 2513 42687
rect 2547 42684 2559 42687
rect 2958 42684 2964 42696
rect 2547 42656 2964 42684
rect 2547 42653 2559 42656
rect 2501 42647 2559 42653
rect 2958 42644 2964 42656
rect 3016 42644 3022 42696
rect 3053 42687 3111 42693
rect 3053 42653 3065 42687
rect 3099 42684 3111 42687
rect 3326 42684 3332 42696
rect 3099 42656 3332 42684
rect 3099 42653 3111 42656
rect 3053 42647 3111 42653
rect 3326 42644 3332 42656
rect 3384 42644 3390 42696
rect 3436 42684 3464 42724
rect 3513 42721 3525 42755
rect 3559 42752 3571 42755
rect 3786 42752 3792 42764
rect 3559 42724 3792 42752
rect 3559 42721 3571 42724
rect 3513 42715 3571 42721
rect 3786 42712 3792 42724
rect 3844 42712 3850 42764
rect 3878 42712 3884 42764
rect 3936 42712 3942 42764
rect 4157 42755 4215 42761
rect 4157 42721 4169 42755
rect 4203 42752 4215 42755
rect 4246 42752 4252 42764
rect 4203 42724 4252 42752
rect 4203 42721 4215 42724
rect 4157 42715 4215 42721
rect 4246 42712 4252 42724
rect 4304 42712 4310 42764
rect 4338 42712 4344 42764
rect 4396 42712 4402 42764
rect 4709 42755 4767 42761
rect 4709 42721 4721 42755
rect 4755 42752 4767 42755
rect 4982 42752 4988 42764
rect 4755 42724 4988 42752
rect 4755 42721 4767 42724
rect 4709 42715 4767 42721
rect 4982 42712 4988 42724
rect 5040 42712 5046 42764
rect 5261 42755 5319 42761
rect 5261 42721 5273 42755
rect 5307 42752 5319 42755
rect 5350 42752 5356 42764
rect 5307 42724 5356 42752
rect 5307 42721 5319 42724
rect 5261 42715 5319 42721
rect 5350 42712 5356 42724
rect 5408 42712 5414 42764
rect 5813 42755 5871 42761
rect 5813 42721 5825 42755
rect 5859 42752 5871 42755
rect 6270 42752 6276 42764
rect 5859 42724 6276 42752
rect 5859 42721 5871 42724
rect 5813 42715 5871 42721
rect 6270 42712 6276 42724
rect 6328 42712 6334 42764
rect 6365 42755 6423 42761
rect 6365 42721 6377 42755
rect 6411 42752 6423 42755
rect 6454 42752 6460 42764
rect 6411 42724 6460 42752
rect 6411 42721 6423 42724
rect 6365 42715 6423 42721
rect 6454 42712 6460 42724
rect 6512 42712 6518 42764
rect 8018 42712 8024 42764
rect 8076 42712 8082 42764
rect 8294 42712 8300 42764
rect 8352 42752 8358 42764
rect 8573 42755 8631 42761
rect 8573 42752 8585 42755
rect 8352 42724 8585 42752
rect 8352 42712 8358 42724
rect 8573 42721 8585 42724
rect 8619 42721 8631 42755
rect 8573 42715 8631 42721
rect 8956 42724 9260 42752
rect 4356 42684 4384 42712
rect 3436 42656 4384 42684
rect 5902 42644 5908 42696
rect 5960 42684 5966 42696
rect 6641 42687 6699 42693
rect 6641 42684 6653 42687
rect 5960 42656 6653 42684
rect 5960 42644 5966 42656
rect 6641 42653 6653 42656
rect 6687 42653 6699 42687
rect 6641 42647 6699 42653
rect 6914 42644 6920 42696
rect 6972 42684 6978 42696
rect 7193 42687 7251 42693
rect 7193 42684 7205 42687
rect 6972 42656 7205 42684
rect 6972 42644 6978 42656
rect 7193 42653 7205 42656
rect 7239 42653 7251 42687
rect 7193 42647 7251 42653
rect 2133 42619 2191 42625
rect 2133 42585 2145 42619
rect 2179 42585 2191 42619
rect 2133 42579 2191 42585
rect 1486 42508 1492 42560
rect 1544 42508 1550 42560
rect 2148 42548 2176 42579
rect 2682 42576 2688 42628
rect 2740 42576 2746 42628
rect 3237 42619 3295 42625
rect 3237 42585 3249 42619
rect 3283 42616 3295 42619
rect 3786 42616 3792 42628
rect 3283 42588 3792 42616
rect 3283 42585 3295 42588
rect 3237 42579 3295 42585
rect 3786 42576 3792 42588
rect 3844 42576 3850 42628
rect 3881 42619 3939 42625
rect 3881 42585 3893 42619
rect 3927 42585 3939 42619
rect 3881 42579 3939 42585
rect 2958 42548 2964 42560
rect 2148 42520 2964 42548
rect 2958 42508 2964 42520
rect 3016 42508 3022 42560
rect 3142 42508 3148 42560
rect 3200 42548 3206 42560
rect 3896 42548 3924 42579
rect 4246 42576 4252 42628
rect 4304 42616 4310 42628
rect 4433 42619 4491 42625
rect 4433 42616 4445 42619
rect 4304 42588 4445 42616
rect 4304 42576 4310 42588
rect 4433 42585 4445 42588
rect 4479 42585 4491 42619
rect 4433 42579 4491 42585
rect 4982 42576 4988 42628
rect 5040 42576 5046 42628
rect 5537 42619 5595 42625
rect 5537 42585 5549 42619
rect 5583 42616 5595 42619
rect 5810 42616 5816 42628
rect 5583 42588 5816 42616
rect 5583 42585 5595 42588
rect 5537 42579 5595 42585
rect 5810 42576 5816 42588
rect 5868 42576 5874 42628
rect 6089 42619 6147 42625
rect 6089 42585 6101 42619
rect 6135 42616 6147 42619
rect 6546 42616 6552 42628
rect 6135 42588 6552 42616
rect 6135 42585 6147 42588
rect 6089 42579 6147 42585
rect 6546 42576 6552 42588
rect 6604 42576 6610 42628
rect 7006 42576 7012 42628
rect 7064 42576 7070 42628
rect 7745 42619 7803 42625
rect 7745 42585 7757 42619
rect 7791 42616 7803 42619
rect 8018 42616 8024 42628
rect 7791 42588 8024 42616
rect 7791 42585 7803 42588
rect 7745 42579 7803 42585
rect 8018 42576 8024 42588
rect 8076 42576 8082 42628
rect 8297 42619 8355 42625
rect 8297 42585 8309 42619
rect 8343 42616 8355 42619
rect 8956 42616 8984 42724
rect 9033 42687 9091 42693
rect 9033 42653 9045 42687
rect 9079 42684 9091 42687
rect 9232 42684 9260 42724
rect 9416 42724 9628 42752
rect 9416 42684 9444 42724
rect 9490 42693 9496 42696
rect 9079 42656 9168 42684
rect 9232 42656 9444 42684
rect 9481 42687 9496 42693
rect 9079 42653 9091 42656
rect 9033 42647 9091 42653
rect 8343 42588 8984 42616
rect 9140 42616 9168 42656
rect 9481 42653 9493 42687
rect 9481 42647 9496 42653
rect 9490 42644 9496 42647
rect 9548 42644 9554 42696
rect 9600 42684 9628 42724
rect 9950 42712 9956 42764
rect 10008 42752 10014 42764
rect 11348 42752 11376 42780
rect 10008 42724 10640 42752
rect 10008 42712 10014 42724
rect 10045 42687 10103 42693
rect 9600 42656 9996 42684
rect 9968 42616 9996 42656
rect 10045 42653 10057 42687
rect 10091 42684 10103 42687
rect 10134 42684 10140 42696
rect 10091 42656 10140 42684
rect 10091 42653 10103 42656
rect 10045 42647 10103 42653
rect 10134 42644 10140 42656
rect 10192 42644 10198 42696
rect 10318 42644 10324 42696
rect 10376 42644 10382 42696
rect 10612 42693 10640 42724
rect 10704 42724 11376 42752
rect 10704 42693 10732 42724
rect 12618 42712 12624 42764
rect 12676 42752 12682 42764
rect 12676 42724 12940 42752
rect 12676 42712 12682 42724
rect 10597 42687 10655 42693
rect 10597 42653 10609 42687
rect 10643 42653 10655 42687
rect 10597 42647 10655 42653
rect 10689 42687 10747 42693
rect 10689 42653 10701 42687
rect 10735 42653 10747 42687
rect 10689 42647 10747 42653
rect 10870 42644 10876 42696
rect 10928 42684 10934 42696
rect 11057 42687 11115 42693
rect 11057 42684 11069 42687
rect 10928 42656 11069 42684
rect 10928 42644 10934 42656
rect 11057 42653 11069 42656
rect 11103 42653 11115 42687
rect 11057 42647 11115 42653
rect 11330 42644 11336 42696
rect 11388 42644 11394 42696
rect 11609 42687 11667 42693
rect 11609 42653 11621 42687
rect 11655 42684 11667 42687
rect 11882 42684 11888 42696
rect 11655 42656 11888 42684
rect 11655 42653 11667 42656
rect 11609 42647 11667 42653
rect 11882 42644 11888 42656
rect 11940 42644 11946 42696
rect 12066 42644 12072 42696
rect 12124 42644 12130 42696
rect 12526 42644 12532 42696
rect 12584 42644 12590 42696
rect 12802 42644 12808 42696
rect 12860 42644 12866 42696
rect 12912 42693 12940 42724
rect 14918 42712 14924 42764
rect 14976 42712 14982 42764
rect 15120 42724 15884 42752
rect 12897 42687 12955 42693
rect 12897 42653 12909 42687
rect 12943 42653 12955 42687
rect 12897 42647 12955 42653
rect 13170 42644 13176 42696
rect 13228 42644 13234 42696
rect 13630 42644 13636 42696
rect 13688 42684 13694 42696
rect 13725 42687 13783 42693
rect 13725 42684 13737 42687
rect 13688 42656 13737 42684
rect 13688 42644 13694 42656
rect 13725 42653 13737 42656
rect 13771 42653 13783 42687
rect 13725 42647 13783 42653
rect 14829 42687 14887 42693
rect 14829 42653 14841 42687
rect 14875 42684 14887 42687
rect 14936 42684 14964 42712
rect 15120 42693 15148 42724
rect 14875 42656 14964 42684
rect 15105 42687 15163 42693
rect 14875 42653 14887 42656
rect 14829 42647 14887 42653
rect 15105 42653 15117 42687
rect 15151 42653 15163 42687
rect 15105 42647 15163 42653
rect 15378 42644 15384 42696
rect 15436 42644 15442 42696
rect 15470 42644 15476 42696
rect 15528 42684 15534 42696
rect 15657 42687 15715 42693
rect 15657 42684 15669 42687
rect 15528 42656 15669 42684
rect 15528 42644 15534 42656
rect 15657 42653 15669 42656
rect 15703 42653 15715 42687
rect 15657 42647 15715 42653
rect 9140 42588 9904 42616
rect 9968 42588 11928 42616
rect 8343 42585 8355 42588
rect 8297 42579 8355 42585
rect 3200 42520 3924 42548
rect 3200 42508 3206 42520
rect 9122 42508 9128 42560
rect 9180 42508 9186 42560
rect 9674 42508 9680 42560
rect 9732 42508 9738 42560
rect 9876 42557 9904 42588
rect 9861 42551 9919 42557
rect 9861 42517 9873 42551
rect 9907 42517 9919 42551
rect 9861 42511 9919 42517
rect 10134 42508 10140 42560
rect 10192 42508 10198 42560
rect 11146 42508 11152 42560
rect 11204 42548 11210 42560
rect 11422 42548 11428 42560
rect 11204 42520 11428 42548
rect 11204 42508 11210 42520
rect 11422 42508 11428 42520
rect 11480 42508 11486 42560
rect 11514 42508 11520 42560
rect 11572 42508 11578 42560
rect 11790 42508 11796 42560
rect 11848 42508 11854 42560
rect 11900 42557 11928 42588
rect 12250 42576 12256 42628
rect 12308 42616 12314 42628
rect 14369 42619 14427 42625
rect 12308 42588 13124 42616
rect 12308 42576 12314 42588
rect 11885 42551 11943 42557
rect 11885 42517 11897 42551
rect 11931 42517 11943 42551
rect 11885 42511 11943 42517
rect 12342 42508 12348 42560
rect 12400 42508 12406 42560
rect 12618 42508 12624 42560
rect 12676 42508 12682 42560
rect 13096 42557 13124 42588
rect 14369 42585 14381 42619
rect 14415 42616 14427 42619
rect 15856 42616 15884 42724
rect 15948 42693 15976 42860
rect 16482 42848 16488 42900
rect 16540 42848 16546 42900
rect 17954 42848 17960 42900
rect 18012 42888 18018 42900
rect 19245 42891 19303 42897
rect 19245 42888 19257 42891
rect 18012 42860 19257 42888
rect 18012 42848 18018 42860
rect 19245 42857 19257 42860
rect 19291 42857 19303 42891
rect 19245 42851 19303 42857
rect 19889 42891 19947 42897
rect 19889 42857 19901 42891
rect 19935 42888 19947 42891
rect 19978 42888 19984 42900
rect 19935 42860 19984 42888
rect 19935 42857 19947 42860
rect 19889 42851 19947 42857
rect 19978 42848 19984 42860
rect 20036 42848 20042 42900
rect 17494 42780 17500 42832
rect 17552 42820 17558 42832
rect 19518 42820 19524 42832
rect 17552 42792 19524 42820
rect 17552 42780 17558 42792
rect 19518 42780 19524 42792
rect 19576 42780 19582 42832
rect 16758 42712 16764 42764
rect 16816 42752 16822 42764
rect 17221 42755 17279 42761
rect 17221 42752 17233 42755
rect 16816 42724 17233 42752
rect 16816 42712 16822 42724
rect 17221 42721 17233 42724
rect 17267 42721 17279 42755
rect 17221 42715 17279 42721
rect 17310 42712 17316 42764
rect 17368 42752 17374 42764
rect 17773 42755 17831 42761
rect 17773 42752 17785 42755
rect 17368 42724 17785 42752
rect 17368 42712 17374 42724
rect 17773 42721 17785 42724
rect 17819 42721 17831 42755
rect 17773 42715 17831 42721
rect 17862 42712 17868 42764
rect 17920 42752 17926 42764
rect 18877 42755 18935 42761
rect 18877 42752 18889 42755
rect 17920 42724 18889 42752
rect 17920 42712 17926 42724
rect 18877 42721 18889 42724
rect 18923 42721 18935 42755
rect 18877 42715 18935 42721
rect 19058 42712 19064 42764
rect 19116 42752 19122 42764
rect 19116 42724 20208 42752
rect 19116 42712 19122 42724
rect 15933 42687 15991 42693
rect 15933 42653 15945 42687
rect 15979 42653 15991 42687
rect 15933 42647 15991 42653
rect 16206 42644 16212 42696
rect 16264 42644 16270 42696
rect 16850 42644 16856 42696
rect 16908 42684 16914 42696
rect 20180 42693 20208 42724
rect 19429 42687 19487 42693
rect 19429 42684 19441 42687
rect 16908 42656 19441 42684
rect 16908 42644 16914 42656
rect 19429 42653 19441 42656
rect 19475 42653 19487 42687
rect 19429 42647 19487 42653
rect 20165 42687 20223 42693
rect 20165 42653 20177 42687
rect 20211 42653 20223 42687
rect 20165 42647 20223 42653
rect 14415 42588 15792 42616
rect 15856 42588 16252 42616
rect 14415 42585 14427 42588
rect 14369 42579 14427 42585
rect 13081 42551 13139 42557
rect 13081 42517 13093 42551
rect 13127 42517 13139 42551
rect 13081 42511 13139 42517
rect 13538 42508 13544 42560
rect 13596 42508 13602 42560
rect 13998 42508 14004 42560
rect 14056 42548 14062 42560
rect 14461 42551 14519 42557
rect 14461 42548 14473 42551
rect 14056 42520 14473 42548
rect 14056 42508 14062 42520
rect 14461 42517 14473 42520
rect 14507 42517 14519 42551
rect 14461 42511 14519 42517
rect 14642 42508 14648 42560
rect 14700 42508 14706 42560
rect 14918 42508 14924 42560
rect 14976 42508 14982 42560
rect 15010 42508 15016 42560
rect 15068 42548 15074 42560
rect 15197 42551 15255 42557
rect 15197 42548 15209 42551
rect 15068 42520 15209 42548
rect 15068 42508 15074 42520
rect 15197 42517 15209 42520
rect 15243 42517 15255 42551
rect 15197 42511 15255 42517
rect 15470 42508 15476 42560
rect 15528 42508 15534 42560
rect 15764 42557 15792 42588
rect 16224 42560 16252 42588
rect 16390 42576 16396 42628
rect 16448 42576 16454 42628
rect 16942 42576 16948 42628
rect 17000 42576 17006 42628
rect 17494 42576 17500 42628
rect 17552 42576 17558 42628
rect 18049 42619 18107 42625
rect 18049 42616 18061 42619
rect 17788 42588 18061 42616
rect 17788 42560 17816 42588
rect 18049 42585 18061 42588
rect 18095 42585 18107 42619
rect 18049 42579 18107 42585
rect 18601 42619 18659 42625
rect 18601 42585 18613 42619
rect 18647 42616 18659 42619
rect 18874 42616 18880 42628
rect 18647 42588 18880 42616
rect 18647 42585 18659 42588
rect 18601 42579 18659 42585
rect 18874 42576 18880 42588
rect 18932 42576 18938 42628
rect 19613 42619 19671 42625
rect 19613 42585 19625 42619
rect 19659 42616 19671 42619
rect 19886 42616 19892 42628
rect 19659 42588 19892 42616
rect 19659 42585 19671 42588
rect 19613 42579 19671 42585
rect 19886 42576 19892 42588
rect 19944 42576 19950 42628
rect 15749 42551 15807 42557
rect 15749 42517 15761 42551
rect 15795 42517 15807 42551
rect 15749 42511 15807 42517
rect 16025 42551 16083 42557
rect 16025 42517 16037 42551
rect 16071 42548 16083 42551
rect 16114 42548 16120 42560
rect 16071 42520 16120 42548
rect 16071 42517 16083 42520
rect 16025 42511 16083 42517
rect 16114 42508 16120 42520
rect 16172 42508 16178 42560
rect 16206 42508 16212 42560
rect 16264 42508 16270 42560
rect 17770 42508 17776 42560
rect 17828 42508 17834 42560
rect 18322 42508 18328 42560
rect 18380 42508 18386 42560
rect 18690 42508 18696 42560
rect 18748 42548 18754 42560
rect 20257 42551 20315 42557
rect 20257 42548 20269 42551
rect 18748 42520 20269 42548
rect 18748 42508 18754 42520
rect 20257 42517 20269 42520
rect 20303 42517 20315 42551
rect 20257 42511 20315 42517
rect 1104 42458 21043 42480
rect 1104 42406 5894 42458
rect 5946 42406 5958 42458
rect 6010 42406 6022 42458
rect 6074 42406 6086 42458
rect 6138 42406 6150 42458
rect 6202 42406 10839 42458
rect 10891 42406 10903 42458
rect 10955 42406 10967 42458
rect 11019 42406 11031 42458
rect 11083 42406 11095 42458
rect 11147 42406 15784 42458
rect 15836 42406 15848 42458
rect 15900 42406 15912 42458
rect 15964 42406 15976 42458
rect 16028 42406 16040 42458
rect 16092 42406 20729 42458
rect 20781 42406 20793 42458
rect 20845 42406 20857 42458
rect 20909 42406 20921 42458
rect 20973 42406 20985 42458
rect 21037 42406 21043 42458
rect 1104 42384 21043 42406
rect 1486 42304 1492 42356
rect 1544 42304 1550 42356
rect 1949 42347 2007 42353
rect 1949 42313 1961 42347
rect 1995 42344 2007 42347
rect 2498 42344 2504 42356
rect 1995 42316 2504 42344
rect 1995 42313 2007 42316
rect 1949 42307 2007 42313
rect 2498 42304 2504 42316
rect 2556 42304 2562 42356
rect 2590 42304 2596 42356
rect 2648 42304 2654 42356
rect 3145 42347 3203 42353
rect 3145 42313 3157 42347
rect 3191 42313 3203 42347
rect 3145 42307 3203 42313
rect 3513 42347 3571 42353
rect 3513 42313 3525 42347
rect 3559 42344 3571 42347
rect 4062 42344 4068 42356
rect 3559 42316 4068 42344
rect 3559 42313 3571 42316
rect 3513 42307 3571 42313
rect 1504 42276 1532 42304
rect 2317 42279 2375 42285
rect 2317 42276 2329 42279
rect 1504 42248 2329 42276
rect 2317 42245 2329 42248
rect 2363 42245 2375 42279
rect 3160 42276 3188 42307
rect 4062 42304 4068 42316
rect 4120 42304 4126 42356
rect 4157 42347 4215 42353
rect 4157 42313 4169 42347
rect 4203 42344 4215 42347
rect 4798 42344 4804 42356
rect 4203 42316 4804 42344
rect 4203 42313 4215 42316
rect 4157 42307 4215 42313
rect 4798 42304 4804 42316
rect 4856 42304 4862 42356
rect 5077 42347 5135 42353
rect 5077 42313 5089 42347
rect 5123 42344 5135 42347
rect 5166 42344 5172 42356
rect 5123 42316 5172 42344
rect 5123 42313 5135 42316
rect 5077 42307 5135 42313
rect 5166 42304 5172 42316
rect 5224 42304 5230 42356
rect 5629 42347 5687 42353
rect 5629 42313 5641 42347
rect 5675 42344 5687 42347
rect 5718 42344 5724 42356
rect 5675 42316 5724 42344
rect 5675 42313 5687 42316
rect 5629 42307 5687 42313
rect 5718 42304 5724 42316
rect 5776 42304 5782 42356
rect 5997 42347 6055 42353
rect 5997 42313 6009 42347
rect 6043 42313 6055 42347
rect 5997 42307 6055 42313
rect 6733 42347 6791 42353
rect 6733 42313 6745 42347
rect 6779 42344 6791 42347
rect 6822 42344 6828 42356
rect 6779 42316 6828 42344
rect 6779 42313 6791 42316
rect 6733 42307 6791 42313
rect 3602 42276 3608 42288
rect 3160 42248 3608 42276
rect 2317 42239 2375 42245
rect 3602 42236 3608 42248
rect 3660 42236 3666 42288
rect 4338 42276 4344 42288
rect 3896 42248 4344 42276
rect 934 42168 940 42220
rect 992 42208 998 42220
rect 2133 42211 2191 42217
rect 2133 42208 2145 42211
rect 992 42180 2145 42208
rect 992 42168 998 42180
rect 2133 42177 2145 42180
rect 2179 42177 2191 42211
rect 2133 42171 2191 42177
rect 2961 42211 3019 42217
rect 2961 42177 2973 42211
rect 3007 42208 3019 42211
rect 3234 42208 3240 42220
rect 3007 42180 3240 42208
rect 3007 42177 3019 42180
rect 2961 42171 3019 42177
rect 3234 42168 3240 42180
rect 3292 42168 3298 42220
rect 3326 42168 3332 42220
rect 3384 42168 3390 42220
rect 3896 42217 3924 42248
rect 4338 42236 4344 42248
rect 4396 42236 4402 42288
rect 6012 42276 6040 42307
rect 6822 42304 6828 42316
rect 6880 42304 6886 42356
rect 7558 42304 7564 42356
rect 7616 42344 7622 42356
rect 7837 42347 7895 42353
rect 7837 42344 7849 42347
rect 7616 42316 7849 42344
rect 7616 42304 7622 42316
rect 7837 42313 7849 42316
rect 7883 42313 7895 42347
rect 7837 42307 7895 42313
rect 8018 42304 8024 42356
rect 8076 42304 8082 42356
rect 8110 42304 8116 42356
rect 8168 42344 8174 42356
rect 8389 42347 8447 42353
rect 8389 42344 8401 42347
rect 8168 42316 8401 42344
rect 8168 42304 8174 42316
rect 8389 42313 8401 42316
rect 8435 42313 8447 42347
rect 8389 42307 8447 42313
rect 8938 42304 8944 42356
rect 8996 42304 9002 42356
rect 9217 42347 9275 42353
rect 9217 42313 9229 42347
rect 9263 42313 9275 42347
rect 9217 42307 9275 42313
rect 7745 42279 7803 42285
rect 7745 42276 7757 42279
rect 4448 42248 5948 42276
rect 6012 42248 7757 42276
rect 4448 42217 4476 42248
rect 3881 42211 3939 42217
rect 3881 42177 3893 42211
rect 3927 42177 3939 42211
rect 3881 42171 3939 42177
rect 3973 42211 4031 42217
rect 3973 42177 3985 42211
rect 4019 42177 4031 42211
rect 3973 42171 4031 42177
rect 4433 42211 4491 42217
rect 4433 42177 4445 42211
rect 4479 42177 4491 42211
rect 4433 42171 4491 42177
rect 1670 42100 1676 42152
rect 1728 42140 1734 42152
rect 2866 42140 2872 42152
rect 1728 42112 2872 42140
rect 1728 42100 1734 42112
rect 2866 42100 2872 42112
rect 2924 42100 2930 42152
rect 3988 42140 4016 42171
rect 4890 42168 4896 42220
rect 4948 42168 4954 42220
rect 5534 42168 5540 42220
rect 5592 42168 5598 42220
rect 4062 42140 4068 42152
rect 3068 42112 3924 42140
rect 3988 42112 4068 42140
rect 842 42032 848 42084
rect 900 42072 906 42084
rect 3068 42072 3096 42112
rect 900 42044 3096 42072
rect 900 42032 906 42044
rect 3694 42032 3700 42084
rect 3752 42032 3758 42084
rect 3896 42004 3924 42112
rect 4062 42100 4068 42112
rect 4120 42100 4126 42152
rect 4522 42100 4528 42152
rect 4580 42140 4586 42152
rect 4709 42143 4767 42149
rect 4709 42140 4721 42143
rect 4580 42112 4721 42140
rect 4580 42100 4586 42112
rect 4709 42109 4721 42112
rect 4755 42109 4767 42143
rect 4709 42103 4767 42109
rect 3970 42032 3976 42084
rect 4028 42072 4034 42084
rect 5920 42072 5948 42248
rect 7745 42245 7757 42248
rect 7791 42245 7803 42279
rect 8036 42276 8064 42304
rect 9232 42276 9260 42307
rect 9582 42304 9588 42356
rect 9640 42344 9646 42356
rect 10873 42347 10931 42353
rect 10873 42344 10885 42347
rect 9640 42316 10885 42344
rect 9640 42304 9646 42316
rect 10873 42313 10885 42316
rect 10919 42313 10931 42347
rect 12342 42344 12348 42356
rect 10873 42307 10931 42313
rect 10980 42316 12348 42344
rect 8036 42248 9260 42276
rect 7745 42239 7803 42245
rect 9766 42236 9772 42288
rect 9824 42276 9830 42288
rect 9824 42248 10732 42276
rect 9824 42236 9830 42248
rect 6181 42211 6239 42217
rect 6181 42177 6193 42211
rect 6227 42177 6239 42211
rect 6181 42171 6239 42177
rect 6196 42140 6224 42171
rect 6270 42168 6276 42220
rect 6328 42208 6334 42220
rect 6641 42211 6699 42217
rect 6641 42208 6653 42211
rect 6328 42180 6653 42208
rect 6328 42168 6334 42180
rect 6641 42177 6653 42180
rect 6687 42177 6699 42211
rect 6641 42171 6699 42177
rect 7098 42168 7104 42220
rect 7156 42168 7162 42220
rect 8202 42168 8208 42220
rect 8260 42168 8266 42220
rect 8846 42168 8852 42220
rect 8904 42168 8910 42220
rect 8938 42168 8944 42220
rect 8996 42208 9002 42220
rect 9125 42211 9183 42217
rect 9125 42208 9137 42211
rect 8996 42180 9137 42208
rect 8996 42168 9002 42180
rect 9125 42177 9137 42180
rect 9171 42177 9183 42211
rect 9125 42171 9183 42177
rect 9401 42211 9459 42217
rect 9401 42177 9413 42211
rect 9447 42177 9459 42211
rect 9401 42171 9459 42177
rect 6914 42140 6920 42152
rect 6196 42112 6920 42140
rect 6914 42100 6920 42112
rect 6972 42100 6978 42152
rect 7742 42100 7748 42152
rect 7800 42100 7806 42152
rect 9416 42140 9444 42171
rect 9490 42168 9496 42220
rect 9548 42208 9554 42220
rect 9677 42211 9735 42217
rect 9677 42208 9689 42211
rect 9548 42180 9689 42208
rect 9548 42168 9554 42180
rect 9677 42177 9689 42180
rect 9723 42177 9735 42211
rect 9677 42171 9735 42177
rect 10042 42168 10048 42220
rect 10100 42168 10106 42220
rect 10594 42168 10600 42220
rect 10652 42168 10658 42220
rect 10704 42217 10732 42248
rect 10689 42211 10747 42217
rect 10689 42177 10701 42211
rect 10735 42177 10747 42211
rect 10689 42171 10747 42177
rect 10980 42140 11008 42316
rect 12342 42304 12348 42316
rect 12400 42304 12406 42356
rect 12713 42347 12771 42353
rect 12713 42313 12725 42347
rect 12759 42344 12771 42347
rect 13446 42344 13452 42356
rect 12759 42316 13452 42344
rect 12759 42313 12771 42316
rect 12713 42307 12771 42313
rect 13446 42304 13452 42316
rect 13504 42304 13510 42356
rect 13538 42304 13544 42356
rect 13596 42304 13602 42356
rect 13722 42344 13728 42356
rect 13648 42316 13728 42344
rect 11606 42236 11612 42288
rect 11664 42276 11670 42288
rect 13556 42276 13584 42304
rect 11664 42248 12940 42276
rect 11664 42236 11670 42248
rect 11330 42168 11336 42220
rect 11388 42168 11394 42220
rect 12342 42168 12348 42220
rect 12400 42168 12406 42220
rect 12912 42217 12940 42248
rect 13004 42248 13584 42276
rect 13004 42217 13032 42248
rect 12621 42211 12679 42217
rect 12621 42177 12633 42211
rect 12667 42177 12679 42211
rect 12621 42171 12679 42177
rect 12897 42211 12955 42217
rect 12897 42177 12909 42211
rect 12943 42177 12955 42211
rect 12897 42171 12955 42177
rect 12989 42211 13047 42217
rect 12989 42177 13001 42211
rect 13035 42177 13047 42211
rect 12989 42171 13047 42177
rect 13357 42211 13415 42217
rect 13357 42177 13369 42211
rect 13403 42208 13415 42211
rect 13648 42208 13676 42316
rect 13722 42304 13728 42316
rect 13780 42304 13786 42356
rect 14642 42304 14648 42356
rect 14700 42304 14706 42356
rect 15286 42344 15292 42356
rect 14752 42316 15292 42344
rect 14660 42276 14688 42304
rect 13740 42248 14688 42276
rect 13740 42217 13768 42248
rect 13403 42180 13676 42208
rect 13725 42211 13783 42217
rect 13403 42177 13415 42180
rect 13357 42171 13415 42177
rect 13725 42177 13737 42211
rect 13771 42177 13783 42211
rect 13725 42171 13783 42177
rect 14185 42211 14243 42217
rect 14185 42177 14197 42211
rect 14231 42177 14243 42211
rect 14185 42171 14243 42177
rect 8680 42112 9444 42140
rect 9508 42112 11008 42140
rect 12636 42140 12664 42171
rect 13630 42140 13636 42152
rect 12636 42112 13636 42140
rect 7006 42072 7012 42084
rect 4028 42044 5304 42072
rect 5920 42044 7012 42072
rect 4028 42032 4034 42044
rect 5166 42004 5172 42016
rect 3896 41976 5172 42004
rect 5166 41964 5172 41976
rect 5224 41964 5230 42016
rect 5276 42004 5304 42044
rect 7006 42032 7012 42044
rect 7064 42032 7070 42084
rect 7285 42075 7343 42081
rect 7285 42041 7297 42075
rect 7331 42072 7343 42075
rect 7760 42072 7788 42100
rect 8680 42081 8708 42112
rect 7331 42044 7788 42072
rect 8665 42075 8723 42081
rect 7331 42041 7343 42044
rect 7285 42035 7343 42041
rect 8665 42041 8677 42075
rect 8711 42041 8723 42075
rect 9508 42072 9536 42112
rect 13630 42100 13636 42112
rect 13688 42100 13694 42152
rect 14200 42140 14228 42171
rect 14458 42168 14464 42220
rect 14516 42168 14522 42220
rect 14642 42168 14648 42220
rect 14700 42208 14706 42220
rect 14752 42208 14780 42316
rect 15286 42304 15292 42316
rect 15344 42304 15350 42356
rect 15470 42304 15476 42356
rect 15528 42304 15534 42356
rect 15933 42347 15991 42353
rect 15933 42344 15945 42347
rect 15672 42316 15945 42344
rect 15488 42276 15516 42304
rect 15672 42285 15700 42316
rect 15933 42313 15945 42316
rect 15979 42313 15991 42347
rect 15933 42307 15991 42313
rect 16114 42304 16120 42356
rect 16172 42304 16178 42356
rect 16206 42304 16212 42356
rect 16264 42344 16270 42356
rect 16669 42347 16727 42353
rect 16669 42344 16681 42347
rect 16264 42316 16681 42344
rect 16264 42304 16270 42316
rect 16669 42313 16681 42316
rect 16715 42313 16727 42347
rect 18966 42344 18972 42356
rect 16669 42307 16727 42313
rect 18064 42316 18972 42344
rect 14844 42248 15516 42276
rect 15657 42279 15715 42285
rect 14844 42217 14872 42248
rect 15657 42245 15669 42279
rect 15703 42245 15715 42279
rect 16132 42276 16160 42304
rect 15657 42239 15715 42245
rect 15764 42248 16160 42276
rect 14700 42180 14780 42208
rect 14829 42211 14887 42217
rect 14700 42168 14706 42180
rect 14829 42177 14841 42211
rect 14875 42177 14887 42211
rect 14829 42171 14887 42177
rect 14918 42168 14924 42220
rect 14976 42168 14982 42220
rect 15197 42211 15255 42217
rect 15197 42177 15209 42211
rect 15243 42208 15255 42211
rect 15764 42208 15792 42248
rect 16482 42236 16488 42288
rect 16540 42276 16546 42288
rect 18064 42285 18092 42316
rect 18966 42304 18972 42316
rect 19024 42304 19030 42356
rect 20257 42347 20315 42353
rect 20257 42313 20269 42347
rect 20303 42344 20315 42347
rect 21174 42344 21180 42356
rect 20303 42316 21180 42344
rect 20303 42313 20315 42316
rect 20257 42307 20315 42313
rect 21174 42304 21180 42316
rect 21232 42304 21238 42356
rect 18049 42279 18107 42285
rect 16540 42248 17816 42276
rect 16540 42236 16546 42248
rect 15243 42180 15792 42208
rect 16117 42211 16175 42217
rect 15243 42177 15255 42180
rect 15197 42171 15255 42177
rect 16117 42177 16129 42211
rect 16163 42177 16175 42211
rect 16117 42171 16175 42177
rect 14936 42140 14964 42168
rect 16132 42140 16160 42171
rect 16298 42168 16304 42220
rect 16356 42208 16362 42220
rect 16393 42211 16451 42217
rect 16393 42208 16405 42211
rect 16356 42180 16405 42208
rect 16356 42168 16362 42180
rect 16393 42177 16405 42180
rect 16439 42177 16451 42211
rect 16393 42171 16451 42177
rect 16574 42168 16580 42220
rect 16632 42208 16638 42220
rect 16853 42211 16911 42217
rect 16853 42208 16865 42211
rect 16632 42180 16865 42208
rect 16632 42168 16638 42180
rect 16853 42177 16865 42180
rect 16899 42177 16911 42211
rect 16853 42171 16911 42177
rect 17126 42168 17132 42220
rect 17184 42168 17190 42220
rect 17310 42168 17316 42220
rect 17368 42208 17374 42220
rect 17681 42211 17739 42217
rect 17681 42208 17693 42211
rect 17368 42180 17693 42208
rect 17368 42168 17374 42180
rect 17681 42177 17693 42180
rect 17727 42177 17739 42211
rect 17788 42208 17816 42248
rect 18049 42245 18061 42279
rect 18095 42245 18107 42279
rect 18049 42239 18107 42245
rect 18230 42236 18236 42288
rect 18288 42236 18294 42288
rect 18598 42236 18604 42288
rect 18656 42236 18662 42288
rect 18877 42211 18935 42217
rect 18877 42208 18889 42211
rect 17788 42180 18889 42208
rect 17681 42171 17739 42177
rect 18877 42177 18889 42180
rect 18923 42177 18935 42211
rect 18877 42171 18935 42177
rect 19061 42211 19119 42217
rect 19061 42177 19073 42211
rect 19107 42177 19119 42211
rect 19061 42171 19119 42177
rect 14200 42112 14964 42140
rect 15212 42112 16160 42140
rect 8665 42035 8723 42041
rect 8772 42044 9536 42072
rect 8772 42004 8800 42044
rect 10318 42032 10324 42084
rect 10376 42072 10382 42084
rect 12437 42075 12495 42081
rect 10376 42044 11192 42072
rect 10376 42032 10382 42044
rect 5276 41976 8800 42004
rect 9490 41964 9496 42016
rect 9548 41964 9554 42016
rect 9766 41964 9772 42016
rect 9824 42004 9830 42016
rect 10229 42007 10287 42013
rect 10229 42004 10241 42007
rect 9824 41976 10241 42004
rect 9824 41964 9830 41976
rect 10229 41973 10241 41976
rect 10275 41973 10287 42007
rect 10229 41967 10287 41973
rect 10410 41964 10416 42016
rect 10468 41964 10474 42016
rect 11164 42013 11192 42044
rect 12437 42041 12449 42075
rect 12483 42072 12495 42075
rect 15212 42072 15240 42112
rect 17862 42100 17868 42152
rect 17920 42140 17926 42152
rect 19076 42140 19104 42171
rect 19610 42168 19616 42220
rect 19668 42208 19674 42220
rect 19797 42211 19855 42217
rect 19797 42208 19809 42211
rect 19668 42180 19809 42208
rect 19668 42168 19674 42180
rect 19797 42177 19809 42180
rect 19843 42177 19855 42211
rect 19797 42171 19855 42177
rect 19981 42211 20039 42217
rect 19981 42177 19993 42211
rect 20027 42208 20039 42211
rect 20622 42208 20628 42220
rect 20027 42180 20628 42208
rect 20027 42177 20039 42180
rect 19981 42171 20039 42177
rect 20622 42168 20628 42180
rect 20680 42168 20686 42220
rect 17920 42112 19104 42140
rect 17920 42100 17926 42112
rect 19150 42100 19156 42152
rect 19208 42100 19214 42152
rect 16209 42075 16267 42081
rect 16209 42072 16221 42075
rect 12483 42044 15240 42072
rect 15304 42044 16221 42072
rect 12483 42041 12495 42044
rect 12437 42035 12495 42041
rect 15304 42016 15332 42044
rect 16209 42041 16221 42044
rect 16255 42041 16267 42075
rect 18693 42075 18751 42081
rect 18693 42072 18705 42075
rect 16209 42035 16267 42041
rect 16776 42044 18705 42072
rect 11149 42007 11207 42013
rect 11149 41973 11161 42007
rect 11195 41973 11207 42007
rect 11149 41967 11207 41973
rect 12158 41964 12164 42016
rect 12216 41964 12222 42016
rect 13170 41964 13176 42016
rect 13228 41964 13234 42016
rect 13262 41964 13268 42016
rect 13320 42004 13326 42016
rect 13541 42007 13599 42013
rect 13541 42004 13553 42007
rect 13320 41976 13553 42004
rect 13320 41964 13326 41976
rect 13541 41973 13553 41976
rect 13587 41973 13599 42007
rect 13541 41967 13599 41973
rect 13906 41964 13912 42016
rect 13964 41964 13970 42016
rect 14274 41964 14280 42016
rect 14332 41964 14338 42016
rect 14366 41964 14372 42016
rect 14424 42004 14430 42016
rect 14645 42007 14703 42013
rect 14645 42004 14657 42007
rect 14424 41976 14657 42004
rect 14424 41964 14430 41976
rect 14645 41973 14657 41976
rect 14691 41973 14703 42007
rect 14645 41967 14703 41973
rect 14826 41964 14832 42016
rect 14884 42004 14890 42016
rect 15013 42007 15071 42013
rect 15013 42004 15025 42007
rect 14884 41976 15025 42004
rect 14884 41964 14890 41976
rect 15013 41973 15025 41976
rect 15059 41973 15071 42007
rect 15013 41967 15071 41973
rect 15286 41964 15292 42016
rect 15344 41964 15350 42016
rect 15378 41964 15384 42016
rect 15436 41964 15442 42016
rect 15470 41964 15476 42016
rect 15528 42004 15534 42016
rect 15749 42007 15807 42013
rect 15749 42004 15761 42007
rect 15528 41976 15761 42004
rect 15528 41964 15534 41976
rect 15749 41973 15761 41976
rect 15795 41973 15807 42007
rect 15749 41967 15807 41973
rect 15838 41964 15844 42016
rect 15896 42004 15902 42016
rect 16776 42004 16804 42044
rect 18693 42041 18705 42044
rect 18739 42041 18751 42075
rect 18693 42035 18751 42041
rect 15896 41976 16804 42004
rect 17405 42007 17463 42013
rect 15896 41964 15902 41976
rect 17405 41973 17417 42007
rect 17451 42004 17463 42007
rect 19168 42004 19196 42100
rect 17451 41976 19196 42004
rect 17451 41973 17463 41976
rect 17405 41967 17463 41973
rect 19334 41964 19340 42016
rect 19392 41964 19398 42016
rect 19613 42007 19671 42013
rect 19613 41973 19625 42007
rect 19659 42004 19671 42007
rect 19886 42004 19892 42016
rect 19659 41976 19892 42004
rect 19659 41973 19671 41976
rect 19613 41967 19671 41973
rect 19886 41964 19892 41976
rect 19944 41964 19950 42016
rect 1104 41914 20884 41936
rect 1104 41862 3422 41914
rect 3474 41862 3486 41914
rect 3538 41862 3550 41914
rect 3602 41862 3614 41914
rect 3666 41862 3678 41914
rect 3730 41862 8367 41914
rect 8419 41862 8431 41914
rect 8483 41862 8495 41914
rect 8547 41862 8559 41914
rect 8611 41862 8623 41914
rect 8675 41862 13312 41914
rect 13364 41862 13376 41914
rect 13428 41862 13440 41914
rect 13492 41862 13504 41914
rect 13556 41862 13568 41914
rect 13620 41862 18257 41914
rect 18309 41862 18321 41914
rect 18373 41862 18385 41914
rect 18437 41862 18449 41914
rect 18501 41862 18513 41914
rect 18565 41862 20884 41914
rect 1104 41840 20884 41862
rect 2130 41760 2136 41812
rect 2188 41760 2194 41812
rect 2317 41803 2375 41809
rect 2317 41769 2329 41803
rect 2363 41800 2375 41803
rect 2682 41800 2688 41812
rect 2363 41772 2688 41800
rect 2363 41769 2375 41772
rect 2317 41763 2375 41769
rect 2682 41760 2688 41772
rect 2740 41760 2746 41812
rect 2869 41803 2927 41809
rect 2869 41769 2881 41803
rect 2915 41800 2927 41803
rect 3050 41800 3056 41812
rect 2915 41772 3056 41800
rect 2915 41769 2927 41772
rect 2869 41763 2927 41769
rect 3050 41760 3056 41772
rect 3108 41760 3114 41812
rect 3142 41760 3148 41812
rect 3200 41760 3206 41812
rect 3234 41760 3240 41812
rect 3292 41800 3298 41812
rect 3421 41803 3479 41809
rect 3421 41800 3433 41803
rect 3292 41772 3433 41800
rect 3292 41760 3298 41772
rect 3421 41769 3433 41772
rect 3467 41769 3479 41803
rect 3970 41800 3976 41812
rect 3421 41763 3479 41769
rect 3528 41772 3976 41800
rect 2148 41732 2176 41760
rect 2593 41735 2651 41741
rect 2593 41732 2605 41735
rect 2148 41704 2605 41732
rect 2593 41701 2605 41704
rect 2639 41701 2651 41735
rect 2593 41695 2651 41701
rect 2958 41692 2964 41744
rect 3016 41732 3022 41744
rect 3528 41732 3556 41772
rect 3970 41760 3976 41772
rect 4028 41760 4034 41812
rect 4154 41760 4160 41812
rect 4212 41760 4218 41812
rect 4246 41760 4252 41812
rect 4304 41760 4310 41812
rect 4709 41803 4767 41809
rect 4709 41769 4721 41803
rect 4755 41800 4767 41803
rect 5534 41800 5540 41812
rect 4755 41772 5540 41800
rect 4755 41769 4767 41772
rect 4709 41763 4767 41769
rect 5534 41760 5540 41772
rect 5592 41760 5598 41812
rect 5997 41803 6055 41809
rect 5997 41769 6009 41803
rect 6043 41800 6055 41803
rect 6638 41800 6644 41812
rect 6043 41772 6644 41800
rect 6043 41769 6055 41772
rect 5997 41763 6055 41769
rect 6638 41760 6644 41772
rect 6696 41760 6702 41812
rect 7006 41760 7012 41812
rect 7064 41760 7070 41812
rect 7098 41760 7104 41812
rect 7156 41800 7162 41812
rect 7929 41803 7987 41809
rect 7929 41800 7941 41803
rect 7156 41772 7941 41800
rect 7156 41760 7162 41772
rect 7929 41769 7941 41772
rect 7975 41769 7987 41803
rect 7929 41763 7987 41769
rect 8202 41760 8208 41812
rect 8260 41800 8266 41812
rect 8297 41803 8355 41809
rect 8297 41800 8309 41803
rect 8260 41772 8309 41800
rect 8260 41760 8266 41772
rect 8297 41769 8309 41772
rect 8343 41769 8355 41803
rect 9490 41800 9496 41812
rect 8297 41763 8355 41769
rect 8404 41772 9496 41800
rect 3016 41704 3556 41732
rect 3881 41735 3939 41741
rect 3016 41692 3022 41704
rect 3881 41701 3893 41735
rect 3927 41732 3939 41735
rect 4264 41732 4292 41760
rect 3927 41704 4292 41732
rect 5261 41735 5319 41741
rect 3927 41701 3939 41704
rect 3881 41695 3939 41701
rect 5261 41701 5273 41735
rect 5307 41701 5319 41735
rect 5261 41695 5319 41701
rect 14 41624 20 41676
rect 72 41664 78 41676
rect 5276 41664 5304 41695
rect 5442 41692 5448 41744
rect 5500 41732 5506 41744
rect 6733 41735 6791 41741
rect 6733 41732 6745 41735
rect 5500 41704 6745 41732
rect 5500 41692 5506 41704
rect 6733 41701 6745 41704
rect 6779 41701 6791 41735
rect 6733 41695 6791 41701
rect 72 41636 4108 41664
rect 72 41624 78 41636
rect 2498 41556 2504 41608
rect 2556 41556 2562 41608
rect 2777 41599 2835 41605
rect 2777 41565 2789 41599
rect 2823 41565 2835 41599
rect 2777 41559 2835 41565
rect 2038 41488 2044 41540
rect 2096 41528 2102 41540
rect 2792 41528 2820 41559
rect 3050 41556 3056 41608
rect 3108 41556 3114 41608
rect 3329 41599 3387 41605
rect 3329 41565 3341 41599
rect 3375 41565 3387 41599
rect 3329 41559 3387 41565
rect 3605 41599 3663 41605
rect 3605 41565 3617 41599
rect 3651 41596 3663 41599
rect 3878 41596 3884 41608
rect 3651 41568 3884 41596
rect 3651 41565 3663 41568
rect 3605 41559 3663 41565
rect 3344 41528 3372 41559
rect 3878 41556 3884 41568
rect 3936 41556 3942 41608
rect 4080 41605 4108 41636
rect 4356 41636 5304 41664
rect 5368 41636 5856 41664
rect 4356 41605 4384 41636
rect 4065 41599 4123 41605
rect 4065 41565 4077 41599
rect 4111 41565 4123 41599
rect 4065 41559 4123 41565
rect 4341 41599 4399 41605
rect 4341 41565 4353 41599
rect 4387 41565 4399 41599
rect 4341 41559 4399 41565
rect 4617 41599 4675 41605
rect 4617 41565 4629 41599
rect 4663 41596 4675 41599
rect 4706 41596 4712 41608
rect 4663 41568 4712 41596
rect 4663 41565 4675 41568
rect 4617 41559 4675 41565
rect 4706 41556 4712 41568
rect 4764 41556 4770 41608
rect 4893 41599 4951 41605
rect 4893 41565 4905 41599
rect 4939 41596 4951 41599
rect 5074 41596 5080 41608
rect 4939 41568 5080 41596
rect 4939 41565 4951 41568
rect 4893 41559 4951 41565
rect 5074 41556 5080 41568
rect 5132 41556 5138 41608
rect 5166 41556 5172 41608
rect 5224 41556 5230 41608
rect 5368 41596 5396 41636
rect 5276 41568 5396 41596
rect 5276 41528 5304 41568
rect 5442 41556 5448 41608
rect 5500 41556 5506 41608
rect 5534 41556 5540 41608
rect 5592 41596 5598 41608
rect 5828 41605 5856 41636
rect 5721 41599 5779 41605
rect 5721 41596 5733 41599
rect 5592 41568 5733 41596
rect 5592 41556 5598 41568
rect 5721 41565 5733 41568
rect 5767 41565 5779 41599
rect 5721 41559 5779 41565
rect 5813 41599 5871 41605
rect 5813 41565 5825 41599
rect 5859 41565 5871 41599
rect 6917 41599 6975 41605
rect 6917 41596 6929 41599
rect 5813 41559 5871 41565
rect 6380 41568 6929 41596
rect 2096 41500 2820 41528
rect 3068 41500 3372 41528
rect 4448 41500 5304 41528
rect 2096 41488 2102 41500
rect 474 41420 480 41472
rect 532 41460 538 41472
rect 3068 41460 3096 41500
rect 4448 41469 4476 41500
rect 532 41432 3096 41460
rect 4433 41463 4491 41469
rect 532 41420 538 41432
rect 4433 41429 4445 41463
rect 4479 41429 4491 41463
rect 4433 41423 4491 41429
rect 4985 41463 5043 41469
rect 4985 41429 4997 41463
rect 5031 41460 5043 41463
rect 5166 41460 5172 41472
rect 5031 41432 5172 41460
rect 5031 41429 5043 41432
rect 4985 41423 5043 41429
rect 5166 41420 5172 41432
rect 5224 41420 5230 41472
rect 5534 41420 5540 41472
rect 5592 41420 5598 41472
rect 5626 41420 5632 41472
rect 5684 41460 5690 41472
rect 6380 41469 6408 41568
rect 6917 41565 6929 41568
rect 6963 41565 6975 41599
rect 6917 41559 6975 41565
rect 7024 41528 7052 41760
rect 7190 41692 7196 41744
rect 7248 41732 7254 41744
rect 7285 41735 7343 41741
rect 7285 41732 7297 41735
rect 7248 41704 7297 41732
rect 7248 41692 7254 41704
rect 7285 41701 7297 41704
rect 7331 41701 7343 41735
rect 7285 41695 7343 41701
rect 7190 41556 7196 41608
rect 7248 41556 7254 41608
rect 7469 41599 7527 41605
rect 7469 41565 7481 41599
rect 7515 41596 7527 41599
rect 7742 41596 7748 41608
rect 7515 41568 7748 41596
rect 7515 41565 7527 41568
rect 7469 41559 7527 41565
rect 7742 41556 7748 41568
rect 7800 41556 7806 41608
rect 8113 41599 8171 41605
rect 8113 41565 8125 41599
rect 8159 41596 8171 41599
rect 8404 41596 8432 41772
rect 9490 41760 9496 41772
rect 9548 41760 9554 41812
rect 12618 41800 12624 41812
rect 9600 41772 12624 41800
rect 8573 41735 8631 41741
rect 8573 41701 8585 41735
rect 8619 41732 8631 41735
rect 8754 41732 8760 41744
rect 8619 41704 8760 41732
rect 8619 41701 8631 41704
rect 8573 41695 8631 41701
rect 8754 41692 8760 41704
rect 8812 41692 8818 41744
rect 8941 41735 8999 41741
rect 8941 41701 8953 41735
rect 8987 41701 8999 41735
rect 8941 41695 8999 41701
rect 8956 41664 8984 41695
rect 8496 41636 8984 41664
rect 8496 41605 8524 41636
rect 8159 41568 8432 41596
rect 8481 41599 8539 41605
rect 8159 41565 8171 41568
rect 8113 41559 8171 41565
rect 8481 41565 8493 41599
rect 8527 41565 8539 41599
rect 8481 41559 8539 41565
rect 8754 41556 8760 41608
rect 8812 41556 8818 41608
rect 9122 41556 9128 41608
rect 9180 41556 9186 41608
rect 9600 41528 9628 41772
rect 12618 41760 12624 41772
rect 12676 41760 12682 41812
rect 13173 41803 13231 41809
rect 13173 41769 13185 41803
rect 13219 41800 13231 41803
rect 14090 41800 14096 41812
rect 13219 41772 14096 41800
rect 13219 41769 13231 41772
rect 13173 41763 13231 41769
rect 14090 41760 14096 41772
rect 14148 41760 14154 41812
rect 15010 41760 15016 41812
rect 15068 41760 15074 41812
rect 17681 41803 17739 41809
rect 17681 41800 17693 41803
rect 15488 41772 17693 41800
rect 12434 41692 12440 41744
rect 12492 41732 12498 41744
rect 13449 41735 13507 41741
rect 13449 41732 13461 41735
rect 12492 41704 13461 41732
rect 12492 41692 12498 41704
rect 13449 41701 13461 41704
rect 13495 41701 13507 41735
rect 13449 41695 13507 41701
rect 13725 41735 13783 41741
rect 13725 41701 13737 41735
rect 13771 41732 13783 41735
rect 13814 41732 13820 41744
rect 13771 41704 13820 41732
rect 13771 41701 13783 41704
rect 13725 41695 13783 41701
rect 13814 41692 13820 41704
rect 13872 41692 13878 41744
rect 14182 41732 14188 41744
rect 13924 41704 14188 41732
rect 13357 41599 13415 41605
rect 13357 41565 13369 41599
rect 13403 41596 13415 41599
rect 13538 41596 13544 41608
rect 13403 41568 13544 41596
rect 13403 41565 13415 41568
rect 13357 41559 13415 41565
rect 13538 41556 13544 41568
rect 13596 41556 13602 41608
rect 13630 41556 13636 41608
rect 13688 41556 13694 41608
rect 13924 41605 13952 41704
rect 14182 41692 14188 41704
rect 14240 41692 14246 41744
rect 14918 41732 14924 41744
rect 14292 41704 14924 41732
rect 14292 41664 14320 41704
rect 14918 41692 14924 41704
rect 14976 41692 14982 41744
rect 15028 41664 15056 41760
rect 15488 41664 15516 41772
rect 17681 41769 17693 41772
rect 17727 41769 17739 41803
rect 17681 41763 17739 41769
rect 18417 41803 18475 41809
rect 18417 41769 18429 41803
rect 18463 41800 18475 41803
rect 18782 41800 18788 41812
rect 18463 41772 18788 41800
rect 18463 41769 18475 41772
rect 18417 41763 18475 41769
rect 18782 41760 18788 41772
rect 18840 41760 18846 41812
rect 18969 41803 19027 41809
rect 18969 41769 18981 41803
rect 19015 41800 19027 41803
rect 19426 41800 19432 41812
rect 19015 41772 19432 41800
rect 19015 41769 19027 41772
rect 18969 41763 19027 41769
rect 19426 41760 19432 41772
rect 19484 41760 19490 41812
rect 15657 41735 15715 41741
rect 15657 41701 15669 41735
rect 15703 41732 15715 41735
rect 15746 41732 15752 41744
rect 15703 41704 15752 41732
rect 15703 41701 15715 41704
rect 15657 41695 15715 41701
rect 15746 41692 15752 41704
rect 15804 41692 15810 41744
rect 16574 41692 16580 41744
rect 16632 41732 16638 41744
rect 17129 41735 17187 41741
rect 17129 41732 17141 41735
rect 16632 41704 17141 41732
rect 16632 41692 16638 41704
rect 17129 41701 17141 41704
rect 17175 41701 17187 41735
rect 17129 41695 17187 41701
rect 17218 41692 17224 41744
rect 17276 41732 17282 41744
rect 18230 41732 18236 41744
rect 17276 41704 18236 41732
rect 17276 41692 17282 41704
rect 18230 41692 18236 41704
rect 18288 41692 18294 41744
rect 19705 41667 19763 41673
rect 14016 41636 14320 41664
rect 14568 41636 15056 41664
rect 15120 41636 15516 41664
rect 16040 41636 19656 41664
rect 13909 41599 13967 41605
rect 13909 41565 13921 41599
rect 13955 41565 13967 41599
rect 13909 41559 13967 41565
rect 7024 41500 9628 41528
rect 9950 41488 9956 41540
rect 10008 41528 10014 41540
rect 10226 41528 10232 41540
rect 10008 41500 10232 41528
rect 10008 41488 10014 41500
rect 10226 41488 10232 41500
rect 10284 41488 10290 41540
rect 11698 41488 11704 41540
rect 11756 41528 11762 41540
rect 12342 41528 12348 41540
rect 11756 41500 12348 41528
rect 11756 41488 11762 41500
rect 12342 41488 12348 41500
rect 12400 41488 12406 41540
rect 12802 41488 12808 41540
rect 12860 41528 12866 41540
rect 14016 41528 14044 41636
rect 14185 41599 14243 41605
rect 14185 41565 14197 41599
rect 14231 41592 14243 41599
rect 14568 41596 14596 41636
rect 15120 41605 15148 41636
rect 14353 41592 14596 41596
rect 14231 41568 14596 41592
rect 14645 41599 14703 41605
rect 14231 41565 14381 41568
rect 14185 41564 14381 41565
rect 14645 41565 14657 41599
rect 14691 41596 14703 41599
rect 15105 41599 15163 41605
rect 14691 41568 15056 41596
rect 14691 41565 14703 41568
rect 14185 41559 14243 41564
rect 14645 41559 14703 41565
rect 12860 41500 14044 41528
rect 12860 41488 12866 41500
rect 6365 41463 6423 41469
rect 6365 41460 6377 41463
rect 5684 41432 6377 41460
rect 5684 41420 5690 41432
rect 6365 41429 6377 41432
rect 6411 41429 6423 41463
rect 6365 41423 6423 41429
rect 7006 41420 7012 41472
rect 7064 41420 7070 41472
rect 14277 41463 14335 41469
rect 14277 41429 14289 41463
rect 14323 41460 14335 41463
rect 14458 41460 14464 41472
rect 14323 41432 14464 41460
rect 14323 41429 14335 41432
rect 14277 41423 14335 41429
rect 14458 41420 14464 41432
rect 14516 41420 14522 41472
rect 14826 41420 14832 41472
rect 14884 41420 14890 41472
rect 15028 41460 15056 41568
rect 15105 41565 15117 41599
rect 15151 41565 15163 41599
rect 15105 41559 15163 41565
rect 15289 41599 15347 41605
rect 15289 41565 15301 41599
rect 15335 41565 15347 41599
rect 15289 41559 15347 41565
rect 15565 41599 15623 41605
rect 15565 41565 15577 41599
rect 15611 41596 15623 41599
rect 15654 41596 15660 41608
rect 15611 41568 15660 41596
rect 15611 41565 15623 41568
rect 15565 41559 15623 41565
rect 15304 41528 15332 41559
rect 15654 41556 15660 41568
rect 15712 41556 15718 41608
rect 15841 41599 15899 41605
rect 15841 41565 15853 41599
rect 15887 41596 15899 41599
rect 15930 41596 15936 41608
rect 15887 41568 15936 41596
rect 15887 41565 15899 41568
rect 15841 41559 15899 41565
rect 15930 41556 15936 41568
rect 15988 41556 15994 41608
rect 16040 41528 16068 41636
rect 16125 41599 16183 41605
rect 16125 41565 16137 41599
rect 16171 41596 16183 41599
rect 16298 41596 16304 41608
rect 16171 41568 16304 41596
rect 16171 41565 16183 41568
rect 16125 41559 16183 41565
rect 16298 41556 16304 41568
rect 16356 41556 16362 41608
rect 16390 41556 16396 41608
rect 16448 41556 16454 41608
rect 16482 41556 16488 41608
rect 16540 41556 16546 41608
rect 16758 41556 16764 41608
rect 16816 41556 16822 41608
rect 16942 41556 16948 41608
rect 17000 41596 17006 41608
rect 17037 41599 17095 41605
rect 17037 41596 17049 41599
rect 17000 41568 17049 41596
rect 17000 41556 17006 41568
rect 17037 41565 17049 41568
rect 17083 41565 17095 41599
rect 17037 41559 17095 41565
rect 17218 41556 17224 41608
rect 17276 41596 17282 41608
rect 17313 41599 17371 41605
rect 17313 41596 17325 41599
rect 17276 41568 17325 41596
rect 17276 41556 17282 41568
rect 17313 41565 17325 41568
rect 17359 41565 17371 41599
rect 17313 41559 17371 41565
rect 17586 41556 17592 41608
rect 17644 41556 17650 41608
rect 17678 41556 17684 41608
rect 17736 41596 17742 41608
rect 17865 41599 17923 41605
rect 17865 41596 17877 41599
rect 17736 41568 17877 41596
rect 17736 41556 17742 41568
rect 17865 41565 17877 41568
rect 17911 41565 17923 41599
rect 17865 41559 17923 41565
rect 18046 41556 18052 41608
rect 18104 41556 18110 41608
rect 19628 41596 19656 41636
rect 19705 41633 19717 41667
rect 19751 41664 19763 41667
rect 21266 41664 21272 41676
rect 19751 41636 21272 41664
rect 19751 41633 19763 41636
rect 19705 41627 19763 41633
rect 21266 41624 21272 41636
rect 21324 41624 21330 41676
rect 20438 41596 20444 41608
rect 19628 41568 20444 41596
rect 20438 41556 20444 41568
rect 20496 41556 20502 41608
rect 16500 41528 16528 41556
rect 18064 41528 18092 41556
rect 15304 41500 16068 41528
rect 16224 41500 16528 41528
rect 16592 41500 18092 41528
rect 15381 41463 15439 41469
rect 15381 41460 15393 41463
rect 15028 41432 15393 41460
rect 15381 41429 15393 41432
rect 15427 41429 15439 41463
rect 15381 41423 15439 41429
rect 15933 41463 15991 41469
rect 15933 41429 15945 41463
rect 15979 41460 15991 41463
rect 16022 41460 16028 41472
rect 15979 41432 16028 41460
rect 15979 41429 15991 41432
rect 15933 41423 15991 41429
rect 16022 41420 16028 41432
rect 16080 41420 16086 41472
rect 16224 41469 16252 41500
rect 16592 41469 16620 41500
rect 18138 41488 18144 41540
rect 18196 41488 18202 41540
rect 18693 41531 18751 41537
rect 18693 41497 18705 41531
rect 18739 41528 18751 41531
rect 18782 41528 18788 41540
rect 18739 41500 18788 41528
rect 18739 41497 18751 41500
rect 18693 41491 18751 41497
rect 18782 41488 18788 41500
rect 18840 41488 18846 41540
rect 19426 41488 19432 41540
rect 19484 41488 19490 41540
rect 20165 41531 20223 41537
rect 20165 41497 20177 41531
rect 20211 41497 20223 41531
rect 20165 41491 20223 41497
rect 16209 41463 16267 41469
rect 16209 41429 16221 41463
rect 16255 41429 16267 41463
rect 16209 41423 16267 41429
rect 16577 41463 16635 41469
rect 16577 41429 16589 41463
rect 16623 41429 16635 41463
rect 16577 41423 16635 41429
rect 16850 41420 16856 41472
rect 16908 41420 16914 41472
rect 17402 41420 17408 41472
rect 17460 41420 17466 41472
rect 17954 41420 17960 41472
rect 18012 41460 18018 41472
rect 19058 41460 19064 41472
rect 18012 41432 19064 41460
rect 18012 41420 18018 41432
rect 19058 41420 19064 41432
rect 19116 41420 19122 41472
rect 19334 41420 19340 41472
rect 19392 41460 19398 41472
rect 20180 41460 20208 41491
rect 20530 41488 20536 41540
rect 20588 41488 20594 41540
rect 19392 41432 20208 41460
rect 19392 41420 19398 41432
rect 1104 41370 21043 41392
rect 1104 41318 5894 41370
rect 5946 41318 5958 41370
rect 6010 41318 6022 41370
rect 6074 41318 6086 41370
rect 6138 41318 6150 41370
rect 6202 41318 10839 41370
rect 10891 41318 10903 41370
rect 10955 41318 10967 41370
rect 11019 41318 11031 41370
rect 11083 41318 11095 41370
rect 11147 41318 15784 41370
rect 15836 41318 15848 41370
rect 15900 41318 15912 41370
rect 15964 41318 15976 41370
rect 16028 41318 16040 41370
rect 16092 41318 20729 41370
rect 20781 41318 20793 41370
rect 20845 41318 20857 41370
rect 20909 41318 20921 41370
rect 20973 41318 20985 41370
rect 21037 41318 21043 41370
rect 1104 41296 21043 41318
rect 3326 41216 3332 41268
rect 3384 41256 3390 41268
rect 3421 41259 3479 41265
rect 3421 41256 3433 41259
rect 3384 41228 3433 41256
rect 3384 41216 3390 41228
rect 3421 41225 3433 41228
rect 3467 41225 3479 41259
rect 3421 41219 3479 41225
rect 3697 41259 3755 41265
rect 3697 41225 3709 41259
rect 3743 41256 3755 41259
rect 3786 41256 3792 41268
rect 3743 41228 3792 41256
rect 3743 41225 3755 41228
rect 3697 41219 3755 41225
rect 3786 41216 3792 41228
rect 3844 41216 3850 41268
rect 3970 41216 3976 41268
rect 4028 41216 4034 41268
rect 4249 41259 4307 41265
rect 4249 41225 4261 41259
rect 4295 41256 4307 41259
rect 4890 41256 4896 41268
rect 4295 41228 4896 41256
rect 4295 41225 4307 41228
rect 4249 41219 4307 41225
rect 4890 41216 4896 41228
rect 4948 41216 4954 41268
rect 4982 41216 4988 41268
rect 5040 41256 5046 41268
rect 5077 41259 5135 41265
rect 5077 41256 5089 41259
rect 5040 41228 5089 41256
rect 5040 41216 5046 41228
rect 5077 41225 5089 41228
rect 5123 41225 5135 41259
rect 5077 41219 5135 41225
rect 5258 41216 5264 41268
rect 5316 41216 5322 41268
rect 5810 41216 5816 41268
rect 5868 41216 5874 41268
rect 6546 41216 6552 41268
rect 6604 41216 6610 41268
rect 6730 41216 6736 41268
rect 6788 41256 6794 41268
rect 6825 41259 6883 41265
rect 6825 41256 6837 41259
rect 6788 41228 6837 41256
rect 6788 41216 6794 41228
rect 6825 41225 6837 41228
rect 6871 41225 6883 41259
rect 6825 41219 6883 41225
rect 7193 41259 7251 41265
rect 7193 41225 7205 41259
rect 7239 41256 7251 41259
rect 7374 41256 7380 41268
rect 7239 41228 7380 41256
rect 7239 41225 7251 41228
rect 7193 41219 7251 41225
rect 7374 41216 7380 41228
rect 7432 41216 7438 41268
rect 14366 41216 14372 41268
rect 14424 41216 14430 41268
rect 14550 41216 14556 41268
rect 14608 41216 14614 41268
rect 14642 41216 14648 41268
rect 14700 41216 14706 41268
rect 14734 41216 14740 41268
rect 14792 41256 14798 41268
rect 14921 41259 14979 41265
rect 14792 41228 14872 41256
rect 14792 41216 14798 41228
rect 1946 41148 1952 41200
rect 2004 41188 2010 41200
rect 2682 41188 2688 41200
rect 2004 41160 2688 41188
rect 2004 41148 2010 41160
rect 2682 41148 2688 41160
rect 2740 41148 2746 41200
rect 5276 41188 5304 41216
rect 6914 41188 6920 41200
rect 5276 41160 6040 41188
rect 1397 41123 1455 41129
rect 1397 41089 1409 41123
rect 1443 41120 1455 41123
rect 2774 41120 2780 41132
rect 1443 41092 2780 41120
rect 1443 41089 1455 41092
rect 1397 41083 1455 41089
rect 2774 41080 2780 41092
rect 2832 41080 2838 41132
rect 3602 41080 3608 41132
rect 3660 41080 3666 41132
rect 3881 41123 3939 41129
rect 3881 41089 3893 41123
rect 3927 41120 3939 41123
rect 4062 41120 4068 41132
rect 3927 41092 4068 41120
rect 3927 41089 3939 41092
rect 3881 41083 3939 41089
rect 4062 41080 4068 41092
rect 4120 41080 4126 41132
rect 4157 41123 4215 41129
rect 4157 41089 4169 41123
rect 4203 41120 4215 41123
rect 4338 41120 4344 41132
rect 4203 41092 4344 41120
rect 4203 41089 4215 41092
rect 4157 41083 4215 41089
rect 4338 41080 4344 41092
rect 4396 41080 4402 41132
rect 4430 41080 4436 41132
rect 4488 41080 4494 41132
rect 4982 41080 4988 41132
rect 5040 41080 5046 41132
rect 5074 41080 5080 41132
rect 5132 41120 5138 41132
rect 6012 41129 6040 41160
rect 6196 41160 6920 41188
rect 5261 41123 5319 41129
rect 5261 41120 5273 41123
rect 5132 41092 5273 41120
rect 5132 41080 5138 41092
rect 5261 41089 5273 41092
rect 5307 41089 5319 41123
rect 5261 41083 5319 41089
rect 5721 41123 5779 41129
rect 5721 41089 5733 41123
rect 5767 41089 5779 41123
rect 5721 41083 5779 41089
rect 5997 41123 6055 41129
rect 5997 41089 6009 41123
rect 6043 41089 6055 41123
rect 5997 41083 6055 41089
rect 2133 41055 2191 41061
rect 2133 41021 2145 41055
rect 2179 41021 2191 41055
rect 2133 41015 2191 41021
rect 2148 40928 2176 41015
rect 5350 41012 5356 41064
rect 5408 41012 5414 41064
rect 5736 41052 5764 41083
rect 6196 41052 6224 41160
rect 6914 41148 6920 41160
rect 6972 41148 6978 41200
rect 14568 41188 14596 41216
rect 14844 41188 14872 41228
rect 14921 41225 14933 41259
rect 14967 41256 14979 41259
rect 15010 41256 15016 41268
rect 14967 41228 15016 41256
rect 14967 41225 14979 41228
rect 14921 41219 14979 41225
rect 15010 41216 15016 41228
rect 15068 41216 15074 41268
rect 15194 41216 15200 41268
rect 15252 41216 15258 41268
rect 15562 41216 15568 41268
rect 15620 41256 15626 41268
rect 15841 41259 15899 41265
rect 15841 41256 15853 41259
rect 15620 41228 15853 41256
rect 15620 41216 15626 41228
rect 15841 41225 15853 41228
rect 15887 41225 15899 41259
rect 15841 41219 15899 41225
rect 16117 41259 16175 41265
rect 16117 41225 16129 41259
rect 16163 41256 16175 41259
rect 16390 41256 16396 41268
rect 16163 41228 16396 41256
rect 16163 41225 16175 41228
rect 16117 41219 16175 41225
rect 16390 41216 16396 41228
rect 16448 41216 16454 41268
rect 16669 41259 16727 41265
rect 16669 41225 16681 41259
rect 16715 41256 16727 41259
rect 16942 41256 16948 41268
rect 16715 41228 16948 41256
rect 16715 41225 16727 41228
rect 16669 41219 16727 41225
rect 16942 41216 16948 41228
rect 17000 41216 17006 41268
rect 17037 41259 17095 41265
rect 17037 41225 17049 41259
rect 17083 41225 17095 41259
rect 17037 41219 17095 41225
rect 14568 41160 14688 41188
rect 14844 41160 15148 41188
rect 6733 41123 6791 41129
rect 6733 41089 6745 41123
rect 6779 41089 6791 41123
rect 6733 41083 6791 41089
rect 7009 41123 7067 41129
rect 7009 41089 7021 41123
rect 7055 41089 7067 41123
rect 7009 41083 7067 41089
rect 7377 41123 7435 41129
rect 7377 41089 7389 41123
rect 7423 41120 7435 41123
rect 7653 41123 7711 41129
rect 7423 41092 7604 41120
rect 7423 41089 7435 41092
rect 7377 41083 7435 41089
rect 5736 41024 6224 41052
rect 6270 41012 6276 41064
rect 6328 41012 6334 41064
rect 4801 40987 4859 40993
rect 4801 40953 4813 40987
rect 4847 40984 4859 40987
rect 5368 40984 5396 41012
rect 4847 40956 5396 40984
rect 5537 40987 5595 40993
rect 4847 40953 4859 40956
rect 4801 40947 4859 40953
rect 5537 40953 5549 40987
rect 5583 40984 5595 40987
rect 6288 40984 6316 41012
rect 5583 40956 6316 40984
rect 5583 40953 5595 40956
rect 5537 40947 5595 40953
rect 2130 40876 2136 40928
rect 2188 40876 2194 40928
rect 5718 40876 5724 40928
rect 5776 40916 5782 40928
rect 6748 40916 6776 41083
rect 7024 41052 7052 41083
rect 7024 41024 7512 41052
rect 7190 40944 7196 40996
rect 7248 40944 7254 40996
rect 7484 40993 7512 41024
rect 7469 40987 7527 40993
rect 7469 40953 7481 40987
rect 7515 40953 7527 40987
rect 7576 40984 7604 41092
rect 7653 41089 7665 41123
rect 7699 41089 7711 41123
rect 7653 41083 7711 41089
rect 7668 41052 7696 41083
rect 7926 41080 7932 41132
rect 7984 41080 7990 41132
rect 14277 41123 14335 41129
rect 14277 41089 14289 41123
rect 14323 41089 14335 41123
rect 14277 41083 14335 41089
rect 8754 41052 8760 41064
rect 7668 41024 8760 41052
rect 8754 41012 8760 41024
rect 8812 41012 8818 41064
rect 14292 41052 14320 41083
rect 14550 41080 14556 41132
rect 14608 41080 14614 41132
rect 14660 41120 14688 41160
rect 15120 41129 15148 41160
rect 15304 41160 16712 41188
rect 14829 41123 14887 41129
rect 14829 41120 14841 41123
rect 14660 41092 14841 41120
rect 14829 41089 14841 41092
rect 14875 41089 14887 41123
rect 14829 41083 14887 41089
rect 15105 41123 15163 41129
rect 15105 41089 15117 41123
rect 15151 41089 15163 41123
rect 15105 41083 15163 41089
rect 15304 41052 15332 41160
rect 16684 41132 16712 41160
rect 16758 41148 16764 41200
rect 16816 41188 16822 41200
rect 17052 41188 17080 41219
rect 17218 41216 17224 41268
rect 17276 41216 17282 41268
rect 17494 41216 17500 41268
rect 17552 41256 17558 41268
rect 17589 41259 17647 41265
rect 17589 41256 17601 41259
rect 17552 41228 17601 41256
rect 17552 41216 17558 41228
rect 17589 41225 17601 41228
rect 17635 41225 17647 41259
rect 17589 41219 17647 41225
rect 18230 41216 18236 41268
rect 18288 41256 18294 41268
rect 18877 41259 18935 41265
rect 18877 41256 18889 41259
rect 18288 41228 18889 41256
rect 18288 41216 18294 41228
rect 18877 41225 18889 41228
rect 18923 41225 18935 41259
rect 18877 41219 18935 41225
rect 19242 41216 19248 41268
rect 19300 41256 19306 41268
rect 20257 41259 20315 41265
rect 20257 41256 20269 41259
rect 19300 41228 20269 41256
rect 19300 41216 19306 41228
rect 20257 41225 20269 41228
rect 20303 41225 20315 41259
rect 20257 41219 20315 41225
rect 17236 41188 17264 41216
rect 16816 41160 17080 41188
rect 17144 41160 17264 41188
rect 16816 41148 16822 41160
rect 15378 41080 15384 41132
rect 15436 41080 15442 41132
rect 15562 41080 15568 41132
rect 15620 41120 15626 41132
rect 15749 41123 15807 41129
rect 15749 41120 15761 41123
rect 15620 41092 15761 41120
rect 15620 41080 15626 41092
rect 15749 41089 15761 41092
rect 15795 41089 15807 41123
rect 15749 41083 15807 41089
rect 16025 41123 16083 41129
rect 16025 41089 16037 41123
rect 16071 41089 16083 41123
rect 16025 41083 16083 41089
rect 14292 41024 15332 41052
rect 15470 41012 15476 41064
rect 15528 41052 15534 41064
rect 16040 41052 16068 41083
rect 16206 41080 16212 41132
rect 16264 41080 16270 41132
rect 16298 41080 16304 41132
rect 16356 41080 16362 41132
rect 16666 41080 16672 41132
rect 16724 41080 16730 41132
rect 16850 41080 16856 41132
rect 16908 41080 16914 41132
rect 16942 41080 16948 41132
rect 17000 41120 17006 41132
rect 17144 41120 17172 41160
rect 17402 41148 17408 41200
rect 17460 41188 17466 41200
rect 20165 41191 20223 41197
rect 20165 41188 20177 41191
rect 17460 41160 20177 41188
rect 17460 41148 17466 41160
rect 20165 41157 20177 41160
rect 20211 41157 20223 41191
rect 20165 41151 20223 41157
rect 17000 41092 17172 41120
rect 17000 41080 17006 41092
rect 17218 41080 17224 41132
rect 17276 41080 17282 41132
rect 17494 41080 17500 41132
rect 17552 41080 17558 41132
rect 17773 41123 17831 41129
rect 17773 41089 17785 41123
rect 17819 41089 17831 41123
rect 17773 41083 17831 41089
rect 15528 41024 16068 41052
rect 15528 41012 15534 41024
rect 12802 40984 12808 40996
rect 7576 40956 12808 40984
rect 7469 40947 7527 40953
rect 12802 40944 12808 40956
rect 12860 40944 12866 40996
rect 15565 40987 15623 40993
rect 15565 40953 15577 40987
rect 15611 40984 15623 40987
rect 16224 40984 16252 41080
rect 17034 41012 17040 41064
rect 17092 41052 17098 41064
rect 17788 41052 17816 41083
rect 18230 41080 18236 41132
rect 18288 41080 18294 41132
rect 18509 41123 18567 41129
rect 18509 41089 18521 41123
rect 18555 41120 18567 41123
rect 18785 41123 18843 41129
rect 18555 41092 18736 41120
rect 18555 41089 18567 41092
rect 18509 41083 18567 41089
rect 18708 41052 18736 41092
rect 18785 41089 18797 41123
rect 18831 41120 18843 41123
rect 18966 41120 18972 41132
rect 18831 41092 18972 41120
rect 18831 41089 18843 41092
rect 18785 41083 18843 41089
rect 18966 41080 18972 41092
rect 19024 41080 19030 41132
rect 19058 41080 19064 41132
rect 19116 41080 19122 41132
rect 19521 41123 19579 41129
rect 19521 41089 19533 41123
rect 19567 41120 19579 41123
rect 19981 41123 20039 41129
rect 19981 41120 19993 41123
rect 19567 41092 19993 41120
rect 19567 41089 19579 41092
rect 19521 41083 19579 41089
rect 19981 41089 19993 41092
rect 20027 41120 20039 41123
rect 21082 41120 21088 41132
rect 20027 41092 21088 41120
rect 20027 41089 20039 41092
rect 19981 41083 20039 41089
rect 21082 41080 21088 41092
rect 21140 41080 21146 41132
rect 19150 41052 19156 41064
rect 17092 41024 17724 41052
rect 17788 41024 18644 41052
rect 18708 41024 19156 41052
rect 17092 41012 17098 41024
rect 15611 40956 16252 40984
rect 15611 40953 15623 40956
rect 15565 40947 15623 40953
rect 16758 40944 16764 40996
rect 16816 40984 16822 40996
rect 17586 40984 17592 40996
rect 16816 40956 17592 40984
rect 16816 40944 16822 40956
rect 17586 40944 17592 40956
rect 17644 40944 17650 40996
rect 5776 40888 6776 40916
rect 7208 40916 7236 40944
rect 7745 40919 7803 40925
rect 7745 40916 7757 40919
rect 7208 40888 7757 40916
rect 5776 40876 5782 40888
rect 7745 40885 7757 40888
rect 7791 40885 7803 40919
rect 7745 40879 7803 40885
rect 14093 40919 14151 40925
rect 14093 40885 14105 40919
rect 14139 40916 14151 40919
rect 14918 40916 14924 40928
rect 14139 40888 14924 40916
rect 14139 40885 14151 40888
rect 14093 40879 14151 40885
rect 14918 40876 14924 40888
rect 14976 40876 14982 40928
rect 15378 40876 15384 40928
rect 15436 40916 15442 40928
rect 16390 40916 16396 40928
rect 15436 40888 16396 40916
rect 15436 40876 15442 40888
rect 16390 40876 16396 40888
rect 16448 40876 16454 40928
rect 16482 40876 16488 40928
rect 16540 40916 16546 40928
rect 17313 40919 17371 40925
rect 17313 40916 17325 40919
rect 16540 40888 17325 40916
rect 16540 40876 16546 40888
rect 17313 40885 17325 40888
rect 17359 40885 17371 40919
rect 17696 40916 17724 41024
rect 17770 40944 17776 40996
rect 17828 40984 17834 40996
rect 18616 40993 18644 41024
rect 19150 41012 19156 41024
rect 19208 41012 19214 41064
rect 18325 40987 18383 40993
rect 18325 40984 18337 40987
rect 17828 40956 18337 40984
rect 17828 40944 17834 40956
rect 18325 40953 18337 40956
rect 18371 40953 18383 40987
rect 18325 40947 18383 40953
rect 18601 40987 18659 40993
rect 18601 40953 18613 40987
rect 18647 40953 18659 40987
rect 18601 40947 18659 40953
rect 17862 40916 17868 40928
rect 17696 40888 17868 40916
rect 17313 40879 17371 40885
rect 17862 40876 17868 40888
rect 17920 40876 17926 40928
rect 18046 40876 18052 40928
rect 18104 40876 18110 40928
rect 19797 40919 19855 40925
rect 19797 40885 19809 40919
rect 19843 40916 19855 40919
rect 20162 40916 20168 40928
rect 19843 40888 20168 40916
rect 19843 40885 19855 40888
rect 19797 40879 19855 40885
rect 20162 40876 20168 40888
rect 20220 40876 20226 40928
rect 1104 40826 20884 40848
rect 1104 40774 3422 40826
rect 3474 40774 3486 40826
rect 3538 40774 3550 40826
rect 3602 40774 3614 40826
rect 3666 40774 3678 40826
rect 3730 40774 8367 40826
rect 8419 40774 8431 40826
rect 8483 40774 8495 40826
rect 8547 40774 8559 40826
rect 8611 40774 8623 40826
rect 8675 40774 13312 40826
rect 13364 40774 13376 40826
rect 13428 40774 13440 40826
rect 13492 40774 13504 40826
rect 13556 40774 13568 40826
rect 13620 40774 18257 40826
rect 18309 40774 18321 40826
rect 18373 40774 18385 40826
rect 18437 40774 18449 40826
rect 18501 40774 18513 40826
rect 18565 40774 20884 40826
rect 1104 40752 20884 40774
rect 5626 40712 5632 40724
rect 2746 40684 5632 40712
rect 750 40536 756 40588
rect 808 40576 814 40588
rect 2746 40576 2774 40684
rect 5626 40672 5632 40684
rect 5684 40672 5690 40724
rect 13078 40712 13084 40724
rect 12406 40684 13084 40712
rect 5258 40604 5264 40656
rect 5316 40644 5322 40656
rect 12406 40644 12434 40684
rect 13078 40672 13084 40684
rect 13136 40672 13142 40724
rect 15194 40672 15200 40724
rect 15252 40672 15258 40724
rect 15470 40672 15476 40724
rect 15528 40672 15534 40724
rect 15654 40672 15660 40724
rect 15712 40712 15718 40724
rect 15749 40715 15807 40721
rect 15749 40712 15761 40715
rect 15712 40684 15761 40712
rect 15712 40672 15718 40684
rect 15749 40681 15761 40684
rect 15795 40681 15807 40715
rect 15749 40675 15807 40681
rect 16206 40672 16212 40724
rect 16264 40672 16270 40724
rect 16393 40715 16451 40721
rect 16393 40681 16405 40715
rect 16439 40712 16451 40715
rect 16758 40712 16764 40724
rect 16439 40684 16764 40712
rect 16439 40681 16451 40684
rect 16393 40675 16451 40681
rect 16758 40672 16764 40684
rect 16816 40672 16822 40724
rect 16853 40715 16911 40721
rect 16853 40681 16865 40715
rect 16899 40712 16911 40715
rect 17218 40712 17224 40724
rect 16899 40684 17224 40712
rect 16899 40681 16911 40684
rect 16853 40675 16911 40681
rect 17218 40672 17224 40684
rect 17276 40672 17282 40724
rect 18601 40715 18659 40721
rect 18601 40681 18613 40715
rect 18647 40712 18659 40715
rect 19426 40712 19432 40724
rect 18647 40684 19432 40712
rect 18647 40681 18659 40684
rect 18601 40675 18659 40681
rect 19426 40672 19432 40684
rect 19484 40672 19490 40724
rect 19518 40672 19524 40724
rect 19576 40672 19582 40724
rect 5316 40616 12434 40644
rect 5316 40604 5322 40616
rect 17034 40604 17040 40656
rect 17092 40644 17098 40656
rect 17313 40647 17371 40653
rect 17313 40644 17325 40647
rect 17092 40616 17325 40644
rect 17092 40604 17098 40616
rect 17313 40613 17325 40616
rect 17359 40613 17371 40647
rect 18141 40647 18199 40653
rect 18141 40644 18153 40647
rect 17313 40607 17371 40613
rect 17420 40616 18153 40644
rect 808 40548 2774 40576
rect 808 40536 814 40548
rect 4062 40536 4068 40588
rect 4120 40576 4126 40588
rect 7558 40576 7564 40588
rect 4120 40548 7564 40576
rect 4120 40536 4126 40548
rect 7558 40536 7564 40548
rect 7616 40536 7622 40588
rect 17420 40576 17448 40616
rect 18141 40613 18153 40616
rect 18187 40613 18199 40647
rect 18141 40607 18199 40613
rect 19245 40647 19303 40653
rect 19245 40613 19257 40647
rect 19291 40613 19303 40647
rect 19245 40607 19303 40613
rect 19260 40576 19288 40607
rect 19794 40576 19800 40588
rect 15120 40548 17448 40576
rect 17980 40548 19288 40576
rect 19720 40548 19800 40576
rect 1394 40468 1400 40520
rect 1452 40468 1458 40520
rect 1673 40511 1731 40517
rect 1673 40477 1685 40511
rect 1719 40508 1731 40511
rect 13538 40508 13544 40520
rect 1719 40480 13544 40508
rect 1719 40477 1731 40480
rect 1673 40471 1731 40477
rect 13538 40468 13544 40480
rect 13596 40468 13602 40520
rect 13630 40468 13636 40520
rect 13688 40468 13694 40520
rect 15120 40517 15148 40548
rect 15105 40511 15163 40517
rect 15105 40477 15117 40511
rect 15151 40477 15163 40511
rect 15105 40471 15163 40477
rect 15378 40468 15384 40520
rect 15436 40468 15442 40520
rect 15654 40468 15660 40520
rect 15712 40468 15718 40520
rect 15933 40511 15991 40517
rect 15933 40477 15945 40511
rect 15979 40477 15991 40511
rect 15933 40471 15991 40477
rect 16025 40511 16083 40517
rect 16025 40477 16037 40511
rect 16071 40508 16083 40511
rect 16114 40508 16120 40520
rect 16071 40480 16120 40508
rect 16071 40477 16083 40480
rect 16025 40471 16083 40477
rect 1946 40400 1952 40452
rect 2004 40400 2010 40452
rect 2682 40400 2688 40452
rect 2740 40400 2746 40452
rect 13648 40440 13676 40468
rect 13648 40412 15240 40440
rect 7650 40332 7656 40384
rect 7708 40372 7714 40384
rect 12434 40372 12440 40384
rect 7708 40344 12440 40372
rect 7708 40332 7714 40344
rect 12434 40332 12440 40344
rect 12492 40332 12498 40384
rect 14918 40332 14924 40384
rect 14976 40332 14982 40384
rect 15212 40372 15240 40412
rect 15286 40400 15292 40452
rect 15344 40440 15350 40452
rect 15948 40440 15976 40471
rect 16114 40468 16120 40480
rect 16172 40468 16178 40520
rect 16577 40511 16635 40517
rect 16577 40477 16589 40511
rect 16623 40508 16635 40511
rect 16758 40508 16764 40520
rect 16623 40480 16764 40508
rect 16623 40477 16635 40480
rect 16577 40471 16635 40477
rect 16758 40468 16764 40480
rect 16816 40468 16822 40520
rect 17037 40511 17095 40517
rect 17037 40477 17049 40511
rect 17083 40477 17095 40511
rect 17037 40471 17095 40477
rect 16482 40440 16488 40452
rect 15344 40412 15976 40440
rect 16040 40412 16488 40440
rect 15344 40400 15350 40412
rect 16040 40372 16068 40412
rect 16482 40400 16488 40412
rect 16540 40400 16546 40452
rect 17052 40384 17080 40471
rect 17402 40468 17408 40520
rect 17460 40468 17466 40520
rect 17497 40511 17555 40517
rect 17497 40477 17509 40511
rect 17543 40477 17555 40511
rect 17497 40471 17555 40477
rect 15212 40344 16068 40372
rect 16206 40332 16212 40384
rect 16264 40372 16270 40384
rect 16942 40372 16948 40384
rect 16264 40344 16948 40372
rect 16264 40332 16270 40344
rect 16942 40332 16948 40344
rect 17000 40332 17006 40384
rect 17034 40332 17040 40384
rect 17092 40332 17098 40384
rect 17420 40372 17448 40468
rect 17512 40440 17540 40471
rect 17770 40468 17776 40520
rect 17828 40468 17834 40520
rect 17980 40440 18008 40548
rect 18049 40511 18107 40517
rect 18049 40477 18061 40511
rect 18095 40508 18107 40511
rect 18138 40508 18144 40520
rect 18095 40480 18144 40508
rect 18095 40477 18107 40480
rect 18049 40471 18107 40477
rect 18138 40468 18144 40480
rect 18196 40468 18202 40520
rect 18325 40511 18383 40517
rect 18325 40477 18337 40511
rect 18371 40508 18383 40511
rect 18785 40511 18843 40517
rect 18371 40480 18460 40508
rect 18371 40477 18383 40480
rect 18325 40471 18383 40477
rect 17512 40412 18008 40440
rect 18432 40384 18460 40480
rect 18785 40477 18797 40511
rect 18831 40508 18843 40511
rect 18831 40480 18920 40508
rect 18831 40477 18843 40480
rect 18785 40471 18843 40477
rect 17589 40375 17647 40381
rect 17589 40372 17601 40375
rect 17420 40344 17601 40372
rect 17589 40341 17601 40344
rect 17635 40341 17647 40375
rect 17589 40335 17647 40341
rect 17770 40332 17776 40384
rect 17828 40372 17834 40384
rect 17865 40375 17923 40381
rect 17865 40372 17877 40375
rect 17828 40344 17877 40372
rect 17828 40332 17834 40344
rect 17865 40341 17877 40344
rect 17911 40341 17923 40375
rect 17865 40335 17923 40341
rect 18414 40332 18420 40384
rect 18472 40332 18478 40384
rect 18892 40381 18920 40480
rect 19058 40468 19064 40520
rect 19116 40468 19122 40520
rect 19426 40468 19432 40520
rect 19484 40468 19490 40520
rect 19720 40517 19748 40548
rect 19794 40536 19800 40548
rect 19852 40536 19858 40588
rect 19705 40511 19763 40517
rect 19705 40477 19717 40511
rect 19751 40477 19763 40511
rect 19705 40471 19763 40477
rect 19978 40468 19984 40520
rect 20036 40468 20042 40520
rect 20165 40443 20223 40449
rect 20165 40409 20177 40443
rect 20211 40440 20223 40443
rect 20346 40440 20352 40452
rect 20211 40412 20352 40440
rect 20211 40409 20223 40412
rect 20165 40403 20223 40409
rect 20346 40400 20352 40412
rect 20404 40400 20410 40452
rect 20533 40443 20591 40449
rect 20533 40409 20545 40443
rect 20579 40440 20591 40443
rect 21266 40440 21272 40452
rect 20579 40412 21272 40440
rect 20579 40409 20591 40412
rect 20533 40403 20591 40409
rect 21266 40400 21272 40412
rect 21324 40400 21330 40452
rect 18877 40375 18935 40381
rect 18877 40341 18889 40375
rect 18923 40341 18935 40375
rect 18877 40335 18935 40341
rect 19794 40332 19800 40384
rect 19852 40332 19858 40384
rect 1104 40282 21043 40304
rect 1104 40230 5894 40282
rect 5946 40230 5958 40282
rect 6010 40230 6022 40282
rect 6074 40230 6086 40282
rect 6138 40230 6150 40282
rect 6202 40230 10839 40282
rect 10891 40230 10903 40282
rect 10955 40230 10967 40282
rect 11019 40230 11031 40282
rect 11083 40230 11095 40282
rect 11147 40230 15784 40282
rect 15836 40230 15848 40282
rect 15900 40230 15912 40282
rect 15964 40230 15976 40282
rect 16028 40230 16040 40282
rect 16092 40230 20729 40282
rect 20781 40230 20793 40282
rect 20845 40230 20857 40282
rect 20909 40230 20921 40282
rect 20973 40230 20985 40282
rect 21037 40230 21043 40282
rect 1104 40208 21043 40230
rect 7650 40128 7656 40180
rect 7708 40128 7714 40180
rect 7760 40140 8064 40168
rect 1302 40060 1308 40112
rect 1360 40100 1366 40112
rect 1397 40103 1455 40109
rect 1397 40100 1409 40103
rect 1360 40072 1409 40100
rect 1360 40060 1366 40072
rect 1397 40069 1409 40072
rect 1443 40069 1455 40103
rect 1397 40063 1455 40069
rect 2682 40060 2688 40112
rect 2740 40060 2746 40112
rect 2777 40103 2835 40109
rect 2777 40069 2789 40103
rect 2823 40100 2835 40103
rect 7668 40100 7696 40128
rect 2823 40072 7696 40100
rect 2823 40069 2835 40072
rect 2777 40063 2835 40069
rect 2501 40035 2559 40041
rect 2501 40032 2513 40035
rect 1504 40004 2513 40032
rect 1302 39924 1308 39976
rect 1360 39964 1366 39976
rect 1504 39964 1532 40004
rect 2501 40001 2513 40004
rect 2547 40001 2559 40035
rect 2700 40032 2728 40060
rect 2700 40004 3004 40032
rect 2501 39995 2559 40001
rect 1360 39936 1532 39964
rect 1360 39924 1366 39936
rect 2038 39924 2044 39976
rect 2096 39964 2102 39976
rect 2133 39967 2191 39973
rect 2133 39964 2145 39967
rect 2096 39936 2145 39964
rect 2096 39924 2102 39936
rect 2133 39933 2145 39936
rect 2179 39964 2191 39967
rect 2976 39964 3004 40004
rect 3050 39992 3056 40044
rect 3108 39992 3114 40044
rect 3329 40035 3387 40041
rect 3329 40001 3341 40035
rect 3375 40032 3387 40035
rect 4799 40035 4857 40041
rect 4799 40032 4811 40035
rect 3375 40004 4811 40032
rect 3375 40001 3387 40004
rect 3329 39995 3387 40001
rect 4799 40001 4811 40004
rect 4845 40032 4857 40035
rect 4890 40032 4896 40044
rect 4845 40004 4896 40032
rect 4845 40001 4857 40004
rect 4799 39995 4857 40001
rect 3344 39964 3372 39995
rect 4890 39992 4896 40004
rect 4948 39992 4954 40044
rect 7760 40032 7788 40140
rect 7668 40004 7788 40032
rect 2179 39936 2774 39964
rect 2976 39936 3372 39964
rect 2179 39933 2191 39936
rect 2133 39927 2191 39933
rect 2746 39896 2774 39936
rect 4062 39924 4068 39976
rect 4120 39924 4126 39976
rect 7668 39973 7696 40004
rect 7834 40002 7840 40054
rect 7892 40041 7898 40054
rect 7892 40035 7953 40041
rect 7892 40002 7907 40035
rect 7895 40001 7907 40002
rect 7941 40001 7953 40035
rect 8036 40032 8064 40140
rect 15562 40128 15568 40180
rect 15620 40128 15626 40180
rect 16114 40128 16120 40180
rect 16172 40128 16178 40180
rect 16666 40128 16672 40180
rect 16724 40168 16730 40180
rect 16853 40171 16911 40177
rect 16853 40168 16865 40171
rect 16724 40140 16865 40168
rect 16724 40128 16730 40140
rect 16853 40137 16865 40140
rect 16899 40137 16911 40171
rect 16853 40131 16911 40137
rect 17129 40171 17187 40177
rect 17129 40137 17141 40171
rect 17175 40168 17187 40171
rect 17310 40168 17316 40180
rect 17175 40140 17316 40168
rect 17175 40137 17187 40140
rect 17129 40131 17187 40137
rect 17310 40128 17316 40140
rect 17368 40128 17374 40180
rect 17405 40171 17463 40177
rect 17405 40137 17417 40171
rect 17451 40168 17463 40171
rect 17678 40168 17684 40180
rect 17451 40140 17684 40168
rect 17451 40137 17463 40140
rect 17405 40131 17463 40137
rect 17678 40128 17684 40140
rect 17736 40128 17742 40180
rect 17957 40171 18015 40177
rect 17957 40137 17969 40171
rect 18003 40168 18015 40171
rect 19058 40168 19064 40180
rect 18003 40140 19064 40168
rect 18003 40137 18015 40140
rect 17957 40131 18015 40137
rect 19058 40128 19064 40140
rect 19116 40128 19122 40180
rect 19794 40128 19800 40180
rect 19852 40168 19858 40180
rect 19852 40140 20208 40168
rect 19852 40128 19858 40140
rect 15580 40100 15608 40128
rect 12452 40072 15608 40100
rect 11330 40032 11336 40044
rect 8036 40004 11336 40032
rect 7895 39995 7953 40001
rect 11330 39992 11336 40004
rect 11388 40032 11394 40044
rect 12452 40032 12480 40072
rect 16942 40060 16948 40112
rect 17000 40100 17006 40112
rect 18046 40100 18052 40112
rect 17000 40072 17080 40100
rect 17000 40060 17006 40072
rect 11388 40004 12480 40032
rect 11388 39992 11394 40004
rect 12802 39992 12808 40044
rect 12860 40032 12866 40044
rect 14182 40032 14188 40044
rect 12860 40004 14188 40032
rect 12860 39992 12866 40004
rect 14182 39992 14188 40004
rect 14240 39992 14246 40044
rect 14642 39992 14648 40044
rect 14700 39992 14706 40044
rect 17052 40041 17080 40072
rect 17328 40072 18052 40100
rect 17328 40041 17356 40072
rect 18046 40060 18052 40072
rect 18104 40060 18110 40112
rect 18230 40060 18236 40112
rect 18288 40100 18294 40112
rect 20180 40109 20208 40140
rect 20254 40128 20260 40180
rect 20312 40168 20318 40180
rect 20312 40140 20392 40168
rect 20312 40128 20318 40140
rect 20165 40103 20223 40109
rect 18288 40072 19104 40100
rect 18288 40060 18294 40072
rect 17037 40035 17095 40041
rect 17037 40001 17049 40035
rect 17083 40001 17095 40035
rect 17037 39995 17095 40001
rect 17313 40035 17371 40041
rect 17313 40001 17325 40035
rect 17359 40001 17371 40035
rect 17313 39995 17371 40001
rect 17586 39992 17592 40044
rect 17644 39992 17650 40044
rect 17862 39992 17868 40044
rect 17920 39992 17926 40044
rect 18141 40035 18199 40041
rect 18141 40001 18153 40035
rect 18187 40032 18199 40035
rect 18322 40032 18328 40044
rect 18187 40004 18328 40032
rect 18187 40001 18199 40004
rect 18141 39995 18199 40001
rect 18322 39992 18328 40004
rect 18380 39992 18386 40044
rect 18601 40035 18659 40041
rect 18601 40001 18613 40035
rect 18647 40032 18659 40035
rect 18874 40032 18880 40044
rect 18647 40004 18880 40032
rect 18647 40001 18659 40004
rect 18601 39995 18659 40001
rect 18874 39992 18880 40004
rect 18932 39992 18938 40044
rect 19076 40041 19104 40072
rect 20165 40069 20177 40103
rect 20211 40069 20223 40103
rect 20165 40063 20223 40069
rect 19061 40035 19119 40041
rect 19061 40001 19073 40035
rect 19107 40001 19119 40035
rect 19061 39995 19119 40001
rect 19242 39992 19248 40044
rect 19300 39992 19306 40044
rect 19334 39992 19340 40044
rect 19392 40032 19398 40044
rect 19429 40035 19487 40041
rect 19429 40032 19441 40035
rect 19392 40004 19441 40032
rect 19392 39992 19398 40004
rect 19429 40001 19441 40004
rect 19475 40001 19487 40035
rect 19429 39995 19487 40001
rect 19705 40035 19763 40041
rect 19705 40001 19717 40035
rect 19751 40032 19763 40035
rect 19886 40032 19892 40044
rect 19751 40004 19892 40032
rect 19751 40001 19763 40004
rect 19705 39995 19763 40001
rect 19886 39992 19892 40004
rect 19944 39992 19950 40044
rect 19981 40035 20039 40041
rect 19981 40001 19993 40035
rect 20027 40032 20039 40035
rect 20254 40032 20260 40044
rect 20027 40004 20260 40032
rect 20027 40001 20039 40004
rect 19981 39995 20039 40001
rect 20254 39992 20260 40004
rect 20312 39992 20318 40044
rect 4525 39967 4583 39973
rect 4525 39933 4537 39967
rect 4571 39933 4583 39967
rect 7653 39967 7711 39973
rect 7653 39964 7665 39967
rect 4525 39927 4583 39933
rect 7576 39936 7665 39964
rect 4080 39896 4108 39924
rect 2746 39868 4108 39896
rect 3786 39788 3792 39840
rect 3844 39828 3850 39840
rect 4540 39828 4568 39927
rect 7576 39840 7604 39936
rect 7653 39933 7665 39936
rect 7699 39933 7711 39967
rect 7653 39927 7711 39933
rect 11422 39924 11428 39976
rect 11480 39964 11486 39976
rect 16482 39964 16488 39976
rect 11480 39936 16488 39964
rect 11480 39924 11486 39936
rect 16482 39924 16488 39936
rect 16540 39924 16546 39976
rect 16574 39924 16580 39976
rect 16632 39924 16638 39976
rect 16666 39924 16672 39976
rect 16724 39964 16730 39976
rect 19260 39964 19288 39992
rect 16724 39936 19288 39964
rect 16724 39924 16730 39936
rect 16592 39896 16620 39924
rect 17681 39899 17739 39905
rect 17681 39896 17693 39899
rect 16592 39868 17693 39896
rect 17681 39865 17693 39868
rect 17727 39865 17739 39899
rect 17681 39859 17739 39865
rect 18046 39856 18052 39908
rect 18104 39896 18110 39908
rect 19245 39899 19303 39905
rect 19245 39896 19257 39899
rect 18104 39868 19257 39896
rect 18104 39856 18110 39868
rect 19245 39865 19257 39868
rect 19291 39865 19303 39899
rect 20364 39896 20392 40140
rect 19245 39859 19303 39865
rect 19352 39868 20392 39896
rect 5442 39828 5448 39840
rect 3844 39800 5448 39828
rect 3844 39788 3850 39800
rect 5442 39788 5448 39800
rect 5500 39788 5506 39840
rect 5534 39788 5540 39840
rect 5592 39788 5598 39840
rect 7558 39788 7564 39840
rect 7616 39788 7622 39840
rect 7926 39788 7932 39840
rect 7984 39828 7990 39840
rect 8665 39831 8723 39837
rect 8665 39828 8677 39831
rect 7984 39800 8677 39828
rect 7984 39788 7990 39800
rect 8665 39797 8677 39800
rect 8711 39797 8723 39831
rect 8665 39791 8723 39797
rect 14918 39788 14924 39840
rect 14976 39828 14982 39840
rect 18138 39828 18144 39840
rect 14976 39800 18144 39828
rect 14976 39788 14982 39800
rect 18138 39788 18144 39800
rect 18196 39788 18202 39840
rect 18417 39831 18475 39837
rect 18417 39797 18429 39831
rect 18463 39828 18475 39831
rect 18690 39828 18696 39840
rect 18463 39800 18696 39828
rect 18463 39797 18475 39800
rect 18417 39791 18475 39797
rect 18690 39788 18696 39800
rect 18748 39788 18754 39840
rect 18874 39788 18880 39840
rect 18932 39788 18938 39840
rect 19058 39788 19064 39840
rect 19116 39828 19122 39840
rect 19352 39828 19380 39868
rect 19116 39800 19380 39828
rect 19116 39788 19122 39800
rect 19518 39788 19524 39840
rect 19576 39788 19582 39840
rect 19794 39788 19800 39840
rect 19852 39788 19858 39840
rect 20441 39831 20499 39837
rect 20441 39797 20453 39831
rect 20487 39828 20499 39831
rect 20990 39828 20996 39840
rect 20487 39800 20996 39828
rect 20487 39797 20499 39800
rect 20441 39791 20499 39797
rect 20990 39788 20996 39800
rect 21048 39788 21054 39840
rect 1104 39738 20884 39760
rect 1104 39686 3422 39738
rect 3474 39686 3486 39738
rect 3538 39686 3550 39738
rect 3602 39686 3614 39738
rect 3666 39686 3678 39738
rect 3730 39686 8367 39738
rect 8419 39686 8431 39738
rect 8483 39686 8495 39738
rect 8547 39686 8559 39738
rect 8611 39686 8623 39738
rect 8675 39686 13312 39738
rect 13364 39686 13376 39738
rect 13428 39686 13440 39738
rect 13492 39686 13504 39738
rect 13556 39686 13568 39738
rect 13620 39686 18257 39738
rect 18309 39686 18321 39738
rect 18373 39686 18385 39738
rect 18437 39686 18449 39738
rect 18501 39686 18513 39738
rect 18565 39686 20884 39738
rect 1104 39664 20884 39686
rect 7558 39624 7564 39636
rect 2746 39596 4476 39624
rect 1394 39380 1400 39432
rect 1452 39380 1458 39432
rect 1949 39423 2007 39429
rect 1949 39389 1961 39423
rect 1995 39420 2007 39423
rect 2130 39420 2136 39432
rect 1995 39392 2136 39420
rect 1995 39389 2007 39392
rect 1949 39383 2007 39389
rect 2130 39380 2136 39392
rect 2188 39380 2194 39432
rect 2223 39423 2281 39429
rect 2223 39389 2235 39423
rect 2269 39420 2281 39423
rect 2746 39420 2774 39596
rect 3786 39516 3792 39568
rect 3844 39516 3850 39568
rect 3804 39429 3832 39516
rect 2269 39392 2774 39420
rect 3789 39423 3847 39429
rect 2269 39389 2281 39392
rect 2223 39383 2281 39389
rect 3789 39389 3801 39423
rect 3835 39389 3847 39423
rect 4062 39420 4068 39432
rect 4023 39392 4068 39420
rect 3789 39383 3847 39389
rect 4062 39380 4068 39392
rect 4120 39380 4126 39432
rect 4448 39420 4476 39596
rect 6380 39596 7564 39624
rect 6380 39497 6408 39596
rect 7558 39584 7564 39596
rect 7616 39584 7622 39636
rect 13722 39584 13728 39636
rect 13780 39584 13786 39636
rect 15289 39627 15347 39633
rect 15289 39593 15301 39627
rect 15335 39624 15347 39627
rect 15654 39624 15660 39636
rect 15335 39596 15660 39624
rect 15335 39593 15347 39596
rect 15289 39587 15347 39593
rect 15654 39584 15660 39596
rect 15712 39584 15718 39636
rect 16945 39627 17003 39633
rect 16945 39624 16957 39627
rect 15764 39596 16957 39624
rect 7374 39516 7380 39568
rect 7432 39516 7438 39568
rect 13740 39556 13768 39584
rect 15764 39556 15792 39596
rect 16945 39593 16957 39596
rect 16991 39593 17003 39627
rect 16945 39587 17003 39593
rect 17221 39627 17279 39633
rect 17221 39593 17233 39627
rect 17267 39624 17279 39627
rect 17586 39624 17592 39636
rect 17267 39596 17592 39624
rect 17267 39593 17279 39596
rect 17221 39587 17279 39593
rect 17586 39584 17592 39596
rect 17644 39584 17650 39636
rect 17678 39584 17684 39636
rect 17736 39624 17742 39636
rect 17773 39627 17831 39633
rect 17773 39624 17785 39627
rect 17736 39596 17785 39624
rect 17736 39584 17742 39596
rect 17773 39593 17785 39596
rect 17819 39593 17831 39627
rect 17773 39587 17831 39593
rect 17862 39584 17868 39636
rect 17920 39584 17926 39636
rect 17954 39584 17960 39636
rect 18012 39624 18018 39636
rect 18325 39627 18383 39633
rect 18325 39624 18337 39627
rect 18012 39596 18337 39624
rect 18012 39584 18018 39596
rect 18325 39593 18337 39596
rect 18371 39593 18383 39627
rect 18325 39587 18383 39593
rect 18877 39627 18935 39633
rect 18877 39593 18889 39627
rect 18923 39624 18935 39627
rect 19334 39624 19340 39636
rect 18923 39596 19340 39624
rect 18923 39593 18935 39596
rect 18877 39587 18935 39593
rect 19334 39584 19340 39596
rect 19392 39584 19398 39636
rect 19426 39584 19432 39636
rect 19484 39624 19490 39636
rect 19613 39627 19671 39633
rect 19613 39624 19625 39627
rect 19484 39596 19625 39624
rect 19484 39584 19490 39596
rect 19613 39593 19625 39596
rect 19659 39593 19671 39627
rect 19613 39587 19671 39593
rect 20162 39584 20168 39636
rect 20220 39584 20226 39636
rect 13740 39528 15792 39556
rect 16206 39516 16212 39568
rect 16264 39516 16270 39568
rect 16393 39559 16451 39565
rect 16393 39525 16405 39559
rect 16439 39556 16451 39559
rect 16574 39556 16580 39568
rect 16439 39528 16580 39556
rect 16439 39525 16451 39528
rect 16393 39519 16451 39525
rect 16574 39516 16580 39528
rect 16632 39516 16638 39568
rect 16669 39559 16727 39565
rect 16669 39525 16681 39559
rect 16715 39556 16727 39559
rect 17880 39556 17908 39584
rect 16715 39528 17908 39556
rect 18049 39559 18107 39565
rect 16715 39525 16727 39528
rect 16669 39519 16727 39525
rect 18049 39525 18061 39559
rect 18095 39556 18107 39559
rect 18506 39556 18512 39568
rect 18095 39528 18512 39556
rect 18095 39525 18107 39528
rect 18049 39519 18107 39525
rect 18506 39516 18512 39528
rect 18564 39516 18570 39568
rect 18601 39559 18659 39565
rect 18601 39525 18613 39559
rect 18647 39525 18659 39559
rect 18601 39519 18659 39525
rect 18708 39528 19334 39556
rect 6365 39491 6423 39497
rect 6365 39457 6377 39491
rect 6411 39457 6423 39491
rect 6365 39451 6423 39457
rect 12618 39448 12624 39500
rect 12676 39488 12682 39500
rect 17586 39488 17592 39500
rect 12676 39460 17592 39488
rect 12676 39448 12682 39460
rect 17586 39448 17592 39460
rect 17644 39448 17650 39500
rect 18616 39488 18644 39519
rect 17696 39460 18644 39488
rect 6638 39420 6644 39432
rect 4448 39392 6644 39420
rect 6638 39380 6644 39392
rect 6696 39380 6702 39432
rect 11422 39420 11428 39432
rect 7392 39392 11428 39420
rect 1673 39355 1731 39361
rect 1673 39321 1685 39355
rect 1719 39352 1731 39355
rect 7392 39352 7420 39392
rect 11422 39380 11428 39392
rect 11480 39380 11486 39432
rect 15286 39420 15292 39432
rect 12406 39392 15292 39420
rect 1719 39324 7420 39352
rect 1719 39321 1731 39324
rect 1673 39315 1731 39321
rect 9582 39312 9588 39364
rect 9640 39352 9646 39364
rect 12406 39352 12434 39392
rect 15286 39380 15292 39392
rect 15344 39380 15350 39432
rect 15470 39380 15476 39432
rect 15528 39380 15534 39432
rect 16577 39423 16635 39429
rect 16577 39389 16589 39423
rect 16623 39389 16635 39423
rect 16577 39383 16635 39389
rect 9640 39324 12434 39352
rect 16592 39352 16620 39383
rect 16850 39380 16856 39432
rect 16908 39380 16914 39432
rect 17126 39380 17132 39432
rect 17184 39380 17190 39432
rect 17402 39380 17408 39432
rect 17460 39380 17466 39432
rect 17696 39429 17724 39460
rect 17681 39423 17739 39429
rect 17681 39389 17693 39423
rect 17727 39389 17739 39423
rect 17681 39383 17739 39389
rect 17957 39423 18015 39429
rect 17957 39389 17969 39423
rect 18003 39420 18015 39423
rect 18003 39392 18184 39420
rect 18003 39389 18015 39392
rect 17957 39383 18015 39389
rect 18156 39364 18184 39392
rect 18230 39380 18236 39432
rect 18288 39380 18294 39432
rect 18509 39423 18567 39429
rect 18509 39389 18521 39423
rect 18555 39420 18567 39423
rect 18708 39420 18736 39528
rect 19306 39488 19334 39528
rect 20180 39488 20208 39584
rect 18892 39460 19196 39488
rect 19306 39460 20208 39488
rect 18555 39392 18736 39420
rect 18785 39423 18843 39429
rect 18555 39389 18567 39392
rect 18509 39383 18567 39389
rect 18785 39389 18797 39423
rect 18831 39416 18843 39423
rect 18892 39416 18920 39460
rect 19168 39436 19196 39460
rect 19168 39432 19288 39436
rect 19061 39423 19119 39429
rect 19061 39420 19073 39423
rect 18831 39389 18920 39416
rect 18785 39388 18920 39389
rect 18984 39392 19073 39420
rect 18785 39383 18843 39388
rect 18046 39352 18052 39364
rect 16592 39324 18052 39352
rect 9640 39312 9646 39324
rect 18046 39312 18052 39324
rect 18104 39312 18110 39364
rect 18138 39312 18144 39364
rect 18196 39312 18202 39364
rect 18322 39312 18328 39364
rect 18380 39352 18386 39364
rect 18984 39352 19012 39392
rect 19061 39389 19073 39392
rect 19107 39389 19119 39423
rect 19168 39408 19248 39432
rect 19061 39383 19119 39389
rect 19242 39380 19248 39408
rect 19300 39380 19306 39432
rect 19426 39380 19432 39432
rect 19484 39420 19490 39432
rect 19521 39423 19579 39429
rect 19521 39420 19533 39423
rect 19484 39392 19533 39420
rect 19484 39380 19490 39392
rect 19521 39389 19533 39392
rect 19567 39389 19579 39423
rect 19521 39383 19579 39389
rect 19702 39380 19708 39432
rect 19760 39420 19766 39432
rect 19797 39423 19855 39429
rect 19797 39420 19809 39423
rect 19760 39392 19809 39420
rect 19760 39380 19766 39392
rect 19797 39389 19809 39392
rect 19843 39389 19855 39423
rect 19797 39383 19855 39389
rect 20165 39355 20223 39361
rect 20165 39352 20177 39355
rect 18380 39324 19012 39352
rect 19076 39324 20177 39352
rect 18380 39312 18386 39324
rect 2961 39287 3019 39293
rect 2961 39253 2973 39287
rect 3007 39284 3019 39287
rect 3786 39284 3792 39296
rect 3007 39256 3792 39284
rect 3007 39253 3019 39256
rect 2961 39247 3019 39253
rect 3786 39244 3792 39256
rect 3844 39244 3850 39296
rect 4706 39244 4712 39296
rect 4764 39284 4770 39296
rect 4801 39287 4859 39293
rect 4801 39284 4813 39287
rect 4764 39256 4813 39284
rect 4764 39244 4770 39256
rect 4801 39253 4813 39256
rect 4847 39253 4859 39287
rect 4801 39247 4859 39253
rect 5442 39244 5448 39296
rect 5500 39284 5506 39296
rect 9600 39284 9628 39312
rect 5500 39256 9628 39284
rect 5500 39244 5506 39256
rect 16850 39244 16856 39296
rect 16908 39284 16914 39296
rect 17310 39284 17316 39296
rect 16908 39256 17316 39284
rect 16908 39244 16914 39256
rect 17310 39244 17316 39256
rect 17368 39244 17374 39296
rect 17497 39287 17555 39293
rect 17497 39253 17509 39287
rect 17543 39284 17555 39287
rect 18782 39284 18788 39296
rect 17543 39256 18788 39284
rect 17543 39253 17555 39256
rect 17497 39247 17555 39253
rect 18782 39244 18788 39256
rect 18840 39244 18846 39296
rect 18966 39244 18972 39296
rect 19024 39284 19030 39296
rect 19076 39284 19104 39324
rect 20165 39321 20177 39324
rect 20211 39321 20223 39355
rect 20165 39315 20223 39321
rect 20533 39355 20591 39361
rect 20533 39321 20545 39355
rect 20579 39352 20591 39355
rect 21266 39352 21272 39364
rect 20579 39324 21272 39352
rect 20579 39321 20591 39324
rect 20533 39315 20591 39321
rect 21266 39312 21272 39324
rect 21324 39312 21330 39364
rect 19024 39256 19104 39284
rect 19337 39287 19395 39293
rect 19024 39244 19030 39256
rect 19337 39253 19349 39287
rect 19383 39284 19395 39287
rect 19978 39284 19984 39296
rect 19383 39256 19984 39284
rect 19383 39253 19395 39256
rect 19337 39247 19395 39253
rect 19978 39244 19984 39256
rect 20036 39244 20042 39296
rect 1104 39194 21043 39216
rect 1104 39142 5894 39194
rect 5946 39142 5958 39194
rect 6010 39142 6022 39194
rect 6074 39142 6086 39194
rect 6138 39142 6150 39194
rect 6202 39142 10839 39194
rect 10891 39142 10903 39194
rect 10955 39142 10967 39194
rect 11019 39142 11031 39194
rect 11083 39142 11095 39194
rect 11147 39142 15784 39194
rect 15836 39142 15848 39194
rect 15900 39142 15912 39194
rect 15964 39142 15976 39194
rect 16028 39142 16040 39194
rect 16092 39142 20729 39194
rect 20781 39142 20793 39194
rect 20845 39142 20857 39194
rect 20909 39142 20921 39194
rect 20973 39142 20985 39194
rect 21037 39142 21043 39194
rect 1104 39120 21043 39142
rect 11238 39080 11244 39092
rect 2240 39052 11244 39080
rect 2240 39021 2268 39052
rect 11238 39040 11244 39052
rect 11296 39080 11302 39092
rect 14550 39080 14556 39092
rect 11296 39052 14556 39080
rect 11296 39040 11302 39052
rect 14550 39040 14556 39052
rect 14608 39080 14614 39092
rect 16390 39080 16396 39092
rect 14608 39052 16396 39080
rect 14608 39040 14614 39052
rect 16390 39040 16396 39052
rect 16448 39040 16454 39092
rect 16485 39083 16543 39089
rect 16485 39049 16497 39083
rect 16531 39049 16543 39083
rect 16485 39043 16543 39049
rect 17037 39083 17095 39089
rect 17037 39049 17049 39083
rect 17083 39080 17095 39083
rect 17402 39080 17408 39092
rect 17083 39052 17408 39080
rect 17083 39049 17095 39052
rect 17037 39043 17095 39049
rect 2225 39015 2283 39021
rect 2225 38981 2237 39015
rect 2271 38981 2283 39015
rect 4246 39012 4252 39024
rect 3068 38984 4252 39012
rect 2225 38975 2283 38981
rect 2943 38977 3001 38983
rect 1397 38947 1455 38953
rect 1397 38913 1409 38947
rect 1443 38944 1455 38947
rect 1486 38944 1492 38956
rect 1443 38916 1492 38944
rect 1443 38913 1455 38916
rect 1397 38907 1455 38913
rect 1486 38904 1492 38916
rect 1544 38904 1550 38956
rect 1946 38904 1952 38956
rect 2004 38904 2010 38956
rect 2943 38943 2955 38977
rect 2989 38974 3001 38977
rect 3068 38974 3096 38984
rect 2989 38946 3096 38974
rect 4246 38972 4252 38984
rect 4304 38972 4310 39024
rect 4525 39015 4583 39021
rect 4525 38981 4537 39015
rect 4571 39012 4583 39015
rect 4614 39012 4620 39024
rect 4571 38984 4620 39012
rect 4571 38981 4583 38984
rect 4525 38975 4583 38981
rect 4614 38972 4620 38984
rect 4672 38972 4678 39024
rect 4798 38972 4804 39024
rect 4856 38972 4862 39024
rect 4893 39015 4951 39021
rect 4893 38981 4905 39015
rect 4939 39012 4951 39015
rect 5534 39012 5540 39024
rect 4939 38984 5540 39012
rect 4939 38981 4951 38984
rect 4893 38975 4951 38981
rect 5534 38972 5540 38984
rect 5592 38972 5598 39024
rect 16500 39012 16528 39043
rect 17402 39040 17408 39052
rect 17460 39040 17466 39092
rect 17681 39083 17739 39089
rect 17681 39049 17693 39083
rect 17727 39080 17739 39083
rect 18230 39080 18236 39092
rect 17727 39052 18236 39080
rect 17727 39049 17739 39052
rect 17681 39043 17739 39049
rect 18230 39040 18236 39052
rect 18288 39040 18294 39092
rect 18322 39040 18328 39092
rect 18380 39080 18386 39092
rect 18509 39083 18567 39089
rect 18509 39080 18521 39083
rect 18380 39052 18521 39080
rect 18380 39040 18386 39052
rect 18509 39049 18521 39052
rect 18555 39049 18567 39083
rect 18509 39043 18567 39049
rect 18785 39083 18843 39089
rect 18785 39049 18797 39083
rect 18831 39080 18843 39083
rect 18966 39080 18972 39092
rect 18831 39052 18972 39080
rect 18831 39049 18843 39052
rect 18785 39043 18843 39049
rect 18966 39040 18972 39052
rect 19024 39040 19030 39092
rect 19061 39083 19119 39089
rect 19061 39049 19073 39083
rect 19107 39080 19119 39083
rect 19107 39052 19196 39080
rect 19107 39049 19119 39052
rect 19061 39043 19119 39049
rect 16500 38984 17540 39012
rect 2989 38943 3001 38946
rect 2943 38937 3001 38943
rect 5166 38904 5172 38956
rect 5224 38944 5230 38956
rect 5261 38947 5319 38953
rect 5261 38944 5273 38947
rect 5224 38916 5273 38944
rect 5224 38904 5230 38916
rect 5261 38913 5273 38916
rect 5307 38913 5319 38947
rect 5261 38907 5319 38913
rect 5626 38904 5632 38956
rect 5684 38953 5690 38956
rect 5684 38947 5701 38953
rect 5689 38913 5701 38947
rect 5684 38907 5701 38913
rect 5684 38904 5690 38907
rect 7926 38904 7932 38956
rect 7984 38904 7990 38956
rect 12434 38904 12440 38956
rect 12492 38944 12498 38956
rect 13078 38944 13084 38956
rect 12492 38916 13084 38944
rect 12492 38904 12498 38916
rect 13078 38904 13084 38916
rect 13136 38904 13142 38956
rect 15194 38904 15200 38956
rect 15252 38944 15258 38956
rect 15361 38947 15419 38953
rect 15361 38944 15373 38947
rect 15252 38916 15373 38944
rect 15252 38904 15258 38916
rect 15361 38913 15373 38916
rect 15407 38913 15419 38947
rect 15361 38907 15419 38913
rect 16850 38904 16856 38956
rect 16908 38944 16914 38956
rect 17512 38953 17540 38984
rect 17770 38972 17776 39024
rect 17828 39012 17834 39024
rect 17828 38984 18736 39012
rect 17828 38972 17834 38984
rect 17221 38947 17279 38953
rect 17221 38944 17233 38947
rect 16908 38916 17233 38944
rect 16908 38904 16914 38916
rect 17221 38913 17233 38916
rect 17267 38913 17279 38947
rect 17221 38907 17279 38913
rect 17497 38947 17555 38953
rect 17497 38913 17509 38947
rect 17543 38913 17555 38947
rect 17497 38907 17555 38913
rect 17865 38947 17923 38953
rect 17865 38913 17877 38947
rect 17911 38944 17923 38947
rect 18046 38944 18052 38956
rect 17911 38916 18052 38944
rect 17911 38913 17923 38916
rect 17865 38907 17923 38913
rect 18046 38904 18052 38916
rect 18104 38904 18110 38956
rect 18141 38947 18199 38953
rect 18141 38913 18153 38947
rect 18187 38944 18199 38947
rect 18322 38944 18328 38956
rect 18187 38916 18328 38944
rect 18187 38913 18199 38916
rect 18141 38907 18199 38913
rect 18322 38904 18328 38916
rect 18380 38904 18386 38956
rect 18414 38904 18420 38956
rect 18472 38953 18478 38956
rect 18708 38953 18736 38984
rect 18472 38944 18483 38953
rect 18693 38947 18751 38953
rect 18472 38916 18517 38944
rect 18472 38907 18483 38916
rect 18693 38913 18705 38947
rect 18739 38913 18751 38947
rect 18693 38907 18751 38913
rect 18969 38947 19027 38953
rect 18969 38913 18981 38947
rect 19015 38944 19027 38947
rect 19168 38944 19196 39052
rect 19242 39040 19248 39092
rect 19300 39040 19306 39092
rect 19429 39083 19487 39089
rect 19429 39049 19441 39083
rect 19475 39080 19487 39083
rect 19610 39080 19616 39092
rect 19475 39052 19616 39080
rect 19475 39049 19487 39052
rect 19429 39043 19487 39049
rect 19610 39040 19616 39052
rect 19668 39040 19674 39092
rect 20622 39080 20628 39092
rect 19720 39052 20628 39080
rect 19260 38953 19288 39040
rect 19015 38916 19196 38944
rect 19245 38947 19303 38953
rect 19015 38913 19027 38916
rect 18969 38907 19027 38913
rect 19245 38913 19257 38947
rect 19291 38913 19303 38947
rect 19245 38907 19303 38913
rect 18472 38904 18478 38907
rect 19334 38904 19340 38956
rect 19392 38944 19398 38956
rect 19613 38947 19671 38953
rect 19613 38944 19625 38947
rect 19392 38916 19625 38944
rect 19392 38904 19398 38916
rect 19613 38913 19625 38916
rect 19659 38913 19671 38947
rect 19613 38907 19671 38913
rect 1673 38879 1731 38885
rect 1673 38845 1685 38879
rect 1719 38845 1731 38879
rect 1673 38839 1731 38845
rect 1688 38740 1716 38839
rect 2314 38836 2320 38888
rect 2372 38876 2378 38888
rect 2685 38879 2743 38885
rect 2685 38876 2697 38879
rect 2372 38848 2697 38876
rect 2372 38836 2378 38848
rect 2685 38845 2697 38848
rect 2731 38845 2743 38879
rect 2685 38839 2743 38845
rect 3878 38836 3884 38888
rect 3936 38876 3942 38888
rect 4249 38879 4307 38885
rect 4249 38876 4261 38879
rect 3936 38848 4261 38876
rect 3936 38836 3942 38848
rect 4249 38845 4261 38848
rect 4295 38845 4307 38879
rect 4249 38839 4307 38845
rect 4706 38836 4712 38888
rect 4764 38836 4770 38888
rect 6546 38836 6552 38888
rect 6604 38876 6610 38888
rect 6733 38879 6791 38885
rect 6733 38876 6745 38879
rect 6604 38848 6745 38876
rect 6604 38836 6610 38848
rect 6733 38845 6745 38848
rect 6779 38845 6791 38879
rect 6733 38839 6791 38845
rect 6914 38836 6920 38888
rect 6972 38836 6978 38888
rect 7374 38836 7380 38888
rect 7432 38836 7438 38888
rect 7834 38885 7840 38888
rect 7653 38879 7711 38885
rect 7653 38876 7665 38879
rect 7484 38848 7665 38876
rect 4062 38808 4068 38820
rect 3620 38780 4068 38808
rect 3620 38740 3648 38780
rect 4062 38768 4068 38780
rect 4120 38768 4126 38820
rect 7484 38808 7512 38848
rect 7653 38845 7665 38848
rect 7699 38845 7711 38879
rect 7653 38839 7711 38845
rect 7791 38879 7840 38885
rect 7791 38845 7803 38879
rect 7837 38845 7840 38879
rect 7791 38839 7840 38845
rect 7834 38836 7840 38839
rect 7892 38836 7898 38888
rect 14090 38836 14096 38888
rect 14148 38876 14154 38888
rect 14642 38876 14648 38888
rect 14148 38848 14648 38876
rect 14148 38836 14154 38848
rect 14642 38836 14648 38848
rect 14700 38876 14706 38888
rect 15105 38879 15163 38885
rect 15105 38876 15117 38879
rect 14700 38848 15117 38876
rect 14700 38836 14706 38848
rect 15105 38845 15117 38848
rect 15151 38845 15163 38879
rect 19720 38876 19748 39052
rect 20622 39040 20628 39052
rect 20680 39040 20686 39092
rect 20070 38972 20076 39024
rect 20128 39012 20134 39024
rect 20165 39015 20223 39021
rect 20165 39012 20177 39015
rect 20128 38984 20177 39012
rect 20128 38972 20134 38984
rect 20165 38981 20177 38984
rect 20211 38981 20223 39015
rect 20165 38975 20223 38981
rect 19886 38904 19892 38956
rect 19944 38944 19950 38956
rect 19981 38947 20039 38953
rect 19981 38944 19993 38947
rect 19944 38916 19993 38944
rect 19944 38904 19950 38916
rect 19981 38913 19993 38916
rect 20027 38913 20039 38947
rect 19981 38907 20039 38913
rect 15105 38839 15163 38845
rect 18248 38848 19748 38876
rect 5828 38780 7512 38808
rect 17313 38811 17371 38817
rect 5828 38752 5856 38780
rect 17313 38777 17325 38811
rect 17359 38808 17371 38811
rect 18138 38808 18144 38820
rect 17359 38780 18144 38808
rect 17359 38777 17371 38780
rect 17313 38771 17371 38777
rect 18138 38768 18144 38780
rect 18196 38768 18202 38820
rect 18248 38817 18276 38848
rect 20346 38836 20352 38888
rect 20404 38836 20410 38888
rect 18233 38811 18291 38817
rect 18233 38777 18245 38811
rect 18279 38777 18291 38811
rect 18233 38771 18291 38777
rect 18414 38768 18420 38820
rect 18472 38808 18478 38820
rect 19518 38808 19524 38820
rect 18472 38780 19524 38808
rect 18472 38768 18478 38780
rect 19518 38768 19524 38780
rect 19576 38768 19582 38820
rect 20364 38808 20392 38836
rect 19628 38780 20392 38808
rect 1688 38712 3648 38740
rect 3697 38743 3755 38749
rect 3697 38709 3709 38743
rect 3743 38740 3755 38743
rect 4154 38740 4160 38752
rect 3743 38712 4160 38740
rect 3743 38709 3755 38712
rect 3697 38703 3755 38709
rect 4154 38700 4160 38712
rect 4212 38700 4218 38752
rect 5810 38700 5816 38752
rect 5868 38700 5874 38752
rect 8573 38743 8631 38749
rect 8573 38709 8585 38743
rect 8619 38740 8631 38743
rect 13814 38740 13820 38752
rect 8619 38712 13820 38740
rect 8619 38709 8631 38712
rect 8573 38703 8631 38709
rect 13814 38700 13820 38712
rect 13872 38700 13878 38752
rect 17957 38743 18015 38749
rect 17957 38709 17969 38743
rect 18003 38740 18015 38743
rect 19628 38740 19656 38780
rect 18003 38712 19656 38740
rect 18003 38709 18015 38712
rect 17957 38703 18015 38709
rect 19702 38700 19708 38752
rect 19760 38740 19766 38752
rect 19797 38743 19855 38749
rect 19797 38740 19809 38743
rect 19760 38712 19809 38740
rect 19760 38700 19766 38712
rect 19797 38709 19809 38712
rect 19843 38709 19855 38743
rect 19797 38703 19855 38709
rect 20438 38700 20444 38752
rect 20496 38700 20502 38752
rect 1104 38650 20884 38672
rect 1104 38598 3422 38650
rect 3474 38598 3486 38650
rect 3538 38598 3550 38650
rect 3602 38598 3614 38650
rect 3666 38598 3678 38650
rect 3730 38598 8367 38650
rect 8419 38598 8431 38650
rect 8483 38598 8495 38650
rect 8547 38598 8559 38650
rect 8611 38598 8623 38650
rect 8675 38598 13312 38650
rect 13364 38598 13376 38650
rect 13428 38598 13440 38650
rect 13492 38598 13504 38650
rect 13556 38598 13568 38650
rect 13620 38598 18257 38650
rect 18309 38598 18321 38650
rect 18373 38598 18385 38650
rect 18437 38598 18449 38650
rect 18501 38598 18513 38650
rect 18565 38598 20884 38650
rect 1104 38576 20884 38598
rect 7282 38496 7288 38548
rect 7340 38536 7346 38548
rect 7340 38508 11192 38536
rect 7340 38496 7346 38508
rect 9674 38468 9680 38480
rect 5276 38440 9680 38468
rect 3792 38412 3844 38418
rect 5276 38412 5304 38440
rect 9674 38428 9680 38440
rect 9732 38428 9738 38480
rect 1578 38360 1584 38412
rect 1636 38400 1642 38412
rect 2314 38400 2320 38412
rect 1636 38372 2320 38400
rect 1636 38360 1642 38372
rect 2314 38360 2320 38372
rect 2372 38360 2378 38412
rect 5258 38360 5264 38412
rect 5316 38360 5322 38412
rect 6270 38360 6276 38412
rect 6328 38400 6334 38412
rect 10318 38400 10324 38412
rect 6328 38372 10324 38400
rect 6328 38360 6334 38372
rect 10318 38360 10324 38372
rect 10376 38360 10382 38412
rect 11164 38400 11192 38508
rect 15212 38508 16252 38536
rect 15212 38480 15240 38508
rect 15194 38428 15200 38480
rect 15252 38428 15258 38480
rect 15473 38471 15531 38477
rect 15473 38437 15485 38471
rect 15519 38437 15531 38471
rect 15473 38431 15531 38437
rect 11164 38372 14228 38400
rect 3792 38354 3844 38360
rect 1118 38292 1124 38344
rect 1176 38332 1182 38344
rect 1397 38335 1455 38341
rect 1397 38332 1409 38335
rect 1176 38304 1409 38332
rect 1176 38292 1182 38304
rect 1397 38301 1409 38304
rect 1443 38301 1455 38335
rect 1397 38295 1455 38301
rect 2591 38335 2649 38341
rect 2591 38301 2603 38335
rect 2637 38332 2649 38335
rect 2682 38332 2688 38344
rect 2637 38304 2688 38332
rect 2637 38301 2649 38304
rect 2591 38295 2649 38301
rect 2682 38292 2688 38304
rect 2740 38292 2746 38344
rect 4154 38292 4160 38344
rect 4212 38332 4218 38344
rect 4341 38335 4399 38341
rect 4341 38332 4353 38335
rect 4212 38304 4353 38332
rect 4212 38292 4218 38304
rect 4341 38301 4353 38304
rect 4387 38301 4399 38335
rect 4798 38332 4804 38344
rect 4341 38295 4399 38301
rect 4448 38304 4804 38332
rect 1670 38224 1676 38276
rect 1728 38224 1734 38276
rect 4249 38267 4307 38273
rect 4249 38233 4261 38267
rect 4295 38264 4307 38267
rect 4448 38264 4476 38304
rect 4798 38292 4804 38304
rect 4856 38292 4862 38344
rect 4890 38292 4896 38344
rect 4948 38332 4954 38344
rect 5626 38332 5632 38344
rect 4948 38304 5632 38332
rect 4948 38292 4954 38304
rect 5626 38292 5632 38304
rect 5684 38292 5690 38344
rect 9766 38292 9772 38344
rect 9824 38332 9830 38344
rect 10502 38332 10508 38344
rect 9824 38304 10508 38332
rect 9824 38292 9830 38304
rect 10502 38292 10508 38304
rect 10560 38292 10566 38344
rect 10778 38332 10784 38344
rect 10739 38304 10784 38332
rect 10778 38292 10784 38304
rect 10836 38292 10842 38344
rect 12250 38332 12256 38344
rect 11992 38304 12256 38332
rect 4295 38236 4476 38264
rect 4709 38267 4767 38273
rect 4295 38233 4307 38236
rect 4249 38227 4307 38233
rect 4709 38233 4721 38267
rect 4755 38264 4767 38267
rect 4982 38264 4988 38276
rect 4755 38236 4988 38264
rect 4755 38233 4767 38236
rect 4709 38227 4767 38233
rect 4982 38224 4988 38236
rect 5040 38264 5046 38276
rect 5166 38264 5172 38276
rect 5040 38236 5172 38264
rect 5040 38224 5046 38236
rect 5166 38224 5172 38236
rect 5224 38224 5230 38276
rect 9950 38224 9956 38276
rect 10008 38264 10014 38276
rect 11992 38273 12020 38304
rect 12250 38292 12256 38304
rect 12308 38292 12314 38344
rect 13814 38292 13820 38344
rect 13872 38332 13878 38344
rect 13909 38335 13967 38341
rect 13909 38332 13921 38335
rect 13872 38304 13921 38332
rect 13872 38292 13878 38304
rect 13909 38301 13921 38304
rect 13955 38301 13967 38335
rect 13909 38295 13967 38301
rect 11977 38267 12035 38273
rect 11977 38264 11989 38267
rect 10008 38236 11989 38264
rect 10008 38224 10014 38236
rect 11977 38233 11989 38236
rect 12023 38233 12035 38267
rect 11977 38227 12035 38233
rect 12158 38224 12164 38276
rect 12216 38224 12222 38276
rect 12434 38224 12440 38276
rect 12492 38264 12498 38276
rect 13924 38264 13952 38295
rect 14090 38292 14096 38344
rect 14148 38292 14154 38344
rect 14200 38332 14228 38372
rect 15488 38332 15516 38431
rect 16224 38341 16252 38508
rect 16390 38496 16396 38548
rect 16448 38536 16454 38548
rect 18322 38536 18328 38548
rect 16448 38508 18328 38536
rect 16448 38496 16454 38508
rect 18322 38496 18328 38508
rect 18380 38496 18386 38548
rect 18509 38539 18567 38545
rect 18509 38505 18521 38539
rect 18555 38536 18567 38539
rect 19242 38536 19248 38548
rect 18555 38508 19248 38536
rect 18555 38505 18567 38508
rect 18509 38499 18567 38505
rect 19242 38496 19248 38508
rect 19300 38496 19306 38548
rect 19352 38508 19564 38536
rect 18233 38471 18291 38477
rect 18233 38437 18245 38471
rect 18279 38437 18291 38471
rect 18233 38431 18291 38437
rect 18877 38471 18935 38477
rect 18877 38437 18889 38471
rect 18923 38468 18935 38471
rect 19352 38468 19380 38508
rect 18923 38440 19380 38468
rect 18923 38437 18935 38440
rect 18877 38431 18935 38437
rect 16853 38403 16911 38409
rect 16853 38369 16865 38403
rect 16899 38400 16911 38403
rect 18248 38400 18276 38431
rect 19426 38428 19432 38480
rect 19484 38428 19490 38480
rect 19536 38468 19564 38508
rect 19794 38496 19800 38548
rect 19852 38536 19858 38548
rect 19852 38508 20208 38536
rect 19852 38496 19858 38508
rect 19978 38468 19984 38480
rect 19536 38440 19984 38468
rect 19978 38428 19984 38440
rect 20036 38428 20042 38480
rect 19444 38400 19472 38428
rect 20070 38400 20076 38412
rect 16899 38372 17540 38400
rect 18248 38372 19472 38400
rect 19812 38372 20076 38400
rect 16899 38369 16911 38372
rect 16853 38363 16911 38369
rect 17512 38341 17540 38372
rect 15749 38335 15807 38341
rect 15749 38332 15761 38335
rect 14200 38304 15056 38332
rect 15488 38304 15761 38332
rect 15028 38276 15056 38304
rect 15749 38301 15761 38304
rect 15795 38301 15807 38335
rect 15749 38295 15807 38301
rect 16209 38335 16267 38341
rect 16209 38301 16221 38335
rect 16255 38301 16267 38335
rect 16209 38295 16267 38301
rect 16761 38335 16819 38341
rect 16761 38301 16773 38335
rect 16807 38301 16819 38335
rect 16761 38295 16819 38301
rect 17497 38335 17555 38341
rect 17497 38301 17509 38335
rect 17543 38301 17555 38335
rect 17497 38295 17555 38301
rect 14338 38267 14396 38273
rect 14338 38264 14350 38267
rect 12492 38236 13860 38264
rect 13924 38236 14350 38264
rect 12492 38224 12498 38236
rect 3326 38156 3332 38208
rect 3384 38156 3390 38208
rect 3973 38199 4031 38205
rect 3973 38165 3985 38199
rect 4019 38196 4031 38199
rect 4154 38196 4160 38208
rect 4019 38168 4160 38196
rect 4019 38165 4031 38168
rect 3973 38159 4031 38165
rect 4154 38156 4160 38168
rect 4212 38196 4218 38208
rect 4614 38196 4620 38208
rect 4212 38168 4620 38196
rect 4212 38156 4218 38168
rect 4614 38156 4620 38168
rect 4672 38156 4678 38208
rect 4890 38156 4896 38208
rect 4948 38196 4954 38208
rect 5077 38199 5135 38205
rect 5077 38196 5089 38199
rect 4948 38168 5089 38196
rect 4948 38156 4954 38168
rect 5077 38165 5089 38168
rect 5123 38165 5135 38199
rect 5077 38159 5135 38165
rect 5258 38156 5264 38208
rect 5316 38156 5322 38208
rect 9122 38156 9128 38208
rect 9180 38196 9186 38208
rect 10410 38196 10416 38208
rect 9180 38168 10416 38196
rect 9180 38156 9186 38168
rect 10410 38156 10416 38168
rect 10468 38156 10474 38208
rect 10502 38156 10508 38208
rect 10560 38196 10566 38208
rect 10778 38196 10784 38208
rect 10560 38168 10784 38196
rect 10560 38156 10566 38168
rect 10778 38156 10784 38168
rect 10836 38156 10842 38208
rect 11514 38156 11520 38208
rect 11572 38156 11578 38208
rect 13722 38156 13728 38208
rect 13780 38156 13786 38208
rect 13832 38196 13860 38236
rect 14338 38233 14350 38236
rect 14384 38233 14396 38267
rect 14338 38227 14396 38233
rect 15010 38224 15016 38276
rect 15068 38224 15074 38276
rect 16776 38264 16804 38295
rect 17678 38292 17684 38344
rect 17736 38332 17742 38344
rect 17957 38335 18015 38341
rect 17957 38332 17969 38335
rect 17736 38304 17969 38332
rect 17736 38292 17742 38304
rect 17957 38301 17969 38304
rect 18003 38301 18015 38335
rect 17957 38295 18015 38301
rect 18138 38292 18144 38344
rect 18196 38292 18202 38344
rect 18322 38292 18328 38344
rect 18380 38332 18386 38344
rect 18417 38335 18475 38341
rect 18417 38332 18429 38335
rect 18380 38304 18429 38332
rect 18380 38292 18386 38304
rect 18417 38301 18429 38304
rect 18463 38301 18475 38335
rect 18417 38295 18475 38301
rect 18693 38335 18751 38341
rect 18693 38301 18705 38335
rect 18739 38301 18751 38335
rect 19061 38335 19119 38341
rect 19061 38332 19073 38335
rect 18693 38295 18751 38301
rect 18984 38304 19073 38332
rect 16040 38236 16804 38264
rect 15470 38196 15476 38208
rect 13832 38168 15476 38196
rect 15470 38156 15476 38168
rect 15528 38156 15534 38208
rect 15562 38156 15568 38208
rect 15620 38156 15626 38208
rect 16040 38205 16068 38236
rect 17770 38224 17776 38276
rect 17828 38224 17834 38276
rect 17865 38267 17923 38273
rect 17865 38233 17877 38267
rect 17911 38264 17923 38267
rect 18049 38267 18107 38273
rect 18049 38264 18061 38267
rect 17911 38236 18061 38264
rect 17911 38233 17923 38236
rect 17865 38227 17923 38233
rect 18049 38233 18061 38236
rect 18095 38233 18107 38267
rect 18049 38227 18107 38233
rect 16025 38199 16083 38205
rect 16025 38165 16037 38199
rect 16071 38165 16083 38199
rect 16025 38159 16083 38165
rect 18138 38156 18144 38208
rect 18196 38196 18202 38208
rect 18708 38196 18736 38295
rect 18984 38208 19012 38304
rect 19061 38301 19073 38304
rect 19107 38301 19119 38335
rect 19061 38295 19119 38301
rect 19426 38292 19432 38344
rect 19484 38292 19490 38344
rect 19518 38292 19524 38344
rect 19576 38292 19582 38344
rect 19812 38341 19840 38372
rect 20070 38360 20076 38372
rect 20128 38360 20134 38412
rect 20180 38341 20208 38508
rect 19797 38335 19855 38341
rect 19797 38301 19809 38335
rect 19843 38301 19855 38335
rect 19797 38295 19855 38301
rect 19981 38335 20039 38341
rect 19981 38301 19993 38335
rect 20027 38301 20039 38335
rect 19981 38295 20039 38301
rect 20165 38335 20223 38341
rect 20165 38301 20177 38335
rect 20211 38301 20223 38335
rect 20165 38295 20223 38301
rect 19996 38264 20024 38295
rect 19260 38236 20024 38264
rect 20533 38267 20591 38273
rect 18196 38168 18736 38196
rect 18196 38156 18202 38168
rect 18966 38156 18972 38208
rect 19024 38156 19030 38208
rect 19260 38205 19288 38236
rect 20533 38233 20545 38267
rect 20579 38264 20591 38267
rect 21266 38264 21272 38276
rect 20579 38236 21272 38264
rect 20579 38233 20591 38236
rect 20533 38227 20591 38233
rect 21266 38224 21272 38236
rect 21324 38224 21330 38276
rect 19245 38199 19303 38205
rect 19245 38165 19257 38199
rect 19291 38165 19303 38199
rect 19245 38159 19303 38165
rect 19610 38156 19616 38208
rect 19668 38156 19674 38208
rect 19978 38156 19984 38208
rect 20036 38156 20042 38208
rect 1104 38106 21043 38128
rect 1104 38054 5894 38106
rect 5946 38054 5958 38106
rect 6010 38054 6022 38106
rect 6074 38054 6086 38106
rect 6138 38054 6150 38106
rect 6202 38054 10839 38106
rect 10891 38054 10903 38106
rect 10955 38054 10967 38106
rect 11019 38054 11031 38106
rect 11083 38054 11095 38106
rect 11147 38054 15784 38106
rect 15836 38054 15848 38106
rect 15900 38054 15912 38106
rect 15964 38054 15976 38106
rect 16028 38054 16040 38106
rect 16092 38054 20729 38106
rect 20781 38054 20793 38106
rect 20845 38054 20857 38106
rect 20909 38054 20921 38106
rect 20973 38054 20985 38106
rect 21037 38054 21043 38106
rect 1104 38032 21043 38054
rect 2869 37995 2927 38001
rect 2869 37961 2881 37995
rect 2915 37992 2927 37995
rect 3973 37995 4031 38001
rect 2915 37964 3924 37992
rect 2915 37961 2927 37964
rect 2869 37955 2927 37961
rect 1673 37927 1731 37933
rect 1673 37893 1685 37927
rect 1719 37924 1731 37927
rect 3237 37927 3295 37933
rect 1719 37896 3004 37924
rect 1719 37893 1731 37896
rect 1673 37887 1731 37893
rect 2976 37868 3004 37896
rect 3237 37893 3249 37927
rect 3283 37924 3295 37927
rect 3326 37924 3332 37936
rect 3283 37896 3332 37924
rect 3283 37893 3295 37896
rect 3237 37887 3295 37893
rect 3326 37884 3332 37896
rect 3384 37884 3390 37936
rect 3786 37924 3792 37936
rect 3528 37896 3792 37924
rect 1397 37859 1455 37865
rect 1397 37825 1409 37859
rect 1443 37825 1455 37859
rect 1397 37819 1455 37825
rect 1412 37732 1440 37819
rect 1854 37816 1860 37868
rect 1912 37856 1918 37868
rect 1949 37859 2007 37865
rect 1949 37856 1961 37859
rect 1912 37828 1961 37856
rect 1912 37816 1918 37828
rect 1949 37825 1961 37828
rect 1995 37825 2007 37859
rect 1949 37819 2007 37825
rect 2958 37816 2964 37868
rect 3016 37816 3022 37868
rect 3145 37859 3203 37865
rect 3145 37825 3157 37859
rect 3191 37856 3203 37859
rect 3528 37856 3556 37896
rect 3786 37884 3792 37896
rect 3844 37884 3850 37936
rect 3896 37924 3924 37964
rect 3973 37961 3985 37995
rect 4019 37992 4031 37995
rect 4019 37964 4476 37992
rect 4019 37961 4031 37964
rect 3973 37955 4031 37961
rect 4154 37924 4160 37936
rect 3896 37896 4160 37924
rect 4154 37884 4160 37896
rect 4212 37884 4218 37936
rect 4448 37924 4476 37964
rect 4522 37952 4528 38004
rect 4580 37992 4586 38004
rect 5353 37995 5411 38001
rect 5353 37992 5365 37995
rect 4580 37964 5365 37992
rect 4580 37952 4586 37964
rect 5353 37961 5365 37964
rect 5399 37961 5411 37995
rect 5353 37955 5411 37961
rect 6454 37952 6460 38004
rect 6512 37992 6518 38004
rect 9674 37992 9680 38004
rect 6512 37964 9680 37992
rect 6512 37952 6518 37964
rect 9674 37952 9680 37964
rect 9732 37952 9738 38004
rect 9950 37952 9956 38004
rect 10008 37952 10014 38004
rect 10318 37952 10324 38004
rect 10376 37952 10382 38004
rect 10594 37952 10600 38004
rect 10652 37992 10658 38004
rect 11514 37992 11520 38004
rect 10652 37964 11520 37992
rect 10652 37952 10658 37964
rect 11514 37952 11520 37964
rect 11572 37952 11578 38004
rect 12529 37995 12587 38001
rect 12529 37961 12541 37995
rect 12575 37961 12587 37995
rect 12529 37955 12587 37961
rect 6270 37924 6276 37936
rect 4448 37896 4936 37924
rect 4908 37868 4936 37896
rect 5552 37896 6276 37924
rect 5552 37868 5580 37896
rect 6270 37884 6276 37896
rect 6328 37884 6334 37936
rect 10226 37884 10232 37936
rect 10284 37884 10290 37936
rect 10336 37924 10364 37952
rect 11057 37927 11115 37933
rect 11057 37924 11069 37927
rect 10336 37896 11069 37924
rect 11057 37893 11069 37896
rect 11103 37893 11115 37927
rect 12544 37924 12572 37955
rect 13722 37952 13728 38004
rect 13780 37952 13786 38004
rect 14366 37952 14372 38004
rect 14424 37992 14430 38004
rect 15470 37992 15476 38004
rect 14424 37964 15476 37992
rect 14424 37952 14430 37964
rect 15470 37952 15476 37964
rect 15528 37952 15534 38004
rect 15562 37952 15568 38004
rect 15620 37952 15626 38004
rect 15764 37964 17356 37992
rect 11057 37887 11115 37893
rect 11624 37896 12572 37924
rect 3191 37828 3556 37856
rect 3605 37859 3663 37865
rect 3191 37825 3203 37828
rect 3145 37819 3203 37825
rect 3605 37825 3617 37859
rect 3651 37856 3663 37859
rect 3651 37828 4844 37856
rect 3651 37825 3663 37828
rect 3605 37819 3663 37825
rect 2225 37791 2283 37797
rect 2225 37757 2237 37791
rect 2271 37788 2283 37791
rect 2314 37788 2320 37800
rect 2271 37760 2320 37788
rect 2271 37757 2283 37760
rect 2225 37751 2283 37757
rect 2314 37748 2320 37760
rect 2372 37748 2378 37800
rect 2774 37748 2780 37800
rect 2832 37748 2838 37800
rect 4816 37788 4844 37828
rect 4890 37816 4896 37868
rect 4948 37816 4954 37868
rect 5534 37816 5540 37868
rect 5592 37816 5598 37868
rect 6638 37816 6644 37868
rect 6696 37856 6702 37868
rect 7283 37859 7341 37865
rect 7283 37856 7295 37859
rect 6696 37828 7295 37856
rect 6696 37816 6702 37828
rect 7283 37825 7295 37828
rect 7329 37825 7341 37859
rect 7283 37819 7341 37825
rect 7374 37816 7380 37868
rect 7432 37856 7438 37868
rect 10042 37856 10048 37868
rect 7432 37828 10048 37856
rect 7432 37816 7438 37828
rect 10042 37816 10048 37828
rect 10100 37816 10106 37868
rect 10321 37859 10379 37865
rect 10321 37825 10333 37859
rect 10367 37856 10379 37859
rect 10594 37856 10600 37868
rect 10367 37828 10600 37856
rect 10367 37825 10379 37828
rect 10321 37819 10379 37825
rect 10594 37816 10600 37828
rect 10652 37816 10658 37868
rect 10689 37859 10747 37865
rect 10689 37825 10701 37859
rect 10735 37856 10747 37859
rect 10778 37856 10784 37868
rect 10735 37828 10784 37856
rect 10735 37825 10747 37828
rect 10689 37819 10747 37825
rect 10778 37816 10784 37828
rect 10836 37816 10842 37868
rect 11624 37856 11652 37896
rect 10980 37828 11652 37856
rect 11791 37859 11849 37865
rect 5350 37788 5356 37800
rect 4816 37760 5356 37788
rect 5350 37748 5356 37760
rect 5408 37748 5414 37800
rect 5902 37748 5908 37800
rect 5960 37788 5966 37800
rect 7009 37791 7067 37797
rect 7009 37788 7021 37791
rect 5960 37760 7021 37788
rect 5960 37748 5966 37760
rect 7009 37757 7021 37760
rect 7055 37757 7067 37791
rect 10980 37774 11008 37828
rect 11791 37825 11803 37859
rect 11837 37856 11849 37859
rect 11882 37856 11888 37868
rect 11837 37828 11888 37856
rect 11837 37825 11849 37828
rect 11791 37819 11849 37825
rect 11882 37816 11888 37828
rect 11940 37856 11946 37868
rect 13740 37856 13768 37952
rect 15212 37896 15516 37924
rect 14461 37859 14519 37865
rect 14461 37856 14473 37859
rect 11940 37828 13124 37856
rect 13740 37828 14473 37856
rect 11940 37816 11946 37828
rect 7009 37751 7067 37757
rect 11514 37748 11520 37800
rect 11572 37748 11578 37800
rect 1394 37680 1400 37732
rect 1452 37680 1458 37732
rect 9030 37720 9036 37732
rect 7668 37692 9036 37720
rect 4154 37612 4160 37664
rect 4212 37612 4218 37664
rect 6362 37612 6368 37664
rect 6420 37652 6426 37664
rect 6730 37652 6736 37664
rect 6420 37624 6736 37652
rect 6420 37612 6426 37624
rect 6730 37612 6736 37624
rect 6788 37612 6794 37664
rect 7466 37612 7472 37664
rect 7524 37652 7530 37664
rect 7668 37652 7696 37692
rect 9030 37680 9036 37692
rect 9088 37720 9094 37732
rect 9582 37720 9588 37732
rect 9088 37692 9588 37720
rect 9088 37680 9094 37692
rect 9582 37680 9588 37692
rect 9640 37680 9646 37732
rect 7524 37624 7696 37652
rect 7524 37612 7530 37624
rect 7926 37612 7932 37664
rect 7984 37652 7990 37664
rect 8021 37655 8079 37661
rect 8021 37652 8033 37655
rect 7984 37624 8033 37652
rect 7984 37612 7990 37624
rect 8021 37621 8033 37624
rect 8067 37621 8079 37655
rect 8021 37615 8079 37621
rect 8754 37612 8760 37664
rect 8812 37652 8818 37664
rect 8941 37655 8999 37661
rect 8941 37652 8953 37655
rect 8812 37624 8953 37652
rect 8812 37612 8818 37624
rect 8941 37621 8953 37624
rect 8987 37621 8999 37655
rect 8941 37615 8999 37621
rect 9214 37612 9220 37664
rect 9272 37652 9278 37664
rect 9490 37652 9496 37664
rect 9272 37624 9496 37652
rect 9272 37612 9278 37624
rect 9490 37612 9496 37624
rect 9548 37612 9554 37664
rect 11241 37655 11299 37661
rect 11241 37621 11253 37655
rect 11287 37652 11299 37655
rect 12986 37652 12992 37664
rect 11287 37624 12992 37652
rect 11287 37621 11299 37624
rect 11241 37615 11299 37621
rect 12986 37612 12992 37624
rect 13044 37612 13050 37664
rect 13096 37652 13124 37828
rect 14461 37825 14473 37828
rect 14507 37825 14519 37859
rect 14461 37819 14519 37825
rect 14553 37859 14611 37865
rect 14553 37825 14565 37859
rect 14599 37856 14611 37859
rect 15013 37859 15071 37865
rect 15013 37856 15025 37859
rect 14599 37828 15025 37856
rect 14599 37825 14611 37828
rect 14553 37819 14611 37825
rect 15013 37825 15025 37828
rect 15059 37825 15071 37859
rect 15013 37819 15071 37825
rect 15102 37816 15108 37868
rect 15160 37856 15166 37868
rect 15212 37865 15240 37896
rect 15197 37859 15255 37865
rect 15197 37856 15209 37859
rect 15160 37828 15209 37856
rect 15160 37816 15166 37828
rect 15197 37825 15209 37828
rect 15243 37825 15255 37859
rect 15197 37819 15255 37825
rect 15286 37816 15292 37868
rect 15344 37816 15350 37868
rect 15488 37865 15516 37896
rect 15381 37859 15439 37865
rect 15381 37825 15393 37859
rect 15427 37825 15439 37859
rect 15381 37819 15439 37825
rect 15473 37859 15531 37865
rect 15473 37825 15485 37859
rect 15519 37825 15531 37859
rect 15580 37856 15608 37952
rect 15657 37859 15715 37865
rect 15657 37856 15669 37859
rect 15580 37828 15669 37856
rect 15473 37819 15531 37825
rect 15657 37825 15669 37828
rect 15703 37825 15715 37859
rect 15657 37819 15715 37825
rect 13906 37748 13912 37800
rect 13964 37788 13970 37800
rect 15396 37788 15424 37819
rect 15565 37791 15623 37797
rect 15565 37788 15577 37791
rect 13964 37760 15332 37788
rect 15396 37760 15577 37788
rect 13964 37748 13970 37760
rect 15304 37720 15332 37760
rect 15565 37757 15577 37760
rect 15611 37757 15623 37791
rect 15565 37751 15623 37757
rect 15764 37720 15792 37964
rect 17328 37924 17356 37964
rect 17678 37952 17684 38004
rect 17736 37952 17742 38004
rect 18693 37995 18751 38001
rect 18693 37961 18705 37995
rect 18739 37961 18751 37995
rect 18693 37955 18751 37961
rect 19245 37995 19303 38001
rect 19245 37961 19257 37995
rect 19291 37992 19303 37995
rect 19518 37992 19524 38004
rect 19291 37964 19524 37992
rect 19291 37961 19303 37964
rect 19245 37955 19303 37961
rect 18138 37924 18144 37936
rect 17328 37896 18144 37924
rect 18138 37884 18144 37896
rect 18196 37884 18202 37936
rect 18708 37924 18736 37955
rect 19518 37952 19524 37964
rect 19576 37952 19582 38004
rect 20254 37952 20260 38004
rect 20312 37952 20318 38004
rect 19334 37924 19340 37936
rect 18708 37896 19340 37924
rect 19334 37884 19340 37896
rect 19392 37884 19398 37936
rect 20272 37924 20300 37952
rect 19812 37896 20300 37924
rect 15838 37816 15844 37868
rect 15896 37856 15902 37868
rect 16943 37859 17001 37865
rect 16943 37856 16955 37859
rect 15896 37828 16955 37856
rect 15896 37816 15902 37828
rect 16943 37825 16955 37828
rect 16989 37856 17001 37859
rect 17862 37856 17868 37868
rect 16989 37828 17868 37856
rect 16989 37825 17001 37828
rect 16943 37819 17001 37825
rect 17862 37816 17868 37828
rect 17920 37816 17926 37868
rect 18877 37859 18935 37865
rect 18877 37825 18889 37859
rect 18923 37825 18935 37859
rect 18877 37819 18935 37825
rect 16482 37748 16488 37800
rect 16540 37788 16546 37800
rect 16666 37788 16672 37800
rect 16540 37760 16672 37788
rect 16540 37748 16546 37760
rect 16666 37748 16672 37760
rect 16724 37748 16730 37800
rect 18892 37720 18920 37819
rect 18966 37816 18972 37868
rect 19024 37856 19030 37868
rect 19153 37859 19211 37865
rect 19153 37856 19165 37859
rect 19024 37828 19165 37856
rect 19024 37816 19030 37828
rect 19153 37825 19165 37828
rect 19199 37825 19211 37859
rect 19153 37819 19211 37825
rect 19242 37816 19248 37868
rect 19300 37856 19306 37868
rect 19429 37859 19487 37865
rect 19429 37856 19441 37859
rect 19300 37828 19441 37856
rect 19300 37816 19306 37828
rect 19429 37825 19441 37828
rect 19475 37825 19487 37859
rect 19429 37819 19487 37825
rect 19518 37816 19524 37868
rect 19576 37856 19582 37868
rect 19705 37859 19763 37865
rect 19705 37856 19717 37859
rect 19576 37828 19717 37856
rect 19576 37816 19582 37828
rect 19705 37825 19717 37828
rect 19751 37825 19763 37859
rect 19705 37819 19763 37825
rect 19812 37788 19840 37896
rect 19981 37859 20039 37865
rect 19981 37825 19993 37859
rect 20027 37825 20039 37859
rect 19981 37819 20039 37825
rect 18984 37760 19840 37788
rect 18984 37729 19012 37760
rect 19886 37748 19892 37800
rect 19944 37748 19950 37800
rect 15304 37692 15792 37720
rect 17328 37692 18920 37720
rect 18969 37723 19027 37729
rect 17328 37652 17356 37692
rect 18969 37689 18981 37723
rect 19015 37689 19027 37723
rect 18969 37683 19027 37689
rect 19521 37723 19579 37729
rect 19521 37689 19533 37723
rect 19567 37720 19579 37723
rect 19904 37720 19932 37748
rect 19567 37692 19932 37720
rect 19567 37689 19579 37692
rect 19521 37683 19579 37689
rect 13096 37624 17356 37652
rect 17770 37612 17776 37664
rect 17828 37652 17834 37664
rect 19334 37652 19340 37664
rect 17828 37624 19340 37652
rect 17828 37612 17834 37624
rect 19334 37612 19340 37624
rect 19392 37612 19398 37664
rect 19794 37612 19800 37664
rect 19852 37612 19858 37664
rect 19886 37612 19892 37664
rect 19944 37652 19950 37664
rect 19996 37652 20024 37819
rect 20162 37816 20168 37868
rect 20220 37816 20226 37868
rect 19944 37624 20024 37652
rect 19944 37612 19950 37624
rect 20438 37612 20444 37664
rect 20496 37612 20502 37664
rect 1104 37562 20884 37584
rect 1104 37510 3422 37562
rect 3474 37510 3486 37562
rect 3538 37510 3550 37562
rect 3602 37510 3614 37562
rect 3666 37510 3678 37562
rect 3730 37510 8367 37562
rect 8419 37510 8431 37562
rect 8483 37510 8495 37562
rect 8547 37510 8559 37562
rect 8611 37510 8623 37562
rect 8675 37510 13312 37562
rect 13364 37510 13376 37562
rect 13428 37510 13440 37562
rect 13492 37510 13504 37562
rect 13556 37510 13568 37562
rect 13620 37510 18257 37562
rect 18309 37510 18321 37562
rect 18373 37510 18385 37562
rect 18437 37510 18449 37562
rect 18501 37510 18513 37562
rect 18565 37510 20884 37562
rect 1104 37488 20884 37510
rect 1026 37408 1032 37460
rect 1084 37448 1090 37460
rect 2685 37451 2743 37457
rect 1084 37420 2360 37448
rect 1084 37408 1090 37420
rect 1578 37272 1584 37324
rect 1636 37312 1642 37324
rect 1673 37315 1731 37321
rect 1673 37312 1685 37315
rect 1636 37284 1685 37312
rect 1636 37272 1642 37284
rect 1673 37281 1685 37284
rect 1719 37281 1731 37315
rect 2332 37312 2360 37420
rect 2685 37417 2697 37451
rect 2731 37448 2743 37451
rect 2774 37448 2780 37460
rect 2731 37420 2780 37448
rect 2731 37417 2743 37420
rect 2685 37411 2743 37417
rect 2774 37408 2780 37420
rect 2832 37408 2838 37460
rect 4062 37408 4068 37460
rect 4120 37448 4126 37460
rect 10594 37448 10600 37460
rect 4120 37420 10600 37448
rect 4120 37408 4126 37420
rect 10594 37408 10600 37420
rect 10652 37408 10658 37460
rect 11514 37448 11520 37460
rect 10704 37420 11520 37448
rect 3786 37340 3792 37392
rect 3844 37380 3850 37392
rect 5258 37380 5264 37392
rect 3844 37352 5264 37380
rect 3844 37340 3850 37352
rect 5258 37340 5264 37352
rect 5316 37340 5322 37392
rect 9674 37340 9680 37392
rect 9732 37380 9738 37392
rect 10704 37380 10732 37420
rect 11514 37408 11520 37420
rect 11572 37408 11578 37460
rect 13998 37408 14004 37460
rect 14056 37448 14062 37460
rect 14056 37420 14780 37448
rect 14056 37408 14062 37420
rect 9732 37352 10732 37380
rect 14752 37380 14780 37420
rect 15102 37408 15108 37460
rect 15160 37408 15166 37460
rect 18785 37451 18843 37457
rect 18785 37417 18797 37451
rect 18831 37448 18843 37451
rect 18966 37448 18972 37460
rect 18831 37420 18972 37448
rect 18831 37417 18843 37420
rect 18785 37411 18843 37417
rect 18966 37408 18972 37420
rect 19024 37408 19030 37460
rect 19150 37408 19156 37460
rect 19208 37448 19214 37460
rect 19208 37420 21864 37448
rect 19208 37408 19214 37420
rect 17586 37380 17592 37392
rect 14752 37352 17592 37380
rect 9732 37340 9738 37352
rect 17586 37340 17592 37352
rect 17644 37340 17650 37392
rect 18233 37383 18291 37389
rect 18233 37380 18245 37383
rect 18064 37352 18245 37380
rect 4062 37312 4068 37324
rect 2332 37284 4068 37312
rect 1673 37275 1731 37281
rect 4062 37272 4068 37284
rect 4120 37272 4126 37324
rect 5902 37272 5908 37324
rect 5960 37272 5966 37324
rect 7466 37272 7472 37324
rect 7524 37272 7530 37324
rect 12066 37272 12072 37324
rect 12124 37312 12130 37324
rect 13630 37312 13636 37324
rect 12124 37284 13636 37312
rect 12124 37272 12130 37284
rect 13630 37272 13636 37284
rect 13688 37272 13694 37324
rect 14093 37315 14151 37321
rect 14093 37281 14105 37315
rect 14139 37281 14151 37315
rect 14093 37275 14151 37281
rect 1947 37247 2005 37253
rect 1947 37213 1959 37247
rect 1993 37244 2005 37247
rect 2038 37244 2044 37256
rect 1993 37216 2044 37244
rect 1993 37213 2005 37216
rect 1947 37207 2005 37213
rect 2038 37204 2044 37216
rect 2096 37244 2102 37256
rect 2682 37244 2688 37256
rect 2096 37216 2688 37244
rect 2096 37204 2102 37216
rect 2682 37204 2688 37216
rect 2740 37204 2746 37256
rect 3053 37247 3111 37253
rect 3053 37213 3065 37247
rect 3099 37213 3111 37247
rect 3789 37247 3847 37253
rect 3789 37244 3801 37247
rect 3053 37207 3111 37213
rect 3252 37216 3801 37244
rect 1210 37136 1216 37188
rect 1268 37176 1274 37188
rect 3068 37176 3096 37207
rect 1268 37148 3096 37176
rect 1268 37136 1274 37148
rect 1302 37068 1308 37120
rect 1360 37108 1366 37120
rect 3252 37108 3280 37216
rect 3789 37213 3801 37216
rect 3835 37213 3847 37247
rect 3789 37207 3847 37213
rect 4246 37204 4252 37256
rect 4304 37244 4310 37256
rect 5258 37244 5264 37256
rect 4304 37216 5264 37244
rect 4304 37204 4310 37216
rect 5258 37204 5264 37216
rect 5316 37204 5322 37256
rect 3329 37179 3387 37185
rect 3329 37145 3341 37179
rect 3375 37145 3387 37179
rect 3329 37139 3387 37145
rect 4065 37179 4123 37185
rect 4065 37145 4077 37179
rect 4111 37176 4123 37179
rect 5442 37176 5448 37188
rect 4111 37148 5448 37176
rect 4111 37145 4123 37148
rect 4065 37139 4123 37145
rect 1360 37080 3280 37108
rect 3344 37108 3372 37139
rect 5442 37136 5448 37148
rect 5500 37136 5506 37188
rect 5534 37136 5540 37188
rect 5592 37176 5598 37188
rect 5920 37176 5948 37272
rect 6179 37247 6237 37253
rect 6179 37213 6191 37247
rect 6225 37244 6237 37247
rect 8941 37247 8999 37253
rect 6225 37216 6316 37244
rect 6225 37213 6237 37216
rect 6179 37207 6237 37213
rect 6288 37188 6316 37216
rect 6380 37234 7604 37244
rect 6380 37216 7650 37234
rect 6380 37188 6408 37216
rect 7576 37214 7650 37216
rect 7727 37217 7785 37223
rect 7727 37214 7739 37217
rect 7576 37206 7739 37214
rect 5592 37148 5948 37176
rect 5592 37136 5598 37148
rect 6270 37136 6276 37188
rect 6328 37136 6334 37188
rect 6362 37136 6368 37188
rect 6420 37136 6426 37188
rect 6730 37136 6736 37188
rect 6788 37136 6794 37188
rect 7622 37186 7739 37206
rect 7727 37183 7739 37186
rect 7773 37183 7785 37217
rect 8941 37213 8953 37247
rect 8987 37244 8999 37247
rect 9215 37247 9273 37253
rect 9030 37244 9036 37246
rect 8987 37216 9036 37244
rect 8987 37213 8999 37216
rect 8941 37207 8999 37213
rect 9030 37194 9036 37216
rect 9088 37194 9094 37246
rect 9215 37213 9227 37247
rect 9261 37244 9273 37247
rect 9261 37216 9444 37244
rect 9261 37213 9273 37216
rect 9215 37207 9273 37213
rect 9416 37188 9444 37216
rect 9950 37204 9956 37256
rect 10008 37244 10014 37256
rect 10778 37244 10784 37256
rect 10008 37216 10784 37244
rect 10008 37204 10014 37216
rect 10778 37204 10784 37216
rect 10836 37204 10842 37256
rect 11057 37247 11115 37253
rect 11057 37213 11069 37247
rect 11103 37213 11115 37247
rect 11057 37207 11115 37213
rect 7727 37177 7785 37183
rect 9398 37136 9404 37188
rect 9456 37136 9462 37188
rect 11072 37176 11100 37207
rect 11238 37204 11244 37256
rect 11296 37244 11302 37256
rect 11331 37247 11389 37253
rect 11331 37244 11343 37247
rect 11296 37216 11343 37244
rect 11296 37204 11302 37216
rect 11331 37213 11343 37216
rect 11377 37213 11389 37247
rect 11331 37207 11389 37213
rect 11072 37148 11836 37176
rect 6748 37108 6776 37136
rect 11808 37120 11836 37148
rect 13446 37136 13452 37188
rect 13504 37176 13510 37188
rect 14108 37176 14136 37275
rect 14367 37247 14425 37253
rect 14367 37213 14379 37247
rect 14413 37244 14425 37247
rect 15562 37244 15568 37256
rect 14413 37216 15568 37244
rect 14413 37213 14425 37216
rect 14367 37207 14425 37213
rect 15562 37204 15568 37216
rect 15620 37204 15626 37256
rect 16482 37204 16488 37256
rect 16540 37204 16546 37256
rect 16500 37176 16528 37204
rect 13504 37148 14136 37176
rect 13504 37136 13510 37148
rect 3344 37080 6776 37108
rect 1360 37068 1366 37080
rect 6914 37068 6920 37120
rect 6972 37068 6978 37120
rect 8478 37068 8484 37120
rect 8536 37068 8542 37120
rect 9030 37068 9036 37120
rect 9088 37108 9094 37120
rect 9953 37111 10011 37117
rect 9953 37108 9965 37111
rect 9088 37080 9965 37108
rect 9088 37068 9094 37080
rect 9953 37077 9965 37080
rect 9999 37077 10011 37111
rect 9953 37071 10011 37077
rect 11790 37068 11796 37120
rect 11848 37068 11854 37120
rect 12066 37068 12072 37120
rect 12124 37068 12130 37120
rect 14108 37108 14136 37148
rect 14658 37148 16528 37176
rect 18064 37176 18092 37352
rect 18233 37349 18245 37352
rect 18279 37349 18291 37383
rect 18509 37383 18567 37389
rect 18509 37380 18521 37383
rect 18233 37343 18291 37349
rect 18340 37352 18521 37380
rect 18340 37312 18368 37352
rect 18509 37349 18521 37352
rect 18555 37349 18567 37383
rect 19794 37380 19800 37392
rect 18509 37343 18567 37349
rect 18616 37352 19800 37380
rect 18616 37312 18644 37352
rect 19794 37340 19800 37352
rect 19852 37340 19858 37392
rect 21542 37380 21548 37392
rect 20180 37352 21548 37380
rect 18156 37284 18368 37312
rect 18432 37284 18644 37312
rect 18156 37253 18184 37284
rect 18432 37253 18460 37284
rect 19334 37272 19340 37324
rect 19392 37312 19398 37324
rect 20180 37312 20208 37352
rect 21542 37340 21548 37352
rect 21600 37340 21606 37392
rect 21836 37324 21864 37420
rect 19392 37284 20208 37312
rect 19392 37272 19398 37284
rect 20254 37272 20260 37324
rect 20312 37272 20318 37324
rect 21818 37272 21824 37324
rect 21876 37272 21882 37324
rect 18141 37247 18199 37253
rect 18141 37213 18153 37247
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 18417 37247 18475 37253
rect 18417 37213 18429 37247
rect 18463 37213 18475 37247
rect 18417 37207 18475 37213
rect 18690 37204 18696 37256
rect 18748 37204 18754 37256
rect 18782 37204 18788 37256
rect 18840 37244 18846 37256
rect 18966 37244 18972 37256
rect 18840 37216 18972 37244
rect 18840 37204 18846 37216
rect 18966 37204 18972 37216
rect 19024 37204 19030 37256
rect 19981 37247 20039 37253
rect 19981 37244 19993 37247
rect 19306 37216 19993 37244
rect 19306 37176 19334 37216
rect 19981 37213 19993 37216
rect 20027 37213 20039 37247
rect 19981 37207 20039 37213
rect 20162 37204 20168 37256
rect 20220 37204 20226 37256
rect 18064 37148 19334 37176
rect 19429 37179 19487 37185
rect 14658 37108 14686 37148
rect 19429 37145 19441 37179
rect 19475 37176 19487 37179
rect 19702 37176 19708 37188
rect 19475 37148 19708 37176
rect 19475 37145 19487 37148
rect 19429 37139 19487 37145
rect 19702 37136 19708 37148
rect 19760 37136 19766 37188
rect 19794 37136 19800 37188
rect 19852 37136 19858 37188
rect 14108 37080 14686 37108
rect 15838 37068 15844 37120
rect 15896 37108 15902 37120
rect 17310 37108 17316 37120
rect 15896 37080 17316 37108
rect 15896 37068 15902 37080
rect 17310 37068 17316 37080
rect 17368 37068 17374 37120
rect 17957 37111 18015 37117
rect 17957 37077 17969 37111
rect 18003 37108 18015 37111
rect 20180 37108 20208 37204
rect 18003 37080 20208 37108
rect 18003 37077 18015 37080
rect 17957 37071 18015 37077
rect 1104 37018 21043 37040
rect 1104 36966 5894 37018
rect 5946 36966 5958 37018
rect 6010 36966 6022 37018
rect 6074 36966 6086 37018
rect 6138 36966 6150 37018
rect 6202 36966 10839 37018
rect 10891 36966 10903 37018
rect 10955 36966 10967 37018
rect 11019 36966 11031 37018
rect 11083 36966 11095 37018
rect 11147 36966 15784 37018
rect 15836 36966 15848 37018
rect 15900 36966 15912 37018
rect 15964 36966 15976 37018
rect 16028 36966 16040 37018
rect 16092 36966 20729 37018
rect 20781 36966 20793 37018
rect 20845 36966 20857 37018
rect 20909 36966 20921 37018
rect 20973 36966 20985 37018
rect 21037 36966 21043 37018
rect 1104 36944 21043 36966
rect 3050 36864 3056 36916
rect 3108 36904 3114 36916
rect 6270 36904 6276 36916
rect 3108 36876 6276 36904
rect 3108 36864 3114 36876
rect 658 36796 664 36848
rect 716 36836 722 36848
rect 1762 36836 1768 36848
rect 716 36808 1768 36836
rect 716 36796 722 36808
rect 1762 36796 1768 36808
rect 1820 36796 1826 36848
rect 3344 36845 3372 36876
rect 6270 36864 6276 36876
rect 6328 36904 6334 36916
rect 9677 36907 9735 36913
rect 6328 36876 9536 36904
rect 6328 36864 6334 36876
rect 3329 36839 3387 36845
rect 3329 36805 3341 36839
rect 3375 36805 3387 36839
rect 6638 36836 6644 36848
rect 3329 36799 3387 36805
rect 3804 36808 6644 36836
rect 1486 36728 1492 36780
rect 1544 36728 1550 36780
rect 1946 36728 1952 36780
rect 2004 36728 2010 36780
rect 3053 36771 3111 36777
rect 3053 36768 3065 36771
rect 2056 36740 3065 36768
rect 1210 36660 1216 36712
rect 1268 36700 1274 36712
rect 2056 36700 2084 36740
rect 3053 36737 3065 36740
rect 3099 36737 3111 36771
rect 3053 36731 3111 36737
rect 3605 36771 3663 36777
rect 3605 36737 3617 36771
rect 3651 36737 3663 36771
rect 3605 36731 3663 36737
rect 1268 36672 2084 36700
rect 2777 36703 2835 36709
rect 1268 36660 1274 36672
rect 2777 36669 2789 36703
rect 2823 36700 2835 36703
rect 3326 36700 3332 36712
rect 2823 36672 3332 36700
rect 2823 36669 2835 36672
rect 2777 36663 2835 36669
rect 3326 36660 3332 36672
rect 3384 36660 3390 36712
rect 1302 36592 1308 36644
rect 1360 36632 1366 36644
rect 3620 36632 3648 36731
rect 3804 36709 3832 36808
rect 6638 36796 6644 36808
rect 6696 36796 6702 36848
rect 9508 36836 9536 36876
rect 9677 36873 9689 36907
rect 9723 36904 9735 36907
rect 17957 36907 18015 36913
rect 9723 36876 15424 36904
rect 9723 36873 9735 36876
rect 9677 36867 9735 36873
rect 10410 36836 10416 36848
rect 9508 36808 10416 36836
rect 10410 36796 10416 36808
rect 10468 36796 10474 36848
rect 13722 36796 13728 36848
rect 13780 36796 13786 36848
rect 13998 36807 14004 36848
rect 13983 36801 14004 36807
rect 4246 36728 4252 36780
rect 4304 36728 4310 36780
rect 5350 36728 5356 36780
rect 5408 36728 5414 36780
rect 5442 36728 5448 36780
rect 5500 36768 5506 36780
rect 7466 36768 7472 36780
rect 5500 36740 7472 36768
rect 5500 36728 5506 36740
rect 7466 36728 7472 36740
rect 7524 36728 7530 36780
rect 8754 36728 8760 36780
rect 8812 36728 8818 36780
rect 9030 36728 9036 36780
rect 9088 36728 9094 36780
rect 9674 36728 9680 36780
rect 9732 36768 9738 36780
rect 10042 36768 10048 36780
rect 9732 36740 10048 36768
rect 9732 36728 9738 36740
rect 10042 36728 10048 36740
rect 10100 36728 10106 36780
rect 11422 36728 11428 36780
rect 11480 36768 11486 36780
rect 11791 36771 11849 36777
rect 11791 36768 11803 36771
rect 11480 36740 11803 36768
rect 11480 36728 11486 36740
rect 11791 36737 11803 36740
rect 11837 36768 11849 36771
rect 13740 36768 13768 36796
rect 11837 36740 13768 36768
rect 13983 36767 13995 36801
rect 14056 36796 14062 36848
rect 15396 36836 15424 36876
rect 17957 36873 17969 36907
rect 18003 36904 18015 36907
rect 18690 36904 18696 36916
rect 18003 36876 18696 36904
rect 18003 36873 18015 36876
rect 17957 36867 18015 36873
rect 18690 36864 18696 36876
rect 18748 36864 18754 36916
rect 18966 36864 18972 36916
rect 19024 36904 19030 36916
rect 19150 36904 19156 36916
rect 19024 36876 19156 36904
rect 19024 36864 19030 36876
rect 19150 36864 19156 36876
rect 19208 36864 19214 36916
rect 19426 36864 19432 36916
rect 19484 36904 19490 36916
rect 19889 36907 19947 36913
rect 19889 36904 19901 36907
rect 19484 36876 19901 36904
rect 19484 36864 19490 36876
rect 19889 36873 19901 36876
rect 19935 36873 19947 36907
rect 19889 36867 19947 36873
rect 18776 36839 18834 36845
rect 18776 36836 18788 36839
rect 15396 36808 18788 36836
rect 18776 36805 18788 36808
rect 18822 36836 18834 36839
rect 19242 36836 19248 36848
rect 18822 36808 19248 36836
rect 18822 36805 18834 36808
rect 18776 36799 18834 36805
rect 19242 36796 19248 36808
rect 19300 36796 19306 36848
rect 14029 36770 14044 36796
rect 15105 36771 15163 36777
rect 14029 36767 14041 36770
rect 15105 36768 15117 36771
rect 13983 36761 14041 36767
rect 14752 36740 15117 36768
rect 11837 36737 11849 36740
rect 11791 36731 11849 36737
rect 3789 36703 3847 36709
rect 3789 36669 3801 36703
rect 3835 36669 3847 36703
rect 3789 36663 3847 36669
rect 1360 36604 3648 36632
rect 1360 36592 1366 36604
rect 1765 36567 1823 36573
rect 1765 36533 1777 36567
rect 1811 36564 1823 36567
rect 2130 36564 2136 36576
rect 1811 36536 2136 36564
rect 1811 36533 1823 36536
rect 1765 36527 1823 36533
rect 2130 36524 2136 36536
rect 2188 36524 2194 36576
rect 3234 36524 3240 36576
rect 3292 36564 3298 36576
rect 3804 36564 3832 36663
rect 5166 36660 5172 36712
rect 5224 36700 5230 36712
rect 5368 36700 5396 36728
rect 14752 36712 14780 36740
rect 15105 36737 15117 36740
rect 15151 36737 15163 36771
rect 15105 36731 15163 36737
rect 15289 36771 15347 36777
rect 15289 36737 15301 36771
rect 15335 36768 15347 36771
rect 15378 36768 15384 36780
rect 15335 36740 15384 36768
rect 15335 36737 15347 36740
rect 15289 36731 15347 36737
rect 15378 36728 15384 36740
rect 15436 36728 15442 36780
rect 15562 36728 15568 36780
rect 15620 36768 15626 36780
rect 15749 36771 15807 36777
rect 15749 36768 15761 36771
rect 15620 36740 15761 36768
rect 15620 36728 15626 36740
rect 15749 36737 15761 36740
rect 15795 36737 15807 36771
rect 15749 36731 15807 36737
rect 18138 36728 18144 36780
rect 18196 36728 18202 36780
rect 18414 36728 18420 36780
rect 18472 36728 18478 36780
rect 20162 36728 20168 36780
rect 20220 36728 20226 36780
rect 7558 36700 7564 36712
rect 5224 36672 7564 36700
rect 5224 36660 5230 36672
rect 7558 36660 7564 36672
rect 7616 36700 7622 36712
rect 7837 36703 7895 36709
rect 7837 36700 7849 36703
rect 7616 36672 7849 36700
rect 7616 36660 7622 36672
rect 7837 36669 7849 36672
rect 7883 36669 7895 36703
rect 7837 36663 7895 36669
rect 8018 36660 8024 36712
rect 8076 36660 8082 36712
rect 8478 36660 8484 36712
rect 8536 36660 8542 36712
rect 8874 36703 8932 36709
rect 8874 36700 8886 36703
rect 8588 36672 8886 36700
rect 4154 36592 4160 36644
rect 4212 36632 4218 36644
rect 7374 36632 7380 36644
rect 4212 36604 7380 36632
rect 4212 36592 4218 36604
rect 7374 36592 7380 36604
rect 7432 36632 7438 36644
rect 8588 36632 8616 36672
rect 8874 36669 8886 36672
rect 8920 36669 8932 36703
rect 9766 36700 9772 36712
rect 8874 36663 8932 36669
rect 9508 36672 9772 36700
rect 7432 36604 8616 36632
rect 7432 36592 7438 36604
rect 3292 36536 3832 36564
rect 4525 36567 4583 36573
rect 3292 36524 3298 36536
rect 4525 36533 4537 36567
rect 4571 36564 4583 36567
rect 7006 36564 7012 36576
rect 4571 36536 7012 36564
rect 4571 36533 4583 36536
rect 4525 36527 4583 36533
rect 7006 36524 7012 36536
rect 7064 36524 7070 36576
rect 9030 36524 9036 36576
rect 9088 36564 9094 36576
rect 9508 36564 9536 36672
rect 9766 36660 9772 36672
rect 9824 36660 9830 36712
rect 11517 36703 11575 36709
rect 11517 36669 11529 36703
rect 11563 36669 11575 36703
rect 11517 36663 11575 36669
rect 9088 36536 9536 36564
rect 9088 36524 9094 36536
rect 9582 36524 9588 36576
rect 9640 36564 9646 36576
rect 10781 36567 10839 36573
rect 10781 36564 10793 36567
rect 9640 36536 10793 36564
rect 9640 36524 9646 36536
rect 10781 36533 10793 36536
rect 10827 36533 10839 36567
rect 10781 36527 10839 36533
rect 11330 36524 11336 36576
rect 11388 36564 11394 36576
rect 11532 36564 11560 36663
rect 13446 36660 13452 36712
rect 13504 36700 13510 36712
rect 13725 36703 13783 36709
rect 13725 36700 13737 36703
rect 13504 36672 13737 36700
rect 13504 36660 13510 36672
rect 13725 36669 13737 36672
rect 13771 36669 13783 36703
rect 13725 36663 13783 36669
rect 14734 36660 14740 36712
rect 14792 36660 14798 36712
rect 16666 36660 16672 36712
rect 16724 36700 16730 36712
rect 18509 36703 18567 36709
rect 18509 36700 18521 36703
rect 16724 36672 18521 36700
rect 16724 36660 16730 36672
rect 18509 36669 18521 36672
rect 18555 36669 18567 36703
rect 18509 36663 18567 36669
rect 17034 36632 17040 36644
rect 12176 36604 13308 36632
rect 11790 36564 11796 36576
rect 11388 36536 11796 36564
rect 11388 36524 11394 36536
rect 11790 36524 11796 36536
rect 11848 36564 11854 36576
rect 12176 36564 12204 36604
rect 11848 36536 12204 36564
rect 12529 36567 12587 36573
rect 11848 36524 11854 36536
rect 12529 36533 12541 36567
rect 12575 36564 12587 36567
rect 12710 36564 12716 36576
rect 12575 36536 12716 36564
rect 12575 36533 12587 36536
rect 12529 36527 12587 36533
rect 12710 36524 12716 36536
rect 12768 36524 12774 36576
rect 12894 36524 12900 36576
rect 12952 36564 12958 36576
rect 13170 36564 13176 36576
rect 12952 36536 13176 36564
rect 12952 36524 12958 36536
rect 13170 36524 13176 36536
rect 13228 36524 13234 36576
rect 13280 36564 13308 36604
rect 14384 36604 17040 36632
rect 14384 36564 14412 36604
rect 17034 36592 17040 36604
rect 17092 36592 17098 36644
rect 13280 36536 14412 36564
rect 14734 36524 14740 36576
rect 14792 36524 14798 36576
rect 15194 36524 15200 36576
rect 15252 36524 15258 36576
rect 15470 36524 15476 36576
rect 15528 36564 15534 36576
rect 15565 36567 15623 36573
rect 15565 36564 15577 36567
rect 15528 36536 15577 36564
rect 15528 36524 15534 36536
rect 15565 36533 15577 36536
rect 15611 36533 15623 36567
rect 15565 36527 15623 36533
rect 18233 36567 18291 36573
rect 18233 36533 18245 36567
rect 18279 36564 18291 36567
rect 19886 36564 19892 36576
rect 18279 36536 19892 36564
rect 18279 36533 18291 36536
rect 18233 36527 18291 36533
rect 19886 36524 19892 36536
rect 19944 36524 19950 36576
rect 20441 36567 20499 36573
rect 20441 36533 20453 36567
rect 20487 36564 20499 36567
rect 21266 36564 21272 36576
rect 20487 36536 21272 36564
rect 20487 36533 20499 36536
rect 20441 36527 20499 36533
rect 21266 36524 21272 36536
rect 21324 36524 21330 36576
rect 1104 36474 20884 36496
rect 1104 36422 3422 36474
rect 3474 36422 3486 36474
rect 3538 36422 3550 36474
rect 3602 36422 3614 36474
rect 3666 36422 3678 36474
rect 3730 36422 8367 36474
rect 8419 36422 8431 36474
rect 8483 36422 8495 36474
rect 8547 36422 8559 36474
rect 8611 36422 8623 36474
rect 8675 36422 13312 36474
rect 13364 36422 13376 36474
rect 13428 36422 13440 36474
rect 13492 36422 13504 36474
rect 13556 36422 13568 36474
rect 13620 36422 18257 36474
rect 18309 36422 18321 36474
rect 18373 36422 18385 36474
rect 18437 36422 18449 36474
rect 18501 36422 18513 36474
rect 18565 36422 20884 36474
rect 1104 36400 20884 36422
rect 382 36320 388 36372
rect 440 36360 446 36372
rect 2590 36360 2596 36372
rect 440 36332 2596 36360
rect 440 36320 446 36332
rect 2590 36320 2596 36332
rect 2648 36320 2654 36372
rect 2866 36320 2872 36372
rect 2924 36360 2930 36372
rect 3421 36363 3479 36369
rect 3421 36360 3433 36363
rect 2924 36332 3433 36360
rect 2924 36320 2930 36332
rect 3421 36329 3433 36332
rect 3467 36329 3479 36363
rect 3421 36323 3479 36329
rect 6914 36320 6920 36372
rect 6972 36360 6978 36372
rect 6972 36332 7236 36360
rect 6972 36320 6978 36332
rect 4154 36292 4160 36304
rect 3804 36264 4160 36292
rect 2222 36184 2228 36236
rect 2280 36184 2286 36236
rect 2501 36227 2559 36233
rect 2501 36193 2513 36227
rect 2547 36224 2559 36227
rect 3804 36224 3832 36264
rect 4154 36252 4160 36264
rect 4212 36252 4218 36304
rect 7208 36301 7236 36332
rect 7466 36320 7472 36372
rect 7524 36360 7530 36372
rect 8389 36363 8447 36369
rect 7524 36332 8340 36360
rect 7524 36320 7530 36332
rect 5537 36295 5595 36301
rect 5537 36261 5549 36295
rect 5583 36261 5595 36295
rect 5537 36255 5595 36261
rect 7193 36295 7251 36301
rect 7193 36261 7205 36295
rect 7239 36261 7251 36295
rect 7193 36255 7251 36261
rect 2547 36196 3832 36224
rect 2547 36193 2559 36196
rect 2501 36187 2559 36193
rect 3878 36184 3884 36236
rect 3936 36224 3942 36236
rect 5552 36224 5580 36255
rect 3936 36196 4094 36224
rect 5552 36196 7512 36224
rect 3936 36184 3942 36196
rect 7484 36168 7512 36196
rect 7558 36184 7564 36236
rect 7616 36233 7622 36236
rect 7616 36227 7644 36233
rect 7632 36193 7644 36227
rect 7616 36187 7644 36193
rect 7745 36227 7803 36233
rect 7745 36193 7757 36227
rect 7791 36224 7803 36227
rect 7926 36224 7932 36236
rect 7791 36196 7932 36224
rect 7791 36193 7803 36196
rect 7745 36187 7803 36193
rect 7616 36184 7622 36187
rect 7926 36184 7932 36196
rect 7984 36184 7990 36236
rect 750 36116 756 36168
rect 808 36156 814 36168
rect 1026 36156 1032 36168
rect 808 36128 1032 36156
rect 808 36116 814 36128
rect 1026 36116 1032 36128
rect 1084 36116 1090 36168
rect 1578 36116 1584 36168
rect 1636 36116 1642 36168
rect 1762 36116 1768 36168
rect 1820 36116 1826 36168
rect 2590 36116 2596 36168
rect 2648 36165 2654 36168
rect 2648 36159 2676 36165
rect 2664 36125 2676 36159
rect 2648 36119 2676 36125
rect 2648 36116 2654 36119
rect 2774 36116 2780 36168
rect 2832 36116 2838 36168
rect 3970 36116 3976 36168
rect 4028 36156 4034 36168
rect 4525 36159 4583 36165
rect 4525 36156 4537 36159
rect 4028 36128 4537 36156
rect 4028 36116 4034 36128
rect 4525 36125 4537 36128
rect 4571 36156 4583 36159
rect 4798 36156 4804 36168
rect 4571 36128 4804 36156
rect 4571 36125 4583 36128
rect 4525 36119 4583 36125
rect 4798 36116 4804 36128
rect 4856 36116 4862 36168
rect 6546 36116 6552 36168
rect 6604 36116 6610 36168
rect 6638 36116 6644 36168
rect 6696 36156 6702 36168
rect 6733 36159 6791 36165
rect 6733 36156 6745 36159
rect 6696 36128 6745 36156
rect 6696 36116 6702 36128
rect 6733 36125 6745 36128
rect 6779 36156 6791 36159
rect 6914 36156 6920 36168
rect 6779 36128 6920 36156
rect 6779 36125 6791 36128
rect 6733 36119 6791 36125
rect 6914 36116 6920 36128
rect 6972 36116 6978 36168
rect 7466 36116 7472 36168
rect 7524 36116 7530 36168
rect 4614 36048 4620 36100
rect 4672 36048 4678 36100
rect 4982 36048 4988 36100
rect 5040 36048 5046 36100
rect 8312 36088 8340 36332
rect 8389 36329 8401 36363
rect 8435 36360 8447 36363
rect 15286 36360 15292 36372
rect 8435 36332 15292 36360
rect 8435 36329 8447 36332
rect 8389 36323 8447 36329
rect 15286 36320 15292 36332
rect 15344 36320 15350 36372
rect 15470 36320 15476 36372
rect 15528 36360 15534 36372
rect 18049 36363 18107 36369
rect 15528 36332 16804 36360
rect 15528 36320 15534 36332
rect 12342 36252 12348 36304
rect 12400 36292 12406 36304
rect 13906 36292 13912 36304
rect 12400 36264 13912 36292
rect 12400 36252 12406 36264
rect 13906 36252 13912 36264
rect 13964 36252 13970 36304
rect 9493 36227 9551 36233
rect 9493 36224 9505 36227
rect 9048 36196 9505 36224
rect 9048 36168 9076 36196
rect 9493 36193 9505 36196
rect 9539 36193 9551 36227
rect 9493 36187 9551 36193
rect 11238 36184 11244 36236
rect 11296 36184 11302 36236
rect 14090 36184 14096 36236
rect 14148 36184 14154 36236
rect 9030 36116 9036 36168
rect 9088 36116 9094 36168
rect 9398 36116 9404 36168
rect 9456 36156 9462 36168
rect 9735 36159 9793 36165
rect 9735 36156 9747 36159
rect 9456 36128 9747 36156
rect 9456 36116 9462 36128
rect 9735 36125 9747 36128
rect 9781 36125 9793 36159
rect 11515 36159 11573 36165
rect 11515 36156 11527 36159
rect 9735 36119 9793 36125
rect 10177 36128 11527 36156
rect 8754 36088 8760 36100
rect 8312 36060 8760 36088
rect 8754 36048 8760 36060
rect 8812 36088 8818 36100
rect 10177 36088 10205 36128
rect 11515 36125 11527 36128
rect 11561 36156 11573 36159
rect 11882 36156 11888 36168
rect 11561 36128 11888 36156
rect 11561 36125 11573 36128
rect 11515 36119 11573 36125
rect 11882 36116 11888 36128
rect 11940 36116 11946 36168
rect 13909 36159 13967 36165
rect 13909 36156 13921 36159
rect 13832 36128 13921 36156
rect 8812 36060 10205 36088
rect 13832 36088 13860 36128
rect 13909 36125 13921 36128
rect 13955 36125 13967 36159
rect 14108 36156 14136 36184
rect 15657 36159 15715 36165
rect 15657 36156 15669 36159
rect 14108 36128 15669 36156
rect 13909 36119 13967 36125
rect 15657 36125 15669 36128
rect 15703 36156 15715 36159
rect 16666 36156 16672 36168
rect 15703 36128 16672 36156
rect 15703 36125 15715 36128
rect 15657 36119 15715 36125
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 16776 36156 16804 36332
rect 18049 36329 18061 36363
rect 18095 36360 18107 36363
rect 18506 36360 18512 36372
rect 18095 36332 18512 36360
rect 18095 36329 18107 36332
rect 18049 36323 18107 36329
rect 18506 36320 18512 36332
rect 18564 36320 18570 36372
rect 18601 36363 18659 36369
rect 18601 36329 18613 36363
rect 18647 36360 18659 36363
rect 20162 36360 20168 36372
rect 18647 36332 20168 36360
rect 18647 36329 18659 36332
rect 18601 36323 18659 36329
rect 20162 36320 20168 36332
rect 20220 36320 20226 36372
rect 17129 36295 17187 36301
rect 17129 36261 17141 36295
rect 17175 36261 17187 36295
rect 17129 36255 17187 36261
rect 17144 36224 17172 36255
rect 18322 36252 18328 36304
rect 18380 36292 18386 36304
rect 18877 36295 18935 36301
rect 18877 36292 18889 36295
rect 18380 36264 18889 36292
rect 18380 36252 18386 36264
rect 18877 36261 18889 36264
rect 18923 36261 18935 36295
rect 18877 36255 18935 36261
rect 18966 36252 18972 36304
rect 19024 36252 19030 36304
rect 20070 36252 20076 36304
rect 20128 36292 20134 36304
rect 20257 36295 20315 36301
rect 20257 36292 20269 36295
rect 20128 36264 20269 36292
rect 20128 36252 20134 36264
rect 20257 36261 20269 36264
rect 20303 36261 20315 36295
rect 20257 36255 20315 36261
rect 18984 36224 19012 36252
rect 19245 36227 19303 36233
rect 19245 36224 19257 36227
rect 17144 36196 18828 36224
rect 18984 36196 19257 36224
rect 17313 36159 17371 36165
rect 17313 36156 17325 36159
rect 16776 36128 17325 36156
rect 17313 36125 17325 36128
rect 17359 36125 17371 36159
rect 17313 36119 17371 36125
rect 17402 36116 17408 36168
rect 17460 36116 17466 36168
rect 17865 36159 17923 36165
rect 17865 36125 17877 36159
rect 17911 36125 17923 36159
rect 18248 36141 18368 36156
rect 17865 36119 17923 36125
rect 18233 36135 18368 36141
rect 14338 36091 14396 36097
rect 14338 36088 14350 36091
rect 13832 36060 14350 36088
rect 8812 36048 8818 36060
rect 13832 36032 13860 36060
rect 14338 36057 14350 36060
rect 14384 36057 14396 36091
rect 14338 36051 14396 36057
rect 15286 36048 15292 36100
rect 15344 36088 15350 36100
rect 15902 36091 15960 36097
rect 15902 36088 15914 36091
rect 15344 36060 15914 36088
rect 15344 36048 15350 36060
rect 15902 36057 15914 36060
rect 15948 36088 15960 36091
rect 16206 36088 16212 36100
rect 15948 36060 16212 36088
rect 15948 36057 15960 36060
rect 15902 36051 15960 36057
rect 16206 36048 16212 36060
rect 16264 36048 16270 36100
rect 17880 36088 17908 36119
rect 18233 36101 18245 36135
rect 18279 36128 18368 36135
rect 18279 36101 18291 36128
rect 18233 36095 18291 36101
rect 17052 36060 17908 36088
rect 18340 36088 18368 36128
rect 18414 36116 18420 36168
rect 18472 36156 18478 36168
rect 18800 36165 18828 36196
rect 19245 36193 19257 36196
rect 19291 36193 19303 36227
rect 19245 36187 19303 36193
rect 18509 36159 18567 36165
rect 18509 36156 18521 36159
rect 18472 36128 18521 36156
rect 18472 36116 18478 36128
rect 18509 36125 18521 36128
rect 18555 36125 18567 36159
rect 18509 36119 18567 36125
rect 18785 36159 18843 36165
rect 18785 36125 18797 36159
rect 18831 36125 18843 36159
rect 18785 36119 18843 36125
rect 18966 36116 18972 36168
rect 19024 36156 19030 36168
rect 19061 36159 19119 36165
rect 19061 36156 19073 36159
rect 19024 36128 19073 36156
rect 19024 36116 19030 36128
rect 19061 36125 19073 36128
rect 19107 36125 19119 36159
rect 19487 36159 19545 36165
rect 19487 36156 19499 36159
rect 19061 36119 19119 36125
rect 19352 36128 19499 36156
rect 19352 36100 19380 36128
rect 19487 36125 19499 36128
rect 19533 36125 19545 36159
rect 19487 36119 19545 36125
rect 19886 36116 19892 36168
rect 19944 36156 19950 36168
rect 20530 36156 20536 36168
rect 19944 36128 20536 36156
rect 19944 36116 19950 36128
rect 20530 36116 20536 36128
rect 20588 36116 20594 36168
rect 18874 36088 18880 36100
rect 18340 36060 18880 36088
rect 2590 35980 2596 36032
rect 2648 36020 2654 36032
rect 2866 36020 2872 36032
rect 2648 35992 2872 36020
rect 2648 35980 2654 35992
rect 2866 35980 2872 35992
rect 2924 36020 2930 36032
rect 3786 36020 3792 36032
rect 2924 35992 3792 36020
rect 2924 35980 2930 35992
rect 3786 35980 3792 35992
rect 3844 35980 3850 36032
rect 4154 35980 4160 36032
rect 4212 36020 4218 36032
rect 4249 36023 4307 36029
rect 4249 36020 4261 36023
rect 4212 35992 4261 36020
rect 4212 35980 4218 35992
rect 4249 35989 4261 35992
rect 4295 35989 4307 36023
rect 4249 35983 4307 35989
rect 4522 35980 4528 36032
rect 4580 36020 4586 36032
rect 4890 36020 4896 36032
rect 4580 35992 4896 36020
rect 4580 35980 4586 35992
rect 4890 35980 4896 35992
rect 4948 36020 4954 36032
rect 5353 36023 5411 36029
rect 5353 36020 5365 36023
rect 4948 35992 5365 36020
rect 4948 35980 4954 35992
rect 5353 35989 5365 35992
rect 5399 35989 5411 36023
rect 5353 35983 5411 35989
rect 6730 35980 6736 36032
rect 6788 36020 6794 36032
rect 9950 36020 9956 36032
rect 6788 35992 9956 36020
rect 6788 35980 6794 35992
rect 9950 35980 9956 35992
rect 10008 35980 10014 36032
rect 10318 35980 10324 36032
rect 10376 36020 10382 36032
rect 10505 36023 10563 36029
rect 10505 36020 10517 36023
rect 10376 35992 10517 36020
rect 10376 35980 10382 35992
rect 10505 35989 10517 35992
rect 10551 35989 10563 36023
rect 10505 35983 10563 35989
rect 11422 35980 11428 36032
rect 11480 36020 11486 36032
rect 11606 36020 11612 36032
rect 11480 35992 11612 36020
rect 11480 35980 11486 35992
rect 11606 35980 11612 35992
rect 11664 35980 11670 36032
rect 11882 35980 11888 36032
rect 11940 36020 11946 36032
rect 12253 36023 12311 36029
rect 12253 36020 12265 36023
rect 11940 35992 12265 36020
rect 11940 35980 11946 35992
rect 12253 35989 12265 35992
rect 12299 35989 12311 36023
rect 12253 35983 12311 35989
rect 13722 35980 13728 36032
rect 13780 35980 13786 36032
rect 13814 35980 13820 36032
rect 13872 35980 13878 36032
rect 15470 35980 15476 36032
rect 15528 35980 15534 36032
rect 17052 36029 17080 36060
rect 18874 36048 18880 36060
rect 18932 36048 18938 36100
rect 19334 36048 19340 36100
rect 19392 36048 19398 36100
rect 17037 36023 17095 36029
rect 17037 35989 17049 36023
rect 17083 35989 17095 36023
rect 17037 35983 17095 35989
rect 17218 35980 17224 36032
rect 17276 36020 17282 36032
rect 17497 36023 17555 36029
rect 17497 36020 17509 36023
rect 17276 35992 17509 36020
rect 17276 35980 17282 35992
rect 17497 35989 17509 35992
rect 17543 35989 17555 36023
rect 17497 35983 17555 35989
rect 17678 35980 17684 36032
rect 17736 35980 17742 36032
rect 18325 36023 18383 36029
rect 18325 35989 18337 36023
rect 18371 36020 18383 36023
rect 19518 36020 19524 36032
rect 18371 35992 19524 36020
rect 18371 35989 18383 35992
rect 18325 35983 18383 35989
rect 19518 35980 19524 35992
rect 19576 35980 19582 36032
rect 1104 35930 21043 35952
rect 1104 35878 5894 35930
rect 5946 35878 5958 35930
rect 6010 35878 6022 35930
rect 6074 35878 6086 35930
rect 6138 35878 6150 35930
rect 6202 35878 10839 35930
rect 10891 35878 10903 35930
rect 10955 35878 10967 35930
rect 11019 35878 11031 35930
rect 11083 35878 11095 35930
rect 11147 35878 15784 35930
rect 15836 35878 15848 35930
rect 15900 35878 15912 35930
rect 15964 35878 15976 35930
rect 16028 35878 16040 35930
rect 16092 35878 20729 35930
rect 20781 35878 20793 35930
rect 20845 35878 20857 35930
rect 20909 35878 20921 35930
rect 20973 35878 20985 35930
rect 21037 35878 21043 35930
rect 1104 35856 21043 35878
rect 2501 35819 2559 35825
rect 2501 35785 2513 35819
rect 2547 35816 2559 35819
rect 2774 35816 2780 35828
rect 2547 35788 2780 35816
rect 2547 35785 2559 35788
rect 2501 35779 2559 35785
rect 2774 35776 2780 35788
rect 2832 35776 2838 35828
rect 3878 35776 3884 35828
rect 3936 35776 3942 35828
rect 4614 35776 4620 35828
rect 4672 35816 4678 35828
rect 5353 35819 5411 35825
rect 5353 35816 5365 35819
rect 4672 35788 5365 35816
rect 4672 35776 4678 35788
rect 5353 35785 5365 35788
rect 5399 35785 5411 35819
rect 10134 35816 10140 35828
rect 5353 35779 5411 35785
rect 9692 35788 10140 35816
rect 1394 35708 1400 35760
rect 1452 35748 1458 35760
rect 1854 35748 1860 35760
rect 1452 35720 1860 35748
rect 1452 35708 1458 35720
rect 1854 35708 1860 35720
rect 1912 35708 1918 35760
rect 5626 35748 5632 35760
rect 2884 35720 5632 35748
rect 1763 35683 1821 35689
rect 1763 35649 1775 35683
rect 1809 35680 1821 35683
rect 2314 35680 2320 35692
rect 1809 35652 2320 35680
rect 1809 35649 1821 35652
rect 1763 35643 1821 35649
rect 2314 35640 2320 35652
rect 2372 35640 2378 35692
rect 2590 35640 2596 35692
rect 2648 35680 2654 35692
rect 2884 35689 2912 35720
rect 2869 35683 2927 35689
rect 2869 35680 2881 35683
rect 2648 35652 2881 35680
rect 2648 35640 2654 35652
rect 2869 35649 2881 35652
rect 2915 35649 2927 35683
rect 3142 35680 3148 35692
rect 3103 35652 3148 35680
rect 2869 35643 2927 35649
rect 3142 35640 3148 35652
rect 3200 35640 3206 35692
rect 4172 35624 4200 35720
rect 5626 35708 5632 35720
rect 5684 35708 5690 35760
rect 9692 35757 9720 35788
rect 10134 35776 10140 35788
rect 10192 35776 10198 35828
rect 10226 35776 10232 35828
rect 10284 35816 10290 35828
rect 10689 35819 10747 35825
rect 10689 35816 10701 35819
rect 10284 35788 10701 35816
rect 10284 35776 10290 35788
rect 10689 35785 10701 35788
rect 10735 35816 10747 35819
rect 10778 35816 10784 35828
rect 10735 35788 10784 35816
rect 10735 35785 10747 35788
rect 10689 35779 10747 35785
rect 10778 35776 10784 35788
rect 10836 35776 10842 35828
rect 13357 35819 13415 35825
rect 13357 35816 13369 35819
rect 11348 35788 13369 35816
rect 9401 35751 9459 35757
rect 9401 35717 9413 35751
rect 9447 35717 9459 35751
rect 9401 35711 9459 35717
rect 9677 35751 9735 35757
rect 9677 35717 9689 35751
rect 9723 35717 9735 35751
rect 9677 35711 9735 35717
rect 4614 35680 4620 35692
rect 4575 35652 4620 35680
rect 4614 35640 4620 35652
rect 4672 35640 4678 35692
rect 9416 35680 9444 35711
rect 9766 35708 9772 35760
rect 9824 35708 9830 35760
rect 9858 35708 9864 35760
rect 9916 35748 9922 35760
rect 9916 35720 10272 35748
rect 9916 35708 9922 35720
rect 9876 35680 9904 35708
rect 9416 35652 9904 35680
rect 10134 35640 10140 35692
rect 10192 35640 10198 35692
rect 10244 35680 10272 35720
rect 10502 35708 10508 35760
rect 10560 35708 10566 35760
rect 10965 35683 11023 35689
rect 10965 35680 10977 35683
rect 10244 35652 10977 35680
rect 10965 35649 10977 35652
rect 11011 35649 11023 35683
rect 10965 35643 11023 35649
rect 1394 35572 1400 35624
rect 1452 35612 1458 35624
rect 1489 35615 1547 35621
rect 1489 35612 1501 35615
rect 1452 35584 1501 35612
rect 1452 35572 1458 35584
rect 1489 35581 1501 35584
rect 1535 35581 1547 35615
rect 1489 35575 1547 35581
rect 4154 35572 4160 35624
rect 4212 35612 4218 35624
rect 4341 35615 4399 35621
rect 4341 35612 4353 35615
rect 4212 35584 4353 35612
rect 4212 35572 4218 35584
rect 4341 35581 4353 35584
rect 4387 35581 4399 35615
rect 4341 35575 4399 35581
rect 5718 35572 5724 35624
rect 5776 35612 5782 35624
rect 6362 35612 6368 35624
rect 5776 35584 6368 35612
rect 5776 35572 5782 35584
rect 6362 35572 6368 35584
rect 6420 35572 6426 35624
rect 9582 35572 9588 35624
rect 9640 35572 9646 35624
rect 10594 35572 10600 35624
rect 10652 35612 10658 35624
rect 11348 35612 11376 35788
rect 13357 35785 13369 35788
rect 13403 35785 13415 35819
rect 13357 35779 13415 35785
rect 13722 35776 13728 35828
rect 13780 35776 13786 35828
rect 15378 35776 15384 35828
rect 15436 35776 15442 35828
rect 15470 35776 15476 35828
rect 15528 35776 15534 35828
rect 16117 35819 16175 35825
rect 16117 35785 16129 35819
rect 16163 35816 16175 35819
rect 17402 35816 17408 35828
rect 16163 35788 17408 35816
rect 16163 35785 16175 35788
rect 16117 35779 16175 35785
rect 17402 35776 17408 35788
rect 17460 35776 17466 35828
rect 17678 35776 17684 35828
rect 17736 35776 17742 35828
rect 18322 35776 18328 35828
rect 18380 35776 18386 35828
rect 18417 35819 18475 35825
rect 18417 35785 18429 35819
rect 18463 35785 18475 35819
rect 18417 35779 18475 35785
rect 12710 35640 12716 35692
rect 12768 35640 12774 35692
rect 13740 35680 13768 35776
rect 15194 35708 15200 35760
rect 15252 35748 15258 35760
rect 15289 35751 15347 35757
rect 15289 35748 15301 35751
rect 15252 35720 15301 35748
rect 15252 35708 15258 35720
rect 15289 35717 15301 35720
rect 15335 35717 15347 35751
rect 15289 35711 15347 35717
rect 14461 35683 14519 35689
rect 14461 35680 14473 35683
rect 13740 35652 14473 35680
rect 14461 35649 14473 35652
rect 14507 35649 14519 35683
rect 14461 35643 14519 35649
rect 14553 35683 14611 35689
rect 14553 35649 14565 35683
rect 14599 35680 14611 35683
rect 14921 35683 14979 35689
rect 14921 35680 14933 35683
rect 14599 35652 14933 35680
rect 14599 35649 14611 35652
rect 14553 35643 14611 35649
rect 14921 35649 14933 35652
rect 14967 35649 14979 35683
rect 15488 35680 15516 35776
rect 16206 35708 16212 35760
rect 16264 35708 16270 35760
rect 15565 35683 15623 35689
rect 15565 35680 15577 35683
rect 15488 35652 15577 35680
rect 14921 35643 14979 35649
rect 15565 35649 15577 35652
rect 15611 35649 15623 35683
rect 16224 35680 16252 35708
rect 16301 35683 16359 35689
rect 16301 35680 16313 35683
rect 16224 35652 16313 35680
rect 15565 35643 15623 35649
rect 16301 35649 16313 35652
rect 16347 35649 16359 35683
rect 16301 35643 16359 35649
rect 17034 35640 17040 35692
rect 17092 35680 17098 35692
rect 17405 35683 17463 35689
rect 17405 35680 17417 35683
rect 17092 35652 17417 35680
rect 17092 35640 17098 35652
rect 17405 35649 17417 35652
rect 17451 35649 17463 35683
rect 17405 35643 17463 35649
rect 17589 35683 17647 35689
rect 17589 35649 17601 35683
rect 17635 35680 17647 35683
rect 17696 35680 17724 35776
rect 18340 35748 18368 35776
rect 17880 35720 18368 35748
rect 18432 35748 18460 35779
rect 18506 35776 18512 35828
rect 18564 35816 18570 35828
rect 19518 35816 19524 35828
rect 18564 35788 19524 35816
rect 18564 35776 18570 35788
rect 19518 35776 19524 35788
rect 19576 35776 19582 35828
rect 19610 35776 19616 35828
rect 19668 35776 19674 35828
rect 19628 35748 19656 35776
rect 18432 35720 18920 35748
rect 17880 35689 17908 35720
rect 17635 35652 17724 35680
rect 17865 35683 17923 35689
rect 17635 35649 17647 35652
rect 17589 35643 17647 35649
rect 17865 35649 17877 35683
rect 17911 35649 17923 35683
rect 17865 35643 17923 35649
rect 17954 35640 17960 35692
rect 18012 35680 18018 35692
rect 18892 35689 18920 35720
rect 19168 35720 19564 35748
rect 19628 35720 19932 35748
rect 19168 35692 19196 35720
rect 18141 35683 18199 35689
rect 18141 35680 18153 35683
rect 18012 35652 18153 35680
rect 18012 35640 18018 35652
rect 18141 35649 18153 35652
rect 18187 35649 18199 35683
rect 18141 35643 18199 35649
rect 18601 35683 18659 35689
rect 18601 35649 18613 35683
rect 18647 35649 18659 35683
rect 18601 35643 18659 35649
rect 18877 35683 18935 35689
rect 18877 35649 18889 35683
rect 18923 35649 18935 35683
rect 18877 35643 18935 35649
rect 10652 35584 11376 35612
rect 11517 35615 11575 35621
rect 10652 35572 10658 35584
rect 11517 35581 11529 35615
rect 11563 35612 11575 35615
rect 11606 35612 11612 35624
rect 11563 35584 11612 35612
rect 11563 35581 11575 35584
rect 11517 35575 11575 35581
rect 11606 35572 11612 35584
rect 11664 35572 11670 35624
rect 11701 35615 11759 35621
rect 11701 35581 11713 35615
rect 11747 35612 11759 35615
rect 11790 35612 11796 35624
rect 11747 35584 11796 35612
rect 11747 35581 11759 35584
rect 11701 35575 11759 35581
rect 11790 35572 11796 35584
rect 11848 35572 11854 35624
rect 12066 35572 12072 35624
rect 12124 35612 12130 35624
rect 12161 35615 12219 35621
rect 12161 35612 12173 35615
rect 12124 35584 12173 35612
rect 12124 35572 12130 35584
rect 12161 35581 12173 35584
rect 12207 35581 12219 35615
rect 12437 35615 12495 35621
rect 12437 35612 12449 35615
rect 12161 35575 12219 35581
rect 12268 35584 12449 35612
rect 10778 35504 10784 35556
rect 10836 35504 10842 35556
rect 10870 35504 10876 35556
rect 10928 35544 10934 35556
rect 11149 35547 11207 35553
rect 11149 35544 11161 35547
rect 10928 35516 11161 35544
rect 10928 35504 10934 35516
rect 11149 35513 11161 35516
rect 11195 35513 11207 35547
rect 11149 35507 11207 35513
rect 3326 35436 3332 35488
rect 3384 35476 3390 35488
rect 6730 35476 6736 35488
rect 3384 35448 6736 35476
rect 3384 35436 3390 35448
rect 6730 35436 6736 35448
rect 6788 35436 6794 35488
rect 10796 35476 10824 35504
rect 12268 35476 12296 35584
rect 12437 35581 12449 35584
rect 12483 35581 12495 35615
rect 12437 35575 12495 35581
rect 12575 35615 12633 35621
rect 12575 35581 12587 35615
rect 12621 35612 12633 35615
rect 14642 35612 14648 35624
rect 12621 35584 14648 35612
rect 12621 35581 12633 35584
rect 12575 35575 12633 35581
rect 14642 35572 14648 35584
rect 14700 35572 14706 35624
rect 14734 35572 14740 35624
rect 14792 35572 14798 35624
rect 15194 35612 15200 35624
rect 14844 35584 15200 35612
rect 13538 35504 13544 35556
rect 13596 35544 13602 35556
rect 14844 35544 14872 35584
rect 15194 35572 15200 35584
rect 15252 35572 15258 35624
rect 17129 35615 17187 35621
rect 17129 35581 17141 35615
rect 17175 35612 17187 35615
rect 17218 35612 17224 35624
rect 17175 35584 17224 35612
rect 17175 35581 17187 35584
rect 17129 35575 17187 35581
rect 17218 35572 17224 35584
rect 17276 35572 17282 35624
rect 17313 35615 17371 35621
rect 17313 35581 17325 35615
rect 17359 35612 17371 35615
rect 17497 35615 17555 35621
rect 17497 35612 17509 35615
rect 17359 35584 17509 35612
rect 17359 35581 17371 35584
rect 17313 35575 17371 35581
rect 17497 35581 17509 35584
rect 17543 35581 17555 35615
rect 18616 35612 18644 35643
rect 19150 35640 19156 35692
rect 19208 35640 19214 35692
rect 19337 35683 19395 35689
rect 19337 35649 19349 35683
rect 19383 35680 19395 35683
rect 19426 35680 19432 35692
rect 19383 35652 19432 35680
rect 19383 35649 19395 35652
rect 19337 35643 19395 35649
rect 19426 35640 19432 35652
rect 19484 35640 19490 35692
rect 17497 35575 17555 35581
rect 17972 35584 18644 35612
rect 17972 35553 18000 35584
rect 18690 35572 18696 35624
rect 18748 35572 18754 35624
rect 19536 35612 19564 35720
rect 19610 35640 19616 35692
rect 19668 35640 19674 35692
rect 19904 35689 19932 35720
rect 19978 35708 19984 35760
rect 20036 35748 20042 35760
rect 20257 35751 20315 35757
rect 20257 35748 20269 35751
rect 20036 35720 20269 35748
rect 20036 35708 20042 35720
rect 20257 35717 20269 35720
rect 20303 35717 20315 35751
rect 20257 35711 20315 35717
rect 19889 35683 19947 35689
rect 19889 35649 19901 35683
rect 19935 35649 19947 35683
rect 19889 35643 19947 35649
rect 20070 35640 20076 35692
rect 20128 35640 20134 35692
rect 20530 35640 20536 35692
rect 20588 35640 20594 35692
rect 20622 35612 20628 35624
rect 19536 35584 20628 35612
rect 20622 35572 20628 35584
rect 20680 35572 20686 35624
rect 13596 35516 14872 35544
rect 15105 35547 15163 35553
rect 13596 35504 13602 35516
rect 15105 35513 15117 35547
rect 15151 35544 15163 35547
rect 17957 35547 18015 35553
rect 15151 35516 17172 35544
rect 15151 35513 15163 35516
rect 15105 35507 15163 35513
rect 17144 35488 17172 35516
rect 17957 35513 17969 35547
rect 18003 35513 18015 35547
rect 17957 35507 18015 35513
rect 10796 35448 12296 35476
rect 12802 35436 12808 35488
rect 12860 35476 12866 35488
rect 13170 35476 13176 35488
rect 12860 35448 13176 35476
rect 12860 35436 12866 35448
rect 13170 35436 13176 35448
rect 13228 35436 13234 35488
rect 14366 35436 14372 35488
rect 14424 35476 14430 35488
rect 16574 35476 16580 35488
rect 14424 35448 16580 35476
rect 14424 35436 14430 35448
rect 16574 35436 16580 35448
rect 16632 35436 16638 35488
rect 17126 35436 17132 35488
rect 17184 35436 17190 35488
rect 17218 35436 17224 35488
rect 17276 35436 17282 35488
rect 17681 35479 17739 35485
rect 17681 35445 17693 35479
rect 17727 35476 17739 35479
rect 18138 35476 18144 35488
rect 17727 35448 18144 35476
rect 17727 35445 17739 35448
rect 17681 35439 17739 35445
rect 18138 35436 18144 35448
rect 18196 35436 18202 35488
rect 18708 35485 18736 35572
rect 19242 35504 19248 35556
rect 19300 35544 19306 35556
rect 19886 35544 19892 35556
rect 19300 35516 19892 35544
rect 19300 35504 19306 35516
rect 19886 35504 19892 35516
rect 19944 35504 19950 35556
rect 20165 35547 20223 35553
rect 20165 35513 20177 35547
rect 20211 35544 20223 35547
rect 20211 35516 21404 35544
rect 20211 35513 20223 35516
rect 20165 35507 20223 35513
rect 21376 35488 21404 35516
rect 18693 35479 18751 35485
rect 18693 35445 18705 35479
rect 18739 35445 18751 35479
rect 18693 35439 18751 35445
rect 19150 35436 19156 35488
rect 19208 35436 19214 35488
rect 19429 35479 19487 35485
rect 19429 35445 19441 35479
rect 19475 35476 19487 35479
rect 19702 35476 19708 35488
rect 19475 35448 19708 35476
rect 19475 35445 19487 35448
rect 19429 35439 19487 35445
rect 19702 35436 19708 35448
rect 19760 35436 19766 35488
rect 19978 35436 19984 35488
rect 20036 35476 20042 35488
rect 20349 35479 20407 35485
rect 20349 35476 20361 35479
rect 20036 35448 20361 35476
rect 20036 35436 20042 35448
rect 20349 35445 20361 35448
rect 20395 35445 20407 35479
rect 20349 35439 20407 35445
rect 21358 35436 21364 35488
rect 21416 35436 21422 35488
rect 1104 35386 20884 35408
rect 1104 35334 3422 35386
rect 3474 35334 3486 35386
rect 3538 35334 3550 35386
rect 3602 35334 3614 35386
rect 3666 35334 3678 35386
rect 3730 35334 8367 35386
rect 8419 35334 8431 35386
rect 8483 35334 8495 35386
rect 8547 35334 8559 35386
rect 8611 35334 8623 35386
rect 8675 35334 13312 35386
rect 13364 35334 13376 35386
rect 13428 35334 13440 35386
rect 13492 35334 13504 35386
rect 13556 35334 13568 35386
rect 13620 35334 18257 35386
rect 18309 35334 18321 35386
rect 18373 35334 18385 35386
rect 18437 35334 18449 35386
rect 18501 35334 18513 35386
rect 18565 35334 20884 35386
rect 1104 35312 20884 35334
rect 2222 35232 2228 35284
rect 2280 35272 2286 35284
rect 2409 35275 2467 35281
rect 2409 35272 2421 35275
rect 2280 35244 2421 35272
rect 2280 35232 2286 35244
rect 2409 35241 2421 35244
rect 2455 35241 2467 35275
rect 2409 35235 2467 35241
rect 4801 35275 4859 35281
rect 4801 35241 4813 35275
rect 4847 35272 4859 35275
rect 5074 35272 5080 35284
rect 4847 35244 5080 35272
rect 4847 35241 4859 35244
rect 4801 35235 4859 35241
rect 5074 35232 5080 35244
rect 5132 35232 5138 35284
rect 6454 35272 6460 35284
rect 5166 35244 6460 35272
rect 2498 35164 2504 35216
rect 2556 35204 2562 35216
rect 5166 35204 5194 35244
rect 6454 35232 6460 35244
rect 6512 35232 6518 35284
rect 7742 35232 7748 35284
rect 7800 35272 7806 35284
rect 10318 35272 10324 35284
rect 7800 35244 10324 35272
rect 7800 35232 7806 35244
rect 10318 35232 10324 35244
rect 10376 35232 10382 35284
rect 10594 35232 10600 35284
rect 10652 35272 10658 35284
rect 11422 35272 11428 35284
rect 10652 35244 11428 35272
rect 10652 35232 10658 35244
rect 11422 35232 11428 35244
rect 11480 35232 11486 35284
rect 11882 35232 11888 35284
rect 11940 35272 11946 35284
rect 11940 35244 12204 35272
rect 11940 35232 11946 35244
rect 2556 35176 5194 35204
rect 2556 35164 2562 35176
rect 8754 35164 8760 35216
rect 8812 35204 8818 35216
rect 9306 35204 9312 35216
rect 8812 35176 9312 35204
rect 8812 35164 8818 35176
rect 9306 35164 9312 35176
rect 9364 35164 9370 35216
rect 9490 35164 9496 35216
rect 9548 35164 9554 35216
rect 12066 35204 12072 35216
rect 10428 35176 12072 35204
rect 1118 35096 1124 35148
rect 1176 35136 1182 35148
rect 1394 35136 1400 35148
rect 1176 35108 1400 35136
rect 1176 35096 1182 35108
rect 1394 35096 1400 35108
rect 1452 35096 1458 35148
rect 3053 35139 3111 35145
rect 3053 35136 3065 35139
rect 2056 35108 3065 35136
rect 1670 35028 1676 35080
rect 1728 35068 1734 35080
rect 2056 35068 2084 35108
rect 3053 35105 3065 35108
rect 3099 35136 3111 35139
rect 3142 35136 3148 35148
rect 3099 35108 3148 35136
rect 3099 35105 3111 35108
rect 3053 35099 3111 35105
rect 3142 35096 3148 35108
rect 3200 35136 3206 35148
rect 9508 35136 9536 35164
rect 3200 35108 4752 35136
rect 3200 35096 3206 35108
rect 1728 35040 2084 35068
rect 1728 35028 1734 35040
rect 2774 35028 2780 35080
rect 2832 35028 2838 35080
rect 3786 35028 3792 35080
rect 3844 35028 3850 35080
rect 4724 35012 4752 35108
rect 8266 35108 9536 35136
rect 4985 35071 5043 35077
rect 4985 35037 4997 35071
rect 5031 35037 5043 35071
rect 4985 35031 5043 35037
rect 5077 35071 5135 35077
rect 5077 35037 5089 35071
rect 5123 35037 5135 35071
rect 5077 35031 5135 35037
rect 4062 34960 4068 35012
rect 4120 34960 4126 35012
rect 4706 34960 4712 35012
rect 4764 34960 4770 35012
rect 2314 34892 2320 34944
rect 2372 34932 2378 34944
rect 4614 34932 4620 34944
rect 2372 34904 4620 34932
rect 2372 34892 2378 34904
rect 4614 34892 4620 34904
rect 4672 34892 4678 34944
rect 5000 34932 5028 35031
rect 5092 35000 5120 35031
rect 5258 35028 5264 35080
rect 5316 35068 5322 35080
rect 5351 35071 5409 35077
rect 5351 35068 5363 35071
rect 5316 35040 5363 35068
rect 5316 35028 5322 35040
rect 5351 35037 5363 35040
rect 5397 35037 5409 35071
rect 5351 35031 5409 35037
rect 6457 35071 6515 35077
rect 6457 35037 6469 35071
rect 6503 35037 6515 35071
rect 6730 35068 6736 35080
rect 6691 35040 6736 35068
rect 6457 35031 6515 35037
rect 6472 35000 6500 35031
rect 6730 35028 6736 35040
rect 6788 35068 6794 35080
rect 7926 35068 7932 35080
rect 6788 35040 7932 35068
rect 6788 35028 6794 35040
rect 7926 35028 7932 35040
rect 7984 35068 7990 35080
rect 8266 35068 8294 35108
rect 7984 35040 8294 35068
rect 8573 35071 8631 35077
rect 7984 35028 7990 35040
rect 8573 35037 8585 35071
rect 8619 35068 8631 35071
rect 8754 35068 8760 35080
rect 8619 35040 8760 35068
rect 8619 35037 8631 35040
rect 8573 35031 8631 35037
rect 8754 35028 8760 35040
rect 8812 35028 8818 35080
rect 9030 35028 9036 35080
rect 9088 35068 9094 35080
rect 9493 35071 9551 35077
rect 9493 35068 9505 35071
rect 9088 35040 9505 35068
rect 9088 35028 9094 35040
rect 9493 35037 9505 35040
rect 9539 35037 9551 35071
rect 10428 35068 10456 35176
rect 12066 35164 12072 35176
rect 12124 35164 12130 35216
rect 12176 35213 12204 35244
rect 12250 35232 12256 35284
rect 12308 35272 12314 35284
rect 13357 35275 13415 35281
rect 12308 35244 13124 35272
rect 12308 35232 12314 35244
rect 12161 35207 12219 35213
rect 12161 35173 12173 35207
rect 12207 35173 12219 35207
rect 12161 35167 12219 35173
rect 11238 35096 11244 35148
rect 11296 35136 11302 35148
rect 11422 35136 11428 35148
rect 11296 35108 11428 35136
rect 11296 35096 11302 35108
rect 11422 35096 11428 35108
rect 11480 35096 11486 35148
rect 11701 35139 11759 35145
rect 11701 35105 11713 35139
rect 11747 35136 11759 35139
rect 11790 35136 11796 35148
rect 11747 35108 11796 35136
rect 11747 35105 11759 35108
rect 11701 35099 11759 35105
rect 11790 35096 11796 35108
rect 11848 35096 11854 35148
rect 13096 35136 13124 35244
rect 13357 35241 13369 35275
rect 13403 35272 13415 35275
rect 13814 35272 13820 35284
rect 13403 35244 13820 35272
rect 13403 35241 13415 35244
rect 13357 35235 13415 35241
rect 13814 35232 13820 35244
rect 13872 35232 13878 35284
rect 15028 35244 16804 35272
rect 13633 35139 13691 35145
rect 13633 35136 13645 35139
rect 13096 35108 13645 35136
rect 13633 35105 13645 35108
rect 13679 35105 13691 35139
rect 13633 35099 13691 35105
rect 9493 35031 9551 35037
rect 9646 35041 10456 35068
rect 9646 35040 9763 35041
rect 6914 35000 6920 35012
rect 5092 34972 6920 35000
rect 6914 34960 6920 34972
rect 6972 34960 6978 35012
rect 7006 34960 7012 35012
rect 7064 35000 7070 35012
rect 9646 35000 9674 35040
rect 9751 35007 9763 35040
rect 9797 35040 10456 35041
rect 11517 35071 11575 35077
rect 9797 35007 9809 35040
rect 11517 35037 11529 35071
rect 11563 35068 11575 35071
rect 11606 35068 11612 35080
rect 11563 35040 11612 35068
rect 11563 35037 11575 35040
rect 11517 35031 11575 35037
rect 11606 35028 11612 35040
rect 11664 35028 11670 35080
rect 12434 35028 12440 35080
rect 12492 35028 12498 35080
rect 12526 35028 12532 35080
rect 12584 35077 12590 35080
rect 12584 35071 12633 35077
rect 12584 35037 12587 35071
rect 12621 35037 12633 35071
rect 12584 35031 12633 35037
rect 12584 35030 12618 35031
rect 12584 35028 12590 35030
rect 12710 35028 12716 35080
rect 12768 35028 12774 35080
rect 13998 35028 14004 35080
rect 14056 35068 14062 35080
rect 14366 35068 14372 35080
rect 14056 35040 14372 35068
rect 14056 35028 14062 35040
rect 14366 35028 14372 35040
rect 14424 35028 14430 35080
rect 14550 35028 14556 35080
rect 14608 35068 14614 35080
rect 14643 35071 14701 35077
rect 14643 35068 14655 35071
rect 14608 35040 14655 35068
rect 14608 35028 14614 35040
rect 14643 35037 14655 35040
rect 14689 35068 14701 35071
rect 15028 35068 15056 35244
rect 15838 35164 15844 35216
rect 15896 35164 15902 35216
rect 16776 35204 16804 35244
rect 17034 35232 17040 35284
rect 17092 35272 17098 35284
rect 17129 35275 17187 35281
rect 17129 35272 17141 35275
rect 17092 35244 17141 35272
rect 17092 35232 17098 35244
rect 17129 35241 17141 35244
rect 17175 35241 17187 35275
rect 17129 35235 17187 35241
rect 17236 35244 18184 35272
rect 17236 35204 17264 35244
rect 16776 35176 17264 35204
rect 18156 35204 18184 35244
rect 18874 35232 18880 35284
rect 18932 35232 18938 35284
rect 19426 35272 19432 35284
rect 19306 35244 19432 35272
rect 19306 35204 19334 35244
rect 19426 35232 19432 35244
rect 19484 35232 19490 35284
rect 20257 35275 20315 35281
rect 20257 35241 20269 35275
rect 20303 35272 20315 35275
rect 20346 35272 20352 35284
rect 20303 35244 20352 35272
rect 20303 35241 20315 35244
rect 20257 35235 20315 35241
rect 20346 35232 20352 35244
rect 20404 35232 20410 35284
rect 18156 35176 19334 35204
rect 18708 35108 19334 35136
rect 18708 35080 18736 35108
rect 14689 35040 15056 35068
rect 16025 35071 16083 35077
rect 14689 35037 14701 35040
rect 14643 35031 14701 35037
rect 16025 35037 16037 35071
rect 16071 35037 16083 35071
rect 16025 35031 16083 35037
rect 16117 35071 16175 35077
rect 16117 35037 16129 35071
rect 16163 35037 16175 35071
rect 16359 35071 16417 35077
rect 16359 35068 16371 35071
rect 16117 35031 16175 35037
rect 16224 35040 16371 35068
rect 9751 35001 9809 35007
rect 7064 34972 9674 35000
rect 7064 34960 7070 34972
rect 10318 34960 10324 35012
rect 10376 35000 10382 35012
rect 10376 34972 11744 35000
rect 10376 34960 10382 34972
rect 5902 34932 5908 34944
rect 5000 34904 5908 34932
rect 5902 34892 5908 34904
rect 5960 34892 5966 34944
rect 6089 34935 6147 34941
rect 6089 34901 6101 34935
rect 6135 34932 6147 34935
rect 6822 34932 6828 34944
rect 6135 34904 6828 34932
rect 6135 34901 6147 34904
rect 6089 34895 6147 34901
rect 6822 34892 6828 34904
rect 6880 34892 6886 34944
rect 7469 34935 7527 34941
rect 7469 34901 7481 34935
rect 7515 34932 7527 34935
rect 7558 34932 7564 34944
rect 7515 34904 7564 34932
rect 7515 34901 7527 34904
rect 7469 34895 7527 34901
rect 7558 34892 7564 34904
rect 7616 34892 7622 34944
rect 8389 34935 8447 34941
rect 8389 34901 8401 34935
rect 8435 34932 8447 34935
rect 9766 34932 9772 34944
rect 8435 34904 9772 34932
rect 8435 34901 8447 34904
rect 8389 34895 8447 34901
rect 9766 34892 9772 34904
rect 9824 34892 9830 34944
rect 9950 34892 9956 34944
rect 10008 34932 10014 34944
rect 10505 34935 10563 34941
rect 10505 34932 10517 34935
rect 10008 34904 10517 34932
rect 10008 34892 10014 34904
rect 10505 34901 10517 34904
rect 10551 34901 10563 34935
rect 10505 34895 10563 34901
rect 10870 34892 10876 34944
rect 10928 34932 10934 34944
rect 11330 34932 11336 34944
rect 10928 34904 11336 34932
rect 10928 34892 10934 34904
rect 11330 34892 11336 34904
rect 11388 34892 11394 34944
rect 11716 34932 11744 34972
rect 13814 34960 13820 35012
rect 13872 35000 13878 35012
rect 14182 35000 14188 35012
rect 13872 34972 14188 35000
rect 13872 34960 13878 34972
rect 14182 34960 14188 34972
rect 14240 35000 14246 35012
rect 16040 35000 16068 35031
rect 14240 34972 16068 35000
rect 14240 34960 14246 34972
rect 14366 34932 14372 34944
rect 11716 34904 14372 34932
rect 14366 34892 14372 34904
rect 14424 34892 14430 34944
rect 15286 34892 15292 34944
rect 15344 34932 15350 34944
rect 15381 34935 15439 34941
rect 15381 34932 15393 34935
rect 15344 34904 15393 34932
rect 15344 34892 15350 34904
rect 15381 34901 15393 34904
rect 15427 34901 15439 34935
rect 16132 34932 16160 35031
rect 16224 35012 16252 35040
rect 16359 35037 16371 35040
rect 16405 35037 16417 35071
rect 16359 35031 16417 35037
rect 16482 35028 16488 35080
rect 16540 35068 16546 35080
rect 17402 35068 17408 35080
rect 16540 35040 17408 35068
rect 16540 35028 16546 35040
rect 17402 35028 17408 35040
rect 17460 35068 17466 35080
rect 17497 35071 17555 35077
rect 17497 35068 17509 35071
rect 17460 35040 17509 35068
rect 17460 35028 17466 35040
rect 17497 35037 17509 35040
rect 17543 35037 17555 35071
rect 17497 35031 17555 35037
rect 17771 35071 17829 35077
rect 17771 35037 17783 35071
rect 17817 35068 17829 35071
rect 17817 35040 18092 35068
rect 17817 35037 17829 35040
rect 17771 35031 17829 35037
rect 18064 35012 18092 35040
rect 18690 35028 18696 35080
rect 18748 35028 18754 35080
rect 19061 35071 19119 35077
rect 19061 35037 19073 35071
rect 19107 35068 19119 35071
rect 19150 35068 19156 35080
rect 19107 35040 19156 35068
rect 19107 35037 19119 35040
rect 19061 35031 19119 35037
rect 19150 35028 19156 35040
rect 19208 35028 19214 35080
rect 19306 35068 19334 35108
rect 19426 35096 19432 35148
rect 19484 35136 19490 35148
rect 20438 35136 20444 35148
rect 19484 35108 20444 35136
rect 19484 35096 19490 35108
rect 20438 35096 20444 35108
rect 20496 35096 20502 35148
rect 19981 35071 20039 35077
rect 19981 35068 19993 35071
rect 19306 35040 19993 35068
rect 19981 35037 19993 35040
rect 20027 35037 20039 35071
rect 19981 35031 20039 35037
rect 16206 34960 16212 35012
rect 16264 34960 16270 35012
rect 18046 34960 18052 35012
rect 18104 34960 18110 35012
rect 18138 34960 18144 35012
rect 18196 35000 18202 35012
rect 19429 35003 19487 35009
rect 19429 35000 19441 35003
rect 18196 34972 19441 35000
rect 18196 34960 18202 34972
rect 19429 34969 19441 34972
rect 19475 34969 19487 35003
rect 19429 34963 19487 34969
rect 19797 35003 19855 35009
rect 19797 34969 19809 35003
rect 19843 34969 19855 35003
rect 19797 34963 19855 34969
rect 16390 34932 16396 34944
rect 16132 34904 16396 34932
rect 15381 34895 15439 34901
rect 16390 34892 16396 34904
rect 16448 34892 16454 34944
rect 18506 34892 18512 34944
rect 18564 34892 18570 34944
rect 18598 34892 18604 34944
rect 18656 34932 18662 34944
rect 18966 34932 18972 34944
rect 18656 34904 18972 34932
rect 18656 34892 18662 34904
rect 18966 34892 18972 34904
rect 19024 34892 19030 34944
rect 19812 34932 19840 34963
rect 21266 34932 21272 34944
rect 19812 34904 21272 34932
rect 21266 34892 21272 34904
rect 21324 34892 21330 34944
rect 1104 34842 21043 34864
rect 1104 34790 5894 34842
rect 5946 34790 5958 34842
rect 6010 34790 6022 34842
rect 6074 34790 6086 34842
rect 6138 34790 6150 34842
rect 6202 34790 10839 34842
rect 10891 34790 10903 34842
rect 10955 34790 10967 34842
rect 11019 34790 11031 34842
rect 11083 34790 11095 34842
rect 11147 34790 15784 34842
rect 15836 34790 15848 34842
rect 15900 34790 15912 34842
rect 15964 34790 15976 34842
rect 16028 34790 16040 34842
rect 16092 34790 20729 34842
rect 20781 34790 20793 34842
rect 20845 34790 20857 34842
rect 20909 34790 20921 34842
rect 20973 34790 20985 34842
rect 21037 34790 21043 34842
rect 1104 34768 21043 34790
rect 1762 34688 1768 34740
rect 1820 34728 1826 34740
rect 1820 34700 3372 34728
rect 1820 34688 1826 34700
rect 2590 34660 2596 34672
rect 2516 34632 2596 34660
rect 1210 34552 1216 34604
rect 1268 34592 1274 34604
rect 1397 34595 1455 34601
rect 1397 34592 1409 34595
rect 1268 34564 1409 34592
rect 1268 34552 1274 34564
rect 1397 34561 1409 34564
rect 1443 34561 1455 34595
rect 1397 34555 1455 34561
rect 1946 34552 1952 34604
rect 2004 34552 2010 34604
rect 2314 34552 2320 34604
rect 2372 34592 2378 34604
rect 2516 34601 2544 34632
rect 2590 34620 2596 34632
rect 2648 34620 2654 34672
rect 3050 34620 3056 34672
rect 3108 34620 3114 34672
rect 3344 34660 3372 34700
rect 3418 34688 3424 34740
rect 3476 34728 3482 34740
rect 5258 34728 5264 34740
rect 3476 34700 5264 34728
rect 3476 34688 3482 34700
rect 5258 34688 5264 34700
rect 5316 34688 5322 34740
rect 5442 34688 5448 34740
rect 5500 34688 5506 34740
rect 6730 34688 6736 34740
rect 6788 34728 6794 34740
rect 8018 34728 8024 34740
rect 6788 34700 8024 34728
rect 6788 34688 6794 34700
rect 8018 34688 8024 34700
rect 8076 34728 8082 34740
rect 8205 34731 8263 34737
rect 8205 34728 8217 34731
rect 8076 34700 8217 34728
rect 8076 34688 8082 34700
rect 8205 34697 8217 34700
rect 8251 34697 8263 34731
rect 8205 34691 8263 34697
rect 8849 34731 8907 34737
rect 8849 34697 8861 34731
rect 8895 34728 8907 34731
rect 8938 34728 8944 34740
rect 8895 34700 8944 34728
rect 8895 34697 8907 34700
rect 8849 34691 8907 34697
rect 8938 34688 8944 34700
rect 8996 34688 9002 34740
rect 9122 34688 9128 34740
rect 9180 34728 9186 34740
rect 9950 34728 9956 34740
rect 9180 34700 9628 34728
rect 9180 34688 9186 34700
rect 4157 34663 4215 34669
rect 3344 34632 4108 34660
rect 2501 34595 2559 34601
rect 2501 34592 2513 34595
rect 2372 34564 2513 34592
rect 2372 34552 2378 34564
rect 2501 34561 2513 34564
rect 2547 34561 2559 34595
rect 2501 34555 2559 34561
rect 2775 34595 2833 34601
rect 2775 34561 2787 34595
rect 2821 34592 2833 34595
rect 3068 34592 3096 34620
rect 2821 34564 3096 34592
rect 2821 34561 2833 34564
rect 2775 34555 2833 34561
rect 3326 34552 3332 34604
rect 3384 34592 3390 34604
rect 3881 34595 3939 34601
rect 3881 34592 3893 34595
rect 3384 34564 3893 34592
rect 3384 34552 3390 34564
rect 3881 34561 3893 34564
rect 3927 34561 3939 34595
rect 4080 34592 4108 34632
rect 4157 34629 4169 34663
rect 4203 34660 4215 34663
rect 4614 34660 4620 34672
rect 4203 34632 4620 34660
rect 4203 34629 4215 34632
rect 4157 34623 4215 34629
rect 4614 34620 4620 34632
rect 4672 34660 4678 34672
rect 7101 34663 7159 34669
rect 4672 34632 5304 34660
rect 4672 34620 4678 34632
rect 5276 34604 5304 34632
rect 7101 34629 7113 34663
rect 7147 34660 7159 34663
rect 7282 34660 7288 34672
rect 7147 34632 7288 34660
rect 7147 34629 7159 34632
rect 7101 34623 7159 34629
rect 7282 34620 7288 34632
rect 7340 34620 7346 34672
rect 7374 34620 7380 34672
rect 7432 34620 7438 34672
rect 7469 34663 7527 34669
rect 7469 34629 7481 34663
rect 7515 34660 7527 34663
rect 8294 34660 8300 34672
rect 7515 34632 8300 34660
rect 7515 34629 7527 34632
rect 7469 34623 7527 34629
rect 8294 34620 8300 34632
rect 8352 34620 8358 34672
rect 9600 34669 9628 34700
rect 9692 34700 9956 34728
rect 9692 34669 9720 34700
rect 9950 34688 9956 34700
rect 10008 34688 10014 34740
rect 10318 34688 10324 34740
rect 10376 34728 10382 34740
rect 10413 34731 10471 34737
rect 10413 34728 10425 34731
rect 10376 34700 10425 34728
rect 10376 34688 10382 34700
rect 10413 34697 10425 34700
rect 10459 34697 10471 34731
rect 11698 34728 11704 34740
rect 10413 34691 10471 34697
rect 10888 34700 11704 34728
rect 10888 34669 10916 34700
rect 11698 34688 11704 34700
rect 11756 34688 11762 34740
rect 12710 34688 12716 34740
rect 12768 34728 12774 34740
rect 12805 34731 12863 34737
rect 12805 34728 12817 34731
rect 12768 34700 12817 34728
rect 12768 34688 12774 34700
rect 12805 34697 12817 34700
rect 12851 34697 12863 34731
rect 12805 34691 12863 34697
rect 18417 34731 18475 34737
rect 18417 34697 18429 34731
rect 18463 34728 18475 34731
rect 19334 34728 19340 34740
rect 18463 34700 19340 34728
rect 18463 34697 18475 34700
rect 18417 34691 18475 34697
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 19429 34731 19487 34737
rect 19429 34697 19441 34731
rect 19475 34728 19487 34731
rect 20530 34728 20536 34740
rect 19475 34700 20536 34728
rect 19475 34697 19487 34700
rect 19429 34691 19487 34697
rect 20530 34688 20536 34700
rect 20588 34688 20594 34740
rect 9309 34663 9367 34669
rect 9309 34629 9321 34663
rect 9355 34629 9367 34663
rect 9309 34623 9367 34629
rect 9585 34663 9643 34669
rect 9585 34629 9597 34663
rect 9631 34629 9643 34663
rect 9585 34623 9643 34629
rect 9677 34663 9735 34669
rect 9677 34629 9689 34663
rect 9723 34629 9735 34663
rect 10873 34663 10931 34669
rect 10873 34660 10885 34663
rect 9677 34623 9735 34629
rect 9766 34632 10885 34660
rect 4433 34595 4491 34601
rect 4433 34592 4445 34595
rect 4080 34564 4445 34592
rect 3881 34555 3939 34561
rect 4433 34561 4445 34564
rect 4479 34561 4491 34595
rect 4433 34555 4491 34561
rect 1673 34527 1731 34533
rect 1673 34493 1685 34527
rect 1719 34524 1731 34527
rect 1762 34524 1768 34536
rect 1719 34496 1768 34524
rect 1719 34493 1731 34496
rect 1673 34487 1731 34493
rect 1762 34484 1768 34496
rect 1820 34484 1826 34536
rect 2225 34527 2283 34533
rect 2225 34493 2237 34527
rect 2271 34524 2283 34527
rect 2406 34524 2412 34536
rect 2271 34496 2412 34524
rect 2271 34493 2283 34496
rect 2225 34487 2283 34493
rect 2406 34484 2412 34496
rect 2464 34484 2470 34536
rect 1486 34348 1492 34400
rect 1544 34388 1550 34400
rect 3418 34388 3424 34400
rect 1544 34360 3424 34388
rect 1544 34348 1550 34360
rect 3418 34348 3424 34360
rect 3476 34348 3482 34400
rect 3513 34391 3571 34397
rect 3513 34357 3525 34391
rect 3559 34388 3571 34391
rect 3878 34388 3884 34400
rect 3559 34360 3884 34388
rect 3559 34357 3571 34360
rect 3513 34351 3571 34357
rect 3878 34348 3884 34360
rect 3936 34348 3942 34400
rect 4448 34388 4476 34555
rect 4706 34552 4712 34604
rect 4764 34592 4770 34604
rect 4764 34564 5194 34592
rect 4764 34552 4770 34564
rect 5166 34524 5194 34564
rect 5258 34552 5264 34604
rect 5316 34592 5322 34604
rect 7742 34592 7748 34604
rect 5316 34564 7748 34592
rect 5316 34552 5322 34564
rect 7742 34552 7748 34564
rect 7800 34552 7806 34604
rect 7834 34552 7840 34604
rect 7892 34552 7898 34604
rect 8573 34595 8631 34601
rect 8573 34561 8585 34595
rect 8619 34592 8631 34595
rect 9324 34592 9352 34623
rect 9766 34592 9794 34632
rect 10873 34629 10885 34632
rect 10919 34629 10931 34663
rect 10873 34623 10931 34629
rect 11422 34620 11428 34672
rect 11480 34620 11486 34672
rect 12526 34660 12532 34672
rect 11716 34632 12532 34660
rect 8619 34564 8984 34592
rect 9324 34564 9794 34592
rect 8619 34561 8631 34564
rect 8573 34555 8631 34561
rect 8956 34536 8984 34564
rect 9858 34552 9864 34604
rect 9916 34592 9922 34604
rect 10045 34595 10103 34601
rect 10045 34592 10057 34595
rect 9916 34564 10057 34592
rect 9916 34552 9922 34564
rect 10045 34561 10057 34564
rect 10091 34561 10103 34595
rect 11440 34592 11468 34620
rect 11716 34592 11744 34632
rect 12526 34620 12532 34632
rect 12584 34620 12590 34672
rect 18046 34660 18052 34672
rect 13004 34632 18052 34660
rect 11781 34595 11839 34601
rect 11781 34592 11793 34595
rect 11440 34564 11793 34592
rect 10045 34555 10103 34561
rect 11781 34561 11793 34564
rect 11827 34561 11839 34595
rect 11781 34555 11839 34561
rect 12067 34595 12125 34601
rect 12067 34561 12079 34595
rect 12113 34592 12125 34595
rect 12158 34592 12164 34604
rect 12113 34564 12164 34592
rect 12113 34561 12125 34564
rect 12067 34555 12125 34561
rect 12158 34552 12164 34564
rect 12216 34592 12222 34604
rect 13004 34592 13032 34632
rect 18046 34620 18052 34632
rect 18104 34620 18110 34672
rect 18506 34660 18512 34672
rect 18156 34632 18512 34660
rect 12216 34564 13032 34592
rect 12216 34552 12222 34564
rect 13814 34552 13820 34604
rect 13872 34592 13878 34604
rect 13909 34595 13967 34601
rect 13909 34592 13921 34595
rect 13872 34564 13921 34592
rect 13872 34552 13878 34564
rect 13909 34561 13921 34564
rect 13955 34561 13967 34595
rect 13909 34555 13967 34561
rect 14183 34595 14241 34601
rect 14183 34561 14195 34595
rect 14229 34592 14241 34595
rect 14274 34592 14280 34604
rect 14229 34564 14280 34592
rect 14229 34561 14241 34564
rect 14183 34555 14241 34561
rect 14274 34552 14280 34564
rect 14332 34552 14338 34604
rect 16666 34552 16672 34604
rect 16724 34552 16730 34604
rect 16942 34601 16948 34604
rect 16936 34592 16948 34601
rect 16903 34564 16948 34592
rect 16936 34555 16948 34564
rect 16942 34552 16948 34555
rect 17000 34552 17006 34604
rect 18156 34601 18184 34632
rect 18506 34620 18512 34632
rect 18564 34660 18570 34672
rect 18564 34632 18828 34660
rect 18564 34620 18570 34632
rect 18800 34601 18828 34632
rect 19518 34620 19524 34672
rect 19576 34660 19582 34672
rect 20165 34663 20223 34669
rect 20165 34660 20177 34663
rect 19576 34632 20177 34660
rect 19576 34620 19582 34632
rect 20165 34629 20177 34632
rect 20211 34629 20223 34663
rect 20165 34623 20223 34629
rect 18141 34595 18199 34601
rect 18141 34561 18153 34595
rect 18187 34561 18199 34595
rect 18693 34595 18751 34601
rect 18693 34592 18705 34595
rect 18141 34555 18199 34561
rect 18340 34564 18705 34592
rect 5902 34524 5908 34536
rect 5166 34496 5908 34524
rect 5902 34484 5908 34496
rect 5960 34484 5966 34536
rect 7558 34484 7564 34536
rect 7616 34484 7622 34536
rect 8846 34484 8852 34536
rect 8904 34484 8910 34536
rect 8938 34484 8944 34536
rect 8996 34484 9002 34536
rect 9950 34484 9956 34536
rect 10008 34484 10014 34536
rect 11054 34484 11060 34536
rect 11112 34484 11118 34536
rect 15010 34484 15016 34536
rect 15068 34524 15074 34536
rect 18340 34524 18368 34564
rect 18693 34561 18705 34564
rect 18739 34561 18751 34595
rect 18693 34555 18751 34561
rect 18785 34595 18843 34601
rect 18785 34561 18797 34595
rect 18831 34561 18843 34595
rect 18785 34555 18843 34561
rect 18969 34595 19027 34601
rect 18969 34561 18981 34595
rect 19015 34561 19027 34595
rect 18969 34555 19027 34561
rect 15068 34496 15792 34524
rect 15068 34484 15074 34496
rect 9030 34456 9036 34468
rect 8404 34428 9036 34456
rect 4890 34388 4896 34400
rect 4448 34360 4896 34388
rect 4890 34348 4896 34360
rect 4948 34348 4954 34400
rect 8404 34397 8432 34428
rect 9030 34416 9036 34428
rect 9088 34416 9094 34468
rect 15764 34456 15792 34496
rect 18064 34496 18368 34524
rect 18417 34527 18475 34533
rect 16574 34456 16580 34468
rect 15764 34428 16580 34456
rect 16574 34416 16580 34428
rect 16632 34416 16638 34468
rect 18064 34465 18092 34496
rect 18417 34493 18429 34527
rect 18463 34524 18475 34527
rect 18877 34527 18935 34533
rect 18877 34524 18889 34527
rect 18463 34496 18889 34524
rect 18463 34493 18475 34496
rect 18417 34487 18475 34493
rect 18877 34493 18889 34496
rect 18923 34493 18935 34527
rect 18877 34487 18935 34493
rect 18049 34459 18107 34465
rect 18049 34425 18061 34459
rect 18095 34425 18107 34459
rect 18049 34419 18107 34425
rect 18509 34459 18567 34465
rect 18509 34425 18521 34459
rect 18555 34456 18567 34459
rect 18984 34456 19012 34555
rect 19334 34552 19340 34604
rect 19392 34552 19398 34604
rect 19426 34552 19432 34604
rect 19484 34592 19490 34604
rect 19613 34595 19671 34601
rect 19613 34592 19625 34595
rect 19484 34564 19625 34592
rect 19484 34552 19490 34564
rect 19613 34561 19625 34564
rect 19659 34561 19671 34595
rect 19613 34555 19671 34561
rect 19886 34552 19892 34604
rect 19944 34552 19950 34604
rect 18555 34428 19012 34456
rect 18555 34425 18567 34428
rect 18509 34419 18567 34425
rect 8389 34391 8447 34397
rect 8389 34357 8401 34391
rect 8435 34357 8447 34391
rect 8389 34351 8447 34357
rect 8665 34391 8723 34397
rect 8665 34357 8677 34391
rect 8711 34388 8723 34391
rect 9306 34388 9312 34400
rect 8711 34360 9312 34388
rect 8711 34357 8723 34360
rect 8665 34351 8723 34357
rect 9306 34348 9312 34360
rect 9364 34348 9370 34400
rect 10594 34348 10600 34400
rect 10652 34388 10658 34400
rect 12250 34388 12256 34400
rect 10652 34360 12256 34388
rect 10652 34348 10658 34360
rect 12250 34348 12256 34360
rect 12308 34348 12314 34400
rect 12710 34348 12716 34400
rect 12768 34388 12774 34400
rect 12986 34388 12992 34400
rect 12768 34360 12992 34388
rect 12768 34348 12774 34360
rect 12986 34348 12992 34360
rect 13044 34388 13050 34400
rect 14274 34388 14280 34400
rect 13044 34360 14280 34388
rect 13044 34348 13050 34360
rect 14274 34348 14280 34360
rect 14332 34348 14338 34400
rect 14921 34391 14979 34397
rect 14921 34357 14933 34391
rect 14967 34388 14979 34391
rect 15010 34388 15016 34400
rect 14967 34360 15016 34388
rect 14967 34357 14979 34360
rect 14921 34351 14979 34357
rect 15010 34348 15016 34360
rect 15068 34348 15074 34400
rect 17586 34348 17592 34400
rect 17644 34388 17650 34400
rect 18233 34391 18291 34397
rect 18233 34388 18245 34391
rect 17644 34360 18245 34388
rect 17644 34348 17650 34360
rect 18233 34357 18245 34360
rect 18279 34357 18291 34391
rect 18233 34351 18291 34357
rect 18690 34348 18696 34400
rect 18748 34388 18754 34400
rect 19153 34391 19211 34397
rect 19153 34388 19165 34391
rect 18748 34360 19165 34388
rect 18748 34348 18754 34360
rect 19153 34357 19165 34360
rect 19199 34357 19211 34391
rect 19153 34351 19211 34357
rect 19705 34391 19763 34397
rect 19705 34357 19717 34391
rect 19751 34388 19763 34391
rect 20346 34388 20352 34400
rect 19751 34360 20352 34388
rect 19751 34357 19763 34360
rect 19705 34351 19763 34357
rect 20346 34348 20352 34360
rect 20404 34348 20410 34400
rect 20438 34348 20444 34400
rect 20496 34348 20502 34400
rect 1104 34298 20884 34320
rect 1104 34246 3422 34298
rect 3474 34246 3486 34298
rect 3538 34246 3550 34298
rect 3602 34246 3614 34298
rect 3666 34246 3678 34298
rect 3730 34246 8367 34298
rect 8419 34246 8431 34298
rect 8483 34246 8495 34298
rect 8547 34246 8559 34298
rect 8611 34246 8623 34298
rect 8675 34246 13312 34298
rect 13364 34246 13376 34298
rect 13428 34246 13440 34298
rect 13492 34246 13504 34298
rect 13556 34246 13568 34298
rect 13620 34246 18257 34298
rect 18309 34246 18321 34298
rect 18373 34246 18385 34298
rect 18437 34246 18449 34298
rect 18501 34246 18513 34298
rect 18565 34246 20884 34298
rect 1104 34224 20884 34246
rect 1688 34156 4292 34184
rect 1688 34057 1716 34156
rect 1673 34051 1731 34057
rect 1673 34017 1685 34051
rect 1719 34017 1731 34051
rect 1673 34011 1731 34017
rect 2314 34008 2320 34060
rect 2372 34008 2378 34060
rect 4264 33992 4292 34156
rect 4430 34144 4436 34196
rect 4488 34184 4494 34196
rect 4617 34187 4675 34193
rect 4617 34184 4629 34187
rect 4488 34156 4629 34184
rect 4488 34144 4494 34156
rect 4617 34153 4629 34156
rect 4663 34153 4675 34187
rect 8570 34184 8576 34196
rect 4617 34147 4675 34153
rect 4816 34156 8576 34184
rect 1394 33940 1400 33992
rect 1452 33940 1458 33992
rect 3234 33980 3240 33992
rect 2606 33959 3240 33980
rect 2575 33953 3240 33959
rect 2575 33950 2587 33953
rect 2038 33872 2044 33924
rect 2096 33912 2102 33924
rect 2516 33922 2587 33950
rect 2516 33912 2544 33922
rect 2575 33919 2587 33922
rect 2621 33952 3240 33953
rect 2621 33922 2634 33952
rect 3234 33940 3240 33952
rect 3292 33940 3298 33992
rect 3789 33983 3847 33989
rect 3789 33949 3801 33983
rect 3835 33949 3847 33983
rect 3789 33943 3847 33949
rect 2621 33919 2633 33922
rect 2575 33913 2633 33919
rect 3804 33912 3832 33943
rect 4246 33940 4252 33992
rect 4304 33940 4310 33992
rect 4614 33940 4620 33992
rect 4672 33980 4678 33992
rect 4816 33989 4844 34156
rect 8570 34144 8576 34156
rect 8628 34144 8634 34196
rect 8665 34187 8723 34193
rect 8665 34153 8677 34187
rect 8711 34184 8723 34187
rect 8846 34184 8852 34196
rect 8711 34156 8852 34184
rect 8711 34153 8723 34156
rect 8665 34147 8723 34153
rect 8846 34144 8852 34156
rect 8904 34144 8910 34196
rect 9306 34144 9312 34196
rect 9364 34184 9370 34196
rect 9364 34156 9720 34184
rect 9364 34144 9370 34156
rect 6546 34076 6552 34128
rect 6604 34076 6610 34128
rect 6822 34076 6828 34128
rect 6880 34116 6886 34128
rect 7098 34116 7104 34128
rect 6880 34088 7104 34116
rect 6880 34076 6886 34088
rect 7098 34076 7104 34088
rect 7156 34116 7162 34128
rect 7193 34119 7251 34125
rect 7193 34116 7205 34119
rect 7156 34088 7205 34116
rect 7156 34076 7162 34088
rect 7193 34085 7205 34088
rect 7239 34085 7251 34119
rect 7193 34079 7251 34085
rect 8389 34119 8447 34125
rect 8389 34085 8401 34119
rect 8435 34116 8447 34119
rect 8754 34116 8760 34128
rect 8435 34088 8760 34116
rect 8435 34085 8447 34088
rect 8389 34079 8447 34085
rect 8754 34076 8760 34088
rect 8812 34076 8818 34128
rect 9692 34116 9720 34156
rect 9950 34144 9956 34196
rect 10008 34184 10014 34196
rect 10045 34187 10103 34193
rect 10045 34184 10057 34187
rect 10008 34156 10057 34184
rect 10008 34144 10014 34156
rect 10045 34153 10057 34156
rect 10091 34153 10103 34187
rect 10045 34147 10103 34153
rect 10134 34144 10140 34196
rect 10192 34184 10198 34196
rect 10410 34184 10416 34196
rect 10192 34156 10416 34184
rect 10192 34144 10198 34156
rect 10410 34144 10416 34156
rect 10468 34144 10474 34196
rect 13725 34187 13783 34193
rect 13725 34153 13737 34187
rect 13771 34184 13783 34187
rect 15378 34184 15384 34196
rect 13771 34156 15384 34184
rect 13771 34153 13783 34156
rect 13725 34147 13783 34153
rect 15378 34144 15384 34156
rect 15436 34144 15442 34196
rect 16574 34144 16580 34196
rect 16632 34184 16638 34196
rect 16850 34184 16856 34196
rect 16632 34156 16856 34184
rect 16632 34144 16638 34156
rect 16850 34144 16856 34156
rect 16908 34144 16914 34196
rect 17586 34144 17592 34196
rect 17644 34144 17650 34196
rect 17773 34187 17831 34193
rect 17773 34153 17785 34187
rect 17819 34184 17831 34187
rect 18506 34184 18512 34196
rect 17819 34156 18512 34184
rect 17819 34153 17831 34156
rect 17773 34147 17831 34153
rect 18506 34144 18512 34156
rect 18564 34144 18570 34196
rect 18601 34187 18659 34193
rect 18601 34153 18613 34187
rect 18647 34184 18659 34187
rect 19334 34184 19340 34196
rect 18647 34156 19340 34184
rect 18647 34153 18659 34156
rect 18601 34147 18659 34153
rect 19334 34144 19340 34156
rect 19392 34144 19398 34196
rect 19518 34144 19524 34196
rect 19576 34144 19582 34196
rect 19610 34144 19616 34196
rect 19668 34144 19674 34196
rect 10505 34119 10563 34125
rect 10505 34116 10517 34119
rect 9692 34088 10517 34116
rect 10505 34085 10517 34088
rect 10551 34085 10563 34119
rect 10505 34079 10563 34085
rect 13814 34076 13820 34128
rect 13872 34076 13878 34128
rect 18049 34119 18107 34125
rect 18049 34085 18061 34119
rect 18095 34116 18107 34119
rect 18095 34088 19012 34116
rect 18095 34085 18107 34088
rect 18049 34079 18107 34085
rect 4890 34008 4896 34060
rect 4948 34048 4954 34060
rect 4985 34051 5043 34057
rect 4985 34048 4997 34051
rect 4948 34020 4997 34048
rect 4948 34008 4954 34020
rect 4985 34017 4997 34020
rect 5031 34017 5043 34051
rect 6564 34048 6592 34076
rect 7466 34048 7472 34060
rect 6564 34020 7472 34048
rect 4985 34011 5043 34017
rect 7466 34008 7472 34020
rect 7524 34008 7530 34060
rect 7650 34057 7656 34060
rect 7607 34051 7656 34057
rect 7607 34017 7619 34051
rect 7653 34017 7656 34051
rect 7607 34011 7656 34017
rect 7650 34008 7656 34011
rect 7708 34008 7714 34060
rect 7926 34048 7932 34060
rect 7760 34020 7932 34048
rect 4801 33983 4859 33989
rect 4801 33980 4813 33983
rect 4672 33952 4813 33980
rect 4672 33940 4678 33952
rect 4801 33949 4813 33952
rect 4847 33949 4859 33983
rect 5258 33980 5264 33992
rect 5219 33952 5264 33980
rect 4801 33943 4859 33949
rect 5258 33940 5264 33952
rect 5316 33940 5322 33992
rect 6549 33983 6607 33989
rect 6549 33949 6561 33983
rect 6595 33980 6607 33983
rect 6638 33980 6644 33992
rect 6595 33952 6644 33980
rect 6595 33949 6607 33952
rect 6549 33943 6607 33949
rect 6638 33940 6644 33952
rect 6696 33940 6702 33992
rect 6730 33940 6736 33992
rect 6788 33940 6794 33992
rect 7760 33989 7788 34020
rect 7926 34008 7932 34020
rect 7984 34008 7990 34060
rect 8110 34008 8116 34060
rect 8168 34048 8174 34060
rect 8662 34048 8668 34060
rect 8168 34020 8668 34048
rect 8168 34008 8174 34020
rect 8662 34008 8668 34020
rect 8720 34048 8726 34060
rect 8720 34020 8890 34048
rect 8720 34008 8726 34020
rect 7745 33983 7803 33989
rect 7745 33949 7757 33983
rect 7791 33949 7803 33983
rect 7745 33943 7803 33949
rect 8573 33983 8631 33989
rect 8573 33949 8585 33983
rect 8619 33949 8631 33983
rect 8573 33943 8631 33949
rect 2096 33884 2544 33912
rect 2746 33884 3832 33912
rect 4065 33915 4123 33921
rect 2096 33872 2102 33884
rect 1302 33804 1308 33856
rect 1360 33844 1366 33856
rect 2746 33844 2774 33884
rect 4065 33881 4077 33915
rect 4111 33912 4123 33915
rect 4111 33884 6776 33912
rect 4111 33881 4123 33884
rect 4065 33875 4123 33881
rect 1360 33816 2774 33844
rect 1360 33804 1366 33816
rect 3326 33804 3332 33856
rect 3384 33804 3390 33856
rect 4154 33804 4160 33856
rect 4212 33844 4218 33856
rect 4614 33844 4620 33856
rect 4212 33816 4620 33844
rect 4212 33804 4218 33816
rect 4614 33804 4620 33816
rect 4672 33804 4678 33856
rect 5534 33804 5540 33856
rect 5592 33844 5598 33856
rect 5997 33847 6055 33853
rect 5997 33844 6009 33847
rect 5592 33816 6009 33844
rect 5592 33804 5598 33816
rect 5997 33813 6009 33816
rect 6043 33813 6055 33847
rect 6748 33844 6776 33884
rect 8478 33844 8484 33856
rect 6748 33816 8484 33844
rect 5997 33807 6055 33813
rect 8478 33804 8484 33816
rect 8536 33804 8542 33856
rect 8588 33844 8616 33943
rect 8754 33940 8760 33992
rect 8812 33940 8818 33992
rect 8862 33980 8890 34020
rect 9766 34008 9772 34060
rect 9824 34048 9830 34060
rect 9824 34020 10456 34048
rect 9824 34008 9830 34020
rect 9033 33983 9091 33989
rect 9033 33980 9045 33983
rect 8862 33952 9045 33980
rect 9033 33949 9045 33952
rect 9079 33949 9091 33983
rect 9033 33943 9091 33949
rect 9307 33973 9365 33979
rect 9307 33939 9319 33973
rect 9353 33939 9365 33973
rect 9398 33940 9404 33992
rect 9456 33980 9462 33992
rect 10318 33980 10324 33992
rect 9456 33952 10324 33980
rect 9456 33940 9462 33952
rect 10318 33940 10324 33952
rect 10376 33940 10382 33992
rect 10428 33989 10456 34020
rect 12526 34008 12532 34060
rect 12584 34048 12590 34060
rect 13722 34048 13728 34060
rect 12584 34020 13728 34048
rect 12584 34008 12590 34020
rect 13722 34008 13728 34020
rect 13780 34008 13786 34060
rect 13906 34008 13912 34060
rect 13964 34008 13970 34060
rect 16758 34048 16764 34060
rect 16132 34020 16764 34048
rect 10413 33983 10471 33989
rect 10413 33949 10425 33983
rect 10459 33949 10471 33983
rect 10413 33943 10471 33949
rect 10781 33983 10839 33989
rect 10781 33949 10793 33983
rect 10827 33949 10839 33983
rect 10781 33943 10839 33949
rect 11055 33983 11113 33989
rect 11055 33949 11067 33983
rect 11101 33980 11113 33983
rect 13633 33983 13691 33989
rect 11101 33952 13308 33980
rect 11101 33949 11113 33952
rect 11055 33943 11113 33949
rect 9307 33933 9365 33939
rect 8938 33844 8944 33856
rect 8588 33816 8944 33844
rect 8938 33804 8944 33816
rect 8996 33804 9002 33856
rect 9324 33844 9352 33933
rect 10796 33912 10824 33943
rect 11238 33912 11244 33924
rect 10796 33884 11244 33912
rect 11238 33872 11244 33884
rect 11296 33872 11302 33924
rect 9490 33844 9496 33856
rect 9324 33816 9496 33844
rect 9490 33804 9496 33816
rect 9548 33844 9554 33856
rect 11346 33844 11374 33952
rect 11606 33872 11612 33924
rect 11664 33912 11670 33924
rect 12158 33912 12164 33924
rect 11664 33884 12164 33912
rect 11664 33872 11670 33884
rect 12158 33872 12164 33884
rect 12216 33872 12222 33924
rect 9548 33816 11374 33844
rect 9548 33804 9554 33816
rect 11790 33804 11796 33856
rect 11848 33804 11854 33856
rect 12618 33804 12624 33856
rect 12676 33844 12682 33856
rect 13170 33844 13176 33856
rect 12676 33816 13176 33844
rect 12676 33804 12682 33816
rect 13170 33804 13176 33816
rect 13228 33804 13234 33856
rect 13280 33844 13308 33952
rect 13633 33949 13645 33983
rect 13679 33949 13691 33983
rect 13740 33980 13768 34008
rect 14093 33983 14151 33989
rect 14093 33980 14105 33983
rect 13740 33952 14105 33980
rect 13633 33943 13691 33949
rect 14093 33949 14105 33952
rect 14139 33949 14151 33983
rect 14093 33943 14151 33949
rect 14367 33983 14425 33989
rect 14367 33949 14379 33983
rect 14413 33980 14425 33983
rect 14413 33952 14596 33980
rect 14413 33949 14425 33952
rect 14367 33943 14425 33949
rect 13648 33912 13676 33943
rect 14568 33924 14596 33952
rect 14734 33940 14740 33992
rect 14792 33980 14798 33992
rect 15473 33983 15531 33989
rect 15473 33980 15485 33983
rect 14792 33952 15485 33980
rect 14792 33940 14798 33952
rect 15473 33949 15485 33952
rect 15519 33949 15531 33983
rect 15473 33943 15531 33949
rect 15654 33940 15660 33992
rect 15712 33980 15718 33992
rect 15747 33983 15805 33989
rect 15747 33980 15759 33983
rect 15712 33952 15759 33980
rect 15712 33940 15718 33952
rect 15747 33949 15759 33952
rect 15793 33980 15805 33983
rect 16132 33980 16160 34020
rect 16758 34008 16764 34020
rect 16816 34048 16822 34060
rect 16816 34020 18000 34048
rect 16816 34008 16822 34020
rect 16942 33980 16948 33992
rect 15793 33952 16160 33980
rect 16592 33952 16948 33980
rect 15793 33949 15805 33952
rect 15747 33943 15805 33949
rect 16592 33924 16620 33952
rect 16942 33940 16948 33952
rect 17000 33980 17006 33992
rect 17972 33989 18000 34020
rect 18598 34008 18604 34060
rect 18656 34048 18662 34060
rect 18984 34048 19012 34088
rect 19150 34076 19156 34128
rect 19208 34116 19214 34128
rect 19628 34116 19656 34144
rect 19208 34088 19656 34116
rect 19208 34076 19214 34088
rect 20070 34048 20076 34060
rect 18656 34020 18828 34048
rect 18984 34020 20076 34048
rect 18656 34008 18662 34020
rect 17037 33983 17095 33989
rect 17037 33980 17049 33983
rect 17000 33952 17049 33980
rect 17000 33940 17006 33952
rect 17037 33949 17049 33952
rect 17083 33949 17095 33983
rect 17037 33943 17095 33949
rect 17497 33983 17555 33989
rect 17497 33949 17509 33983
rect 17543 33949 17555 33983
rect 17497 33943 17555 33949
rect 17957 33983 18015 33989
rect 17957 33949 17969 33983
rect 18003 33949 18015 33983
rect 17957 33943 18015 33949
rect 13814 33912 13820 33924
rect 13648 33884 13820 33912
rect 13814 33872 13820 33884
rect 13872 33872 13878 33924
rect 14550 33872 14556 33924
rect 14608 33872 14614 33924
rect 16574 33872 16580 33924
rect 16632 33872 16638 33924
rect 17512 33912 17540 33943
rect 18230 33940 18236 33992
rect 18288 33940 18294 33992
rect 18509 33983 18567 33989
rect 18509 33949 18521 33983
rect 18555 33980 18567 33983
rect 18690 33980 18696 33992
rect 18555 33952 18696 33980
rect 18555 33949 18567 33952
rect 18509 33943 18567 33949
rect 18690 33940 18696 33952
rect 18748 33940 18754 33992
rect 18800 33989 18828 34020
rect 20070 34008 20076 34020
rect 20128 34008 20134 34060
rect 18785 33983 18843 33989
rect 18785 33949 18797 33983
rect 18831 33949 18843 33983
rect 18785 33943 18843 33949
rect 18874 33940 18880 33992
rect 18932 33980 18938 33992
rect 19061 33983 19119 33989
rect 19061 33980 19073 33983
rect 18932 33952 19073 33980
rect 18932 33940 18938 33952
rect 19061 33949 19073 33952
rect 19107 33949 19119 33983
rect 19061 33943 19119 33949
rect 19426 33940 19432 33992
rect 19484 33940 19490 33992
rect 19610 33940 19616 33992
rect 19668 33940 19674 33992
rect 19981 33983 20039 33989
rect 19981 33949 19993 33983
rect 20027 33980 20039 33983
rect 20162 33980 20168 33992
rect 20027 33952 20168 33980
rect 20027 33949 20039 33952
rect 19981 33943 20039 33949
rect 20162 33940 20168 33952
rect 20220 33940 20226 33992
rect 20257 33983 20315 33989
rect 20257 33949 20269 33983
rect 20303 33949 20315 33983
rect 20257 33943 20315 33949
rect 20272 33912 20300 33943
rect 16868 33884 17540 33912
rect 18340 33884 19380 33912
rect 14568 33844 14596 33872
rect 13280 33816 14596 33844
rect 14734 33804 14740 33856
rect 14792 33844 14798 33856
rect 15105 33847 15163 33853
rect 15105 33844 15117 33847
rect 14792 33816 15117 33844
rect 14792 33804 14798 33816
rect 15105 33813 15117 33816
rect 15151 33813 15163 33847
rect 15105 33807 15163 33813
rect 15194 33804 15200 33856
rect 15252 33844 15258 33856
rect 16868 33853 16896 33884
rect 16485 33847 16543 33853
rect 16485 33844 16497 33847
rect 15252 33816 16497 33844
rect 15252 33804 15258 33816
rect 16485 33813 16497 33816
rect 16531 33813 16543 33847
rect 16485 33807 16543 33813
rect 16853 33847 16911 33853
rect 16853 33813 16865 33847
rect 16899 33813 16911 33847
rect 16853 33807 16911 33813
rect 17126 33804 17132 33856
rect 17184 33844 17190 33856
rect 17586 33844 17592 33856
rect 17184 33816 17592 33844
rect 17184 33804 17190 33816
rect 17586 33804 17592 33816
rect 17644 33804 17650 33856
rect 18340 33853 18368 33884
rect 18325 33847 18383 33853
rect 18325 33813 18337 33847
rect 18371 33813 18383 33847
rect 18325 33807 18383 33813
rect 18877 33847 18935 33853
rect 18877 33813 18889 33847
rect 18923 33844 18935 33847
rect 19150 33844 19156 33856
rect 18923 33816 19156 33844
rect 18923 33813 18935 33816
rect 18877 33807 18935 33813
rect 19150 33804 19156 33816
rect 19208 33804 19214 33856
rect 19352 33844 19380 33884
rect 19628 33884 20300 33912
rect 19628 33844 19656 33884
rect 19352 33816 19656 33844
rect 19794 33804 19800 33856
rect 19852 33804 19858 33856
rect 20441 33847 20499 33853
rect 20441 33813 20453 33847
rect 20487 33844 20499 33847
rect 21174 33844 21180 33856
rect 20487 33816 21180 33844
rect 20487 33813 20499 33816
rect 20441 33807 20499 33813
rect 21174 33804 21180 33816
rect 21232 33804 21238 33856
rect 1104 33754 21043 33776
rect 1104 33702 5894 33754
rect 5946 33702 5958 33754
rect 6010 33702 6022 33754
rect 6074 33702 6086 33754
rect 6138 33702 6150 33754
rect 6202 33702 10839 33754
rect 10891 33702 10903 33754
rect 10955 33702 10967 33754
rect 11019 33702 11031 33754
rect 11083 33702 11095 33754
rect 11147 33702 15784 33754
rect 15836 33702 15848 33754
rect 15900 33702 15912 33754
rect 15964 33702 15976 33754
rect 16028 33702 16040 33754
rect 16092 33702 20729 33754
rect 20781 33702 20793 33754
rect 20845 33702 20857 33754
rect 20909 33702 20921 33754
rect 20973 33702 20985 33754
rect 21037 33702 21043 33754
rect 1104 33680 21043 33702
rect 1670 33640 1676 33652
rect 1654 33600 1676 33640
rect 1728 33600 1734 33652
rect 3326 33600 3332 33652
rect 3384 33640 3390 33652
rect 7190 33640 7196 33652
rect 3384 33612 4108 33640
rect 3384 33600 3390 33612
rect 1654 33543 1682 33600
rect 1654 33537 1713 33543
rect 1654 33506 1667 33537
rect 1655 33503 1667 33506
rect 1701 33503 1713 33537
rect 1854 33532 1860 33584
rect 1912 33572 1918 33584
rect 3234 33572 3240 33584
rect 1912 33544 3240 33572
rect 1912 33532 1918 33544
rect 3234 33532 3240 33544
rect 3292 33532 3298 33584
rect 3694 33532 3700 33584
rect 3752 33532 3758 33584
rect 3970 33532 3976 33584
rect 4028 33532 4034 33584
rect 4080 33581 4108 33612
rect 4356 33612 7196 33640
rect 4065 33575 4123 33581
rect 4065 33541 4077 33575
rect 4111 33541 4123 33575
rect 4065 33535 4123 33541
rect 1655 33497 1713 33503
rect 2774 33464 2780 33516
rect 2832 33464 2838 33516
rect 3053 33507 3111 33513
rect 3053 33473 3065 33507
rect 3099 33504 3111 33507
rect 4356 33504 4384 33612
rect 7190 33600 7196 33612
rect 7248 33600 7254 33652
rect 7650 33600 7656 33652
rect 7708 33640 7714 33652
rect 7834 33640 7840 33652
rect 7708 33612 7840 33640
rect 7708 33600 7714 33612
rect 7834 33600 7840 33612
rect 7892 33600 7898 33652
rect 8754 33600 8760 33652
rect 8812 33640 8818 33652
rect 9953 33643 10011 33649
rect 9953 33640 9965 33643
rect 8812 33612 9965 33640
rect 8812 33600 8818 33612
rect 9953 33609 9965 33612
rect 9999 33609 10011 33643
rect 14734 33640 14740 33652
rect 9953 33603 10011 33609
rect 14200 33612 14740 33640
rect 4522 33532 4528 33584
rect 4580 33572 4586 33584
rect 4801 33575 4859 33581
rect 4801 33572 4813 33575
rect 4580 33544 4813 33572
rect 4580 33532 4586 33544
rect 4801 33541 4813 33544
rect 4847 33541 4859 33575
rect 4801 33535 4859 33541
rect 6270 33532 6276 33584
rect 6328 33572 6334 33584
rect 6822 33572 6828 33584
rect 6328 33544 6828 33572
rect 6328 33532 6334 33544
rect 3099 33476 4384 33504
rect 3099 33473 3111 33476
rect 3053 33467 3111 33473
rect 4430 33464 4436 33516
rect 4488 33504 4494 33516
rect 4982 33504 4988 33516
rect 4488 33476 4988 33504
rect 4488 33464 4494 33476
rect 4982 33464 4988 33476
rect 5040 33464 5046 33516
rect 6656 33513 6684 33544
rect 6822 33532 6828 33544
rect 6880 33532 6886 33584
rect 8481 33575 8539 33581
rect 8481 33541 8493 33575
rect 8527 33572 8539 33575
rect 12066 33572 12072 33584
rect 8527 33544 10180 33572
rect 8527 33541 8539 33544
rect 8481 33535 8539 33541
rect 6641 33507 6699 33513
rect 6641 33473 6653 33507
rect 6687 33473 6699 33507
rect 6641 33467 6699 33473
rect 7558 33464 7564 33516
rect 7616 33464 7622 33516
rect 7678 33507 7736 33513
rect 7678 33473 7690 33507
rect 7724 33473 7736 33507
rect 7678 33467 7736 33473
rect 8573 33507 8631 33513
rect 8573 33473 8585 33507
rect 8619 33473 8631 33507
rect 8846 33504 8852 33516
rect 8807 33476 8852 33504
rect 8573 33467 8631 33473
rect 1302 33396 1308 33448
rect 1360 33436 1366 33448
rect 1397 33439 1455 33445
rect 1397 33436 1409 33439
rect 1360 33408 1409 33436
rect 1360 33396 1366 33408
rect 1397 33405 1409 33408
rect 1443 33405 1455 33439
rect 1397 33399 1455 33405
rect 3878 33396 3884 33448
rect 3936 33396 3942 33448
rect 5258 33396 5264 33448
rect 5316 33436 5322 33448
rect 6825 33439 6883 33445
rect 6825 33436 6837 33439
rect 5316 33408 6837 33436
rect 5316 33396 5322 33408
rect 6825 33405 6837 33408
rect 6871 33405 6883 33439
rect 6825 33399 6883 33405
rect 7374 33396 7380 33448
rect 7432 33436 7438 33448
rect 7693 33436 7721 33467
rect 7432 33408 7721 33436
rect 7837 33439 7895 33445
rect 7432 33396 7438 33408
rect 7837 33405 7849 33439
rect 7883 33436 7895 33439
rect 8018 33436 8024 33448
rect 7883 33408 8024 33436
rect 7883 33405 7895 33408
rect 7837 33399 7895 33405
rect 8018 33396 8024 33408
rect 8076 33396 8082 33448
rect 8588 33436 8616 33467
rect 8846 33464 8852 33476
rect 8904 33464 8910 33516
rect 8938 33464 8944 33516
rect 8996 33504 9002 33516
rect 10152 33513 10180 33544
rect 11806 33544 12072 33572
rect 10137 33507 10195 33513
rect 8996 33476 9628 33504
rect 8996 33464 9002 33476
rect 8220 33408 8616 33436
rect 4985 33371 5043 33377
rect 4985 33337 4997 33371
rect 5031 33368 5043 33371
rect 5276 33368 5304 33396
rect 5031 33340 5304 33368
rect 5031 33337 5043 33340
rect 4985 33331 5043 33337
rect 7098 33328 7104 33380
rect 7156 33368 7162 33380
rect 7285 33371 7343 33377
rect 7285 33368 7297 33371
rect 7156 33340 7297 33368
rect 7156 33328 7162 33340
rect 7285 33337 7297 33340
rect 7331 33337 7343 33371
rect 7285 33331 7343 33337
rect 2406 33260 2412 33312
rect 2464 33260 2470 33312
rect 6730 33260 6736 33312
rect 6788 33300 6794 33312
rect 7558 33300 7564 33312
rect 6788 33272 7564 33300
rect 6788 33260 6794 33272
rect 7558 33260 7564 33272
rect 7616 33260 7622 33312
rect 7650 33260 7656 33312
rect 7708 33300 7714 33312
rect 8220 33300 8248 33408
rect 9600 33377 9628 33476
rect 10137 33473 10149 33507
rect 10183 33473 10195 33507
rect 10137 33467 10195 33473
rect 11238 33464 11244 33516
rect 11296 33504 11302 33516
rect 11806 33513 11834 33544
rect 12066 33532 12072 33544
rect 12124 33572 12130 33584
rect 13814 33572 13820 33584
rect 12124 33544 13820 33572
rect 12124 33532 12130 33544
rect 13814 33532 13820 33544
rect 13872 33532 13878 33584
rect 11517 33507 11575 33513
rect 11517 33504 11529 33507
rect 11296 33476 11529 33504
rect 11296 33464 11302 33476
rect 11517 33473 11529 33476
rect 11563 33473 11575 33507
rect 11517 33467 11575 33473
rect 11791 33507 11849 33513
rect 11791 33473 11803 33507
rect 11837 33473 11849 33507
rect 11791 33467 11849 33473
rect 12986 33464 12992 33516
rect 13044 33504 13050 33516
rect 14200 33504 14228 33612
rect 14734 33600 14740 33612
rect 14792 33600 14798 33652
rect 15010 33600 15016 33652
rect 15068 33640 15074 33652
rect 15841 33643 15899 33649
rect 15068 33612 15700 33640
rect 15068 33600 15074 33612
rect 15672 33572 15700 33612
rect 15841 33609 15853 33643
rect 15887 33640 15899 33643
rect 16574 33640 16580 33652
rect 15887 33612 16580 33640
rect 15887 33609 15899 33612
rect 15841 33603 15899 33609
rect 16574 33600 16580 33612
rect 16632 33600 16638 33652
rect 18230 33600 18236 33652
rect 18288 33600 18294 33652
rect 18506 33600 18512 33652
rect 18564 33600 18570 33652
rect 18601 33643 18659 33649
rect 18601 33609 18613 33643
rect 18647 33609 18659 33643
rect 18601 33603 18659 33609
rect 19153 33643 19211 33649
rect 19153 33609 19165 33643
rect 19199 33640 19211 33643
rect 19610 33640 19616 33652
rect 19199 33612 19616 33640
rect 19199 33609 19211 33612
rect 19153 33603 19211 33609
rect 15672 33544 15976 33572
rect 13044 33476 14136 33504
rect 14200 33476 14412 33504
rect 13044 33464 13050 33476
rect 13906 33396 13912 33448
rect 13964 33396 13970 33448
rect 14001 33439 14059 33445
rect 14001 33405 14013 33439
rect 14047 33405 14059 33439
rect 14108 33436 14136 33476
rect 14185 33439 14243 33445
rect 14185 33436 14197 33439
rect 14108 33408 14197 33436
rect 14001 33399 14059 33405
rect 14185 33405 14197 33408
rect 14231 33405 14243 33439
rect 14384 33436 14412 33476
rect 15194 33464 15200 33516
rect 15252 33464 15258 33516
rect 15948 33513 15976 33544
rect 15933 33507 15991 33513
rect 15933 33473 15945 33507
rect 15979 33473 15991 33507
rect 15933 33467 15991 33473
rect 16114 33464 16120 33516
rect 16172 33464 16178 33516
rect 14645 33439 14703 33445
rect 14645 33436 14657 33439
rect 14384 33408 14657 33436
rect 14185 33399 14243 33405
rect 14645 33405 14657 33408
rect 14691 33405 14703 33439
rect 14645 33399 14703 33405
rect 9585 33371 9643 33377
rect 9585 33337 9597 33371
rect 9631 33337 9643 33371
rect 9585 33331 9643 33337
rect 12176 33340 13216 33368
rect 7708 33272 8248 33300
rect 7708 33260 7714 33272
rect 8478 33260 8484 33312
rect 8536 33300 8542 33312
rect 9490 33300 9496 33312
rect 8536 33272 9496 33300
rect 8536 33260 8542 33272
rect 9490 33260 9496 33272
rect 9548 33300 9554 33312
rect 12176 33300 12204 33340
rect 13188 33312 13216 33340
rect 9548 33272 12204 33300
rect 9548 33260 9554 33272
rect 12342 33260 12348 33312
rect 12400 33300 12406 33312
rect 12529 33303 12587 33309
rect 12529 33300 12541 33303
rect 12400 33272 12541 33300
rect 12400 33260 12406 33272
rect 12529 33269 12541 33272
rect 12575 33269 12587 33303
rect 12529 33263 12587 33269
rect 13170 33260 13176 33312
rect 13228 33260 13234 33312
rect 13924 33300 13952 33396
rect 14016 33368 14044 33399
rect 14734 33396 14740 33448
rect 14792 33436 14798 33448
rect 14921 33439 14979 33445
rect 14921 33436 14933 33439
rect 14792 33408 14933 33436
rect 14792 33396 14798 33408
rect 14921 33405 14933 33408
rect 14967 33405 14979 33439
rect 14921 33399 14979 33405
rect 15010 33396 15016 33448
rect 15068 33445 15074 33448
rect 15068 33439 15096 33445
rect 15084 33405 15096 33439
rect 15068 33399 15096 33405
rect 15068 33396 15074 33399
rect 14366 33368 14372 33380
rect 14016 33340 14372 33368
rect 14366 33328 14372 33340
rect 14424 33328 14430 33380
rect 18248 33368 18276 33600
rect 18524 33504 18552 33600
rect 18616 33572 18644 33603
rect 19610 33600 19616 33612
rect 19668 33600 19674 33652
rect 19720 33612 20208 33640
rect 19720 33572 19748 33612
rect 20180 33581 20208 33612
rect 18616 33544 19748 33572
rect 20165 33575 20223 33581
rect 20165 33541 20177 33575
rect 20211 33541 20223 33575
rect 20165 33535 20223 33541
rect 18785 33507 18843 33513
rect 18785 33504 18797 33507
rect 18524 33476 18797 33504
rect 18785 33473 18797 33476
rect 18831 33473 18843 33507
rect 18785 33467 18843 33473
rect 18966 33464 18972 33516
rect 19024 33504 19030 33516
rect 19061 33507 19119 33513
rect 19061 33504 19073 33507
rect 19024 33476 19073 33504
rect 19024 33464 19030 33476
rect 19061 33473 19073 33476
rect 19107 33473 19119 33507
rect 19061 33467 19119 33473
rect 19337 33507 19395 33513
rect 19337 33473 19349 33507
rect 19383 33504 19395 33507
rect 19518 33504 19524 33516
rect 19383 33476 19524 33504
rect 19383 33473 19395 33476
rect 19337 33467 19395 33473
rect 19518 33464 19524 33476
rect 19576 33464 19582 33516
rect 19812 33513 19932 33528
rect 19797 33507 19932 33513
rect 19797 33473 19809 33507
rect 19843 33504 19932 33507
rect 20254 33504 20260 33516
rect 19843 33500 20260 33504
rect 19843 33473 19855 33500
rect 19904 33476 20260 33500
rect 19797 33467 19855 33473
rect 20254 33464 20260 33476
rect 20312 33464 20318 33516
rect 19613 33371 19671 33377
rect 19613 33368 19625 33371
rect 18248 33340 19625 33368
rect 19613 33337 19625 33340
rect 19659 33337 19671 33371
rect 19613 33331 19671 33337
rect 16025 33303 16083 33309
rect 16025 33300 16037 33303
rect 13924 33272 16037 33300
rect 16025 33269 16037 33272
rect 16071 33269 16083 33303
rect 16025 33263 16083 33269
rect 18877 33303 18935 33309
rect 18877 33269 18889 33303
rect 18923 33300 18935 33303
rect 19334 33300 19340 33312
rect 18923 33272 19340 33300
rect 18923 33269 18935 33272
rect 18877 33263 18935 33269
rect 19334 33260 19340 33272
rect 19392 33260 19398 33312
rect 20438 33260 20444 33312
rect 20496 33260 20502 33312
rect 1104 33210 20884 33232
rect 1104 33158 3422 33210
rect 3474 33158 3486 33210
rect 3538 33158 3550 33210
rect 3602 33158 3614 33210
rect 3666 33158 3678 33210
rect 3730 33158 8367 33210
rect 8419 33158 8431 33210
rect 8483 33158 8495 33210
rect 8547 33158 8559 33210
rect 8611 33158 8623 33210
rect 8675 33158 13312 33210
rect 13364 33158 13376 33210
rect 13428 33158 13440 33210
rect 13492 33158 13504 33210
rect 13556 33158 13568 33210
rect 13620 33158 18257 33210
rect 18309 33158 18321 33210
rect 18373 33158 18385 33210
rect 18437 33158 18449 33210
rect 18501 33158 18513 33210
rect 18565 33158 20884 33210
rect 1104 33136 20884 33158
rect 1946 33056 1952 33108
rect 2004 33096 2010 33108
rect 3050 33096 3056 33108
rect 2004 33068 3056 33096
rect 2004 33056 2010 33068
rect 3050 33056 3056 33068
rect 3108 33056 3114 33108
rect 4338 33056 4344 33108
rect 4396 33096 4402 33108
rect 4709 33099 4767 33105
rect 4709 33096 4721 33099
rect 4396 33068 4721 33096
rect 4396 33056 4402 33068
rect 4709 33065 4721 33068
rect 4755 33065 4767 33099
rect 4709 33059 4767 33065
rect 4982 33056 4988 33108
rect 5040 33096 5046 33108
rect 5166 33096 5172 33108
rect 5040 33068 5172 33096
rect 5040 33056 5046 33068
rect 5166 33056 5172 33068
rect 5224 33056 5230 33108
rect 7558 33056 7564 33108
rect 7616 33096 7622 33108
rect 7742 33096 7748 33108
rect 7616 33068 7748 33096
rect 7616 33056 7622 33068
rect 7742 33056 7748 33068
rect 7800 33056 7806 33108
rect 8202 33056 8208 33108
rect 8260 33096 8266 33108
rect 8297 33099 8355 33105
rect 8297 33096 8309 33099
rect 8260 33068 8309 33096
rect 8260 33056 8266 33068
rect 8297 33065 8309 33068
rect 8343 33065 8355 33099
rect 9306 33096 9312 33108
rect 8297 33059 8355 33065
rect 8588 33068 9312 33096
rect 8588 33040 8616 33068
rect 9306 33056 9312 33068
rect 9364 33096 9370 33108
rect 10502 33096 10508 33108
rect 9364 33068 10508 33096
rect 9364 33056 9370 33068
rect 10502 33056 10508 33068
rect 10560 33056 10566 33108
rect 12434 33096 12440 33108
rect 11716 33068 12440 33096
rect 6638 32988 6644 33040
rect 6696 33028 6702 33040
rect 7282 33028 7288 33040
rect 6696 33000 7288 33028
rect 6696 32988 6702 33000
rect 7282 32988 7288 33000
rect 7340 32988 7346 33040
rect 8570 32988 8576 33040
rect 8628 32988 8634 33040
rect 11716 33028 11744 33068
rect 12434 33056 12440 33068
rect 12492 33056 12498 33108
rect 12526 33056 12532 33108
rect 12584 33096 12590 33108
rect 12989 33099 13047 33105
rect 12989 33096 13001 33099
rect 12584 33068 13001 33096
rect 12584 33056 12590 33068
rect 12989 33065 13001 33068
rect 13035 33065 13047 33099
rect 12989 33059 13047 33065
rect 15378 33056 15384 33108
rect 15436 33056 15442 33108
rect 15473 33099 15531 33105
rect 15473 33065 15485 33099
rect 15519 33096 15531 33099
rect 16114 33096 16120 33108
rect 15519 33068 16120 33096
rect 15519 33065 15531 33068
rect 15473 33059 15531 33065
rect 16114 33056 16120 33068
rect 16172 33056 16178 33108
rect 17218 33056 17224 33108
rect 17276 33096 17282 33108
rect 18046 33096 18052 33108
rect 17276 33068 18052 33096
rect 17276 33056 17282 33068
rect 18046 33056 18052 33068
rect 18104 33056 18110 33108
rect 18785 33099 18843 33105
rect 18785 33065 18797 33099
rect 18831 33096 18843 33099
rect 19426 33096 19432 33108
rect 18831 33068 19432 33096
rect 18831 33065 18843 33068
rect 18785 33059 18843 33065
rect 9646 33000 11744 33028
rect 1302 32920 1308 32972
rect 1360 32960 1366 32972
rect 1949 32963 2007 32969
rect 1949 32960 1961 32963
rect 1360 32932 1961 32960
rect 1360 32920 1366 32932
rect 1949 32929 1961 32932
rect 1995 32929 2007 32963
rect 1949 32923 2007 32929
rect 750 32852 756 32904
rect 808 32892 814 32904
rect 1397 32895 1455 32901
rect 1397 32892 1409 32895
rect 808 32864 1409 32892
rect 808 32852 814 32864
rect 1397 32861 1409 32864
rect 1443 32861 1455 32895
rect 1397 32855 1455 32861
rect 1486 32784 1492 32836
rect 1544 32824 1550 32836
rect 1673 32827 1731 32833
rect 1673 32824 1685 32827
rect 1544 32796 1685 32824
rect 1544 32784 1550 32796
rect 1673 32793 1685 32796
rect 1719 32793 1731 32827
rect 1964 32824 1992 32923
rect 2958 32920 2964 32972
rect 3016 32960 3022 32972
rect 4798 32960 4804 32972
rect 3016 32932 4804 32960
rect 3016 32920 3022 32932
rect 4798 32920 4804 32932
rect 4856 32920 4862 32972
rect 5442 32920 5448 32972
rect 5500 32920 5506 32972
rect 6914 32920 6920 32972
rect 6972 32960 6978 32972
rect 7098 32960 7104 32972
rect 6972 32932 7104 32960
rect 6972 32920 6978 32932
rect 7098 32920 7104 32932
rect 7156 32960 7162 32972
rect 8846 32960 8852 32972
rect 7156 32932 7328 32960
rect 7156 32920 7162 32932
rect 2222 32892 2228 32904
rect 2183 32864 2228 32892
rect 2222 32852 2228 32864
rect 2280 32852 2286 32904
rect 2866 32852 2872 32904
rect 2924 32892 2930 32904
rect 3789 32895 3847 32901
rect 3789 32892 3801 32895
rect 2924 32864 3801 32892
rect 2924 32852 2930 32864
rect 3789 32861 3801 32864
rect 3835 32861 3847 32895
rect 3789 32855 3847 32861
rect 4062 32852 4068 32904
rect 4120 32852 4126 32904
rect 4893 32895 4951 32901
rect 4893 32861 4905 32895
rect 4939 32861 4951 32895
rect 4893 32855 4951 32861
rect 2682 32824 2688 32836
rect 1964 32796 2688 32824
rect 1673 32787 1731 32793
rect 2682 32784 2688 32796
rect 2740 32784 2746 32836
rect 2884 32796 3280 32824
rect 1210 32716 1216 32768
rect 1268 32756 1274 32768
rect 2884 32756 2912 32796
rect 1268 32728 2912 32756
rect 2961 32759 3019 32765
rect 1268 32716 1274 32728
rect 2961 32725 2973 32759
rect 3007 32756 3019 32759
rect 3050 32756 3056 32768
rect 3007 32728 3056 32756
rect 3007 32725 3019 32728
rect 2961 32719 3019 32725
rect 3050 32716 3056 32728
rect 3108 32716 3114 32768
rect 3252 32756 3280 32796
rect 3326 32784 3332 32836
rect 3384 32824 3390 32836
rect 3878 32824 3884 32836
rect 3384 32796 3884 32824
rect 3384 32784 3390 32796
rect 3878 32784 3884 32796
rect 3936 32784 3942 32836
rect 4908 32824 4936 32855
rect 5534 32852 5540 32904
rect 5592 32852 5598 32904
rect 6454 32852 6460 32904
rect 6512 32892 6518 32904
rect 6638 32892 6644 32904
rect 6512 32864 6644 32892
rect 6512 32852 6518 32864
rect 6638 32852 6644 32864
rect 6696 32852 6702 32904
rect 7006 32852 7012 32904
rect 7064 32852 7070 32904
rect 7300 32901 7328 32932
rect 8128 32932 8852 32960
rect 8128 32904 8156 32932
rect 8846 32920 8852 32932
rect 8904 32960 8910 32972
rect 8941 32963 8999 32969
rect 8941 32960 8953 32963
rect 8904 32932 8953 32960
rect 8904 32920 8910 32932
rect 8941 32929 8953 32932
rect 8987 32929 8999 32963
rect 8941 32923 8999 32929
rect 7285 32895 7343 32901
rect 7285 32861 7297 32895
rect 7331 32861 7343 32895
rect 7527 32895 7585 32901
rect 7527 32892 7539 32895
rect 7285 32855 7343 32861
rect 7374 32864 7539 32892
rect 5445 32827 5503 32833
rect 4908 32796 5302 32824
rect 4908 32756 4936 32796
rect 3252 32728 4936 32756
rect 5166 32716 5172 32768
rect 5224 32716 5230 32768
rect 5274 32756 5302 32796
rect 5445 32793 5457 32827
rect 5491 32824 5503 32827
rect 5626 32824 5632 32836
rect 5491 32796 5632 32824
rect 5491 32793 5503 32796
rect 5445 32787 5503 32793
rect 5626 32784 5632 32796
rect 5684 32784 5690 32836
rect 5905 32827 5963 32833
rect 5905 32793 5917 32827
rect 5951 32824 5963 32827
rect 6362 32824 6368 32836
rect 5951 32796 6368 32824
rect 5951 32793 5963 32796
rect 5905 32787 5963 32793
rect 6362 32784 6368 32796
rect 6420 32784 6426 32836
rect 7024 32824 7052 32852
rect 7374 32824 7402 32864
rect 7527 32861 7539 32864
rect 7573 32861 7585 32895
rect 7527 32855 7585 32861
rect 8110 32852 8116 32904
rect 8168 32852 8174 32904
rect 9183 32895 9241 32901
rect 9183 32892 9195 32895
rect 8956 32864 9195 32892
rect 8956 32836 8984 32864
rect 9183 32861 9195 32864
rect 9229 32861 9241 32895
rect 9646 32892 9674 33000
rect 11790 32988 11796 33040
rect 11848 32988 11854 33040
rect 15396 33028 15424 33056
rect 15841 33031 15899 33037
rect 15841 33028 15853 33031
rect 15396 33000 15853 33028
rect 15841 32997 15853 33000
rect 15887 32997 15899 33031
rect 15841 32991 15899 32997
rect 11698 32920 11704 32972
rect 11756 32960 11762 32972
rect 12069 32963 12127 32969
rect 12069 32960 12081 32963
rect 11756 32932 12081 32960
rect 11756 32920 11762 32932
rect 12069 32929 12081 32932
rect 12115 32929 12127 32963
rect 12069 32923 12127 32929
rect 12342 32920 12348 32972
rect 12400 32920 12406 32972
rect 12526 32920 12532 32972
rect 12584 32960 12590 32972
rect 12584 32932 13952 32960
rect 12584 32920 12590 32932
rect 9183 32855 9241 32861
rect 9322 32864 9674 32892
rect 7024 32796 7402 32824
rect 8938 32784 8944 32836
rect 8996 32784 9002 32836
rect 6273 32759 6331 32765
rect 6273 32756 6285 32759
rect 5274 32728 6285 32756
rect 6273 32725 6285 32728
rect 6319 32725 6331 32759
rect 6273 32719 6331 32725
rect 6457 32759 6515 32765
rect 6457 32725 6469 32759
rect 6503 32756 6515 32759
rect 6730 32756 6736 32768
rect 6503 32728 6736 32756
rect 6503 32725 6515 32728
rect 6457 32719 6515 32725
rect 6730 32716 6736 32728
rect 6788 32716 6794 32768
rect 6914 32716 6920 32768
rect 6972 32756 6978 32768
rect 9322 32756 9350 32864
rect 11146 32852 11152 32904
rect 11204 32852 11210 32904
rect 11333 32895 11391 32901
rect 11333 32861 11345 32895
rect 11379 32861 11391 32895
rect 11333 32855 11391 32861
rect 6972 32728 9350 32756
rect 6972 32716 6978 32728
rect 9858 32716 9864 32768
rect 9916 32756 9922 32768
rect 9953 32759 10011 32765
rect 9953 32756 9965 32759
rect 9916 32728 9965 32756
rect 9916 32716 9922 32728
rect 9953 32725 9965 32728
rect 9999 32725 10011 32759
rect 11348 32756 11376 32855
rect 12158 32852 12164 32904
rect 12216 32901 12222 32904
rect 12216 32895 12244 32901
rect 12232 32861 12244 32895
rect 13924 32892 13952 32932
rect 13998 32920 14004 32972
rect 14056 32960 14062 32972
rect 14093 32963 14151 32969
rect 14093 32960 14105 32963
rect 14056 32932 14105 32960
rect 14056 32920 14062 32932
rect 14093 32929 14105 32932
rect 14139 32929 14151 32963
rect 14093 32923 14151 32929
rect 15580 32932 15884 32960
rect 14335 32895 14393 32901
rect 14335 32892 14347 32895
rect 13924 32864 14347 32892
rect 12216 32855 12244 32861
rect 14335 32861 14347 32864
rect 14381 32892 14393 32895
rect 15580 32892 15608 32932
rect 14381 32864 15608 32892
rect 14381 32861 14393 32864
rect 14335 32855 14393 32861
rect 12216 32852 12222 32855
rect 15654 32852 15660 32904
rect 15712 32852 15718 32904
rect 15749 32895 15807 32901
rect 15749 32861 15761 32895
rect 15795 32861 15807 32895
rect 15749 32855 15807 32861
rect 13814 32784 13820 32836
rect 13872 32824 13878 32836
rect 15764 32824 15792 32855
rect 13872 32796 15792 32824
rect 15856 32824 15884 32932
rect 17402 32852 17408 32904
rect 17460 32892 17466 32904
rect 17773 32895 17831 32901
rect 17773 32892 17785 32895
rect 17460 32864 17785 32892
rect 17460 32852 17466 32864
rect 17773 32861 17785 32864
rect 17819 32861 17831 32895
rect 18015 32895 18073 32901
rect 18015 32892 18027 32895
rect 17773 32855 17831 32861
rect 17880 32864 18027 32892
rect 17880 32824 17908 32864
rect 18015 32861 18027 32864
rect 18061 32892 18073 32895
rect 18598 32892 18604 32904
rect 18061 32864 18604 32892
rect 18061 32861 18073 32864
rect 18015 32855 18073 32861
rect 18598 32852 18604 32864
rect 18656 32852 18662 32904
rect 19260 32901 19288 33068
rect 19426 33056 19432 33068
rect 19484 33056 19490 33108
rect 19702 33056 19708 33108
rect 19760 33056 19766 33108
rect 19720 33028 19748 33056
rect 19536 33000 19748 33028
rect 19889 33031 19947 33037
rect 19536 32969 19564 33000
rect 19889 32997 19901 33031
rect 19935 33028 19947 33031
rect 21266 33028 21272 33040
rect 19935 33000 21272 33028
rect 19935 32997 19947 33000
rect 19889 32991 19947 32997
rect 21266 32988 21272 33000
rect 21324 32988 21330 33040
rect 19521 32963 19579 32969
rect 19521 32929 19533 32963
rect 19567 32929 19579 32963
rect 19521 32923 19579 32929
rect 19245 32895 19303 32901
rect 19245 32861 19257 32895
rect 19291 32861 19303 32895
rect 19245 32855 19303 32861
rect 19334 32852 19340 32904
rect 19392 32852 19398 32904
rect 19705 32895 19763 32901
rect 19705 32861 19717 32895
rect 19751 32861 19763 32895
rect 19705 32855 19763 32861
rect 15856 32796 17908 32824
rect 13872 32784 13878 32796
rect 18782 32784 18788 32836
rect 18840 32824 18846 32836
rect 19610 32824 19616 32836
rect 18840 32796 19616 32824
rect 18840 32784 18846 32796
rect 19610 32784 19616 32796
rect 19668 32784 19674 32836
rect 19720 32824 19748 32855
rect 19978 32852 19984 32904
rect 20036 32852 20042 32904
rect 20070 32852 20076 32904
rect 20128 32892 20134 32904
rect 20165 32895 20223 32901
rect 20165 32892 20177 32895
rect 20128 32864 20177 32892
rect 20128 32852 20134 32864
rect 20165 32861 20177 32864
rect 20211 32861 20223 32895
rect 20165 32855 20223 32861
rect 19996 32824 20024 32852
rect 19720 32796 20024 32824
rect 20530 32784 20536 32836
rect 20588 32784 20594 32836
rect 12434 32756 12440 32768
rect 11348 32728 12440 32756
rect 9953 32719 10011 32725
rect 12434 32716 12440 32728
rect 12492 32756 12498 32768
rect 12986 32756 12992 32768
rect 12492 32728 12992 32756
rect 12492 32716 12498 32728
rect 12986 32716 12992 32728
rect 13044 32716 13050 32768
rect 13722 32716 13728 32768
rect 13780 32756 13786 32768
rect 13998 32756 14004 32768
rect 13780 32728 14004 32756
rect 13780 32716 13786 32728
rect 13998 32716 14004 32728
rect 14056 32756 14062 32768
rect 14550 32756 14556 32768
rect 14056 32728 14556 32756
rect 14056 32716 14062 32728
rect 14550 32716 14556 32728
rect 14608 32716 14614 32768
rect 14826 32716 14832 32768
rect 14884 32756 14890 32768
rect 15105 32759 15163 32765
rect 15105 32756 15117 32759
rect 14884 32728 15117 32756
rect 14884 32716 14890 32728
rect 15105 32725 15117 32728
rect 15151 32725 15163 32759
rect 15105 32719 15163 32725
rect 16206 32716 16212 32768
rect 16264 32756 16270 32768
rect 16850 32756 16856 32768
rect 16264 32728 16856 32756
rect 16264 32716 16270 32728
rect 16850 32716 16856 32728
rect 16908 32716 16914 32768
rect 17310 32716 17316 32768
rect 17368 32756 17374 32768
rect 19426 32756 19432 32768
rect 17368 32728 19432 32756
rect 17368 32716 17374 32728
rect 19426 32716 19432 32728
rect 19484 32716 19490 32768
rect 19521 32759 19579 32765
rect 19521 32725 19533 32759
rect 19567 32756 19579 32759
rect 21634 32756 21640 32768
rect 19567 32728 21640 32756
rect 19567 32725 19579 32728
rect 19521 32719 19579 32725
rect 21634 32716 21640 32728
rect 21692 32716 21698 32768
rect 1104 32666 21043 32688
rect 1104 32614 5894 32666
rect 5946 32614 5958 32666
rect 6010 32614 6022 32666
rect 6074 32614 6086 32666
rect 6138 32614 6150 32666
rect 6202 32614 10839 32666
rect 10891 32614 10903 32666
rect 10955 32614 10967 32666
rect 11019 32614 11031 32666
rect 11083 32614 11095 32666
rect 11147 32614 15784 32666
rect 15836 32614 15848 32666
rect 15900 32614 15912 32666
rect 15964 32614 15976 32666
rect 16028 32614 16040 32666
rect 16092 32614 20729 32666
rect 20781 32614 20793 32666
rect 20845 32614 20857 32666
rect 20909 32614 20921 32666
rect 20973 32614 20985 32666
rect 21037 32614 21043 32666
rect 1104 32592 21043 32614
rect 1302 32512 1308 32564
rect 1360 32552 1366 32564
rect 1360 32524 3740 32552
rect 1360 32512 1366 32524
rect 1854 32444 1860 32496
rect 1912 32484 1918 32496
rect 2225 32487 2283 32493
rect 2225 32484 2237 32487
rect 1912 32456 2237 32484
rect 1912 32444 1918 32456
rect 2225 32453 2237 32456
rect 2271 32453 2283 32487
rect 2225 32447 2283 32453
rect 2501 32487 2559 32493
rect 2501 32453 2513 32487
rect 2547 32453 2559 32487
rect 2501 32447 2559 32453
rect 2593 32487 2651 32493
rect 2593 32453 2605 32487
rect 2639 32484 2651 32487
rect 3050 32484 3056 32496
rect 2639 32456 3056 32484
rect 2639 32453 2651 32456
rect 2593 32447 2651 32453
rect 1394 32376 1400 32428
rect 1452 32376 1458 32428
rect 2516 32416 2544 32447
rect 3050 32444 3056 32456
rect 3108 32444 3114 32496
rect 3326 32444 3332 32496
rect 3384 32444 3390 32496
rect 2774 32416 2780 32428
rect 2516 32388 2780 32416
rect 2774 32376 2780 32388
rect 2832 32376 2838 32428
rect 2958 32376 2964 32428
rect 3016 32376 3022 32428
rect 3712 32425 3740 32524
rect 4062 32512 4068 32564
rect 4120 32552 4126 32564
rect 4120 32524 7586 32552
rect 4120 32512 4126 32524
rect 5442 32444 5448 32496
rect 5500 32484 5506 32496
rect 7466 32484 7472 32496
rect 5500 32456 7472 32484
rect 5500 32444 5506 32456
rect 7466 32444 7472 32456
rect 7524 32444 7530 32496
rect 3697 32419 3755 32425
rect 3697 32385 3709 32419
rect 3743 32385 3755 32419
rect 3697 32379 3755 32385
rect 3878 32376 3884 32428
rect 3936 32416 3942 32428
rect 3973 32419 4031 32425
rect 3973 32416 3985 32419
rect 3936 32388 3985 32416
rect 3936 32376 3942 32388
rect 3973 32385 3985 32388
rect 4019 32416 4031 32419
rect 4338 32416 4344 32428
rect 4019 32388 4344 32416
rect 4019 32385 4031 32388
rect 3973 32379 4031 32385
rect 4338 32376 4344 32388
rect 4396 32376 4402 32428
rect 4707 32419 4765 32425
rect 4707 32385 4719 32419
rect 4753 32416 4765 32419
rect 4798 32416 4804 32428
rect 4753 32388 4804 32416
rect 4753 32385 4765 32388
rect 4707 32379 4765 32385
rect 4798 32376 4804 32388
rect 4856 32376 4862 32428
rect 5534 32376 5540 32428
rect 5592 32416 5598 32428
rect 6914 32416 6920 32428
rect 5592 32388 6920 32416
rect 5592 32376 5598 32388
rect 6914 32376 6920 32388
rect 6972 32376 6978 32428
rect 7098 32376 7104 32428
rect 7156 32376 7162 32428
rect 7374 32416 7380 32428
rect 7335 32388 7380 32416
rect 7374 32376 7380 32388
rect 7432 32376 7438 32428
rect 7558 32416 7586 32524
rect 8018 32512 8024 32564
rect 8076 32552 8082 32564
rect 8113 32555 8171 32561
rect 8113 32552 8125 32555
rect 8076 32524 8125 32552
rect 8076 32512 8082 32524
rect 8113 32521 8125 32524
rect 8159 32521 8171 32555
rect 9306 32552 9312 32564
rect 8113 32515 8171 32521
rect 9232 32524 9312 32552
rect 9232 32425 9260 32524
rect 9306 32512 9312 32524
rect 9364 32512 9370 32564
rect 13814 32512 13820 32564
rect 13872 32512 13878 32564
rect 16025 32555 16083 32561
rect 13970 32524 15790 32552
rect 9398 32444 9404 32496
rect 9456 32484 9462 32496
rect 13970 32484 13998 32524
rect 9456 32456 13998 32484
rect 9456 32444 9462 32456
rect 14274 32444 14280 32496
rect 14332 32444 14338 32496
rect 15762 32484 15790 32524
rect 16025 32521 16037 32555
rect 16071 32521 16083 32555
rect 16025 32515 16083 32521
rect 16040 32484 16068 32515
rect 16666 32512 16672 32564
rect 16724 32512 16730 32564
rect 17126 32512 17132 32564
rect 17184 32512 17190 32564
rect 18785 32555 18843 32561
rect 18785 32521 18797 32555
rect 18831 32552 18843 32555
rect 18831 32524 19104 32552
rect 18831 32521 18843 32524
rect 18785 32515 18843 32521
rect 16684 32484 16712 32512
rect 19076 32484 19104 32524
rect 19334 32512 19340 32564
rect 19392 32552 19398 32564
rect 20349 32555 20407 32561
rect 20349 32552 20361 32555
rect 19392 32524 20361 32552
rect 19392 32512 19398 32524
rect 20349 32521 20361 32524
rect 20395 32521 20407 32555
rect 20349 32515 20407 32521
rect 19518 32484 19524 32496
rect 15762 32456 15884 32484
rect 16040 32456 16344 32484
rect 16684 32456 18920 32484
rect 19076 32456 19524 32484
rect 9217 32419 9275 32425
rect 7558 32388 9168 32416
rect 1673 32351 1731 32357
rect 1673 32317 1685 32351
rect 1719 32317 1731 32351
rect 1673 32311 1731 32317
rect 1688 32280 1716 32311
rect 2406 32308 2412 32360
rect 2464 32308 2470 32360
rect 4433 32351 4491 32357
rect 4433 32317 4445 32351
rect 4479 32317 4491 32351
rect 4433 32311 4491 32317
rect 2130 32280 2136 32292
rect 1688 32252 2136 32280
rect 2130 32240 2136 32252
rect 2188 32240 2194 32292
rect 3510 32240 3516 32292
rect 3568 32240 3574 32292
rect 4448 32212 4476 32311
rect 8938 32308 8944 32360
rect 8996 32308 9002 32360
rect 9140 32348 9168 32388
rect 9217 32385 9229 32419
rect 9263 32385 9275 32419
rect 9674 32416 9680 32428
rect 9217 32379 9275 32385
rect 9324 32388 9680 32416
rect 9324 32348 9352 32388
rect 9674 32376 9680 32388
rect 9732 32376 9738 32428
rect 9767 32419 9825 32425
rect 9767 32385 9779 32419
rect 9813 32416 9825 32419
rect 10778 32416 10784 32428
rect 9813 32388 10784 32416
rect 9813 32385 9825 32388
rect 9767 32379 9825 32385
rect 10778 32376 10784 32388
rect 10836 32416 10842 32428
rect 11606 32416 11612 32428
rect 10836 32388 11612 32416
rect 10836 32376 10842 32388
rect 11606 32376 11612 32388
rect 11664 32376 11670 32428
rect 12619 32419 12677 32425
rect 12619 32385 12631 32419
rect 12665 32416 12677 32419
rect 13170 32416 13176 32428
rect 12665 32388 13176 32416
rect 12665 32385 12677 32388
rect 12619 32379 12677 32385
rect 13170 32376 13176 32388
rect 13228 32376 13234 32428
rect 13814 32376 13820 32428
rect 13872 32416 13878 32428
rect 14001 32420 14059 32425
rect 13924 32419 14059 32420
rect 13924 32416 14013 32419
rect 13872 32392 14013 32416
rect 13872 32388 13952 32392
rect 13998 32388 14013 32392
rect 13872 32376 13878 32388
rect 14001 32385 14013 32388
rect 14047 32385 14059 32419
rect 14292 32416 14320 32444
rect 14292 32388 14394 32416
rect 14001 32379 14059 32385
rect 9140 32320 9352 32348
rect 9493 32351 9551 32357
rect 9493 32317 9505 32351
rect 9539 32317 9551 32351
rect 9493 32311 9551 32317
rect 12345 32351 12403 32357
rect 12345 32317 12357 32351
rect 12391 32317 12403 32351
rect 12345 32311 12403 32317
rect 14093 32351 14151 32357
rect 14093 32317 14105 32351
rect 14139 32317 14151 32351
rect 14093 32311 14151 32317
rect 8956 32280 8984 32308
rect 9508 32280 9536 32311
rect 8956 32252 9536 32280
rect 4890 32212 4896 32224
rect 4448 32184 4896 32212
rect 4890 32172 4896 32184
rect 4948 32212 4954 32224
rect 5350 32212 5356 32224
rect 4948 32184 5356 32212
rect 4948 32172 4954 32184
rect 5350 32172 5356 32184
rect 5408 32172 5414 32224
rect 5442 32172 5448 32224
rect 5500 32172 5506 32224
rect 6546 32172 6552 32224
rect 6604 32212 6610 32224
rect 9309 32215 9367 32221
rect 9309 32212 9321 32215
rect 6604 32184 9321 32212
rect 6604 32172 6610 32184
rect 9309 32181 9321 32184
rect 9355 32181 9367 32215
rect 9309 32175 9367 32181
rect 9490 32172 9496 32224
rect 9548 32212 9554 32224
rect 10226 32212 10232 32224
rect 9548 32184 10232 32212
rect 9548 32172 9554 32184
rect 10226 32172 10232 32184
rect 10284 32172 10290 32224
rect 10502 32172 10508 32224
rect 10560 32172 10566 32224
rect 11054 32172 11060 32224
rect 11112 32212 11118 32224
rect 11974 32212 11980 32224
rect 11112 32184 11980 32212
rect 11112 32172 11118 32184
rect 11974 32172 11980 32184
rect 12032 32172 12038 32224
rect 12158 32172 12164 32224
rect 12216 32212 12222 32224
rect 12360 32212 12388 32311
rect 14108 32280 14136 32311
rect 14274 32308 14280 32360
rect 14332 32308 14338 32360
rect 14366 32348 14394 32388
rect 15286 32376 15292 32428
rect 15344 32376 15350 32428
rect 15013 32351 15071 32357
rect 15013 32348 15025 32351
rect 14366 32320 15025 32348
rect 15013 32317 15025 32320
rect 15059 32317 15071 32351
rect 15013 32311 15071 32317
rect 15102 32308 15108 32360
rect 15160 32357 15166 32360
rect 15160 32351 15188 32357
rect 15176 32317 15188 32351
rect 15856 32348 15884 32456
rect 16206 32376 16212 32428
rect 16264 32376 16270 32428
rect 16316 32425 16344 32456
rect 16301 32419 16359 32425
rect 16301 32385 16313 32419
rect 16347 32385 16359 32419
rect 16301 32379 16359 32385
rect 16574 32376 16580 32428
rect 16632 32416 16638 32428
rect 17420 32425 17448 32456
rect 17313 32419 17371 32425
rect 17313 32416 17325 32419
rect 16632 32388 17325 32416
rect 16632 32376 16638 32388
rect 17313 32385 17325 32388
rect 17359 32385 17371 32419
rect 17313 32379 17371 32385
rect 17405 32419 17463 32425
rect 17405 32385 17417 32419
rect 17451 32385 17463 32419
rect 17661 32419 17719 32425
rect 17661 32416 17673 32419
rect 17405 32379 17463 32385
rect 17512 32388 17673 32416
rect 17512 32348 17540 32388
rect 17661 32385 17673 32388
rect 17707 32416 17719 32419
rect 17954 32416 17960 32428
rect 17707 32388 17960 32416
rect 17707 32385 17719 32388
rect 17661 32379 17719 32385
rect 17954 32376 17960 32388
rect 18012 32376 18018 32428
rect 18230 32376 18236 32428
rect 18288 32416 18294 32428
rect 18892 32425 18920 32456
rect 19518 32444 19524 32456
rect 19576 32444 19582 32496
rect 18877 32419 18935 32425
rect 18288 32388 18828 32416
rect 18288 32376 18294 32388
rect 15856 32320 17540 32348
rect 18800 32348 18828 32388
rect 18877 32385 18889 32419
rect 18923 32385 18935 32419
rect 19133 32419 19191 32425
rect 19133 32416 19145 32419
rect 18877 32379 18935 32385
rect 18984 32388 19145 32416
rect 18984 32348 19012 32388
rect 19133 32385 19145 32388
rect 19179 32416 19191 32419
rect 20533 32419 20591 32425
rect 20533 32416 20545 32419
rect 19179 32388 20545 32416
rect 19179 32385 19191 32388
rect 19133 32379 19191 32385
rect 20533 32385 20545 32388
rect 20579 32385 20591 32419
rect 20533 32379 20591 32385
rect 18800 32320 19012 32348
rect 15160 32311 15188 32317
rect 15160 32308 15166 32311
rect 14041 32252 14136 32280
rect 14041 32224 14069 32252
rect 14550 32240 14556 32292
rect 14608 32240 14614 32292
rect 14737 32283 14795 32289
rect 14737 32249 14749 32283
rect 14783 32280 14795 32283
rect 14826 32280 14832 32292
rect 14783 32252 14832 32280
rect 14783 32249 14795 32252
rect 14737 32243 14795 32249
rect 14826 32240 14832 32252
rect 14884 32240 14890 32292
rect 15746 32240 15752 32292
rect 15804 32280 15810 32292
rect 16574 32280 16580 32292
rect 15804 32252 16580 32280
rect 15804 32240 15810 32252
rect 16574 32240 16580 32252
rect 16632 32240 16638 32292
rect 19886 32240 19892 32292
rect 19944 32280 19950 32292
rect 20257 32283 20315 32289
rect 20257 32280 20269 32283
rect 19944 32252 20269 32280
rect 19944 32240 19950 32252
rect 20257 32249 20269 32252
rect 20303 32249 20315 32283
rect 20257 32243 20315 32249
rect 13078 32212 13084 32224
rect 12216 32184 13084 32212
rect 12216 32172 12222 32184
rect 13078 32172 13084 32184
rect 13136 32172 13142 32224
rect 13170 32172 13176 32224
rect 13228 32212 13234 32224
rect 13357 32215 13415 32221
rect 13357 32212 13369 32215
rect 13228 32184 13369 32212
rect 13228 32172 13234 32184
rect 13357 32181 13369 32184
rect 13403 32181 13415 32215
rect 13357 32175 13415 32181
rect 13998 32172 14004 32224
rect 14056 32184 14069 32224
rect 14568 32212 14596 32240
rect 15838 32212 15844 32224
rect 14568 32184 15844 32212
rect 14056 32172 14062 32184
rect 15838 32172 15844 32184
rect 15896 32172 15902 32224
rect 15930 32172 15936 32224
rect 15988 32172 15994 32224
rect 16390 32172 16396 32224
rect 16448 32172 16454 32224
rect 18598 32172 18604 32224
rect 18656 32212 18662 32224
rect 20162 32212 20168 32224
rect 18656 32184 20168 32212
rect 18656 32172 18662 32184
rect 20162 32172 20168 32184
rect 20220 32172 20226 32224
rect 1104 32122 20884 32144
rect 1104 32070 3422 32122
rect 3474 32070 3486 32122
rect 3538 32070 3550 32122
rect 3602 32070 3614 32122
rect 3666 32070 3678 32122
rect 3730 32070 8367 32122
rect 8419 32070 8431 32122
rect 8483 32070 8495 32122
rect 8547 32070 8559 32122
rect 8611 32070 8623 32122
rect 8675 32070 13312 32122
rect 13364 32070 13376 32122
rect 13428 32070 13440 32122
rect 13492 32070 13504 32122
rect 13556 32070 13568 32122
rect 13620 32070 18257 32122
rect 18309 32070 18321 32122
rect 18373 32070 18385 32122
rect 18437 32070 18449 32122
rect 18501 32070 18513 32122
rect 18565 32070 20884 32122
rect 1104 32048 20884 32070
rect 1854 31968 1860 32020
rect 1912 32008 1918 32020
rect 4062 32008 4068 32020
rect 1912 31980 4068 32008
rect 1912 31968 1918 31980
rect 4062 31968 4068 31980
rect 4120 31968 4126 32020
rect 6457 32011 6515 32017
rect 6457 31977 6469 32011
rect 6503 32008 6515 32011
rect 6914 32008 6920 32020
rect 6503 31980 6920 32008
rect 6503 31977 6515 31980
rect 6457 31971 6515 31977
rect 6914 31968 6920 31980
rect 6972 31968 6978 32020
rect 7024 31980 8248 32008
rect 2590 31900 2596 31952
rect 2648 31940 2654 31952
rect 3237 31943 3295 31949
rect 3237 31940 3249 31943
rect 2648 31912 3249 31940
rect 2648 31900 2654 31912
rect 3237 31909 3249 31912
rect 3283 31909 3295 31943
rect 3237 31903 3295 31909
rect 1118 31832 1124 31884
rect 1176 31872 1182 31884
rect 1489 31875 1547 31881
rect 1489 31872 1501 31875
rect 1176 31844 1501 31872
rect 1176 31832 1182 31844
rect 1489 31841 1501 31844
rect 1535 31841 1547 31875
rect 4080 31872 4108 31968
rect 7024 31940 7052 31980
rect 6288 31912 7052 31940
rect 6288 31884 6316 31912
rect 4080 31844 4936 31872
rect 1489 31835 1547 31841
rect 1504 31668 1532 31835
rect 1747 31777 1805 31783
rect 1747 31743 1759 31777
rect 1793 31774 1805 31777
rect 1793 31743 1806 31774
rect 1854 31764 1860 31816
rect 1912 31804 1918 31816
rect 1912 31776 2268 31804
rect 1912 31764 1918 31776
rect 1747 31737 1806 31743
rect 1778 31736 1806 31737
rect 2130 31736 2136 31748
rect 1778 31708 2136 31736
rect 2130 31696 2136 31708
rect 2188 31696 2194 31748
rect 2240 31736 2268 31776
rect 3050 31764 3056 31816
rect 3108 31764 3114 31816
rect 4614 31764 4620 31816
rect 4672 31764 4678 31816
rect 4908 31804 4936 31844
rect 5442 31832 5448 31884
rect 5500 31832 5506 31884
rect 6270 31832 6276 31884
rect 6328 31832 6334 31884
rect 4908 31776 5304 31804
rect 3421 31739 3479 31745
rect 3421 31736 3433 31739
rect 2240 31708 3433 31736
rect 3421 31705 3433 31708
rect 3467 31705 3479 31739
rect 3421 31699 3479 31705
rect 3602 31696 3608 31748
rect 3660 31696 3666 31748
rect 3786 31696 3792 31748
rect 3844 31696 3850 31748
rect 5166 31696 5172 31748
rect 5224 31696 5230 31748
rect 1670 31668 1676 31680
rect 1504 31640 1676 31668
rect 1670 31628 1676 31640
rect 1728 31668 1734 31680
rect 2222 31668 2228 31680
rect 1728 31640 2228 31668
rect 1728 31628 1734 31640
rect 2222 31628 2228 31640
rect 2280 31628 2286 31680
rect 2501 31671 2559 31677
rect 2501 31637 2513 31671
rect 2547 31668 2559 31671
rect 2682 31668 2688 31680
rect 2547 31640 2688 31668
rect 2547 31637 2559 31640
rect 2501 31631 2559 31637
rect 2682 31628 2688 31640
rect 2740 31628 2746 31680
rect 5276 31668 5304 31776
rect 5350 31764 5356 31816
rect 5408 31804 5414 31816
rect 5537 31807 5595 31813
rect 5537 31804 5549 31807
rect 5408 31776 5549 31804
rect 5408 31764 5414 31776
rect 5537 31773 5549 31776
rect 5583 31773 5595 31807
rect 5905 31807 5963 31813
rect 5905 31804 5917 31807
rect 5537 31767 5595 31773
rect 5644 31776 5917 31804
rect 5442 31696 5448 31748
rect 5500 31696 5506 31748
rect 5644 31668 5672 31776
rect 5905 31773 5917 31776
rect 5951 31773 5963 31807
rect 5905 31767 5963 31773
rect 6917 31807 6975 31813
rect 6917 31773 6929 31807
rect 6963 31804 6975 31807
rect 7098 31804 7104 31816
rect 6963 31776 7104 31804
rect 6963 31773 6975 31776
rect 6917 31767 6975 31773
rect 7098 31764 7104 31776
rect 7156 31764 7162 31816
rect 7191 31807 7249 31813
rect 7191 31773 7203 31807
rect 7237 31804 7249 31807
rect 8220 31804 8248 31980
rect 13078 31968 13084 32020
rect 13136 32008 13142 32020
rect 14182 32008 14188 32020
rect 13136 31980 14188 32008
rect 13136 31968 13142 31980
rect 14182 31968 14188 31980
rect 14240 31968 14246 32020
rect 14274 31968 14280 32020
rect 14332 31968 14338 32020
rect 15194 32008 15200 32020
rect 14844 31980 15200 32008
rect 10781 31943 10839 31949
rect 10781 31909 10793 31943
rect 10827 31909 10839 31943
rect 10781 31903 10839 31909
rect 14292 31940 14320 31968
rect 14458 31940 14464 31952
rect 14292 31912 14464 31940
rect 9306 31832 9312 31884
rect 9364 31872 9370 31884
rect 9769 31875 9827 31881
rect 9769 31872 9781 31875
rect 9364 31844 9781 31872
rect 9364 31832 9370 31844
rect 9769 31841 9781 31844
rect 9815 31841 9827 31875
rect 10796 31872 10824 31903
rect 14292 31881 14320 31912
rect 14458 31900 14464 31912
rect 14516 31900 14522 31952
rect 14734 31900 14740 31952
rect 14792 31900 14798 31952
rect 14277 31875 14335 31881
rect 10796 31844 11178 31872
rect 9769 31835 9827 31841
rect 14277 31841 14289 31875
rect 14323 31841 14335 31875
rect 14844 31872 14872 31980
rect 15194 31968 15200 31980
rect 15252 31968 15258 32020
rect 15654 31968 15660 32020
rect 15712 32008 15718 32020
rect 15933 32011 15991 32017
rect 15933 32008 15945 32011
rect 15712 31980 15945 32008
rect 15712 31968 15718 31980
rect 15933 31977 15945 31980
rect 15979 31977 15991 32011
rect 18325 32011 18383 32017
rect 15933 31971 15991 31977
rect 17604 31980 18276 32008
rect 17604 31949 17632 31980
rect 17589 31943 17647 31949
rect 17589 31909 17601 31943
rect 17635 31909 17647 31943
rect 17589 31903 17647 31909
rect 17954 31900 17960 31952
rect 18012 31900 18018 31952
rect 15013 31875 15071 31881
rect 15013 31872 15025 31875
rect 14844 31844 15025 31872
rect 14277 31835 14335 31841
rect 15013 31841 15025 31844
rect 15059 31841 15071 31875
rect 15013 31835 15071 31841
rect 15102 31832 15108 31884
rect 15160 31881 15166 31884
rect 15160 31875 15188 31881
rect 15176 31841 15188 31875
rect 15160 31835 15188 31841
rect 15289 31875 15347 31881
rect 15289 31841 15301 31875
rect 15335 31872 15347 31875
rect 15470 31872 15476 31884
rect 15335 31844 15476 31872
rect 15335 31841 15347 31844
rect 15289 31835 15347 31841
rect 15160 31832 15166 31835
rect 15470 31832 15476 31844
rect 15528 31832 15534 31884
rect 15838 31832 15844 31884
rect 15896 31872 15902 31884
rect 16025 31875 16083 31881
rect 16025 31872 16037 31875
rect 15896 31844 16037 31872
rect 15896 31832 15902 31844
rect 16025 31841 16037 31844
rect 16071 31841 16083 31875
rect 16025 31835 16083 31841
rect 16850 31832 16856 31884
rect 16908 31832 16914 31884
rect 10011 31807 10069 31813
rect 7237 31776 8156 31804
rect 8220 31776 9904 31804
rect 7237 31773 7249 31776
rect 7191 31767 7249 31773
rect 7392 31748 7420 31776
rect 6270 31696 6276 31748
rect 6328 31696 6334 31748
rect 7374 31696 7380 31748
rect 7432 31696 7438 31748
rect 8128 31736 8156 31776
rect 8846 31736 8852 31748
rect 7760 31708 8064 31736
rect 8128 31708 8852 31736
rect 5276 31640 5672 31668
rect 5810 31628 5816 31680
rect 5868 31668 5874 31680
rect 7760 31668 7788 31708
rect 5868 31640 7788 31668
rect 5868 31628 5874 31640
rect 7834 31628 7840 31680
rect 7892 31668 7898 31680
rect 7929 31671 7987 31677
rect 7929 31668 7941 31671
rect 7892 31640 7941 31668
rect 7892 31628 7898 31640
rect 7929 31637 7941 31640
rect 7975 31637 7987 31671
rect 8036 31668 8064 31708
rect 8846 31696 8852 31708
rect 8904 31696 8910 31748
rect 9398 31696 9404 31748
rect 9456 31736 9462 31748
rect 9876 31736 9904 31776
rect 10011 31773 10023 31807
rect 10057 31804 10069 31807
rect 10134 31804 10140 31816
rect 10057 31776 10140 31804
rect 10057 31773 10069 31776
rect 10011 31767 10069 31773
rect 10134 31764 10140 31776
rect 10192 31764 10198 31816
rect 11606 31764 11612 31816
rect 11664 31764 11670 31816
rect 11701 31807 11759 31813
rect 11701 31773 11713 31807
rect 11747 31804 11759 31807
rect 12526 31804 12532 31816
rect 11747 31776 12532 31804
rect 11747 31773 11759 31776
rect 11701 31767 11759 31773
rect 12526 31764 12532 31776
rect 12584 31764 12590 31816
rect 13906 31764 13912 31816
rect 13964 31804 13970 31816
rect 14093 31807 14151 31813
rect 14093 31804 14105 31807
rect 13964 31776 14105 31804
rect 13964 31764 13970 31776
rect 14093 31773 14105 31776
rect 14139 31773 14151 31807
rect 16868 31804 16896 31832
rect 17773 31807 17831 31813
rect 17773 31804 17785 31807
rect 14093 31767 14151 31773
rect 16283 31777 16341 31783
rect 9456 31708 9904 31736
rect 11256 31708 11928 31736
rect 9456 31696 9462 31708
rect 11256 31668 11284 31708
rect 8036 31640 11284 31668
rect 11333 31671 11391 31677
rect 7929 31631 7987 31637
rect 11333 31637 11345 31671
rect 11379 31668 11391 31671
rect 11790 31668 11796 31680
rect 11379 31640 11796 31668
rect 11379 31637 11391 31640
rect 11333 31631 11391 31637
rect 11790 31628 11796 31640
rect 11848 31628 11854 31680
rect 11900 31668 11928 31708
rect 11974 31696 11980 31748
rect 12032 31736 12038 31748
rect 12069 31739 12127 31745
rect 12069 31736 12081 31739
rect 12032 31708 12081 31736
rect 12032 31696 12038 31708
rect 12069 31705 12081 31708
rect 12115 31705 12127 31739
rect 16283 31743 16295 31777
rect 16329 31774 16341 31777
rect 16868 31776 17785 31804
rect 16329 31743 16344 31774
rect 17773 31773 17785 31776
rect 17819 31773 17831 31807
rect 17972 31804 18000 31900
rect 18248 31872 18276 31980
rect 18325 31977 18337 32011
rect 18371 32008 18383 32011
rect 18598 32008 18604 32020
rect 18371 31980 18604 32008
rect 18371 31977 18383 31980
rect 18325 31971 18383 31977
rect 18598 31968 18604 31980
rect 18656 31968 18662 32020
rect 19702 32008 19708 32020
rect 18708 31980 19708 32008
rect 18248 31844 18552 31872
rect 18524 31813 18552 31844
rect 18708 31813 18736 31980
rect 19702 31968 19708 31980
rect 19760 31968 19766 32020
rect 19058 31832 19064 31884
rect 19116 31872 19122 31884
rect 19245 31875 19303 31881
rect 19245 31872 19257 31875
rect 19116 31844 19257 31872
rect 19116 31832 19122 31844
rect 19245 31841 19257 31844
rect 19291 31841 19303 31875
rect 19245 31835 19303 31841
rect 18233 31807 18291 31813
rect 18233 31804 18245 31807
rect 17972 31776 18245 31804
rect 17773 31767 17831 31773
rect 18233 31773 18245 31776
rect 18279 31773 18291 31807
rect 18233 31767 18291 31773
rect 18509 31807 18567 31813
rect 18509 31773 18521 31807
rect 18555 31773 18567 31807
rect 18509 31767 18567 31773
rect 18693 31807 18751 31813
rect 18693 31773 18705 31807
rect 18739 31773 18751 31807
rect 19519 31807 19577 31813
rect 18693 31767 18751 31773
rect 18800 31776 19472 31804
rect 18800 31748 18828 31776
rect 16283 31737 16344 31743
rect 16316 31736 16344 31737
rect 16850 31736 16856 31748
rect 12069 31699 12127 31705
rect 12360 31708 14320 31736
rect 16316 31708 16856 31736
rect 12360 31668 12388 31708
rect 11900 31640 12388 31668
rect 12434 31628 12440 31680
rect 12492 31628 12498 31680
rect 12621 31671 12679 31677
rect 12621 31637 12633 31671
rect 12667 31668 12679 31671
rect 13078 31668 13084 31680
rect 12667 31640 13084 31668
rect 12667 31637 12679 31640
rect 12621 31631 12679 31637
rect 13078 31628 13084 31640
rect 13136 31628 13142 31680
rect 14292 31668 14320 31708
rect 16850 31696 16856 31708
rect 16908 31696 16914 31748
rect 17586 31696 17592 31748
rect 17644 31736 17650 31748
rect 17862 31736 17868 31748
rect 17644 31708 17868 31736
rect 17644 31696 17650 31708
rect 17862 31696 17868 31708
rect 17920 31696 17926 31748
rect 18414 31696 18420 31748
rect 18472 31736 18478 31748
rect 18472 31708 18727 31736
rect 18472 31696 18478 31708
rect 14918 31668 14924 31680
rect 14292 31640 14924 31668
rect 14918 31628 14924 31640
rect 14976 31668 14982 31680
rect 15746 31668 15752 31680
rect 14976 31640 15752 31668
rect 14976 31628 14982 31640
rect 15746 31628 15752 31640
rect 15804 31628 15810 31680
rect 15930 31628 15936 31680
rect 15988 31668 15994 31680
rect 16298 31668 16304 31680
rect 15988 31640 16304 31668
rect 15988 31628 15994 31640
rect 16298 31628 16304 31640
rect 16356 31628 16362 31680
rect 16574 31628 16580 31680
rect 16632 31668 16638 31680
rect 17037 31671 17095 31677
rect 17037 31668 17049 31671
rect 16632 31640 17049 31668
rect 16632 31628 16638 31640
rect 17037 31637 17049 31640
rect 17083 31637 17095 31671
rect 17037 31631 17095 31637
rect 18049 31671 18107 31677
rect 18049 31637 18061 31671
rect 18095 31668 18107 31671
rect 18598 31668 18604 31680
rect 18095 31640 18604 31668
rect 18095 31637 18107 31640
rect 18049 31631 18107 31637
rect 18598 31628 18604 31640
rect 18656 31628 18662 31680
rect 18699 31668 18727 31708
rect 18782 31696 18788 31748
rect 18840 31696 18846 31748
rect 19058 31696 19064 31748
rect 19116 31736 19122 31748
rect 19334 31736 19340 31748
rect 19116 31708 19340 31736
rect 19116 31696 19122 31708
rect 19334 31696 19340 31708
rect 19392 31696 19398 31748
rect 18969 31671 19027 31677
rect 18969 31668 18981 31671
rect 18699 31640 18981 31668
rect 18969 31637 18981 31640
rect 19015 31637 19027 31671
rect 19444 31668 19472 31776
rect 19519 31773 19531 31807
rect 19565 31804 19577 31807
rect 20622 31804 20628 31816
rect 19565 31776 20628 31804
rect 19565 31773 19577 31776
rect 19519 31767 19577 31773
rect 20622 31764 20628 31776
rect 20680 31764 20686 31816
rect 19610 31696 19616 31748
rect 19668 31736 19674 31748
rect 21910 31736 21916 31748
rect 19668 31708 21916 31736
rect 19668 31696 19674 31708
rect 21910 31696 21916 31708
rect 21968 31696 21974 31748
rect 19978 31668 19984 31680
rect 19444 31640 19984 31668
rect 18969 31631 19027 31637
rect 19978 31628 19984 31640
rect 20036 31628 20042 31680
rect 20254 31628 20260 31680
rect 20312 31628 20318 31680
rect 1104 31578 21043 31600
rect 1104 31526 5894 31578
rect 5946 31526 5958 31578
rect 6010 31526 6022 31578
rect 6074 31526 6086 31578
rect 6138 31526 6150 31578
rect 6202 31526 10839 31578
rect 10891 31526 10903 31578
rect 10955 31526 10967 31578
rect 11019 31526 11031 31578
rect 11083 31526 11095 31578
rect 11147 31526 15784 31578
rect 15836 31526 15848 31578
rect 15900 31526 15912 31578
rect 15964 31526 15976 31578
rect 16028 31526 16040 31578
rect 16092 31526 20729 31578
rect 20781 31526 20793 31578
rect 20845 31526 20857 31578
rect 20909 31526 20921 31578
rect 20973 31526 20985 31578
rect 21037 31526 21043 31578
rect 1104 31504 21043 31526
rect 1578 31424 1584 31476
rect 1636 31424 1642 31476
rect 5092 31436 5304 31464
rect 1596 31328 1624 31424
rect 3050 31396 3056 31408
rect 2056 31368 3056 31396
rect 1673 31331 1731 31337
rect 1673 31328 1685 31331
rect 1596 31300 1685 31328
rect 1673 31297 1685 31300
rect 1719 31328 1731 31331
rect 1946 31328 1952 31340
rect 1719 31300 1952 31328
rect 1719 31297 1731 31300
rect 1673 31291 1731 31297
rect 1946 31288 1952 31300
rect 2004 31288 2010 31340
rect 1397 31263 1455 31269
rect 1397 31229 1409 31263
rect 1443 31260 1455 31263
rect 1578 31260 1584 31272
rect 1443 31232 1584 31260
rect 1443 31229 1455 31232
rect 1397 31223 1455 31229
rect 1578 31220 1584 31232
rect 1636 31220 1642 31272
rect 566 31152 572 31204
rect 624 31192 630 31204
rect 2056 31192 2084 31368
rect 3050 31356 3056 31368
rect 3108 31356 3114 31408
rect 5092 31396 5120 31436
rect 3344 31368 5120 31396
rect 5276 31396 5304 31436
rect 5350 31424 5356 31476
rect 5408 31464 5414 31476
rect 5905 31467 5963 31473
rect 5905 31464 5917 31467
rect 5408 31436 5917 31464
rect 5408 31424 5414 31436
rect 5905 31433 5917 31436
rect 5951 31433 5963 31467
rect 7650 31464 7656 31476
rect 5905 31427 5963 31433
rect 7300 31436 7656 31464
rect 5534 31396 5540 31408
rect 5276 31368 5540 31396
rect 3344 31340 3372 31368
rect 5534 31356 5540 31368
rect 5592 31356 5598 31408
rect 2222 31288 2228 31340
rect 2280 31288 2286 31340
rect 2406 31288 2412 31340
rect 2464 31328 2470 31340
rect 2743 31331 2801 31337
rect 2743 31328 2755 31331
rect 2464 31300 2755 31328
rect 2464 31288 2470 31300
rect 2743 31297 2755 31300
rect 2789 31328 2801 31331
rect 3326 31328 3332 31340
rect 2789 31300 3332 31328
rect 2789 31297 2801 31300
rect 2743 31291 2801 31297
rect 3326 31288 3332 31300
rect 3384 31288 3390 31340
rect 3881 31331 3939 31337
rect 3881 31297 3893 31331
rect 3927 31328 3939 31331
rect 4798 31328 4804 31340
rect 3927 31300 4804 31328
rect 3927 31297 3939 31300
rect 3881 31291 3939 31297
rect 4798 31288 4804 31300
rect 4856 31288 4862 31340
rect 5074 31288 5080 31340
rect 5132 31328 5138 31340
rect 5167 31331 5225 31337
rect 5167 31328 5179 31331
rect 5132 31300 5179 31328
rect 5132 31288 5138 31300
rect 5167 31297 5179 31300
rect 5213 31328 5225 31331
rect 5213 31300 5672 31328
rect 5213 31297 5225 31300
rect 5167 31291 5225 31297
rect 2240 31260 2268 31288
rect 2501 31263 2559 31269
rect 2501 31260 2513 31263
rect 2240 31232 2513 31260
rect 2501 31229 2513 31232
rect 2547 31229 2559 31263
rect 2501 31223 2559 31229
rect 4157 31263 4215 31269
rect 4157 31229 4169 31263
rect 4203 31229 4215 31263
rect 4157 31223 4215 31229
rect 4172 31192 4200 31223
rect 4890 31220 4896 31272
rect 4948 31220 4954 31272
rect 5644 31260 5672 31300
rect 7098 31288 7104 31340
rect 7156 31328 7162 31340
rect 7300 31337 7328 31436
rect 7650 31424 7656 31436
rect 7708 31424 7714 31476
rect 10410 31424 10416 31476
rect 10468 31464 10474 31476
rect 10965 31467 11023 31473
rect 10965 31464 10977 31467
rect 10468 31436 10977 31464
rect 10468 31424 10474 31436
rect 10965 31433 10977 31436
rect 11011 31433 11023 31467
rect 10965 31427 11023 31433
rect 11790 31424 11796 31476
rect 11848 31464 11854 31476
rect 12066 31464 12072 31476
rect 11848 31436 12072 31464
rect 11848 31424 11854 31436
rect 12066 31424 12072 31436
rect 12124 31424 12130 31476
rect 12158 31424 12164 31476
rect 12216 31424 12222 31476
rect 12526 31424 12532 31476
rect 12584 31424 12590 31476
rect 13814 31424 13820 31476
rect 13872 31464 13878 31476
rect 14737 31467 14795 31473
rect 14737 31464 14749 31467
rect 13872 31436 14749 31464
rect 13872 31424 13878 31436
rect 14737 31433 14749 31436
rect 14783 31433 14795 31467
rect 15470 31464 15476 31476
rect 14737 31427 14795 31433
rect 14844 31436 15476 31464
rect 12176 31396 12204 31424
rect 11532 31368 12204 31396
rect 7543 31361 7601 31367
rect 7285 31331 7343 31337
rect 7285 31328 7297 31331
rect 7156 31300 7297 31328
rect 7156 31288 7162 31300
rect 7285 31297 7297 31300
rect 7331 31297 7343 31331
rect 7543 31327 7555 31361
rect 7589 31358 7601 31361
rect 7589 31328 7604 31358
rect 8202 31328 8208 31340
rect 7589 31327 8208 31328
rect 7543 31321 8208 31327
rect 7576 31300 8208 31321
rect 7285 31291 7343 31297
rect 8202 31288 8208 31300
rect 8260 31288 8266 31340
rect 9140 31300 9444 31328
rect 9140 31269 9168 31300
rect 9416 31272 9444 31300
rect 10042 31288 10048 31340
rect 10100 31288 10106 31340
rect 10318 31288 10324 31340
rect 10376 31288 10382 31340
rect 11146 31288 11152 31340
rect 11204 31328 11210 31340
rect 11532 31337 11560 31368
rect 12342 31356 12348 31408
rect 12400 31396 12406 31408
rect 12434 31396 12440 31408
rect 12400 31368 12440 31396
rect 12400 31356 12406 31368
rect 12434 31356 12440 31368
rect 12492 31396 12498 31408
rect 14844 31396 14872 31436
rect 15470 31424 15476 31436
rect 15528 31464 15534 31476
rect 15841 31467 15899 31473
rect 15841 31464 15853 31467
rect 15528 31436 15853 31464
rect 15528 31424 15534 31436
rect 15841 31433 15853 31436
rect 15887 31433 15899 31467
rect 15841 31427 15899 31433
rect 16209 31467 16267 31473
rect 16209 31433 16221 31467
rect 16255 31433 16267 31467
rect 16209 31427 16267 31433
rect 18141 31467 18199 31473
rect 18141 31433 18153 31467
rect 18187 31433 18199 31467
rect 18141 31427 18199 31433
rect 18601 31467 18659 31473
rect 18601 31433 18613 31467
rect 18647 31464 18659 31467
rect 18782 31464 18788 31476
rect 18647 31436 18788 31464
rect 18647 31433 18659 31436
rect 18601 31427 18659 31433
rect 12492 31368 13124 31396
rect 12492 31356 12498 31368
rect 11517 31331 11575 31337
rect 11517 31328 11529 31331
rect 11204 31300 11529 31328
rect 11204 31288 11210 31300
rect 11517 31297 11529 31300
rect 11563 31297 11575 31331
rect 11790 31328 11796 31340
rect 11751 31300 11796 31328
rect 11517 31291 11575 31297
rect 11790 31288 11796 31300
rect 11848 31288 11854 31340
rect 12526 31288 12532 31340
rect 12584 31328 12590 31340
rect 12710 31328 12716 31340
rect 12584 31300 12716 31328
rect 12584 31288 12590 31300
rect 12710 31288 12716 31300
rect 12768 31288 12774 31340
rect 13096 31337 13124 31368
rect 14752 31368 14872 31396
rect 13081 31331 13139 31337
rect 13081 31297 13093 31331
rect 13127 31297 13139 31331
rect 13081 31291 13139 31297
rect 9125 31263 9183 31269
rect 5644 31232 7144 31260
rect 7116 31204 7144 31232
rect 9125 31229 9137 31263
rect 9171 31229 9183 31263
rect 9125 31223 9183 31229
rect 9309 31263 9367 31269
rect 9309 31229 9321 31263
rect 9355 31229 9367 31263
rect 9309 31223 9367 31229
rect 624 31164 2084 31192
rect 3160 31164 4200 31192
rect 624 31152 630 31164
rect 2406 31084 2412 31136
rect 2464 31124 2470 31136
rect 3160 31124 3188 31164
rect 7098 31152 7104 31204
rect 7156 31152 7162 31204
rect 2464 31096 3188 31124
rect 2464 31084 2470 31096
rect 3234 31084 3240 31136
rect 3292 31124 3298 31136
rect 3513 31127 3571 31133
rect 3513 31124 3525 31127
rect 3292 31096 3525 31124
rect 3292 31084 3298 31096
rect 3513 31093 3525 31096
rect 3559 31093 3571 31127
rect 3513 31087 3571 31093
rect 3602 31084 3608 31136
rect 3660 31124 3666 31136
rect 5350 31124 5356 31136
rect 3660 31096 5356 31124
rect 3660 31084 3666 31096
rect 5350 31084 5356 31096
rect 5408 31084 5414 31136
rect 7190 31084 7196 31136
rect 7248 31124 7254 31136
rect 7374 31124 7380 31136
rect 7248 31096 7380 31124
rect 7248 31084 7254 31096
rect 7374 31084 7380 31096
rect 7432 31084 7438 31136
rect 8202 31084 8208 31136
rect 8260 31124 8266 31136
rect 8297 31127 8355 31133
rect 8297 31124 8309 31127
rect 8260 31096 8309 31124
rect 8260 31084 8266 31096
rect 8297 31093 8309 31096
rect 8343 31093 8355 31127
rect 9324 31124 9352 31223
rect 9398 31220 9404 31272
rect 9456 31220 9462 31272
rect 10183 31263 10241 31269
rect 10183 31260 10195 31263
rect 9876 31232 10195 31260
rect 9876 31204 9904 31232
rect 10183 31229 10195 31232
rect 10229 31229 10241 31263
rect 10183 31223 10241 31229
rect 12897 31263 12955 31269
rect 12897 31229 12909 31263
rect 12943 31260 12955 31263
rect 12986 31260 12992 31272
rect 12943 31232 12992 31260
rect 12943 31229 12955 31232
rect 12897 31223 12955 31229
rect 12986 31220 12992 31232
rect 13044 31220 13050 31272
rect 13170 31220 13176 31272
rect 13228 31260 13234 31272
rect 13541 31263 13599 31269
rect 13541 31260 13553 31263
rect 13228 31232 13553 31260
rect 13228 31220 13234 31232
rect 13541 31229 13553 31232
rect 13587 31229 13599 31263
rect 13541 31223 13599 31229
rect 13814 31220 13820 31272
rect 13872 31220 13878 31272
rect 13998 31269 14004 31272
rect 13955 31263 14004 31269
rect 13955 31229 13967 31263
rect 14001 31229 14004 31263
rect 13955 31223 14004 31229
rect 13998 31220 14004 31223
rect 14056 31220 14062 31272
rect 14093 31263 14151 31269
rect 14093 31229 14105 31263
rect 14139 31260 14151 31263
rect 14752 31260 14780 31368
rect 14918 31356 14924 31408
rect 14976 31356 14982 31408
rect 16224 31396 16252 31427
rect 18156 31396 18184 31427
rect 18782 31424 18788 31436
rect 18840 31424 18846 31476
rect 19076 31436 20208 31464
rect 19076 31396 19104 31436
rect 20180 31405 20208 31436
rect 20254 31424 20260 31476
rect 20312 31424 20318 31476
rect 20622 31424 20628 31476
rect 20680 31464 20686 31476
rect 21818 31464 21824 31476
rect 20680 31436 21824 31464
rect 20680 31424 20686 31436
rect 21818 31424 21824 31436
rect 21876 31424 21882 31476
rect 16224 31368 16896 31396
rect 18156 31368 19104 31396
rect 20165 31399 20223 31405
rect 14936 31328 14964 31356
rect 15071 31331 15129 31337
rect 15071 31328 15083 31331
rect 14936 31300 15083 31328
rect 15071 31297 15083 31300
rect 15117 31297 15129 31331
rect 15071 31291 15129 31297
rect 16298 31288 16304 31340
rect 16356 31328 16362 31340
rect 16868 31337 16896 31368
rect 20165 31365 20177 31399
rect 20211 31365 20223 31399
rect 20165 31359 20223 31365
rect 16393 31331 16451 31337
rect 16393 31328 16405 31331
rect 16356 31300 16405 31328
rect 16356 31288 16362 31300
rect 16393 31297 16405 31300
rect 16439 31297 16451 31331
rect 16669 31331 16727 31337
rect 16669 31328 16681 31331
rect 16393 31291 16451 31297
rect 16592 31300 16681 31328
rect 16592 31272 16620 31300
rect 16669 31297 16681 31300
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 16853 31331 16911 31337
rect 16853 31297 16865 31331
rect 16899 31297 16911 31331
rect 16853 31291 16911 31297
rect 17586 31288 17592 31340
rect 17644 31328 17650 31340
rect 18049 31331 18107 31337
rect 18049 31328 18061 31331
rect 17644 31300 18061 31328
rect 17644 31288 17650 31300
rect 18049 31297 18061 31300
rect 18095 31297 18107 31331
rect 18049 31291 18107 31297
rect 18325 31331 18383 31337
rect 18325 31297 18337 31331
rect 18371 31297 18383 31331
rect 18325 31291 18383 31297
rect 18417 31331 18475 31337
rect 18417 31297 18429 31331
rect 18463 31297 18475 31331
rect 18417 31291 18475 31297
rect 14139 31232 14780 31260
rect 14829 31263 14887 31269
rect 14139 31229 14151 31232
rect 14093 31223 14151 31229
rect 14829 31229 14841 31263
rect 14875 31229 14887 31263
rect 14829 31223 14887 31229
rect 9766 31152 9772 31204
rect 9824 31152 9830 31204
rect 9858 31152 9864 31204
rect 9916 31152 9922 31204
rect 14844 31192 14872 31223
rect 16574 31220 16580 31272
rect 16632 31220 16638 31272
rect 18230 31220 18236 31272
rect 18288 31260 18294 31272
rect 18340 31260 18368 31291
rect 18288 31232 18368 31260
rect 18432 31260 18460 31291
rect 18506 31288 18512 31340
rect 18564 31328 18570 31340
rect 18601 31331 18659 31337
rect 18601 31328 18613 31331
rect 18564 31300 18613 31328
rect 18564 31288 18570 31300
rect 18601 31297 18613 31300
rect 18647 31297 18659 31331
rect 18601 31291 18659 31297
rect 18690 31288 18696 31340
rect 18748 31288 18754 31340
rect 19153 31337 19211 31343
rect 19153 31332 19165 31337
rect 19076 31328 19165 31332
rect 18984 31304 19165 31328
rect 18984 31300 19104 31304
rect 19153 31303 19165 31304
rect 19199 31303 19211 31337
rect 18782 31260 18788 31272
rect 18432 31232 18788 31260
rect 18288 31220 18294 31232
rect 18782 31220 18788 31232
rect 18840 31220 18846 31272
rect 18984 31252 19012 31300
rect 19153 31297 19211 31303
rect 19242 31288 19248 31340
rect 19300 31332 19306 31340
rect 19300 31304 19380 31332
rect 19300 31288 19306 31304
rect 19058 31252 19064 31272
rect 18984 31224 19064 31252
rect 19058 31220 19064 31224
rect 19116 31220 19122 31272
rect 14752 31164 14872 31192
rect 10502 31124 10508 31136
rect 9324 31096 10508 31124
rect 8297 31087 8355 31093
rect 10502 31084 10508 31096
rect 10560 31084 10566 31136
rect 14182 31084 14188 31136
rect 14240 31124 14246 31136
rect 14752 31124 14780 31164
rect 15562 31152 15568 31204
rect 15620 31192 15626 31204
rect 16942 31192 16948 31204
rect 15620 31164 16948 31192
rect 15620 31152 15626 31164
rect 16942 31152 16948 31164
rect 17000 31152 17006 31204
rect 19242 31152 19248 31204
rect 19300 31152 19306 31204
rect 19352 31192 19380 31304
rect 19610 31288 19616 31340
rect 19668 31288 19674 31340
rect 19705 31331 19763 31337
rect 19705 31297 19717 31331
rect 19751 31328 19763 31331
rect 19794 31328 19800 31340
rect 19751 31300 19800 31328
rect 19751 31297 19763 31300
rect 19705 31291 19763 31297
rect 19794 31288 19800 31300
rect 19852 31328 19858 31340
rect 20272 31328 20300 31424
rect 19852 31300 20300 31328
rect 19852 31288 19858 31300
rect 19978 31220 19984 31272
rect 20036 31220 20042 31272
rect 19797 31195 19855 31201
rect 19797 31192 19809 31195
rect 19352 31164 19809 31192
rect 19797 31161 19809 31164
rect 19843 31161 19855 31195
rect 21726 31192 21732 31204
rect 19797 31155 19855 31161
rect 19904 31164 21732 31192
rect 14240 31096 14780 31124
rect 14240 31084 14246 31096
rect 16758 31084 16764 31136
rect 16816 31084 16822 31136
rect 17865 31127 17923 31133
rect 17865 31093 17877 31127
rect 17911 31124 17923 31127
rect 18414 31124 18420 31136
rect 17911 31096 18420 31124
rect 17911 31093 17923 31096
rect 17865 31087 17923 31093
rect 18414 31084 18420 31096
rect 18472 31084 18478 31136
rect 18690 31084 18696 31136
rect 18748 31124 18754 31136
rect 18785 31127 18843 31133
rect 18785 31124 18797 31127
rect 18748 31096 18797 31124
rect 18748 31084 18754 31096
rect 18785 31093 18797 31096
rect 18831 31093 18843 31127
rect 18785 31087 18843 31093
rect 19429 31127 19487 31133
rect 19429 31093 19441 31127
rect 19475 31124 19487 31127
rect 19702 31124 19708 31136
rect 19475 31096 19708 31124
rect 19475 31093 19487 31096
rect 19429 31087 19487 31093
rect 19702 31084 19708 31096
rect 19760 31084 19766 31136
rect 19904 31133 19932 31164
rect 21726 31152 21732 31164
rect 21784 31152 21790 31204
rect 19889 31127 19947 31133
rect 19889 31093 19901 31127
rect 19935 31093 19947 31127
rect 19889 31087 19947 31093
rect 20438 31084 20444 31136
rect 20496 31084 20502 31136
rect 1104 31034 20884 31056
rect 1104 30982 3422 31034
rect 3474 30982 3486 31034
rect 3538 30982 3550 31034
rect 3602 30982 3614 31034
rect 3666 30982 3678 31034
rect 3730 30982 8367 31034
rect 8419 30982 8431 31034
rect 8483 30982 8495 31034
rect 8547 30982 8559 31034
rect 8611 30982 8623 31034
rect 8675 30982 13312 31034
rect 13364 30982 13376 31034
rect 13428 30982 13440 31034
rect 13492 30982 13504 31034
rect 13556 30982 13568 31034
rect 13620 30982 18257 31034
rect 18309 30982 18321 31034
rect 18373 30982 18385 31034
rect 18437 30982 18449 31034
rect 18501 30982 18513 31034
rect 18565 30982 20884 31034
rect 1104 30960 20884 30982
rect 658 30880 664 30932
rect 716 30920 722 30932
rect 3421 30923 3479 30929
rect 3421 30920 3433 30923
rect 716 30892 3433 30920
rect 716 30880 722 30892
rect 3421 30889 3433 30892
rect 3467 30889 3479 30923
rect 3421 30883 3479 30889
rect 4154 30880 4160 30932
rect 4212 30920 4218 30932
rect 5626 30920 5632 30932
rect 4212 30892 5632 30920
rect 4212 30880 4218 30892
rect 5626 30880 5632 30892
rect 5684 30880 5690 30932
rect 8202 30880 8208 30932
rect 8260 30880 8266 30932
rect 9398 30880 9404 30932
rect 9456 30920 9462 30932
rect 10318 30920 10324 30932
rect 9456 30892 10324 30920
rect 9456 30880 9462 30892
rect 10318 30880 10324 30892
rect 10376 30880 10382 30932
rect 11146 30920 11152 30932
rect 10796 30892 11152 30920
rect 1854 30852 1860 30864
rect 1596 30824 1860 30852
rect 1596 30725 1624 30824
rect 1854 30812 1860 30824
rect 1912 30812 1918 30864
rect 2225 30787 2283 30793
rect 2225 30784 2237 30787
rect 1688 30756 2237 30784
rect 1581 30719 1639 30725
rect 1581 30685 1593 30719
rect 1627 30685 1639 30719
rect 1581 30679 1639 30685
rect 1302 30608 1308 30660
rect 1360 30648 1366 30660
rect 1688 30648 1716 30756
rect 2225 30753 2237 30756
rect 2271 30753 2283 30787
rect 2225 30747 2283 30753
rect 2590 30744 2596 30796
rect 2648 30793 2654 30796
rect 2648 30787 2676 30793
rect 2664 30753 2676 30787
rect 2648 30747 2676 30753
rect 2648 30744 2654 30747
rect 7834 30744 7840 30796
rect 7892 30744 7898 30796
rect 1765 30719 1823 30725
rect 1765 30685 1777 30719
rect 1811 30685 1823 30719
rect 1765 30679 1823 30685
rect 1360 30620 1716 30648
rect 1360 30608 1366 30620
rect 1780 30580 1808 30679
rect 2498 30676 2504 30728
rect 2556 30676 2562 30728
rect 2774 30676 2780 30728
rect 2832 30676 2838 30728
rect 3418 30676 3424 30728
rect 3476 30716 3482 30728
rect 3789 30719 3847 30725
rect 3789 30716 3801 30719
rect 3476 30688 3801 30716
rect 3476 30676 3482 30688
rect 3789 30685 3801 30688
rect 3835 30685 3847 30719
rect 3789 30679 3847 30685
rect 4065 30719 4123 30725
rect 4065 30685 4077 30719
rect 4111 30685 4123 30719
rect 4065 30679 4123 30685
rect 4339 30719 4397 30725
rect 4339 30685 4351 30719
rect 4385 30716 4397 30719
rect 5074 30716 5080 30728
rect 4385 30688 5080 30716
rect 4385 30685 4397 30688
rect 4339 30679 4397 30685
rect 4080 30648 4108 30679
rect 5074 30676 5080 30688
rect 5132 30676 5138 30728
rect 5350 30676 5356 30728
rect 5408 30716 5414 30728
rect 6730 30716 6736 30728
rect 5408 30688 6736 30716
rect 5408 30676 5414 30688
rect 6730 30676 6736 30688
rect 6788 30716 6794 30728
rect 7285 30719 7343 30725
rect 7285 30716 7297 30719
rect 6788 30688 7297 30716
rect 6788 30676 6794 30688
rect 7285 30685 7297 30688
rect 7331 30685 7343 30719
rect 7285 30679 7343 30685
rect 7377 30719 7435 30725
rect 7377 30685 7389 30719
rect 7423 30716 7435 30719
rect 8220 30716 8248 30880
rect 8297 30855 8355 30861
rect 8297 30821 8309 30855
rect 8343 30852 8355 30855
rect 8846 30852 8852 30864
rect 8343 30824 8852 30852
rect 8343 30821 8355 30824
rect 8297 30815 8355 30821
rect 8846 30812 8852 30824
rect 8904 30812 8910 30864
rect 9306 30784 9312 30796
rect 8312 30756 9312 30784
rect 8312 30728 8340 30756
rect 9306 30744 9312 30756
rect 9364 30784 9370 30796
rect 10796 30793 10824 30892
rect 11146 30880 11152 30892
rect 11204 30880 11210 30932
rect 11238 30880 11244 30932
rect 11296 30920 11302 30932
rect 11296 30892 12434 30920
rect 11296 30880 11302 30892
rect 9401 30787 9459 30793
rect 9401 30784 9413 30787
rect 9364 30756 9413 30784
rect 9364 30744 9370 30756
rect 9401 30753 9413 30756
rect 9447 30753 9459 30787
rect 9401 30747 9459 30753
rect 10781 30787 10839 30793
rect 10781 30753 10793 30787
rect 10827 30753 10839 30787
rect 10781 30747 10839 30753
rect 7423 30688 8248 30716
rect 7423 30685 7435 30688
rect 7377 30679 7435 30685
rect 8294 30676 8300 30728
rect 8352 30676 8358 30728
rect 8478 30676 8484 30728
rect 8536 30676 8542 30728
rect 8665 30719 8723 30725
rect 8665 30685 8677 30719
rect 8711 30685 8723 30719
rect 8665 30679 8723 30685
rect 7009 30651 7067 30657
rect 7009 30648 7021 30651
rect 3804 30620 4108 30648
rect 5000 30620 7021 30648
rect 3804 30592 3832 30620
rect 3602 30580 3608 30592
rect 1780 30552 3608 30580
rect 3602 30540 3608 30552
rect 3660 30540 3666 30592
rect 3786 30540 3792 30592
rect 3844 30540 3850 30592
rect 3973 30583 4031 30589
rect 3973 30549 3985 30583
rect 4019 30580 4031 30583
rect 5000 30580 5028 30620
rect 7009 30617 7021 30620
rect 7055 30617 7067 30651
rect 7009 30611 7067 30617
rect 4019 30552 5028 30580
rect 5077 30583 5135 30589
rect 4019 30549 4031 30552
rect 3973 30543 4031 30549
rect 5077 30549 5089 30583
rect 5123 30580 5135 30583
rect 5166 30580 5172 30592
rect 5123 30552 5172 30580
rect 5123 30549 5135 30552
rect 5077 30543 5135 30549
rect 5166 30540 5172 30552
rect 5224 30540 5230 30592
rect 7024 30580 7052 30611
rect 7190 30608 7196 30660
rect 7248 30648 7254 30660
rect 7745 30651 7803 30657
rect 7745 30648 7757 30651
rect 7248 30620 7757 30648
rect 7248 30608 7254 30620
rect 7745 30617 7757 30620
rect 7791 30648 7803 30651
rect 7834 30648 7840 30660
rect 7791 30620 7840 30648
rect 7791 30617 7803 30620
rect 7745 30611 7803 30617
rect 7834 30608 7840 30620
rect 7892 30608 7898 30660
rect 7926 30608 7932 30660
rect 7984 30648 7990 30660
rect 8680 30648 8708 30679
rect 7984 30620 8708 30648
rect 9416 30648 9444 30747
rect 9675 30719 9733 30725
rect 9675 30685 9687 30719
rect 9721 30716 9733 30719
rect 9766 30716 9772 30728
rect 9721 30688 9772 30716
rect 9721 30685 9733 30688
rect 9675 30679 9733 30685
rect 9766 30676 9772 30688
rect 9824 30676 9830 30728
rect 10042 30676 10048 30728
rect 10100 30716 10106 30728
rect 10594 30716 10600 30728
rect 10100 30688 10600 30716
rect 10100 30676 10106 30688
rect 10594 30676 10600 30688
rect 10652 30676 10658 30728
rect 10796 30648 10824 30747
rect 11882 30744 11888 30796
rect 11940 30784 11946 30796
rect 12250 30784 12256 30796
rect 11940 30756 12256 30784
rect 11940 30744 11946 30756
rect 12250 30744 12256 30756
rect 12308 30744 12314 30796
rect 12406 30784 12434 30892
rect 13354 30880 13360 30932
rect 13412 30920 13418 30932
rect 13722 30920 13728 30932
rect 13412 30892 13728 30920
rect 13412 30880 13418 30892
rect 13722 30880 13728 30892
rect 13780 30880 13786 30932
rect 13814 30880 13820 30932
rect 13872 30920 13878 30932
rect 15010 30920 15016 30932
rect 13872 30892 15016 30920
rect 13872 30880 13878 30892
rect 15010 30880 15016 30892
rect 15068 30880 15074 30932
rect 15933 30923 15991 30929
rect 15933 30889 15945 30923
rect 15979 30920 15991 30923
rect 16206 30920 16212 30932
rect 15979 30892 16212 30920
rect 15979 30889 15991 30892
rect 15933 30883 15991 30889
rect 16206 30880 16212 30892
rect 16264 30880 16270 30932
rect 16758 30880 16764 30932
rect 16816 30880 16822 30932
rect 17972 30892 19196 30920
rect 14734 30812 14740 30864
rect 14792 30812 14798 30864
rect 12406 30756 15148 30784
rect 15120 30728 15148 30756
rect 15286 30744 15292 30796
rect 15344 30744 15350 30796
rect 15654 30744 15660 30796
rect 15712 30784 15718 30796
rect 16114 30784 16120 30796
rect 15712 30756 16120 30784
rect 15712 30744 15718 30756
rect 16114 30744 16120 30756
rect 16172 30744 16178 30796
rect 16209 30787 16267 30793
rect 16209 30753 16221 30787
rect 16255 30784 16267 30787
rect 16574 30784 16580 30796
rect 16255 30756 16580 30784
rect 16255 30753 16267 30756
rect 16209 30747 16267 30753
rect 16574 30744 16580 30756
rect 16632 30744 16638 30796
rect 11054 30725 11060 30728
rect 11023 30719 11060 30725
rect 11023 30685 11035 30719
rect 11023 30679 11060 30685
rect 11054 30676 11060 30679
rect 11112 30676 11118 30728
rect 12342 30676 12348 30728
rect 12400 30676 12406 30728
rect 14093 30719 14151 30725
rect 14093 30685 14105 30719
rect 14139 30716 14151 30719
rect 14182 30716 14188 30728
rect 14139 30688 14188 30716
rect 14139 30685 14151 30688
rect 14093 30679 14151 30685
rect 14182 30676 14188 30688
rect 14240 30676 14246 30728
rect 14277 30719 14335 30725
rect 14277 30685 14289 30719
rect 14323 30685 14335 30719
rect 14277 30679 14335 30685
rect 9416 30620 10824 30648
rect 7984 30608 7990 30620
rect 11882 30608 11888 30660
rect 11940 30648 11946 30660
rect 12360 30648 12388 30676
rect 14292 30648 14320 30679
rect 15010 30676 15016 30728
rect 15068 30676 15074 30728
rect 15102 30676 15108 30728
rect 15160 30725 15166 30728
rect 15160 30719 15188 30725
rect 15176 30685 15188 30719
rect 15160 30679 15188 30685
rect 15160 30676 15166 30679
rect 16390 30676 16396 30728
rect 16448 30676 16454 30728
rect 16776 30716 16804 30880
rect 17972 30861 18000 30892
rect 17957 30855 18015 30861
rect 17957 30821 17969 30855
rect 18003 30821 18015 30855
rect 17957 30815 18015 30821
rect 18601 30855 18659 30861
rect 18601 30821 18613 30855
rect 18647 30821 18659 30855
rect 18601 30815 18659 30821
rect 18877 30855 18935 30861
rect 18877 30821 18889 30855
rect 18923 30852 18935 30855
rect 19168 30852 19196 30892
rect 19242 30880 19248 30932
rect 19300 30880 19306 30932
rect 18923 30824 19104 30852
rect 19168 30824 19334 30852
rect 18923 30821 18935 30824
rect 18877 30815 18935 30821
rect 17678 30744 17684 30796
rect 17736 30784 17742 30796
rect 18616 30784 18644 30815
rect 19076 30784 19104 30824
rect 17736 30756 18000 30784
rect 18616 30756 19012 30784
rect 19076 30756 19176 30784
rect 17736 30744 17742 30756
rect 17972 30728 18000 30756
rect 16853 30719 16911 30725
rect 16853 30716 16865 30719
rect 16776 30688 16865 30716
rect 16853 30685 16865 30688
rect 16899 30685 16911 30719
rect 17221 30719 17279 30725
rect 17221 30716 17233 30719
rect 16853 30679 16911 30685
rect 16960 30688 17233 30716
rect 11940 30620 14320 30648
rect 11940 30608 11946 30620
rect 16298 30608 16304 30660
rect 16356 30648 16362 30660
rect 16960 30648 16988 30688
rect 17221 30685 17233 30688
rect 17267 30685 17279 30719
rect 17221 30679 17279 30685
rect 17770 30676 17776 30728
rect 17828 30676 17834 30728
rect 17954 30676 17960 30728
rect 18012 30676 18018 30728
rect 18138 30676 18144 30728
rect 18196 30676 18202 30728
rect 18782 30676 18788 30728
rect 18840 30676 18846 30728
rect 18984 30718 19012 30756
rect 19061 30719 19119 30725
rect 19061 30718 19073 30719
rect 18984 30690 19073 30718
rect 19061 30685 19073 30690
rect 19107 30685 19119 30719
rect 19061 30679 19119 30685
rect 16356 30620 16988 30648
rect 17129 30651 17187 30657
rect 16356 30608 16362 30620
rect 17129 30617 17141 30651
rect 17175 30648 17187 30651
rect 18230 30648 18236 30660
rect 17175 30620 18236 30648
rect 17175 30617 17187 30620
rect 17129 30611 17187 30617
rect 18230 30608 18236 30620
rect 18288 30608 18294 30660
rect 19148 30648 19176 30756
rect 19306 30716 19334 30824
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 19306 30688 19441 30716
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19518 30676 19524 30728
rect 19576 30716 19582 30728
rect 19705 30719 19763 30725
rect 19705 30716 19717 30719
rect 19576 30688 19717 30716
rect 19576 30676 19582 30688
rect 19705 30685 19717 30688
rect 19751 30685 19763 30719
rect 19705 30679 19763 30685
rect 19794 30676 19800 30728
rect 19852 30716 19858 30728
rect 19981 30719 20039 30725
rect 19981 30716 19993 30719
rect 19852 30688 19993 30716
rect 19852 30676 19858 30688
rect 19981 30685 19993 30688
rect 20027 30685 20039 30719
rect 19981 30679 20039 30685
rect 20165 30651 20223 30657
rect 20165 30648 20177 30651
rect 19148 30620 20177 30648
rect 20165 30617 20177 30620
rect 20211 30617 20223 30651
rect 20165 30611 20223 30617
rect 20533 30651 20591 30657
rect 20533 30617 20545 30651
rect 20579 30648 20591 30651
rect 21266 30648 21272 30660
rect 20579 30620 21272 30648
rect 20579 30617 20591 30620
rect 20533 30611 20591 30617
rect 21266 30608 21272 30620
rect 21324 30608 21330 30660
rect 7558 30580 7564 30592
rect 7024 30552 7564 30580
rect 7558 30540 7564 30552
rect 7616 30540 7622 30592
rect 8110 30540 8116 30592
rect 8168 30540 8174 30592
rect 8570 30540 8576 30592
rect 8628 30540 8634 30592
rect 10410 30540 10416 30592
rect 10468 30540 10474 30592
rect 10594 30540 10600 30592
rect 10652 30580 10658 30592
rect 11330 30580 11336 30592
rect 10652 30552 11336 30580
rect 10652 30540 10658 30552
rect 11330 30540 11336 30552
rect 11388 30540 11394 30592
rect 11790 30540 11796 30592
rect 11848 30540 11854 30592
rect 13078 30540 13084 30592
rect 13136 30580 13142 30592
rect 16758 30580 16764 30592
rect 13136 30552 16764 30580
rect 13136 30540 13142 30552
rect 16758 30540 16764 30552
rect 16816 30540 16822 30592
rect 17310 30540 17316 30592
rect 17368 30540 17374 30592
rect 17586 30540 17592 30592
rect 17644 30540 17650 30592
rect 17678 30540 17684 30592
rect 17736 30580 17742 30592
rect 19521 30583 19579 30589
rect 19521 30580 19533 30583
rect 17736 30552 19533 30580
rect 17736 30540 17742 30552
rect 19521 30549 19533 30552
rect 19567 30549 19579 30583
rect 19521 30543 19579 30549
rect 19797 30583 19855 30589
rect 19797 30549 19809 30583
rect 19843 30580 19855 30583
rect 19978 30580 19984 30592
rect 19843 30552 19984 30580
rect 19843 30549 19855 30552
rect 19797 30543 19855 30549
rect 19978 30540 19984 30552
rect 20036 30540 20042 30592
rect 1104 30490 21043 30512
rect 1104 30438 5894 30490
rect 5946 30438 5958 30490
rect 6010 30438 6022 30490
rect 6074 30438 6086 30490
rect 6138 30438 6150 30490
rect 6202 30438 10839 30490
rect 10891 30438 10903 30490
rect 10955 30438 10967 30490
rect 11019 30438 11031 30490
rect 11083 30438 11095 30490
rect 11147 30438 15784 30490
rect 15836 30438 15848 30490
rect 15900 30438 15912 30490
rect 15964 30438 15976 30490
rect 16028 30438 16040 30490
rect 16092 30438 20729 30490
rect 20781 30438 20793 30490
rect 20845 30438 20857 30490
rect 20909 30438 20921 30490
rect 20973 30438 20985 30490
rect 21037 30438 21043 30490
rect 1104 30416 21043 30438
rect 2240 30348 4016 30376
rect 1394 30268 1400 30320
rect 1452 30308 1458 30320
rect 1489 30311 1547 30317
rect 1489 30308 1501 30311
rect 1452 30280 1501 30308
rect 1452 30268 1458 30280
rect 1489 30277 1501 30280
rect 1535 30277 1547 30311
rect 1489 30271 1547 30277
rect 750 30200 756 30252
rect 808 30240 814 30252
rect 2240 30240 2268 30348
rect 3988 30308 4016 30348
rect 4798 30336 4804 30388
rect 4856 30376 4862 30388
rect 7190 30376 7196 30388
rect 4856 30348 5672 30376
rect 4856 30336 4862 30348
rect 5644 30308 5672 30348
rect 6840 30348 7196 30376
rect 5813 30311 5871 30317
rect 5813 30308 5825 30311
rect 3988 30280 4108 30308
rect 5644 30280 5825 30308
rect 808 30212 2268 30240
rect 808 30200 814 30212
rect 2972 30200 2978 30252
rect 3030 30249 3036 30252
rect 3030 30203 3037 30249
rect 3030 30200 3036 30203
rect 3970 30200 3976 30252
rect 4028 30200 4034 30252
rect 4080 30240 4108 30280
rect 5813 30277 5825 30280
rect 5859 30277 5871 30311
rect 5813 30271 5871 30277
rect 4338 30240 4344 30252
rect 4080 30212 4344 30240
rect 4338 30200 4344 30212
rect 4396 30200 4402 30252
rect 5166 30200 5172 30252
rect 5224 30200 5230 30252
rect 2041 30175 2099 30181
rect 2041 30172 2053 30175
rect 1412 30144 2053 30172
rect 1412 30048 1440 30144
rect 2041 30141 2053 30144
rect 2087 30141 2099 30175
rect 2041 30135 2099 30141
rect 2056 30104 2084 30135
rect 2222 30132 2228 30184
rect 2280 30132 2286 30184
rect 3078 30175 3136 30181
rect 3078 30172 3090 30175
rect 2792 30144 3090 30172
rect 2590 30104 2596 30116
rect 2056 30076 2596 30104
rect 2590 30064 2596 30076
rect 2648 30064 2654 30116
rect 2682 30064 2688 30116
rect 2740 30064 2746 30116
rect 1394 29996 1400 30048
rect 1452 29996 1458 30048
rect 1762 29996 1768 30048
rect 1820 29996 1826 30048
rect 2792 30036 2820 30144
rect 3078 30141 3090 30144
rect 3124 30141 3136 30175
rect 3216 30172 3222 30184
rect 3274 30181 3280 30184
rect 3181 30144 3222 30172
rect 3078 30135 3136 30141
rect 3216 30132 3222 30144
rect 3274 30135 3281 30181
rect 3274 30132 3280 30135
rect 4154 30132 4160 30184
rect 4212 30132 4218 30184
rect 4893 30175 4951 30181
rect 4893 30172 4905 30175
rect 4724 30144 4905 30172
rect 3881 30107 3939 30113
rect 3881 30073 3893 30107
rect 3927 30104 3939 30107
rect 3970 30104 3976 30116
rect 3927 30076 3976 30104
rect 3927 30073 3939 30076
rect 3881 30067 3939 30073
rect 3970 30064 3976 30076
rect 4028 30064 4034 30116
rect 4614 30064 4620 30116
rect 4672 30064 4678 30116
rect 4724 30036 4752 30144
rect 4893 30141 4905 30144
rect 4939 30141 4951 30175
rect 4893 30135 4951 30141
rect 5031 30175 5089 30181
rect 5031 30141 5043 30175
rect 5077 30172 5089 30175
rect 5350 30172 5356 30184
rect 5077 30144 5356 30172
rect 5077 30141 5089 30144
rect 5031 30135 5089 30141
rect 5350 30132 5356 30144
rect 5408 30132 5414 30184
rect 6840 30172 6868 30348
rect 7190 30336 7196 30348
rect 7248 30376 7254 30388
rect 7650 30376 7656 30388
rect 7248 30348 7656 30376
rect 7248 30336 7254 30348
rect 7650 30336 7656 30348
rect 7708 30376 7714 30388
rect 8294 30376 8300 30388
rect 7708 30348 8300 30376
rect 7708 30336 7714 30348
rect 8294 30336 8300 30348
rect 8352 30336 8358 30388
rect 9582 30336 9588 30388
rect 9640 30336 9646 30388
rect 11606 30336 11612 30388
rect 11664 30376 11670 30388
rect 11974 30376 11980 30388
rect 11664 30348 11980 30376
rect 11664 30336 11670 30348
rect 11974 30336 11980 30348
rect 12032 30376 12038 30388
rect 13998 30376 14004 30388
rect 12032 30348 14004 30376
rect 12032 30336 12038 30348
rect 13998 30336 14004 30348
rect 14056 30336 14062 30388
rect 14642 30336 14648 30388
rect 14700 30336 14706 30388
rect 16298 30336 16304 30388
rect 16356 30336 16362 30388
rect 17126 30336 17132 30388
rect 17184 30376 17190 30388
rect 17402 30376 17408 30388
rect 17184 30348 17408 30376
rect 17184 30336 17190 30348
rect 17402 30336 17408 30348
rect 17460 30336 17466 30388
rect 17586 30336 17592 30388
rect 17644 30336 17650 30388
rect 17770 30336 17776 30388
rect 17828 30376 17834 30388
rect 18049 30379 18107 30385
rect 18049 30376 18061 30379
rect 17828 30348 18061 30376
rect 17828 30336 17834 30348
rect 18049 30345 18061 30348
rect 18095 30345 18107 30379
rect 18049 30339 18107 30345
rect 18782 30336 18788 30388
rect 18840 30376 18846 30388
rect 19061 30379 19119 30385
rect 19061 30376 19073 30379
rect 18840 30348 19073 30376
rect 18840 30336 18846 30348
rect 19061 30345 19073 30348
rect 19107 30345 19119 30379
rect 19061 30339 19119 30345
rect 19429 30379 19487 30385
rect 19429 30345 19441 30379
rect 19475 30376 19487 30379
rect 19610 30376 19616 30388
rect 19475 30348 19616 30376
rect 19475 30345 19487 30348
rect 19429 30339 19487 30345
rect 19610 30336 19616 30348
rect 19668 30336 19674 30388
rect 19702 30336 19708 30388
rect 19760 30376 19766 30388
rect 20162 30376 20168 30388
rect 19760 30348 20168 30376
rect 19760 30336 19766 30348
rect 20162 30336 20168 30348
rect 20220 30336 20226 30388
rect 6914 30268 6920 30320
rect 6972 30268 6978 30320
rect 7006 30268 7012 30320
rect 7064 30308 7070 30320
rect 8573 30311 8631 30317
rect 7064 30280 8432 30308
rect 7064 30268 7070 30280
rect 6932 30240 6960 30268
rect 7159 30243 7217 30249
rect 7159 30240 7171 30243
rect 6932 30212 7171 30240
rect 7159 30209 7171 30212
rect 7205 30240 7217 30243
rect 7558 30240 7564 30252
rect 7205 30212 7564 30240
rect 7205 30209 7217 30212
rect 7159 30203 7217 30209
rect 7558 30200 7564 30212
rect 7616 30200 7622 30252
rect 8297 30243 8355 30249
rect 8297 30209 8309 30243
rect 8343 30209 8355 30243
rect 8404 30240 8432 30280
rect 8573 30277 8585 30311
rect 8619 30308 8631 30311
rect 9122 30308 9128 30320
rect 8619 30280 9128 30308
rect 8619 30277 8631 30280
rect 8573 30271 8631 30277
rect 9122 30268 9128 30280
rect 9180 30268 9186 30320
rect 8662 30240 8668 30252
rect 8404 30212 8668 30240
rect 8297 30203 8355 30209
rect 6917 30175 6975 30181
rect 6917 30172 6929 30175
rect 6840 30144 6929 30172
rect 6917 30141 6929 30144
rect 6963 30141 6975 30175
rect 6917 30135 6975 30141
rect 8312 30172 8340 30203
rect 8662 30200 8668 30212
rect 8720 30200 8726 30252
rect 8939 30243 8997 30249
rect 8939 30209 8951 30243
rect 8985 30240 8997 30243
rect 9600 30240 9628 30336
rect 14660 30308 14688 30336
rect 14829 30311 14887 30317
rect 14660 30280 14780 30308
rect 8985 30212 9628 30240
rect 8985 30209 8997 30212
rect 8939 30203 8997 30209
rect 11974 30200 11980 30252
rect 12032 30240 12038 30252
rect 13354 30240 13360 30252
rect 12032 30212 13360 30240
rect 12032 30200 12038 30212
rect 13354 30200 13360 30212
rect 13412 30200 13418 30252
rect 13998 30200 14004 30252
rect 14056 30249 14062 30252
rect 14056 30243 14084 30249
rect 14072 30209 14084 30243
rect 14752 30240 14780 30280
rect 14829 30277 14841 30311
rect 14875 30308 14887 30311
rect 16914 30311 16972 30317
rect 16914 30308 16926 30311
rect 14875 30280 16926 30308
rect 14875 30277 14887 30280
rect 14829 30271 14887 30277
rect 14921 30243 14979 30249
rect 14921 30240 14933 30243
rect 14752 30212 14933 30240
rect 14056 30203 14084 30209
rect 14921 30209 14933 30212
rect 14967 30209 14979 30243
rect 14921 30203 14979 30209
rect 14056 30200 14062 30203
rect 15102 30200 15108 30252
rect 15160 30240 15166 30252
rect 16500 30249 16528 30280
rect 16914 30277 16926 30280
rect 16960 30277 16972 30311
rect 17604 30308 17632 30336
rect 17604 30280 18736 30308
rect 16914 30271 16972 30277
rect 15195 30243 15253 30249
rect 15195 30240 15207 30243
rect 15160 30212 15207 30240
rect 15160 30200 15166 30212
rect 15195 30209 15207 30212
rect 15241 30240 15253 30243
rect 16485 30243 16543 30249
rect 15241 30212 16068 30240
rect 15241 30209 15253 30212
rect 15195 30203 15253 30209
rect 8478 30172 8484 30184
rect 8312 30144 8484 30172
rect 6638 30064 6644 30116
rect 6696 30064 6702 30116
rect 7929 30107 7987 30113
rect 7929 30073 7941 30107
rect 7975 30104 7987 30107
rect 8312 30104 8340 30144
rect 8478 30132 8484 30144
rect 8536 30132 8542 30184
rect 8570 30132 8576 30184
rect 8628 30132 8634 30184
rect 12989 30175 13047 30181
rect 12989 30141 13001 30175
rect 13035 30172 13047 30175
rect 13078 30172 13084 30184
rect 13035 30144 13084 30172
rect 13035 30141 13047 30144
rect 12989 30135 13047 30141
rect 13078 30132 13084 30144
rect 13136 30132 13142 30184
rect 13170 30132 13176 30184
rect 13228 30132 13234 30184
rect 13906 30132 13912 30184
rect 13964 30132 13970 30184
rect 14185 30175 14243 30181
rect 14185 30141 14197 30175
rect 14231 30172 14243 30175
rect 14231 30144 14872 30172
rect 14231 30141 14243 30144
rect 14185 30135 14243 30141
rect 7975 30076 8340 30104
rect 8389 30107 8447 30113
rect 7975 30073 7987 30076
rect 7929 30067 7987 30073
rect 8389 30073 8401 30107
rect 8435 30104 8447 30107
rect 8435 30076 8800 30104
rect 8435 30073 8447 30076
rect 8389 30067 8447 30073
rect 5074 30036 5080 30048
rect 2792 30008 5080 30036
rect 5074 29996 5080 30008
rect 5132 29996 5138 30048
rect 5258 29996 5264 30048
rect 5316 30036 5322 30048
rect 6546 30036 6552 30048
rect 5316 30008 6552 30036
rect 5316 29996 5322 30008
rect 6546 29996 6552 30008
rect 6604 29996 6610 30048
rect 6656 30036 6684 30064
rect 8772 30048 8800 30076
rect 13630 30064 13636 30116
rect 13688 30064 13694 30116
rect 14844 30104 14872 30144
rect 14844 30076 14964 30104
rect 8110 30036 8116 30048
rect 6656 30008 8116 30036
rect 8110 29996 8116 30008
rect 8168 29996 8174 30048
rect 8754 29996 8760 30048
rect 8812 29996 8818 30048
rect 9674 29996 9680 30048
rect 9732 29996 9738 30048
rect 10042 29996 10048 30048
rect 10100 30036 10106 30048
rect 10870 30036 10876 30048
rect 10100 30008 10876 30036
rect 10100 29996 10106 30008
rect 10870 29996 10876 30008
rect 10928 30036 10934 30048
rect 14826 30036 14832 30048
rect 10928 30008 14832 30036
rect 10928 29996 10934 30008
rect 14826 29996 14832 30008
rect 14884 29996 14890 30048
rect 14936 30036 14964 30076
rect 15933 30039 15991 30045
rect 15933 30036 15945 30039
rect 14936 30008 15945 30036
rect 15933 30005 15945 30008
rect 15979 30005 15991 30039
rect 16040 30036 16068 30212
rect 16485 30209 16497 30243
rect 16531 30209 16543 30243
rect 16485 30203 16543 30209
rect 16666 30200 16672 30252
rect 16724 30200 16730 30252
rect 17310 30200 17316 30252
rect 17368 30240 17374 30252
rect 17368 30212 17816 30240
rect 17368 30200 17374 30212
rect 17788 30172 17816 30212
rect 18138 30200 18144 30252
rect 18196 30240 18202 30252
rect 18708 30249 18736 30280
rect 18791 30280 19288 30308
rect 18509 30243 18567 30249
rect 18509 30240 18521 30243
rect 18196 30212 18521 30240
rect 18196 30200 18202 30212
rect 18509 30209 18521 30212
rect 18555 30209 18567 30243
rect 18509 30203 18567 30209
rect 18693 30243 18751 30249
rect 18693 30209 18705 30243
rect 18739 30209 18751 30243
rect 18693 30203 18751 30209
rect 18233 30175 18291 30181
rect 18233 30172 18245 30175
rect 17788 30144 18245 30172
rect 18233 30141 18245 30144
rect 18279 30141 18291 30175
rect 18233 30135 18291 30141
rect 18417 30175 18475 30181
rect 18417 30141 18429 30175
rect 18463 30172 18475 30175
rect 18601 30175 18659 30181
rect 18601 30172 18613 30175
rect 18463 30144 18613 30172
rect 18463 30141 18475 30144
rect 18417 30135 18475 30141
rect 18601 30141 18613 30144
rect 18647 30141 18659 30175
rect 18791 30172 18819 30280
rect 18966 30200 18972 30252
rect 19024 30200 19030 30252
rect 19260 30249 19288 30280
rect 19534 30280 20208 30308
rect 19245 30243 19303 30249
rect 19245 30209 19257 30243
rect 19291 30209 19303 30243
rect 19245 30203 19303 30209
rect 19534 30172 19562 30280
rect 19610 30200 19616 30252
rect 19668 30200 19674 30252
rect 19702 30200 19708 30252
rect 19760 30200 19766 30252
rect 20180 30249 20208 30280
rect 19889 30243 19947 30249
rect 19889 30209 19901 30243
rect 19935 30209 19947 30243
rect 19889 30203 19947 30209
rect 20165 30243 20223 30249
rect 20165 30209 20177 30243
rect 20211 30209 20223 30243
rect 20165 30203 20223 30209
rect 18601 30135 18659 30141
rect 18699 30144 18819 30172
rect 18892 30144 19562 30172
rect 18699 30104 18727 30144
rect 17604 30076 18727 30104
rect 18785 30107 18843 30113
rect 17604 30036 17632 30076
rect 18785 30073 18797 30107
rect 18831 30104 18843 30107
rect 18892 30104 18920 30144
rect 19904 30104 19932 30203
rect 20070 30132 20076 30184
rect 20128 30172 20134 30184
rect 20128 30144 20392 30172
rect 20128 30132 20134 30144
rect 18831 30076 18920 30104
rect 19306 30076 19932 30104
rect 18831 30073 18843 30076
rect 18785 30067 18843 30073
rect 16040 30008 17632 30036
rect 18325 30039 18383 30045
rect 15933 29999 15991 30005
rect 18325 30005 18337 30039
rect 18371 30036 18383 30039
rect 18690 30036 18696 30048
rect 18371 30008 18696 30036
rect 18371 30005 18383 30008
rect 18325 29999 18383 30005
rect 18690 29996 18696 30008
rect 18748 29996 18754 30048
rect 18874 29996 18880 30048
rect 18932 30036 18938 30048
rect 19306 30036 19334 30076
rect 20364 30048 20392 30144
rect 18932 30008 19334 30036
rect 19797 30039 19855 30045
rect 18932 29996 18938 30008
rect 19797 30005 19809 30039
rect 19843 30036 19855 30039
rect 20070 30036 20076 30048
rect 19843 30008 20076 30036
rect 19843 30005 19855 30008
rect 19797 29999 19855 30005
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 20346 29996 20352 30048
rect 20404 29996 20410 30048
rect 20438 29996 20444 30048
rect 20496 29996 20502 30048
rect 1104 29946 20884 29968
rect 1104 29894 3422 29946
rect 3474 29894 3486 29946
rect 3538 29894 3550 29946
rect 3602 29894 3614 29946
rect 3666 29894 3678 29946
rect 3730 29894 8367 29946
rect 8419 29894 8431 29946
rect 8483 29894 8495 29946
rect 8547 29894 8559 29946
rect 8611 29894 8623 29946
rect 8675 29894 13312 29946
rect 13364 29894 13376 29946
rect 13428 29894 13440 29946
rect 13492 29894 13504 29946
rect 13556 29894 13568 29946
rect 13620 29894 18257 29946
rect 18309 29894 18321 29946
rect 18373 29894 18385 29946
rect 18437 29894 18449 29946
rect 18501 29894 18513 29946
rect 18565 29894 20884 29946
rect 1104 29872 20884 29894
rect 2222 29792 2228 29844
rect 2280 29832 2286 29844
rect 2280 29804 2544 29832
rect 2280 29792 2286 29804
rect 1026 29724 1032 29776
rect 1084 29764 1090 29776
rect 1084 29736 1716 29764
rect 1084 29724 1090 29736
rect 1688 29708 1716 29736
rect 1486 29656 1492 29708
rect 1544 29656 1550 29708
rect 1670 29656 1676 29708
rect 1728 29696 1734 29708
rect 1857 29699 1915 29705
rect 1857 29696 1869 29699
rect 1728 29668 1869 29696
rect 1728 29656 1734 29668
rect 1857 29665 1869 29668
rect 1903 29665 1915 29699
rect 2516 29696 2544 29804
rect 2682 29792 2688 29844
rect 2740 29832 2746 29844
rect 2869 29835 2927 29841
rect 2869 29832 2881 29835
rect 2740 29804 2881 29832
rect 2740 29792 2746 29804
rect 2869 29801 2881 29804
rect 2915 29801 2927 29835
rect 4522 29832 4528 29844
rect 2869 29795 2927 29801
rect 2976 29804 4528 29832
rect 2976 29764 3004 29804
rect 4522 29792 4528 29804
rect 4580 29792 4586 29844
rect 4614 29792 4620 29844
rect 4672 29832 4678 29844
rect 4801 29835 4859 29841
rect 4801 29832 4813 29835
rect 4672 29804 4813 29832
rect 4672 29792 4678 29804
rect 4801 29801 4813 29804
rect 4847 29801 4859 29835
rect 6914 29832 6920 29844
rect 4801 29795 4859 29801
rect 6012 29804 6920 29832
rect 6012 29773 6040 29804
rect 6914 29792 6920 29804
rect 6972 29832 6978 29844
rect 8297 29835 8355 29841
rect 8297 29832 8309 29835
rect 6972 29804 8309 29832
rect 6972 29792 6978 29804
rect 8297 29801 8309 29804
rect 8343 29801 8355 29835
rect 13449 29835 13507 29841
rect 8297 29795 8355 29801
rect 12544 29804 13124 29832
rect 2746 29736 3004 29764
rect 5997 29767 6055 29773
rect 2746 29696 2774 29736
rect 5997 29733 6009 29767
rect 6043 29733 6055 29767
rect 12544 29764 12572 29804
rect 5997 29727 6055 29733
rect 12452 29736 12572 29764
rect 13096 29764 13124 29804
rect 13449 29801 13461 29835
rect 13495 29832 13507 29835
rect 13630 29832 13636 29844
rect 13495 29804 13636 29832
rect 13495 29801 13507 29804
rect 13449 29795 13507 29801
rect 13630 29792 13636 29804
rect 13688 29792 13694 29844
rect 14550 29832 14556 29844
rect 13740 29804 14556 29832
rect 13538 29764 13544 29776
rect 13096 29736 13544 29764
rect 10416 29708 10468 29714
rect 3786 29696 3792 29708
rect 2516 29668 2774 29696
rect 3160 29668 3792 29696
rect 1857 29659 1915 29665
rect 1504 29628 1532 29656
rect 3160 29640 3188 29668
rect 3786 29656 3792 29668
rect 3844 29656 3850 29708
rect 6390 29699 6448 29705
rect 6390 29696 6402 29699
rect 4722 29668 6402 29696
rect 2131 29631 2189 29637
rect 1504 29600 1808 29628
rect 1780 29598 1808 29600
rect 1486 29520 1492 29572
rect 1544 29520 1550 29572
rect 1670 29520 1676 29572
rect 1728 29520 1734 29572
rect 1780 29570 1990 29598
rect 2131 29597 2143 29631
rect 2177 29628 2189 29631
rect 2774 29628 2780 29640
rect 2177 29600 2780 29628
rect 2177 29597 2189 29600
rect 2131 29591 2189 29597
rect 2774 29588 2780 29600
rect 2832 29588 2838 29640
rect 3142 29588 3148 29640
rect 3200 29588 3206 29640
rect 3326 29588 3332 29640
rect 3384 29588 3390 29640
rect 3970 29628 3976 29640
rect 3436 29600 3976 29628
rect 1962 29560 1990 29570
rect 2222 29560 2228 29572
rect 1962 29532 2228 29560
rect 2222 29520 2228 29532
rect 2280 29520 2286 29572
rect 3234 29520 3240 29572
rect 3292 29560 3298 29572
rect 3436 29560 3464 29600
rect 3970 29588 3976 29600
rect 4028 29628 4034 29640
rect 4063 29631 4121 29637
rect 4063 29628 4075 29631
rect 4028 29600 4075 29628
rect 4028 29588 4034 29600
rect 4063 29597 4075 29600
rect 4109 29597 4121 29631
rect 4722 29628 4750 29668
rect 6390 29665 6402 29668
rect 6436 29665 6448 29699
rect 6390 29659 6448 29665
rect 6549 29699 6607 29705
rect 6549 29665 6561 29699
rect 6595 29696 6607 29699
rect 6730 29696 6736 29708
rect 6595 29668 6736 29696
rect 6595 29665 6607 29668
rect 6549 29659 6607 29665
rect 6730 29656 6736 29668
rect 6788 29656 6794 29708
rect 7190 29656 7196 29708
rect 7248 29696 7254 29708
rect 7285 29699 7343 29705
rect 7285 29696 7297 29699
rect 7248 29668 7297 29696
rect 7248 29656 7254 29668
rect 7285 29665 7297 29668
rect 7331 29665 7343 29699
rect 7285 29659 7343 29665
rect 4063 29591 4121 29597
rect 4448 29600 4750 29628
rect 3292 29532 3464 29560
rect 3513 29563 3571 29569
rect 3292 29520 3298 29532
rect 3513 29529 3525 29563
rect 3559 29560 3571 29563
rect 4154 29560 4160 29572
rect 3559 29532 4160 29560
rect 3559 29529 3571 29532
rect 3513 29523 3571 29529
rect 4154 29520 4160 29532
rect 4212 29560 4218 29572
rect 4448 29560 4476 29600
rect 5258 29588 5264 29640
rect 5316 29628 5322 29640
rect 5353 29631 5411 29637
rect 5353 29628 5365 29631
rect 5316 29600 5365 29628
rect 5316 29588 5322 29600
rect 5353 29597 5365 29600
rect 5399 29597 5411 29631
rect 5353 29591 5411 29597
rect 5537 29631 5595 29637
rect 5537 29597 5549 29631
rect 5583 29597 5595 29631
rect 5537 29591 5595 29597
rect 4212 29532 4476 29560
rect 4212 29520 4218 29532
rect 4522 29520 4528 29572
rect 4580 29560 4586 29572
rect 5166 29560 5172 29572
rect 4580 29532 5172 29560
rect 4580 29520 4586 29532
rect 5166 29520 5172 29532
rect 5224 29560 5230 29572
rect 5552 29560 5580 29591
rect 6270 29588 6276 29640
rect 6328 29588 6334 29640
rect 5224 29532 5580 29560
rect 5224 29520 5230 29532
rect 1026 29452 1032 29504
rect 1084 29492 1090 29504
rect 2590 29492 2596 29504
rect 1084 29464 2596 29492
rect 1084 29452 1090 29464
rect 2590 29452 2596 29464
rect 2648 29452 2654 29504
rect 3326 29452 3332 29504
rect 3384 29492 3390 29504
rect 4798 29492 4804 29504
rect 3384 29464 4804 29492
rect 3384 29452 3390 29464
rect 4798 29452 4804 29464
rect 4856 29452 4862 29504
rect 7190 29452 7196 29504
rect 7248 29452 7254 29504
rect 7300 29492 7328 29659
rect 8938 29656 8944 29708
rect 8996 29696 9002 29708
rect 9033 29699 9091 29705
rect 9033 29696 9045 29699
rect 8996 29668 9045 29696
rect 8996 29656 9002 29668
rect 9033 29665 9045 29668
rect 9079 29665 9091 29699
rect 9033 29659 9091 29665
rect 11698 29656 11704 29708
rect 11756 29696 11762 29708
rect 12452 29705 12480 29736
rect 13538 29724 13544 29736
rect 13596 29764 13602 29776
rect 13740 29764 13768 29804
rect 14550 29792 14556 29804
rect 14608 29792 14614 29844
rect 17126 29832 17132 29844
rect 16776 29804 17132 29832
rect 13596 29736 13768 29764
rect 13596 29724 13602 29736
rect 12437 29699 12495 29705
rect 11756 29668 11928 29696
rect 11756 29656 11762 29668
rect 10416 29650 10468 29656
rect 7527 29631 7585 29637
rect 7527 29628 7539 29631
rect 7392 29600 7539 29628
rect 7392 29572 7420 29600
rect 7527 29597 7539 29600
rect 7573 29597 7585 29631
rect 7527 29591 7585 29597
rect 8202 29588 8208 29640
rect 8260 29628 8266 29640
rect 9306 29628 9312 29640
rect 8260 29600 9312 29628
rect 8260 29588 8266 29600
rect 9306 29588 9312 29600
rect 9364 29588 9370 29640
rect 10870 29588 10876 29640
rect 10928 29588 10934 29640
rect 10965 29631 11023 29637
rect 10965 29597 10977 29631
rect 11011 29628 11023 29631
rect 11790 29628 11796 29640
rect 11011 29600 11796 29628
rect 11011 29597 11023 29600
rect 10965 29591 11023 29597
rect 11790 29588 11796 29600
rect 11848 29588 11854 29640
rect 11900 29628 11928 29668
rect 12437 29665 12449 29699
rect 12483 29665 12495 29699
rect 12437 29659 12495 29665
rect 15562 29656 15568 29708
rect 15620 29656 15626 29708
rect 16776 29705 16804 29804
rect 17126 29792 17132 29804
rect 17184 29792 17190 29844
rect 17773 29835 17831 29841
rect 17773 29801 17785 29835
rect 17819 29832 17831 29835
rect 18138 29832 18144 29844
rect 17819 29804 18144 29832
rect 17819 29801 17831 29804
rect 17773 29795 17831 29801
rect 18138 29792 18144 29804
rect 18196 29792 18202 29844
rect 18601 29835 18659 29841
rect 18601 29801 18613 29835
rect 18647 29832 18659 29835
rect 18966 29832 18972 29844
rect 18647 29804 18972 29832
rect 18647 29801 18659 29804
rect 18601 29795 18659 29801
rect 18966 29792 18972 29804
rect 19024 29792 19030 29844
rect 19797 29835 19855 29841
rect 19797 29801 19809 29835
rect 19843 29832 19855 29835
rect 19886 29832 19892 29844
rect 19843 29804 19892 29832
rect 19843 29801 19855 29804
rect 19797 29795 19855 29801
rect 17586 29724 17592 29776
rect 17644 29764 17650 29776
rect 19245 29767 19303 29773
rect 17644 29736 19104 29764
rect 17644 29724 17650 29736
rect 16761 29699 16819 29705
rect 16761 29665 16773 29699
rect 16807 29665 16819 29699
rect 16761 29659 16819 29665
rect 18598 29656 18604 29708
rect 18656 29696 18662 29708
rect 18656 29668 19012 29696
rect 18656 29656 18662 29668
rect 12679 29631 12737 29637
rect 12679 29628 12691 29631
rect 11900 29600 12691 29628
rect 12679 29597 12691 29600
rect 12725 29628 12737 29631
rect 13170 29628 13176 29640
rect 12725 29600 13176 29628
rect 12725 29597 12737 29600
rect 12679 29591 12737 29597
rect 13170 29588 13176 29600
rect 13228 29588 13234 29640
rect 14277 29631 14335 29637
rect 14277 29597 14289 29631
rect 14323 29597 14335 29631
rect 14550 29628 14556 29640
rect 14511 29600 14556 29628
rect 14277 29591 14335 29597
rect 7374 29520 7380 29572
rect 7432 29520 7438 29572
rect 8294 29520 8300 29572
rect 8352 29560 8358 29572
rect 8352 29532 9904 29560
rect 8352 29520 8358 29532
rect 9876 29504 9904 29532
rect 11238 29520 11244 29572
rect 11296 29560 11302 29572
rect 11333 29563 11391 29569
rect 11333 29560 11345 29563
rect 11296 29532 11345 29560
rect 11296 29520 11302 29532
rect 11333 29529 11345 29532
rect 11379 29529 11391 29563
rect 14292 29560 14320 29591
rect 14550 29588 14556 29600
rect 14608 29588 14614 29640
rect 14642 29560 14648 29572
rect 14292 29532 14648 29560
rect 11333 29523 11391 29529
rect 14642 29520 14648 29532
rect 14700 29560 14706 29572
rect 15580 29560 15608 29656
rect 16942 29588 16948 29640
rect 17000 29628 17006 29640
rect 17035 29631 17093 29637
rect 17035 29628 17047 29631
rect 17000 29600 17047 29628
rect 17000 29588 17006 29600
rect 17035 29597 17047 29600
rect 17081 29597 17093 29631
rect 17035 29591 17093 29597
rect 18785 29631 18843 29637
rect 18785 29597 18797 29631
rect 18831 29628 18843 29631
rect 18831 29600 18920 29628
rect 18831 29597 18843 29600
rect 18785 29591 18843 29597
rect 14700 29532 15608 29560
rect 14700 29520 14706 29532
rect 7650 29492 7656 29504
rect 7300 29464 7656 29492
rect 7650 29452 7656 29464
rect 7708 29452 7714 29504
rect 9858 29452 9864 29504
rect 9916 29452 9922 29504
rect 10042 29452 10048 29504
rect 10100 29452 10106 29504
rect 10597 29495 10655 29501
rect 10597 29461 10609 29495
rect 10643 29492 10655 29495
rect 11606 29492 11612 29504
rect 10643 29464 11612 29492
rect 10643 29461 10655 29464
rect 10597 29455 10655 29461
rect 11606 29452 11612 29464
rect 11664 29452 11670 29504
rect 11698 29452 11704 29504
rect 11756 29452 11762 29504
rect 11885 29495 11943 29501
rect 11885 29461 11897 29495
rect 11931 29492 11943 29495
rect 12434 29492 12440 29504
rect 11931 29464 12440 29492
rect 11931 29461 11943 29464
rect 11885 29455 11943 29461
rect 12434 29452 12440 29464
rect 12492 29452 12498 29504
rect 12710 29452 12716 29504
rect 12768 29492 12774 29504
rect 14550 29492 14556 29504
rect 12768 29464 14556 29492
rect 12768 29452 12774 29464
rect 14550 29452 14556 29464
rect 14608 29452 14614 29504
rect 15010 29452 15016 29504
rect 15068 29492 15074 29504
rect 15289 29495 15347 29501
rect 15289 29492 15301 29495
rect 15068 29464 15301 29492
rect 15068 29452 15074 29464
rect 15289 29461 15301 29464
rect 15335 29461 15347 29495
rect 15289 29455 15347 29461
rect 15470 29452 15476 29504
rect 15528 29492 15534 29504
rect 18598 29492 18604 29504
rect 15528 29464 18604 29492
rect 15528 29452 15534 29464
rect 18598 29452 18604 29464
rect 18656 29452 18662 29504
rect 18892 29501 18920 29600
rect 18984 29560 19012 29668
rect 19076 29637 19104 29736
rect 19245 29733 19257 29767
rect 19291 29764 19303 29767
rect 19518 29764 19524 29776
rect 19291 29736 19524 29764
rect 19291 29733 19303 29736
rect 19245 29727 19303 29733
rect 19518 29724 19524 29736
rect 19576 29724 19582 29776
rect 19061 29631 19119 29637
rect 19061 29597 19073 29631
rect 19107 29597 19119 29631
rect 19061 29591 19119 29597
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29628 19487 29631
rect 19812 29628 19840 29795
rect 19886 29792 19892 29804
rect 19944 29792 19950 29844
rect 19475 29600 19840 29628
rect 19475 29597 19487 29600
rect 19429 29591 19487 29597
rect 20165 29563 20223 29569
rect 20165 29560 20177 29563
rect 18984 29532 20177 29560
rect 20165 29529 20177 29532
rect 20211 29529 20223 29563
rect 20165 29523 20223 29529
rect 20533 29563 20591 29569
rect 20533 29529 20545 29563
rect 20579 29560 20591 29563
rect 21266 29560 21272 29572
rect 20579 29532 21272 29560
rect 20579 29529 20591 29532
rect 20533 29523 20591 29529
rect 21266 29520 21272 29532
rect 21324 29520 21330 29572
rect 18877 29495 18935 29501
rect 18877 29461 18889 29495
rect 18923 29461 18935 29495
rect 18877 29455 18935 29461
rect 1104 29402 21043 29424
rect 1104 29350 5894 29402
rect 5946 29350 5958 29402
rect 6010 29350 6022 29402
rect 6074 29350 6086 29402
rect 6138 29350 6150 29402
rect 6202 29350 10839 29402
rect 10891 29350 10903 29402
rect 10955 29350 10967 29402
rect 11019 29350 11031 29402
rect 11083 29350 11095 29402
rect 11147 29350 15784 29402
rect 15836 29350 15848 29402
rect 15900 29350 15912 29402
rect 15964 29350 15976 29402
rect 16028 29350 16040 29402
rect 16092 29350 20729 29402
rect 20781 29350 20793 29402
rect 20845 29350 20857 29402
rect 20909 29350 20921 29402
rect 20973 29350 20985 29402
rect 21037 29350 21043 29402
rect 1104 29328 21043 29350
rect 1302 29248 1308 29300
rect 1360 29288 1366 29300
rect 2409 29291 2467 29297
rect 2409 29288 2421 29291
rect 1360 29260 2421 29288
rect 1360 29248 1366 29260
rect 2409 29257 2421 29260
rect 2455 29257 2467 29291
rect 3878 29288 3884 29300
rect 2409 29251 2467 29257
rect 2976 29260 3884 29288
rect 2976 29232 3004 29260
rect 3878 29248 3884 29260
rect 3936 29248 3942 29300
rect 3970 29248 3976 29300
rect 4028 29288 4034 29300
rect 4246 29288 4252 29300
rect 4028 29260 4252 29288
rect 4028 29248 4034 29260
rect 4246 29248 4252 29260
rect 4304 29248 4310 29300
rect 4430 29248 4436 29300
rect 4488 29248 4494 29300
rect 4706 29248 4712 29300
rect 4764 29288 4770 29300
rect 4982 29288 4988 29300
rect 4764 29260 4988 29288
rect 4764 29248 4770 29260
rect 4982 29248 4988 29260
rect 5040 29248 5046 29300
rect 7650 29288 7656 29300
rect 5092 29260 7656 29288
rect 2038 29220 2044 29232
rect 1962 29192 2044 29220
rect 1671 29165 1729 29171
rect 1026 29112 1032 29164
rect 1084 29152 1090 29164
rect 1397 29155 1455 29161
rect 1397 29152 1409 29155
rect 1084 29124 1409 29152
rect 1084 29112 1090 29124
rect 1397 29121 1409 29124
rect 1443 29121 1455 29155
rect 1671 29131 1683 29165
rect 1717 29162 1729 29165
rect 1962 29162 1990 29192
rect 2038 29180 2044 29192
rect 2096 29220 2102 29232
rect 2096 29192 2728 29220
rect 2096 29180 2102 29192
rect 1717 29134 1990 29162
rect 2590 29152 2596 29164
rect 1717 29131 1729 29134
rect 1671 29125 1729 29131
rect 2056 29130 2596 29152
rect 1397 29115 1455 29121
rect 2038 29078 2044 29130
rect 2096 29124 2596 29130
rect 2096 29078 2102 29124
rect 2590 29112 2596 29124
rect 2648 29112 2654 29164
rect 2700 29084 2728 29192
rect 2958 29180 2964 29232
rect 3016 29180 3022 29232
rect 5092 29220 5120 29260
rect 7650 29248 7656 29260
rect 7708 29288 7714 29300
rect 8202 29288 8208 29300
rect 7708 29260 8208 29288
rect 7708 29248 7714 29260
rect 8202 29248 8208 29260
rect 8260 29248 8266 29300
rect 9214 29288 9220 29300
rect 8956 29260 9220 29288
rect 4264 29192 4844 29220
rect 2866 29112 2872 29164
rect 2924 29112 2930 29164
rect 2976 29152 3004 29180
rect 4264 29164 4292 29192
rect 3111 29155 3169 29161
rect 3111 29152 3123 29155
rect 2976 29124 3123 29152
rect 3111 29121 3123 29124
rect 3157 29121 3169 29155
rect 3111 29115 3169 29121
rect 4246 29112 4252 29164
rect 4304 29112 4310 29164
rect 4525 29155 4583 29161
rect 4525 29121 4537 29155
rect 4571 29121 4583 29155
rect 4525 29115 4583 29121
rect 2700 29056 2774 29084
rect 566 28908 572 28960
rect 624 28948 630 28960
rect 2498 28948 2504 28960
rect 624 28920 2504 28948
rect 624 28908 630 28920
rect 2498 28908 2504 28920
rect 2556 28908 2562 28960
rect 2746 28948 2774 29056
rect 3786 29044 3792 29096
rect 3844 29084 3850 29096
rect 4540 29084 4568 29115
rect 4816 29096 4844 29192
rect 4908 29192 5120 29220
rect 4908 29161 4936 29192
rect 5442 29180 5448 29232
rect 5500 29180 5506 29232
rect 7098 29220 7104 29232
rect 5570 29192 7104 29220
rect 4893 29155 4951 29161
rect 4893 29121 4905 29155
rect 4939 29121 4951 29155
rect 4893 29115 4951 29121
rect 5167 29155 5225 29161
rect 5167 29121 5179 29155
rect 5213 29152 5225 29155
rect 5460 29152 5488 29180
rect 5213 29124 5488 29152
rect 5213 29121 5225 29124
rect 5167 29115 5225 29121
rect 3844 29056 4568 29084
rect 3844 29044 3850 29056
rect 4798 29044 4804 29096
rect 4856 29044 4862 29096
rect 3878 28976 3884 29028
rect 3936 28976 3942 29028
rect 5570 29016 5598 29192
rect 7098 29180 7104 29192
rect 7156 29180 7162 29232
rect 7190 29180 7196 29232
rect 7248 29180 7254 29232
rect 7374 29191 7380 29232
rect 7359 29185 7380 29191
rect 7432 29220 7438 29232
rect 7558 29220 7564 29232
rect 7432 29192 7564 29220
rect 7009 29155 7067 29161
rect 7009 29121 7021 29155
rect 7055 29152 7067 29155
rect 7208 29152 7236 29180
rect 7055 29124 7236 29152
rect 7359 29151 7371 29185
rect 7432 29180 7438 29192
rect 7558 29180 7564 29192
rect 7616 29180 7622 29232
rect 8956 29229 8984 29260
rect 9214 29248 9220 29260
rect 9272 29248 9278 29300
rect 9674 29288 9680 29300
rect 9324 29260 9680 29288
rect 8665 29223 8723 29229
rect 8665 29189 8677 29223
rect 8711 29189 8723 29223
rect 8665 29183 8723 29189
rect 8941 29223 8999 29229
rect 8941 29189 8953 29223
rect 8987 29189 8999 29223
rect 8941 29183 8999 29189
rect 9033 29223 9091 29229
rect 9033 29189 9045 29223
rect 9079 29220 9091 29223
rect 9324 29220 9352 29260
rect 9674 29248 9680 29260
rect 9732 29248 9738 29300
rect 9769 29291 9827 29297
rect 9769 29257 9781 29291
rect 9815 29288 9827 29291
rect 9858 29288 9864 29300
rect 9815 29260 9864 29288
rect 9815 29257 9827 29260
rect 9769 29251 9827 29257
rect 9858 29248 9864 29260
rect 9916 29248 9922 29300
rect 10502 29248 10508 29300
rect 10560 29288 10566 29300
rect 11698 29288 11704 29300
rect 10560 29260 11704 29288
rect 10560 29248 10566 29260
rect 11348 29232 11376 29260
rect 11698 29248 11704 29260
rect 11756 29248 11762 29300
rect 12250 29248 12256 29300
rect 12308 29248 12314 29300
rect 13170 29248 13176 29300
rect 13228 29288 13234 29300
rect 14734 29288 14740 29300
rect 13228 29260 14740 29288
rect 13228 29248 13234 29260
rect 14734 29248 14740 29260
rect 14792 29288 14798 29300
rect 17586 29288 17592 29300
rect 14792 29260 17592 29288
rect 14792 29248 14798 29260
rect 17586 29248 17592 29260
rect 17644 29248 17650 29300
rect 18417 29291 18475 29297
rect 18417 29257 18429 29291
rect 18463 29257 18475 29291
rect 18417 29251 18475 29257
rect 18693 29291 18751 29297
rect 18693 29257 18705 29291
rect 18739 29288 18751 29291
rect 18874 29288 18880 29300
rect 18739 29260 18880 29288
rect 18739 29257 18751 29260
rect 18693 29251 18751 29257
rect 9079 29192 9352 29220
rect 9079 29189 9091 29192
rect 9033 29183 9091 29189
rect 7405 29154 7420 29180
rect 7405 29151 7417 29154
rect 7359 29145 7417 29151
rect 8680 29152 8708 29183
rect 9398 29180 9404 29232
rect 9456 29180 9462 29232
rect 10229 29223 10287 29229
rect 10229 29220 10241 29223
rect 9646 29192 10241 29220
rect 9646 29152 9674 29192
rect 10229 29189 10241 29192
rect 10275 29220 10287 29223
rect 10686 29220 10692 29232
rect 10275 29192 10692 29220
rect 10275 29189 10287 29192
rect 10229 29183 10287 29189
rect 10686 29180 10692 29192
rect 10744 29180 10750 29232
rect 11330 29180 11336 29232
rect 11388 29180 11394 29232
rect 8680 29124 9674 29152
rect 11791 29155 11849 29161
rect 7055 29121 7067 29124
rect 7009 29115 7067 29121
rect 11791 29121 11803 29155
rect 11837 29152 11849 29155
rect 12268 29152 12296 29248
rect 17310 29220 17316 29232
rect 14016 29192 17316 29220
rect 13415 29155 13473 29161
rect 13415 29152 13427 29155
rect 11837 29124 12204 29152
rect 12268 29124 13427 29152
rect 11837 29121 11849 29124
rect 11791 29115 11849 29121
rect 7101 29087 7159 29093
rect 7101 29084 7113 29087
rect 7024 29056 7113 29084
rect 7024 29028 7052 29056
rect 7101 29053 7113 29056
rect 7147 29053 7159 29087
rect 11517 29087 11575 29093
rect 7101 29047 7159 29053
rect 5552 28988 5598 29016
rect 6825 29019 6883 29025
rect 2866 28948 2872 28960
rect 2746 28920 2872 28948
rect 2866 28908 2872 28920
rect 2924 28908 2930 28960
rect 4798 28908 4804 28960
rect 4856 28948 4862 28960
rect 5552 28948 5580 28988
rect 6825 28985 6837 29019
rect 6871 29016 6883 29019
rect 6914 29016 6920 29028
rect 6871 28988 6920 29016
rect 6871 28985 6883 28988
rect 6825 28979 6883 28985
rect 6914 28976 6920 28988
rect 6972 28976 6978 29028
rect 7006 28976 7012 29028
rect 7064 28976 7070 29028
rect 8113 29019 8171 29025
rect 8113 28985 8125 29019
rect 8159 29016 8171 29019
rect 8496 29016 8524 29070
rect 11517 29053 11529 29087
rect 11563 29053 11575 29087
rect 12176 29084 12204 29124
rect 13415 29121 13427 29124
rect 13461 29152 13473 29155
rect 14016 29152 14044 29192
rect 17310 29180 17316 29192
rect 17368 29180 17374 29232
rect 18432 29220 18460 29251
rect 18874 29248 18880 29260
rect 18932 29248 18938 29300
rect 18969 29291 19027 29297
rect 18969 29257 18981 29291
rect 19015 29288 19027 29291
rect 19610 29288 19616 29300
rect 19015 29260 19616 29288
rect 19015 29257 19027 29260
rect 18969 29251 19027 29257
rect 19610 29248 19616 29260
rect 19668 29248 19674 29300
rect 18432 29192 19472 29220
rect 13461 29124 14044 29152
rect 13461 29121 13473 29124
rect 13415 29115 13473 29121
rect 14090 29112 14096 29164
rect 14148 29152 14154 29164
rect 14795 29155 14853 29161
rect 14795 29152 14807 29155
rect 14148 29124 14807 29152
rect 14148 29112 14154 29124
rect 14795 29121 14807 29124
rect 14841 29121 14853 29155
rect 14795 29115 14853 29121
rect 17770 29112 17776 29164
rect 17828 29152 17834 29164
rect 18601 29155 18659 29161
rect 18601 29152 18613 29155
rect 17828 29124 18613 29152
rect 17828 29112 17834 29124
rect 18601 29121 18613 29124
rect 18647 29121 18659 29155
rect 18601 29115 18659 29121
rect 18874 29112 18880 29164
rect 18932 29112 18938 29164
rect 19150 29112 19156 29164
rect 19208 29112 19214 29164
rect 19444 29161 19472 29192
rect 20162 29180 20168 29232
rect 20220 29180 20226 29232
rect 19429 29155 19487 29161
rect 19429 29121 19441 29155
rect 19475 29121 19487 29155
rect 19429 29115 19487 29121
rect 19521 29155 19579 29161
rect 19521 29121 19533 29155
rect 19567 29121 19579 29155
rect 19521 29115 19579 29121
rect 12710 29084 12716 29096
rect 12176 29056 12716 29084
rect 11517 29047 11575 29053
rect 8159 28988 8524 29016
rect 8159 28985 8171 28988
rect 8113 28979 8171 28985
rect 10410 28976 10416 29028
rect 10468 28976 10474 29028
rect 11532 29016 11560 29047
rect 12710 29044 12716 29056
rect 12768 29044 12774 29096
rect 13173 29087 13231 29093
rect 13173 29053 13185 29087
rect 13219 29053 13231 29087
rect 14550 29084 14556 29096
rect 13173 29047 13231 29053
rect 13832 29056 14556 29084
rect 11532 28988 11652 29016
rect 11624 28960 11652 28988
rect 12250 28976 12256 29028
rect 12308 29016 12314 29028
rect 12529 29019 12587 29025
rect 12529 29016 12541 29019
rect 12308 28988 12541 29016
rect 12308 28976 12314 28988
rect 12529 28985 12541 28988
rect 12575 28985 12587 29019
rect 12529 28979 12587 28985
rect 4856 28920 5580 28948
rect 5905 28951 5963 28957
rect 4856 28908 4862 28920
rect 5905 28917 5917 28951
rect 5951 28948 5963 28951
rect 6730 28948 6736 28960
rect 5951 28920 6736 28948
rect 5951 28917 5963 28920
rect 5905 28911 5963 28917
rect 6730 28908 6736 28920
rect 6788 28948 6794 28960
rect 7098 28948 7104 28960
rect 6788 28920 7104 28948
rect 6788 28908 6794 28920
rect 7098 28908 7104 28920
rect 7156 28908 7162 28960
rect 9953 28951 10011 28957
rect 9953 28917 9965 28951
rect 9999 28948 10011 28951
rect 10318 28948 10324 28960
rect 9999 28920 10324 28948
rect 9999 28917 10011 28920
rect 9953 28911 10011 28917
rect 10318 28908 10324 28920
rect 10376 28948 10382 28960
rect 11238 28948 11244 28960
rect 10376 28920 11244 28948
rect 10376 28908 10382 28920
rect 11238 28908 11244 28920
rect 11296 28908 11302 28960
rect 11606 28908 11612 28960
rect 11664 28908 11670 28960
rect 13188 28948 13216 29047
rect 13832 28948 13860 29056
rect 14550 29044 14556 29056
rect 14608 29044 14614 29096
rect 19242 29044 19248 29096
rect 19300 29084 19306 29096
rect 19536 29084 19564 29115
rect 19886 29112 19892 29164
rect 19944 29152 19950 29164
rect 19981 29155 20039 29161
rect 19981 29152 19993 29155
rect 19944 29124 19993 29152
rect 19944 29112 19950 29124
rect 19981 29121 19993 29124
rect 20027 29121 20039 29155
rect 19981 29115 20039 29121
rect 19300 29056 19564 29084
rect 19300 29044 19306 29056
rect 19794 29044 19800 29096
rect 19852 29044 19858 29096
rect 17862 28976 17868 29028
rect 17920 29016 17926 29028
rect 19150 29016 19156 29028
rect 17920 28988 19156 29016
rect 17920 28976 17926 28988
rect 19150 28976 19156 28988
rect 19208 28976 19214 29028
rect 19812 29016 19840 29044
rect 19260 28988 19840 29016
rect 13188 28920 13860 28948
rect 14182 28908 14188 28960
rect 14240 28908 14246 28960
rect 15470 28908 15476 28960
rect 15528 28948 15534 28960
rect 19260 28957 19288 28988
rect 20438 28976 20444 29028
rect 20496 28976 20502 29028
rect 15565 28951 15623 28957
rect 15565 28948 15577 28951
rect 15528 28920 15577 28948
rect 15528 28908 15534 28920
rect 15565 28917 15577 28920
rect 15611 28917 15623 28951
rect 15565 28911 15623 28917
rect 19245 28951 19303 28957
rect 19245 28917 19257 28951
rect 19291 28917 19303 28951
rect 19245 28911 19303 28917
rect 19610 28908 19616 28960
rect 19668 28908 19674 28960
rect 19794 28908 19800 28960
rect 19852 28908 19858 28960
rect 1104 28858 20884 28880
rect 1104 28806 3422 28858
rect 3474 28806 3486 28858
rect 3538 28806 3550 28858
rect 3602 28806 3614 28858
rect 3666 28806 3678 28858
rect 3730 28806 8367 28858
rect 8419 28806 8431 28858
rect 8483 28806 8495 28858
rect 8547 28806 8559 28858
rect 8611 28806 8623 28858
rect 8675 28806 13312 28858
rect 13364 28806 13376 28858
rect 13428 28806 13440 28858
rect 13492 28806 13504 28858
rect 13556 28806 13568 28858
rect 13620 28806 18257 28858
rect 18309 28806 18321 28858
rect 18373 28806 18385 28858
rect 18437 28806 18449 28858
rect 18501 28806 18513 28858
rect 18565 28806 20884 28858
rect 1104 28784 20884 28806
rect 4430 28744 4436 28756
rect 3988 28716 4436 28744
rect 1210 28568 1216 28620
rect 1268 28608 1274 28620
rect 2317 28611 2375 28617
rect 2317 28608 2329 28611
rect 1268 28580 2329 28608
rect 1268 28568 1274 28580
rect 2317 28577 2329 28580
rect 2363 28577 2375 28611
rect 2317 28571 2375 28577
rect 2590 28568 2596 28620
rect 2648 28568 2654 28620
rect 3988 28617 4016 28716
rect 4430 28704 4436 28716
rect 4488 28744 4494 28756
rect 4890 28744 4896 28756
rect 4488 28716 4896 28744
rect 4488 28704 4494 28716
rect 4890 28704 4896 28716
rect 4948 28704 4954 28756
rect 6822 28744 6828 28756
rect 6196 28716 6828 28744
rect 5534 28636 5540 28688
rect 5592 28676 5598 28688
rect 5718 28676 5724 28688
rect 5592 28648 5724 28676
rect 5592 28636 5598 28648
rect 5718 28636 5724 28648
rect 5776 28636 5782 28688
rect 6196 28685 6224 28716
rect 6822 28704 6828 28716
rect 6880 28704 6886 28756
rect 6914 28704 6920 28756
rect 6972 28744 6978 28756
rect 8113 28747 8171 28753
rect 6972 28716 8064 28744
rect 6972 28704 6978 28716
rect 6181 28679 6239 28685
rect 6181 28645 6193 28679
rect 6227 28645 6239 28679
rect 6181 28639 6239 28645
rect 7745 28679 7803 28685
rect 7745 28645 7757 28679
rect 7791 28676 7803 28679
rect 7926 28676 7932 28688
rect 7791 28648 7932 28676
rect 7791 28645 7803 28648
rect 7745 28639 7803 28645
rect 7926 28636 7932 28648
rect 7984 28636 7990 28688
rect 3973 28611 4031 28617
rect 3973 28577 3985 28611
rect 4019 28577 4031 28611
rect 7098 28608 7104 28620
rect 3973 28571 4031 28577
rect 6746 28580 7104 28608
rect 750 28500 756 28552
rect 808 28540 814 28552
rect 1489 28543 1547 28549
rect 1489 28540 1501 28543
rect 808 28512 1501 28540
rect 808 28500 814 28512
rect 1489 28509 1501 28512
rect 1535 28509 1547 28543
rect 1489 28503 1547 28509
rect 3234 28500 3240 28552
rect 3292 28500 3298 28552
rect 4247 28543 4305 28549
rect 4247 28509 4259 28543
rect 4293 28540 4305 28543
rect 4614 28540 4620 28552
rect 4293 28512 4620 28540
rect 4293 28509 4305 28512
rect 4247 28503 4305 28509
rect 4614 28500 4620 28512
rect 4672 28540 4678 28552
rect 5350 28540 5356 28552
rect 4672 28512 5356 28540
rect 4672 28500 4678 28512
rect 5350 28500 5356 28512
rect 5408 28500 5414 28552
rect 5442 28500 5448 28552
rect 5500 28540 5506 28552
rect 5537 28543 5595 28549
rect 5537 28540 5549 28543
rect 5500 28512 5549 28540
rect 5500 28500 5506 28512
rect 5537 28509 5549 28512
rect 5583 28509 5595 28543
rect 5537 28503 5595 28509
rect 5718 28500 5724 28552
rect 5776 28500 5782 28552
rect 6454 28500 6460 28552
rect 6512 28500 6518 28552
rect 6546 28500 6552 28552
rect 6604 28549 6610 28552
rect 6746 28549 6774 28580
rect 7098 28568 7104 28580
rect 7156 28568 7162 28620
rect 8036 28549 8064 28716
rect 8113 28713 8125 28747
rect 8159 28744 8171 28747
rect 8754 28744 8760 28756
rect 8159 28716 8760 28744
rect 8159 28713 8171 28716
rect 8113 28707 8171 28713
rect 8754 28704 8760 28716
rect 8812 28704 8818 28756
rect 12894 28704 12900 28756
rect 12952 28744 12958 28756
rect 13538 28744 13544 28756
rect 12952 28716 13544 28744
rect 12952 28704 12958 28716
rect 13538 28704 13544 28716
rect 13596 28704 13602 28756
rect 14182 28704 14188 28756
rect 14240 28704 14246 28756
rect 15933 28747 15991 28753
rect 15933 28713 15945 28747
rect 15979 28744 15991 28747
rect 15979 28716 17724 28744
rect 15979 28713 15991 28716
rect 15933 28707 15991 28713
rect 14200 28676 14228 28704
rect 14737 28679 14795 28685
rect 14737 28676 14749 28679
rect 14200 28648 14749 28676
rect 14737 28645 14749 28648
rect 14783 28645 14795 28679
rect 14737 28639 14795 28645
rect 14277 28611 14335 28617
rect 14277 28608 14289 28611
rect 8680 28580 9246 28608
rect 13004 28580 14289 28608
rect 8680 28552 8708 28580
rect 13004 28552 13032 28580
rect 14277 28577 14289 28580
rect 14323 28577 14335 28611
rect 14277 28571 14335 28577
rect 14826 28568 14832 28620
rect 14884 28608 14890 28620
rect 15013 28611 15071 28617
rect 15013 28608 15025 28611
rect 14884 28580 15025 28608
rect 14884 28568 14890 28580
rect 15013 28577 15025 28580
rect 15059 28577 15071 28611
rect 15013 28571 15071 28577
rect 15289 28611 15347 28617
rect 15289 28577 15301 28611
rect 15335 28608 15347 28611
rect 15470 28608 15476 28620
rect 15335 28580 15476 28608
rect 15335 28577 15347 28580
rect 15289 28571 15347 28577
rect 15470 28568 15476 28580
rect 15528 28568 15534 28620
rect 17696 28608 17724 28716
rect 18874 28704 18880 28756
rect 18932 28744 18938 28756
rect 19061 28747 19119 28753
rect 19061 28744 19073 28747
rect 18932 28716 19073 28744
rect 18932 28704 18938 28716
rect 19061 28713 19073 28716
rect 19107 28713 19119 28747
rect 19061 28707 19119 28713
rect 19242 28704 19248 28756
rect 19300 28704 19306 28756
rect 19610 28704 19616 28756
rect 19668 28744 19674 28756
rect 19981 28747 20039 28753
rect 19981 28744 19993 28747
rect 19668 28716 19993 28744
rect 19668 28704 19674 28716
rect 19981 28713 19993 28716
rect 20027 28713 20039 28747
rect 19981 28707 20039 28713
rect 20070 28704 20076 28756
rect 20128 28704 20134 28756
rect 19702 28636 19708 28688
rect 19760 28636 19766 28688
rect 19720 28608 19748 28636
rect 20088 28608 20116 28704
rect 20165 28611 20223 28617
rect 20165 28608 20177 28611
rect 17696 28580 17816 28608
rect 19720 28580 19932 28608
rect 20088 28580 20177 28608
rect 6604 28543 6632 28549
rect 6620 28509 6632 28543
rect 6604 28503 6632 28509
rect 6733 28543 6791 28549
rect 6733 28509 6745 28543
rect 6779 28509 6791 28543
rect 6733 28503 6791 28509
rect 7377 28543 7435 28549
rect 7377 28509 7389 28543
rect 7423 28540 7435 28543
rect 7929 28543 7987 28549
rect 7929 28540 7941 28543
rect 7423 28512 7941 28540
rect 7423 28509 7435 28512
rect 7377 28503 7435 28509
rect 7929 28509 7941 28512
rect 7975 28509 7987 28543
rect 7929 28503 7987 28509
rect 8021 28543 8079 28549
rect 8021 28509 8033 28543
rect 8067 28509 8079 28543
rect 8021 28503 8079 28509
rect 6604 28500 6610 28503
rect 8662 28500 8668 28552
rect 8720 28500 8726 28552
rect 9582 28500 9588 28552
rect 9640 28540 9646 28552
rect 9677 28543 9735 28549
rect 9677 28540 9689 28543
rect 9640 28512 9689 28540
rect 9640 28500 9646 28512
rect 9677 28509 9689 28512
rect 9723 28509 9735 28543
rect 9677 28503 9735 28509
rect 10042 28500 10048 28552
rect 10100 28500 10106 28552
rect 10137 28543 10195 28549
rect 10137 28509 10149 28543
rect 10183 28540 10195 28543
rect 10318 28540 10324 28552
rect 10183 28512 10324 28540
rect 10183 28509 10195 28512
rect 10137 28503 10195 28509
rect 10318 28500 10324 28512
rect 10376 28500 10382 28552
rect 11517 28543 11575 28549
rect 11517 28509 11529 28543
rect 11563 28540 11575 28543
rect 11698 28540 11704 28552
rect 11563 28512 11704 28540
rect 11563 28509 11575 28512
rect 11517 28503 11575 28509
rect 11698 28500 11704 28512
rect 11756 28500 11762 28552
rect 11791 28543 11849 28549
rect 11791 28509 11803 28543
rect 11837 28540 11849 28543
rect 11882 28540 11888 28552
rect 11837 28512 11888 28540
rect 11837 28509 11849 28512
rect 11791 28503 11849 28509
rect 11882 28500 11888 28512
rect 11940 28540 11946 28552
rect 12710 28540 12716 28552
rect 11940 28512 12716 28540
rect 11940 28500 11946 28512
rect 12710 28500 12716 28512
rect 12768 28500 12774 28552
rect 12986 28500 12992 28552
rect 13044 28500 13050 28552
rect 13078 28500 13084 28552
rect 13136 28540 13142 28552
rect 15194 28549 15200 28552
rect 14093 28543 14151 28549
rect 14093 28540 14105 28543
rect 13136 28512 14105 28540
rect 13136 28500 13142 28512
rect 14093 28509 14105 28512
rect 14139 28509 14151 28543
rect 14093 28503 14151 28509
rect 15151 28543 15200 28549
rect 15151 28509 15163 28543
rect 15197 28509 15200 28543
rect 15151 28503 15200 28509
rect 15194 28500 15200 28503
rect 15252 28500 15258 28552
rect 16025 28543 16083 28549
rect 16025 28509 16037 28543
rect 16071 28540 16083 28543
rect 16666 28540 16672 28552
rect 16071 28512 16672 28540
rect 16071 28509 16083 28512
rect 16025 28503 16083 28509
rect 1670 28432 1676 28484
rect 1728 28432 1734 28484
rect 9769 28475 9827 28481
rect 3436 28444 5764 28472
rect 934 28364 940 28416
rect 992 28404 998 28416
rect 2590 28404 2596 28416
rect 992 28376 2596 28404
rect 992 28364 998 28376
rect 2590 28364 2596 28376
rect 2648 28364 2654 28416
rect 3436 28413 3464 28444
rect 3421 28407 3479 28413
rect 3421 28373 3433 28407
rect 3467 28373 3479 28407
rect 3421 28367 3479 28373
rect 4982 28364 4988 28416
rect 5040 28364 5046 28416
rect 5736 28404 5764 28444
rect 7944 28444 9628 28472
rect 7944 28404 7972 28444
rect 5736 28376 7972 28404
rect 8294 28364 8300 28416
rect 8352 28404 8358 28416
rect 9398 28404 9404 28416
rect 8352 28376 9404 28404
rect 8352 28364 8358 28376
rect 9398 28364 9404 28376
rect 9456 28364 9462 28416
rect 9600 28404 9628 28444
rect 9769 28441 9781 28475
rect 9815 28472 9827 28475
rect 10060 28472 10088 28500
rect 14274 28472 14280 28484
rect 9815 28444 10088 28472
rect 10428 28444 14280 28472
rect 9815 28441 9827 28444
rect 9769 28435 9827 28441
rect 10428 28404 10456 28444
rect 14274 28432 14280 28444
rect 14332 28432 14338 28484
rect 9600 28376 10456 28404
rect 10502 28364 10508 28416
rect 10560 28364 10566 28416
rect 10686 28364 10692 28416
rect 10744 28364 10750 28416
rect 11606 28364 11612 28416
rect 11664 28404 11670 28416
rect 11974 28404 11980 28416
rect 11664 28376 11980 28404
rect 11664 28364 11670 28376
rect 11974 28364 11980 28376
rect 12032 28364 12038 28416
rect 12529 28407 12587 28413
rect 12529 28373 12541 28407
rect 12575 28404 12587 28407
rect 12710 28404 12716 28416
rect 12575 28376 12716 28404
rect 12575 28373 12587 28376
rect 12529 28367 12587 28373
rect 12710 28364 12716 28376
rect 12768 28364 12774 28416
rect 14642 28364 14648 28416
rect 14700 28404 14706 28416
rect 15010 28404 15016 28416
rect 14700 28376 15016 28404
rect 14700 28364 14706 28376
rect 15010 28364 15016 28376
rect 15068 28364 15074 28416
rect 15194 28364 15200 28416
rect 15252 28404 15258 28416
rect 16040 28404 16068 28503
rect 16666 28500 16672 28512
rect 16724 28540 16730 28552
rect 17681 28543 17739 28549
rect 17681 28540 17693 28543
rect 16724 28512 17693 28540
rect 16724 28500 16730 28512
rect 17681 28509 17693 28512
rect 17727 28509 17739 28543
rect 17788 28540 17816 28580
rect 19904 28549 19932 28580
rect 20165 28577 20177 28580
rect 20211 28577 20223 28611
rect 20165 28571 20223 28577
rect 17937 28543 17995 28549
rect 17937 28540 17949 28543
rect 17788 28512 17949 28540
rect 17681 28503 17739 28509
rect 17937 28509 17949 28512
rect 17983 28540 17995 28543
rect 19429 28543 19487 28549
rect 19429 28540 19441 28543
rect 17983 28512 19441 28540
rect 17983 28509 17995 28512
rect 17937 28503 17995 28509
rect 19429 28509 19441 28512
rect 19475 28509 19487 28543
rect 19429 28503 19487 28509
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 19889 28543 19947 28549
rect 19889 28509 19901 28543
rect 19935 28509 19947 28543
rect 19889 28503 19947 28509
rect 16298 28481 16304 28484
rect 16281 28475 16304 28481
rect 16281 28441 16293 28475
rect 16281 28435 16304 28441
rect 16298 28432 16304 28435
rect 16356 28432 16362 28484
rect 19150 28432 19156 28484
rect 19208 28472 19214 28484
rect 19812 28472 19840 28503
rect 19978 28500 19984 28552
rect 20036 28540 20042 28552
rect 20257 28543 20315 28549
rect 20257 28540 20269 28543
rect 20036 28512 20269 28540
rect 20036 28500 20042 28512
rect 20257 28509 20269 28512
rect 20303 28509 20315 28543
rect 20257 28503 20315 28509
rect 19208 28444 19840 28472
rect 19208 28432 19214 28444
rect 15252 28376 16068 28404
rect 17405 28407 17463 28413
rect 15252 28364 15258 28376
rect 17405 28373 17417 28407
rect 17451 28404 17463 28407
rect 18046 28404 18052 28416
rect 17451 28376 18052 28404
rect 17451 28373 17463 28376
rect 17405 28367 17463 28373
rect 18046 28364 18052 28376
rect 18104 28364 18110 28416
rect 19613 28407 19671 28413
rect 19613 28373 19625 28407
rect 19659 28404 19671 28407
rect 19978 28404 19984 28416
rect 19659 28376 19984 28404
rect 19659 28373 19671 28376
rect 19613 28367 19671 28373
rect 19978 28364 19984 28376
rect 20036 28364 20042 28416
rect 20070 28364 20076 28416
rect 20128 28404 20134 28416
rect 20165 28407 20223 28413
rect 20165 28404 20177 28407
rect 20128 28376 20177 28404
rect 20128 28364 20134 28376
rect 20165 28373 20177 28376
rect 20211 28373 20223 28407
rect 20165 28367 20223 28373
rect 20438 28364 20444 28416
rect 20496 28364 20502 28416
rect 1104 28314 21043 28336
rect 1104 28262 5894 28314
rect 5946 28262 5958 28314
rect 6010 28262 6022 28314
rect 6074 28262 6086 28314
rect 6138 28262 6150 28314
rect 6202 28262 10839 28314
rect 10891 28262 10903 28314
rect 10955 28262 10967 28314
rect 11019 28262 11031 28314
rect 11083 28262 11095 28314
rect 11147 28262 15784 28314
rect 15836 28262 15848 28314
rect 15900 28262 15912 28314
rect 15964 28262 15976 28314
rect 16028 28262 16040 28314
rect 16092 28262 20729 28314
rect 20781 28262 20793 28314
rect 20845 28262 20857 28314
rect 20909 28262 20921 28314
rect 20973 28262 20985 28314
rect 21037 28262 21043 28314
rect 1104 28240 21043 28262
rect 1394 28160 1400 28212
rect 1452 28200 1458 28212
rect 2038 28200 2044 28212
rect 1452 28172 2044 28200
rect 1452 28160 1458 28172
rect 2038 28160 2044 28172
rect 2096 28160 2102 28212
rect 2406 28160 2412 28212
rect 2464 28200 2470 28212
rect 4246 28200 4252 28212
rect 2464 28172 4252 28200
rect 2464 28160 2470 28172
rect 4246 28160 4252 28172
rect 4304 28160 4310 28212
rect 5902 28160 5908 28212
rect 5960 28200 5966 28212
rect 6546 28200 6552 28212
rect 5960 28172 6552 28200
rect 5960 28160 5966 28172
rect 6546 28160 6552 28172
rect 6604 28160 6610 28212
rect 8662 28160 8668 28212
rect 8720 28200 8726 28212
rect 9953 28203 10011 28209
rect 9953 28200 9965 28203
rect 8720 28172 9965 28200
rect 8720 28160 8726 28172
rect 9953 28169 9965 28172
rect 9999 28169 10011 28203
rect 15286 28200 15292 28212
rect 9953 28163 10011 28169
rect 10058 28172 13216 28200
rect 290 28092 296 28144
rect 348 28092 354 28144
rect 1302 28092 1308 28144
rect 1360 28132 1366 28144
rect 2869 28135 2927 28141
rect 2869 28132 2881 28135
rect 1360 28104 2881 28132
rect 1360 28092 1366 28104
rect 2869 28101 2881 28104
rect 2915 28101 2927 28135
rect 2869 28095 2927 28101
rect 3970 28092 3976 28144
rect 4028 28092 4034 28144
rect 5074 28092 5080 28144
rect 5132 28092 5138 28144
rect 5350 28092 5356 28144
rect 5408 28132 5414 28144
rect 8202 28132 8208 28144
rect 5408 28104 8208 28132
rect 5408 28092 5414 28104
rect 8202 28092 8208 28104
rect 8260 28092 8266 28144
rect 8956 28104 9352 28132
rect 308 28064 336 28092
rect 1639 28067 1697 28073
rect 1639 28064 1651 28067
rect 308 28036 1651 28064
rect 1639 28033 1651 28036
rect 1685 28064 1697 28067
rect 2038 28064 2044 28076
rect 1685 28036 2044 28064
rect 1685 28033 1697 28036
rect 1639 28027 1697 28033
rect 2038 28024 2044 28036
rect 2096 28024 2102 28076
rect 3050 28024 3056 28076
rect 3108 28064 3114 28076
rect 3419 28067 3477 28073
rect 3108 28036 3188 28064
rect 3108 28024 3114 28036
rect 750 27956 756 28008
rect 808 27996 814 28008
rect 1394 27996 1400 28008
rect 808 27968 1400 27996
rect 808 27956 814 27968
rect 1394 27956 1400 27968
rect 1452 27956 1458 28008
rect 3160 28005 3188 28036
rect 3419 28033 3431 28067
rect 3465 28064 3477 28067
rect 3988 28064 4016 28092
rect 4798 28064 4804 28076
rect 3465 28036 4016 28064
rect 4759 28036 4804 28064
rect 3465 28033 3477 28036
rect 3419 28027 3477 28033
rect 4798 28024 4804 28036
rect 4856 28024 4862 28076
rect 5092 28064 5120 28092
rect 5092 28036 5580 28064
rect 3145 27999 3203 28005
rect 3145 27965 3157 27999
rect 3191 27965 3203 27999
rect 3145 27959 3203 27965
rect 3050 27888 3056 27940
rect 3108 27888 3114 27940
rect 1026 27820 1032 27872
rect 1084 27820 1090 27872
rect 2406 27820 2412 27872
rect 2464 27820 2470 27872
rect 3160 27860 3188 27959
rect 4522 27956 4528 28008
rect 4580 27956 4586 28008
rect 5552 27937 5580 28036
rect 8956 28008 8984 28104
rect 9122 28024 9128 28076
rect 9180 28064 9186 28076
rect 9215 28067 9273 28073
rect 9215 28064 9227 28067
rect 9180 28036 9227 28064
rect 9180 28024 9186 28036
rect 9215 28033 9227 28036
rect 9261 28033 9273 28067
rect 9324 28064 9352 28104
rect 9398 28092 9404 28144
rect 9456 28132 9462 28144
rect 10058 28132 10086 28172
rect 9456 28104 10086 28132
rect 9456 28092 9462 28104
rect 10318 28092 10324 28144
rect 10376 28132 10382 28144
rect 10778 28132 10784 28144
rect 10376 28104 10784 28132
rect 10376 28092 10382 28104
rect 10778 28092 10784 28104
rect 10836 28092 10842 28144
rect 10870 28092 10876 28144
rect 10928 28132 10934 28144
rect 11606 28132 11612 28144
rect 10928 28104 11612 28132
rect 10928 28092 10934 28104
rect 11606 28092 11612 28104
rect 11664 28092 11670 28144
rect 11698 28092 11704 28144
rect 11756 28092 11762 28144
rect 13188 28132 13216 28172
rect 13464 28172 15292 28200
rect 13464 28132 13492 28172
rect 15286 28160 15292 28172
rect 15344 28160 15350 28212
rect 16301 28203 16359 28209
rect 16301 28169 16313 28203
rect 16347 28169 16359 28203
rect 16301 28163 16359 28169
rect 13188 28104 13492 28132
rect 16316 28132 16344 28163
rect 17954 28160 17960 28212
rect 18012 28200 18018 28212
rect 19426 28200 19432 28212
rect 18012 28172 19432 28200
rect 18012 28160 18018 28172
rect 19426 28160 19432 28172
rect 19484 28160 19490 28212
rect 19521 28203 19579 28209
rect 19521 28169 19533 28203
rect 19567 28200 19579 28203
rect 19702 28200 19708 28212
rect 19567 28172 19708 28200
rect 19567 28169 19579 28172
rect 19521 28163 19579 28169
rect 19702 28160 19708 28172
rect 19760 28160 19766 28212
rect 16316 28104 18092 28132
rect 11716 28064 11744 28092
rect 9324 28036 11744 28064
rect 9215 28027 9273 28033
rect 12710 28024 12716 28076
rect 12768 28024 12774 28076
rect 14182 28064 14188 28076
rect 13280 28036 14188 28064
rect 7282 27956 7288 28008
rect 7340 27996 7346 28008
rect 7650 27996 7656 28008
rect 7340 27968 7656 27996
rect 7340 27956 7346 27968
rect 7650 27956 7656 27968
rect 7708 27956 7714 28008
rect 8938 27956 8944 28008
rect 8996 27956 9002 28008
rect 11517 27999 11575 28005
rect 11517 27965 11529 27999
rect 11563 27996 11575 27999
rect 11606 27996 11612 28008
rect 11563 27968 11612 27996
rect 11563 27965 11575 27968
rect 11517 27959 11575 27965
rect 11606 27956 11612 27968
rect 11664 27956 11670 28008
rect 11698 27956 11704 28008
rect 11756 27956 11762 28008
rect 12161 27999 12219 28005
rect 12161 27965 12173 27999
rect 12207 27996 12219 27999
rect 12250 27996 12256 28008
rect 12207 27968 12256 27996
rect 12207 27965 12219 27968
rect 12161 27959 12219 27965
rect 12250 27956 12256 27968
rect 12308 27956 12314 28008
rect 12434 27956 12440 28008
rect 12492 27956 12498 28008
rect 12575 27999 12633 28005
rect 12575 27965 12587 27999
rect 12621 27996 12633 27999
rect 12894 27996 12900 28008
rect 12621 27968 12900 27996
rect 12621 27965 12633 27968
rect 12575 27959 12633 27965
rect 12894 27956 12900 27968
rect 12952 27996 12958 28008
rect 13280 27996 13308 28036
rect 14182 28024 14188 28036
rect 14240 28024 14246 28076
rect 14274 28024 14280 28076
rect 14332 28024 14338 28076
rect 15286 28024 15292 28076
rect 15344 28073 15350 28076
rect 15344 28067 15372 28073
rect 15360 28033 15372 28067
rect 15344 28027 15372 28033
rect 16117 28067 16175 28073
rect 16117 28033 16129 28067
rect 16163 28064 16175 28067
rect 16298 28064 16304 28076
rect 16163 28036 16304 28064
rect 16163 28033 16175 28036
rect 16117 28027 16175 28033
rect 15344 28024 15350 28027
rect 16298 28024 16304 28036
rect 16356 28064 16362 28076
rect 16485 28067 16543 28073
rect 16485 28064 16497 28067
rect 16356 28036 16497 28064
rect 16356 28024 16362 28036
rect 16485 28033 16497 28036
rect 16531 28033 16543 28067
rect 16485 28027 16543 28033
rect 16850 28024 16856 28076
rect 16908 28064 16914 28076
rect 18064 28073 18092 28104
rect 18782 28103 18788 28144
rect 18767 28097 18788 28103
rect 16943 28067 17001 28073
rect 16943 28064 16955 28067
rect 16908 28036 16955 28064
rect 16908 28024 16914 28036
rect 16943 28033 16955 28036
rect 16989 28064 17001 28067
rect 18049 28067 18107 28073
rect 16989 28036 17908 28064
rect 16989 28033 17001 28036
rect 16943 28027 17001 28033
rect 17880 28008 17908 28036
rect 18049 28033 18061 28067
rect 18095 28033 18107 28067
rect 18767 28063 18779 28097
rect 18840 28092 18846 28144
rect 19058 28092 19064 28144
rect 19116 28132 19122 28144
rect 19610 28132 19616 28144
rect 19116 28104 19616 28132
rect 19116 28092 19122 28104
rect 19610 28092 19616 28104
rect 19668 28092 19674 28144
rect 19794 28092 19800 28144
rect 19852 28132 19858 28144
rect 20165 28135 20223 28141
rect 20165 28132 20177 28135
rect 19852 28104 20177 28132
rect 19852 28092 19858 28104
rect 20165 28101 20177 28104
rect 20211 28101 20223 28135
rect 20165 28095 20223 28101
rect 18813 28066 18828 28092
rect 18813 28063 18825 28066
rect 18767 28057 18825 28063
rect 18049 28027 18107 28033
rect 18874 28024 18880 28076
rect 18932 28064 18938 28076
rect 20622 28064 20628 28076
rect 18932 28036 20628 28064
rect 18932 28024 18938 28036
rect 20622 28024 20628 28036
rect 20680 28024 20686 28076
rect 14366 27996 14372 28008
rect 12952 27968 13308 27996
rect 13924 27968 14372 27996
rect 12952 27956 12958 27968
rect 5537 27931 5595 27937
rect 3802 27900 4288 27928
rect 3802 27860 3830 27900
rect 3160 27832 3830 27860
rect 4154 27820 4160 27872
rect 4212 27820 4218 27872
rect 4260 27860 4288 27900
rect 5537 27897 5549 27931
rect 5583 27897 5595 27931
rect 5537 27891 5595 27897
rect 13170 27888 13176 27940
rect 13228 27928 13234 27940
rect 13357 27931 13415 27937
rect 13357 27928 13369 27931
rect 13228 27900 13369 27928
rect 13228 27888 13234 27900
rect 13357 27897 13369 27900
rect 13403 27897 13415 27931
rect 13357 27891 13415 27897
rect 13924 27872 13952 27968
rect 14366 27956 14372 27968
rect 14424 27996 14430 28008
rect 14461 27999 14519 28005
rect 14461 27996 14473 27999
rect 14424 27968 14473 27996
rect 14424 27956 14430 27968
rect 14461 27965 14473 27968
rect 14507 27965 14519 27999
rect 14461 27959 14519 27965
rect 14642 27956 14648 28008
rect 14700 27996 14706 28008
rect 14921 27999 14979 28005
rect 14921 27996 14933 27999
rect 14700 27968 14933 27996
rect 14700 27956 14706 27968
rect 14921 27965 14933 27968
rect 14967 27965 14979 27999
rect 15197 27999 15255 28005
rect 15197 27996 15209 27999
rect 14921 27959 14979 27965
rect 15028 27968 15209 27996
rect 15028 27928 15056 27968
rect 15197 27965 15209 27968
rect 15243 27965 15255 27999
rect 15197 27959 15255 27965
rect 15470 27956 15476 28008
rect 15528 27956 15534 28008
rect 16669 27999 16727 28005
rect 16669 27965 16681 27999
rect 16715 27965 16727 27999
rect 16669 27959 16727 27965
rect 14476 27900 15056 27928
rect 14476 27872 14504 27900
rect 6822 27860 6828 27872
rect 4260 27832 6828 27860
rect 6822 27820 6828 27832
rect 6880 27820 6886 27872
rect 7282 27820 7288 27872
rect 7340 27860 7346 27872
rect 13078 27860 13084 27872
rect 7340 27832 13084 27860
rect 7340 27820 7346 27832
rect 13078 27820 13084 27832
rect 13136 27820 13142 27872
rect 13906 27820 13912 27872
rect 13964 27820 13970 27872
rect 14458 27820 14464 27872
rect 14516 27820 14522 27872
rect 16684 27860 16712 27959
rect 17862 27956 17868 28008
rect 17920 27956 17926 28008
rect 18509 27999 18567 28005
rect 18509 27965 18521 27999
rect 18555 27965 18567 27999
rect 18509 27959 18567 27965
rect 18524 27928 18552 27959
rect 17512 27900 18552 27928
rect 17126 27860 17132 27872
rect 16684 27832 17132 27860
rect 17126 27820 17132 27832
rect 17184 27860 17190 27872
rect 17512 27860 17540 27900
rect 17184 27832 17540 27860
rect 17184 27820 17190 27832
rect 17586 27820 17592 27872
rect 17644 27860 17650 27872
rect 17681 27863 17739 27869
rect 17681 27860 17693 27863
rect 17644 27832 17693 27860
rect 17644 27820 17650 27832
rect 17681 27829 17693 27832
rect 17727 27829 17739 27863
rect 17681 27823 17739 27829
rect 17770 27820 17776 27872
rect 17828 27860 17834 27872
rect 18141 27863 18199 27869
rect 18141 27860 18153 27863
rect 17828 27832 18153 27860
rect 17828 27820 17834 27832
rect 18141 27829 18153 27832
rect 18187 27829 18199 27863
rect 18141 27823 18199 27829
rect 20438 27820 20444 27872
rect 20496 27820 20502 27872
rect 1044 27600 1072 27820
rect 1104 27770 20884 27792
rect 1104 27718 3422 27770
rect 3474 27718 3486 27770
rect 3538 27718 3550 27770
rect 3602 27718 3614 27770
rect 3666 27718 3678 27770
rect 3730 27718 8367 27770
rect 8419 27718 8431 27770
rect 8483 27718 8495 27770
rect 8547 27718 8559 27770
rect 8611 27718 8623 27770
rect 8675 27718 13312 27770
rect 13364 27718 13376 27770
rect 13428 27718 13440 27770
rect 13492 27718 13504 27770
rect 13556 27718 13568 27770
rect 13620 27718 18257 27770
rect 18309 27718 18321 27770
rect 18373 27718 18385 27770
rect 18437 27718 18449 27770
rect 18501 27718 18513 27770
rect 18565 27718 20884 27770
rect 1104 27696 20884 27718
rect 3050 27616 3056 27668
rect 3108 27656 3114 27668
rect 3145 27659 3203 27665
rect 3145 27656 3157 27659
rect 3108 27628 3157 27656
rect 3108 27616 3114 27628
rect 3145 27625 3157 27628
rect 3191 27625 3203 27659
rect 3145 27619 3203 27625
rect 6840 27628 7510 27656
rect 1026 27548 1032 27600
rect 1084 27548 1090 27600
rect 2406 27480 2412 27532
rect 2464 27480 2470 27532
rect 2958 27480 2964 27532
rect 3016 27520 3022 27532
rect 3694 27520 3700 27532
rect 3016 27492 3700 27520
rect 3016 27480 3022 27492
rect 3694 27480 3700 27492
rect 3752 27480 3758 27532
rect 4982 27480 4988 27532
rect 5040 27480 5046 27532
rect 6840 27464 6868 27628
rect 7482 27588 7510 27628
rect 7834 27616 7840 27668
rect 7892 27616 7898 27668
rect 7944 27628 9674 27656
rect 7944 27588 7972 27628
rect 7482 27560 7972 27588
rect 8110 27480 8116 27532
rect 8168 27520 8174 27532
rect 9646 27520 9674 27628
rect 10318 27616 10324 27668
rect 10376 27656 10382 27668
rect 11514 27656 11520 27668
rect 10376 27628 11520 27656
rect 10376 27616 10382 27628
rect 11514 27616 11520 27628
rect 11572 27616 11578 27668
rect 12250 27616 12256 27668
rect 12308 27656 12314 27668
rect 13170 27656 13176 27668
rect 12308 27628 13176 27656
rect 12308 27616 12314 27628
rect 13170 27616 13176 27628
rect 13228 27616 13234 27668
rect 14182 27616 14188 27668
rect 14240 27616 14246 27668
rect 15470 27616 15476 27668
rect 15528 27656 15534 27668
rect 16485 27659 16543 27665
rect 16485 27656 16497 27659
rect 15528 27628 16497 27656
rect 15528 27616 15534 27628
rect 16485 27625 16497 27628
rect 16531 27625 16543 27659
rect 16485 27619 16543 27625
rect 17770 27616 17776 27668
rect 17828 27616 17834 27668
rect 19886 27656 19892 27668
rect 18524 27628 18736 27656
rect 10502 27548 10508 27600
rect 10560 27588 10566 27600
rect 12710 27588 12716 27600
rect 10560 27560 12716 27588
rect 10560 27548 10566 27560
rect 12710 27548 12716 27560
rect 12768 27548 12774 27600
rect 13909 27591 13967 27597
rect 13909 27557 13921 27591
rect 13955 27588 13967 27591
rect 14200 27588 14228 27616
rect 13955 27560 14228 27588
rect 17313 27591 17371 27597
rect 13955 27557 13967 27560
rect 13909 27551 13967 27557
rect 17313 27557 17325 27591
rect 17359 27588 17371 27591
rect 17788 27588 17816 27616
rect 17359 27560 17816 27588
rect 17359 27557 17371 27560
rect 17313 27551 17371 27557
rect 18046 27548 18052 27600
rect 18104 27548 18110 27600
rect 18141 27591 18199 27597
rect 18141 27557 18153 27591
rect 18187 27588 18199 27591
rect 18524 27588 18552 27628
rect 18187 27560 18552 27588
rect 18601 27591 18659 27597
rect 18187 27557 18199 27560
rect 18141 27551 18199 27557
rect 18601 27557 18613 27591
rect 18647 27557 18659 27591
rect 18708 27588 18736 27628
rect 19260 27628 19892 27656
rect 19260 27597 19288 27628
rect 19886 27616 19892 27628
rect 19944 27616 19950 27668
rect 21266 27616 21272 27668
rect 21324 27656 21330 27668
rect 21818 27656 21824 27668
rect 21324 27628 21824 27656
rect 21324 27616 21330 27628
rect 21818 27616 21824 27628
rect 21876 27616 21882 27668
rect 19245 27591 19303 27597
rect 18708 27560 19196 27588
rect 18601 27551 18659 27557
rect 13630 27520 13636 27532
rect 8168 27492 8708 27520
rect 9646 27492 13636 27520
rect 8168 27480 8174 27492
rect 8680 27464 8708 27492
rect 12544 27464 12572 27492
rect 13630 27480 13636 27492
rect 13688 27520 13694 27532
rect 14093 27523 14151 27529
rect 14093 27520 14105 27523
rect 13688 27492 14105 27520
rect 13688 27480 13694 27492
rect 14093 27489 14105 27492
rect 14139 27489 14151 27523
rect 14093 27483 14151 27489
rect 15470 27480 15476 27532
rect 15528 27480 15534 27532
rect 17497 27523 17555 27529
rect 17497 27489 17509 27523
rect 17543 27520 17555 27523
rect 17681 27523 17739 27529
rect 17681 27520 17693 27523
rect 17543 27492 17693 27520
rect 17543 27489 17555 27492
rect 17497 27483 17555 27489
rect 17681 27489 17693 27492
rect 17727 27489 17739 27523
rect 17681 27483 17739 27489
rect 1394 27412 1400 27464
rect 1452 27412 1458 27464
rect 3789 27455 3847 27461
rect 3789 27452 3801 27455
rect 1504 27424 3801 27452
rect 1118 27344 1124 27396
rect 1176 27384 1182 27396
rect 1504 27384 1532 27424
rect 3789 27421 3801 27424
rect 3835 27421 3847 27455
rect 3789 27415 3847 27421
rect 4065 27455 4123 27461
rect 4065 27421 4077 27455
rect 4111 27452 4123 27455
rect 4614 27452 4620 27464
rect 4111 27424 4620 27452
rect 4111 27421 4123 27424
rect 4065 27415 4123 27421
rect 4614 27412 4620 27424
rect 4672 27412 4678 27464
rect 4893 27455 4951 27461
rect 4893 27421 4905 27455
rect 4939 27452 4951 27455
rect 5074 27452 5080 27464
rect 4939 27424 5080 27452
rect 4939 27421 4951 27424
rect 4893 27415 4951 27421
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 5810 27452 5816 27464
rect 5184 27424 5816 27452
rect 1176 27356 1532 27384
rect 1176 27344 1182 27356
rect 1946 27344 1952 27396
rect 2004 27384 2010 27396
rect 2133 27387 2191 27393
rect 2133 27384 2145 27387
rect 2004 27356 2145 27384
rect 2004 27344 2010 27356
rect 2133 27353 2145 27356
rect 2179 27353 2191 27387
rect 2133 27347 2191 27353
rect 2222 27344 2228 27396
rect 2280 27344 2286 27396
rect 2314 27344 2320 27396
rect 2372 27384 2378 27396
rect 2593 27387 2651 27393
rect 2593 27384 2605 27387
rect 2372 27356 2605 27384
rect 2372 27344 2378 27356
rect 2593 27353 2605 27356
rect 2639 27353 2651 27387
rect 4801 27387 4859 27393
rect 2593 27347 2651 27353
rect 2746 27356 4752 27384
rect 1578 27276 1584 27328
rect 1636 27276 1642 27328
rect 1857 27319 1915 27325
rect 1857 27285 1869 27319
rect 1903 27316 1915 27319
rect 2746 27316 2774 27356
rect 4724 27328 4752 27356
rect 4801 27353 4813 27387
rect 4847 27384 4859 27387
rect 5184 27384 5212 27424
rect 5810 27412 5816 27424
rect 5868 27452 5874 27464
rect 6362 27452 6368 27464
rect 5868 27424 6368 27452
rect 5868 27412 5874 27424
rect 6362 27412 6368 27424
rect 6420 27412 6426 27464
rect 6822 27412 6828 27464
rect 6880 27412 6886 27464
rect 7098 27452 7104 27464
rect 7059 27424 7104 27452
rect 7098 27412 7104 27424
rect 7156 27412 7162 27464
rect 8386 27412 8392 27464
rect 8444 27412 8450 27464
rect 8662 27412 8668 27464
rect 8720 27452 8726 27464
rect 8941 27455 8999 27461
rect 8941 27452 8953 27455
rect 8720 27424 8953 27452
rect 8720 27412 8726 27424
rect 8941 27421 8953 27424
rect 8987 27421 8999 27455
rect 8941 27415 8999 27421
rect 9122 27412 9128 27464
rect 9180 27452 9186 27464
rect 9215 27455 9273 27461
rect 9215 27452 9227 27455
rect 9180 27424 9227 27452
rect 9180 27412 9186 27424
rect 9215 27421 9227 27424
rect 9261 27421 9273 27455
rect 9215 27415 9273 27421
rect 9324 27424 10456 27452
rect 4847 27356 5212 27384
rect 5261 27387 5319 27393
rect 4847 27353 4859 27356
rect 4801 27347 4859 27353
rect 5261 27353 5273 27387
rect 5307 27353 5319 27387
rect 9324 27384 9352 27424
rect 5261 27347 5319 27353
rect 5828 27356 9352 27384
rect 10428 27384 10456 27424
rect 10778 27412 10784 27464
rect 10836 27452 10842 27464
rect 11514 27452 11520 27464
rect 10836 27424 11520 27452
rect 10836 27412 10842 27424
rect 11514 27412 11520 27424
rect 11572 27452 11578 27464
rect 12066 27452 12072 27464
rect 11572 27424 12072 27452
rect 11572 27412 11578 27424
rect 12066 27412 12072 27424
rect 12124 27412 12130 27464
rect 12526 27412 12532 27464
rect 12584 27412 12590 27464
rect 14335 27455 14393 27461
rect 14335 27452 14347 27455
rect 12634 27424 14347 27452
rect 12250 27384 12256 27396
rect 10428 27356 12256 27384
rect 1903 27288 2774 27316
rect 1903 27285 1915 27288
rect 1857 27279 1915 27285
rect 2958 27276 2964 27328
rect 3016 27276 3022 27328
rect 3973 27319 4031 27325
rect 3973 27285 3985 27319
rect 4019 27316 4031 27319
rect 4062 27316 4068 27328
rect 4019 27288 4068 27316
rect 4019 27285 4031 27288
rect 3973 27279 4031 27285
rect 4062 27276 4068 27288
rect 4120 27276 4126 27328
rect 4249 27319 4307 27325
rect 4249 27285 4261 27319
rect 4295 27316 4307 27319
rect 4430 27316 4436 27328
rect 4295 27288 4436 27316
rect 4295 27285 4307 27288
rect 4249 27279 4307 27285
rect 4430 27276 4436 27288
rect 4488 27316 4494 27328
rect 4525 27319 4583 27325
rect 4525 27316 4537 27319
rect 4488 27288 4537 27316
rect 4488 27276 4494 27288
rect 4525 27285 4537 27288
rect 4571 27285 4583 27319
rect 4525 27279 4583 27285
rect 4706 27276 4712 27328
rect 4764 27276 4770 27328
rect 4890 27276 4896 27328
rect 4948 27316 4954 27328
rect 5276 27316 5304 27347
rect 4948 27288 5304 27316
rect 4948 27276 4954 27288
rect 5350 27276 5356 27328
rect 5408 27316 5414 27328
rect 5828 27325 5856 27356
rect 12250 27344 12256 27356
rect 12308 27344 12314 27396
rect 5629 27319 5687 27325
rect 5629 27316 5641 27319
rect 5408 27288 5641 27316
rect 5408 27276 5414 27288
rect 5629 27285 5641 27288
rect 5675 27285 5687 27319
rect 5629 27279 5687 27285
rect 5813 27319 5871 27325
rect 5813 27285 5825 27319
rect 5859 27285 5871 27319
rect 5813 27279 5871 27285
rect 8294 27276 8300 27328
rect 8352 27316 8358 27328
rect 9953 27319 10011 27325
rect 9953 27316 9965 27319
rect 8352 27288 9965 27316
rect 8352 27276 8358 27288
rect 9953 27285 9965 27288
rect 9999 27285 10011 27319
rect 9953 27279 10011 27285
rect 11974 27276 11980 27328
rect 12032 27316 12038 27328
rect 12158 27316 12164 27328
rect 12032 27288 12164 27316
rect 12032 27276 12038 27288
rect 12158 27276 12164 27288
rect 12216 27316 12222 27328
rect 12634 27316 12662 27424
rect 14335 27421 14347 27424
rect 14381 27421 14393 27455
rect 14335 27415 14393 27421
rect 15715 27455 15773 27461
rect 15715 27421 15727 27455
rect 15761 27421 15773 27455
rect 15715 27415 15773 27421
rect 14350 27384 14378 27415
rect 15730 27384 15758 27415
rect 16942 27412 16948 27464
rect 17000 27412 17006 27464
rect 17221 27455 17279 27461
rect 17221 27421 17233 27455
rect 17267 27421 17279 27455
rect 17221 27415 17279 27421
rect 16298 27384 16304 27396
rect 14350 27356 16304 27384
rect 16298 27344 16304 27356
rect 16356 27344 16362 27396
rect 17236 27384 17264 27415
rect 17586 27412 17592 27464
rect 17644 27412 17650 27464
rect 18064 27461 18092 27548
rect 18616 27520 18644 27551
rect 18616 27492 19104 27520
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27452 17831 27455
rect 18049 27455 18107 27461
rect 17819 27424 17908 27452
rect 17819 27421 17831 27424
rect 17773 27415 17831 27421
rect 17604 27384 17632 27412
rect 17236 27356 17632 27384
rect 12216 27288 12662 27316
rect 12216 27276 12222 27288
rect 14182 27276 14188 27328
rect 14240 27316 14246 27328
rect 15105 27319 15163 27325
rect 15105 27316 15117 27319
rect 14240 27288 15117 27316
rect 14240 27276 14246 27288
rect 15105 27285 15117 27288
rect 15151 27285 15163 27319
rect 15105 27279 15163 27285
rect 17034 27276 17040 27328
rect 17092 27276 17098 27328
rect 17497 27319 17555 27325
rect 17497 27285 17509 27319
rect 17543 27316 17555 27319
rect 17770 27316 17776 27328
rect 17543 27288 17776 27316
rect 17543 27285 17555 27288
rect 17497 27279 17555 27285
rect 17770 27276 17776 27288
rect 17828 27276 17834 27328
rect 17880 27325 17908 27424
rect 18049 27421 18061 27455
rect 18095 27421 18107 27455
rect 18049 27415 18107 27421
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 17865 27319 17923 27325
rect 17865 27285 17877 27319
rect 17911 27285 17923 27319
rect 17865 27279 17923 27285
rect 18046 27276 18052 27328
rect 18104 27316 18110 27328
rect 18340 27316 18368 27415
rect 18782 27412 18788 27464
rect 18840 27412 18846 27464
rect 19076 27461 19104 27492
rect 19061 27455 19119 27461
rect 19061 27421 19073 27455
rect 19107 27421 19119 27455
rect 19168 27452 19196 27560
rect 19245 27557 19257 27591
rect 19291 27557 19303 27591
rect 19245 27551 19303 27557
rect 19889 27523 19947 27529
rect 19889 27489 19901 27523
rect 19935 27520 19947 27523
rect 21266 27520 21272 27532
rect 19935 27492 21272 27520
rect 19935 27489 19947 27492
rect 19889 27483 19947 27489
rect 21266 27480 21272 27492
rect 21324 27480 21330 27532
rect 19429 27455 19487 27461
rect 19429 27452 19441 27455
rect 19168 27424 19441 27452
rect 19061 27415 19119 27421
rect 19429 27421 19441 27424
rect 19475 27421 19487 27455
rect 19429 27415 19487 27421
rect 19978 27412 19984 27464
rect 20036 27452 20042 27464
rect 20165 27455 20223 27461
rect 20165 27452 20177 27455
rect 20036 27424 20177 27452
rect 20036 27412 20042 27424
rect 20165 27421 20177 27424
rect 20211 27421 20223 27455
rect 20165 27415 20223 27421
rect 19613 27387 19671 27393
rect 19613 27384 19625 27387
rect 18892 27356 19625 27384
rect 18892 27325 18920 27356
rect 19613 27353 19625 27356
rect 19659 27353 19671 27387
rect 19613 27347 19671 27353
rect 20530 27344 20536 27396
rect 20588 27344 20594 27396
rect 18104 27288 18368 27316
rect 18877 27319 18935 27325
rect 18104 27276 18110 27288
rect 18877 27285 18889 27319
rect 18923 27285 18935 27319
rect 18877 27279 18935 27285
rect 1104 27226 21043 27248
rect 1104 27174 5894 27226
rect 5946 27174 5958 27226
rect 6010 27174 6022 27226
rect 6074 27174 6086 27226
rect 6138 27174 6150 27226
rect 6202 27174 10839 27226
rect 10891 27174 10903 27226
rect 10955 27174 10967 27226
rect 11019 27174 11031 27226
rect 11083 27174 11095 27226
rect 11147 27174 15784 27226
rect 15836 27174 15848 27226
rect 15900 27174 15912 27226
rect 15964 27174 15976 27226
rect 16028 27174 16040 27226
rect 16092 27174 20729 27226
rect 20781 27174 20793 27226
rect 20845 27174 20857 27226
rect 20909 27174 20921 27226
rect 20973 27174 20985 27226
rect 21037 27174 21043 27226
rect 1104 27152 21043 27174
rect 2222 27072 2228 27124
rect 2280 27112 2286 27124
rect 2593 27115 2651 27121
rect 2593 27112 2605 27115
rect 2280 27084 2605 27112
rect 2280 27072 2286 27084
rect 2593 27081 2605 27084
rect 2639 27081 2651 27115
rect 2593 27075 2651 27081
rect 3421 27115 3479 27121
rect 3421 27081 3433 27115
rect 3467 27112 3479 27115
rect 6730 27112 6736 27124
rect 3467 27084 6736 27112
rect 3467 27081 3479 27084
rect 3421 27075 3479 27081
rect 6730 27072 6736 27084
rect 6788 27072 6794 27124
rect 8386 27112 8392 27124
rect 7484 27084 8392 27112
rect 1302 27004 1308 27056
rect 1360 27044 1366 27056
rect 1360 27016 3556 27044
rect 1360 27004 1366 27016
rect 750 26936 756 26988
rect 808 26936 814 26988
rect 1855 26979 1913 26985
rect 1855 26945 1867 26979
rect 1901 26976 1913 26979
rect 2406 26976 2412 26988
rect 1901 26948 2412 26976
rect 1901 26945 1913 26948
rect 1855 26939 1913 26945
rect 2406 26936 2412 26948
rect 2464 26936 2470 26988
rect 2961 26979 3019 26985
rect 2961 26976 2973 26979
rect 2746 26948 2973 26976
rect 768 26908 796 26936
rect 1581 26911 1639 26917
rect 1581 26908 1593 26911
rect 768 26880 1593 26908
rect 1581 26877 1593 26880
rect 1627 26877 1639 26911
rect 1581 26871 1639 26877
rect 1210 26732 1216 26784
rect 1268 26772 1274 26784
rect 2746 26772 2774 26948
rect 2961 26945 2973 26948
rect 3007 26945 3019 26979
rect 2961 26939 3019 26945
rect 3234 26936 3240 26988
rect 3292 26936 3298 26988
rect 3528 26985 3556 27016
rect 3602 27004 3608 27056
rect 3660 27044 3666 27056
rect 4065 27047 4123 27053
rect 4065 27044 4077 27047
rect 3660 27016 4077 27044
rect 3660 27004 3666 27016
rect 4065 27013 4077 27016
rect 4111 27013 4123 27047
rect 4065 27007 4123 27013
rect 4154 27004 4160 27056
rect 4212 27044 4218 27056
rect 4433 27047 4491 27053
rect 4433 27044 4445 27047
rect 4212 27016 4445 27044
rect 4212 27004 4218 27016
rect 4433 27013 4445 27016
rect 4479 27013 4491 27047
rect 5442 27044 5448 27056
rect 4433 27007 4491 27013
rect 4724 27016 5448 27044
rect 3513 26979 3571 26985
rect 3513 26945 3525 26979
rect 3559 26945 3571 26979
rect 3513 26939 3571 26945
rect 4341 26979 4399 26985
rect 4341 26945 4353 26979
rect 4387 26976 4399 26979
rect 4724 26976 4752 27016
rect 5442 27004 5448 27016
rect 5500 27044 5506 27056
rect 5500 27016 5856 27044
rect 5500 27004 5506 27016
rect 5828 26988 5856 27016
rect 6914 27004 6920 27056
rect 6972 27044 6978 27056
rect 7193 27047 7251 27053
rect 7193 27044 7205 27047
rect 6972 27016 7205 27044
rect 6972 27004 6978 27016
rect 7193 27013 7205 27016
rect 7239 27013 7251 27047
rect 7193 27007 7251 27013
rect 4387 26948 4752 26976
rect 4387 26945 4399 26948
rect 4341 26939 4399 26945
rect 4798 26936 4804 26988
rect 4856 26936 4862 26988
rect 5166 26936 5172 26988
rect 5224 26985 5230 26988
rect 5224 26979 5241 26985
rect 5229 26976 5241 26979
rect 5350 26976 5356 26988
rect 5229 26948 5356 26976
rect 5229 26945 5241 26948
rect 5224 26939 5241 26945
rect 5224 26936 5230 26939
rect 5350 26936 5356 26948
rect 5408 26936 5414 26988
rect 5810 26936 5816 26988
rect 5868 26936 5874 26988
rect 7484 26985 7512 27084
rect 8386 27072 8392 27084
rect 8444 27072 8450 27124
rect 9950 27072 9956 27124
rect 10008 27112 10014 27124
rect 10594 27112 10600 27124
rect 10008 27084 10600 27112
rect 10008 27072 10014 27084
rect 10594 27072 10600 27084
rect 10652 27072 10658 27124
rect 13814 27112 13820 27124
rect 11790 27084 13820 27112
rect 8110 27004 8116 27056
rect 8168 27044 8174 27056
rect 8297 27047 8355 27053
rect 8297 27044 8309 27047
rect 8168 27016 8309 27044
rect 8168 27004 8174 27016
rect 8297 27013 8309 27016
rect 8343 27044 8355 27047
rect 8754 27044 8760 27056
rect 8343 27016 8760 27044
rect 8343 27013 8355 27016
rect 8297 27007 8355 27013
rect 8754 27004 8760 27016
rect 8812 27004 8818 27056
rect 10686 27044 10692 27056
rect 10060 27016 10692 27044
rect 7469 26979 7527 26985
rect 7469 26945 7481 26979
rect 7515 26945 7527 26979
rect 7469 26939 7527 26945
rect 7558 26936 7564 26988
rect 7616 26936 7622 26988
rect 7926 26936 7932 26988
rect 7984 26936 7990 26988
rect 3884 26920 3936 26926
rect 3050 26868 3056 26920
rect 3108 26908 3114 26920
rect 3694 26908 3700 26920
rect 3108 26880 3700 26908
rect 3108 26868 3114 26880
rect 3694 26868 3700 26880
rect 3752 26868 3758 26920
rect 7834 26868 7840 26920
rect 7892 26868 7898 26920
rect 9398 26868 9404 26920
rect 9456 26908 9462 26920
rect 10060 26917 10088 27016
rect 10686 27004 10692 27016
rect 10744 27044 10750 27056
rect 10744 27016 11560 27044
rect 10744 27004 10750 27016
rect 11532 26985 11560 27016
rect 11790 27015 11818 27084
rect 13814 27072 13820 27084
rect 13872 27072 13878 27124
rect 13906 27072 13912 27124
rect 13964 27112 13970 27124
rect 14090 27112 14096 27124
rect 13964 27084 14096 27112
rect 13964 27072 13970 27084
rect 14090 27072 14096 27084
rect 14148 27072 14154 27124
rect 16298 27072 16304 27124
rect 16356 27072 16362 27124
rect 16669 27115 16727 27121
rect 16669 27081 16681 27115
rect 16715 27112 16727 27115
rect 16942 27112 16948 27124
rect 16715 27084 16948 27112
rect 16715 27081 16727 27084
rect 16669 27075 16727 27081
rect 16942 27072 16948 27084
rect 17000 27072 17006 27124
rect 17052 27084 18368 27112
rect 11775 27009 11833 27015
rect 10319 26979 10377 26985
rect 10319 26945 10331 26979
rect 10365 26976 10377 26979
rect 11517 26979 11575 26985
rect 10365 26948 10732 26976
rect 10365 26945 10377 26948
rect 10319 26939 10377 26945
rect 10045 26911 10103 26917
rect 10045 26908 10057 26911
rect 9456 26880 10057 26908
rect 9456 26868 9462 26880
rect 10045 26877 10057 26880
rect 10091 26877 10103 26911
rect 10704 26908 10732 26948
rect 11517 26945 11529 26979
rect 11563 26945 11575 26979
rect 11775 26975 11787 27009
rect 11821 26975 11833 27009
rect 12066 27004 12072 27056
rect 12124 27044 12130 27056
rect 12124 27016 12278 27044
rect 12124 27004 12130 27016
rect 11775 26969 11833 26975
rect 12250 26976 12278 27016
rect 12710 27004 12716 27056
rect 12768 27044 12774 27056
rect 14829 27047 14887 27053
rect 12768 27016 13216 27044
rect 12768 27004 12774 27016
rect 13188 26985 13216 27016
rect 14829 27013 14841 27047
rect 14875 27044 14887 27047
rect 16316 27044 16344 27072
rect 17052 27056 17080 27084
rect 14875 27016 15332 27044
rect 16316 27016 16968 27044
rect 14875 27013 14887 27016
rect 14829 27007 14887 27013
rect 12989 26979 13047 26985
rect 12989 26976 13001 26979
rect 12250 26948 13001 26976
rect 11517 26939 11575 26945
rect 12989 26945 13001 26948
rect 13035 26945 13047 26979
rect 12989 26939 13047 26945
rect 13173 26979 13231 26985
rect 13173 26945 13185 26979
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 13906 26936 13912 26988
rect 13964 26936 13970 26988
rect 14182 26936 14188 26988
rect 14240 26936 14246 26988
rect 15105 26979 15163 26985
rect 15105 26945 15117 26979
rect 15151 26976 15163 26979
rect 15194 26976 15200 26988
rect 15151 26948 15200 26976
rect 15151 26945 15163 26948
rect 15105 26939 15163 26945
rect 15194 26936 15200 26948
rect 15252 26936 15258 26988
rect 15304 26976 15332 27016
rect 15372 26979 15430 26985
rect 15372 26976 15384 26979
rect 15304 26948 15384 26976
rect 15372 26945 15384 26948
rect 15418 26976 15430 26979
rect 16853 26979 16911 26985
rect 16853 26976 16865 26979
rect 15418 26948 16865 26976
rect 15418 26945 15430 26948
rect 15372 26939 15430 26945
rect 16853 26945 16865 26948
rect 16899 26945 16911 26979
rect 16940 26976 16968 27016
rect 17034 27004 17040 27056
rect 17092 27004 17098 27056
rect 18340 27044 18368 27084
rect 18782 27072 18788 27124
rect 18840 27112 18846 27124
rect 18877 27115 18935 27121
rect 18877 27112 18889 27115
rect 18840 27084 18889 27112
rect 18840 27072 18846 27084
rect 18877 27081 18889 27084
rect 18923 27081 18935 27115
rect 18877 27075 18935 27081
rect 18966 27072 18972 27124
rect 19024 27072 19030 27124
rect 19150 27072 19156 27124
rect 19208 27072 19214 27124
rect 19334 27072 19340 27124
rect 19392 27072 19398 27124
rect 19978 27072 19984 27124
rect 20036 27112 20042 27124
rect 21542 27112 21548 27124
rect 20036 27084 21548 27112
rect 20036 27072 20042 27084
rect 21542 27072 21548 27084
rect 21600 27072 21606 27124
rect 18340 27016 18460 27044
rect 17187 26979 17245 26985
rect 17187 26976 17199 26979
rect 16940 26948 17199 26976
rect 16853 26939 16911 26945
rect 17187 26945 17199 26948
rect 17233 26945 17245 26979
rect 17187 26939 17245 26945
rect 17862 26936 17868 26988
rect 17920 26976 17926 26988
rect 18432 26985 18460 27016
rect 18325 26979 18383 26985
rect 18325 26976 18337 26979
rect 17920 26948 18337 26976
rect 17920 26936 17926 26948
rect 18325 26945 18337 26948
rect 18371 26945 18383 26979
rect 18325 26939 18383 26945
rect 18417 26979 18475 26985
rect 18417 26945 18429 26979
rect 18463 26945 18475 26979
rect 18984 26976 19012 27072
rect 19352 27044 19380 27072
rect 20165 27047 20223 27053
rect 20165 27044 20177 27047
rect 19352 27016 20177 27044
rect 20165 27013 20177 27016
rect 20211 27013 20223 27047
rect 20165 27007 20223 27013
rect 19061 26979 19119 26985
rect 19061 26976 19073 26979
rect 18417 26939 18475 26945
rect 18504 26948 19073 26976
rect 10962 26908 10968 26920
rect 10704 26880 10968 26908
rect 10045 26871 10103 26877
rect 10962 26868 10968 26880
rect 11020 26868 11026 26920
rect 12434 26908 12440 26920
rect 12176 26880 12440 26908
rect 3884 26862 3936 26868
rect 3142 26800 3148 26852
rect 3200 26800 3206 26852
rect 5350 26800 5356 26852
rect 5408 26800 5414 26852
rect 10980 26812 11652 26840
rect 10980 26784 11008 26812
rect 1268 26744 2774 26772
rect 3697 26775 3755 26781
rect 1268 26732 1274 26744
rect 3697 26741 3709 26775
rect 3743 26772 3755 26775
rect 4062 26772 4068 26784
rect 3743 26744 4068 26772
rect 3743 26741 3755 26744
rect 3697 26735 3755 26741
rect 4062 26732 4068 26744
rect 4120 26732 4126 26784
rect 8481 26775 8539 26781
rect 8481 26741 8493 26775
rect 8527 26772 8539 26775
rect 10502 26772 10508 26784
rect 8527 26744 10508 26772
rect 8527 26741 8539 26744
rect 8481 26735 8539 26741
rect 10502 26732 10508 26744
rect 10560 26732 10566 26784
rect 10962 26732 10968 26784
rect 11020 26732 11026 26784
rect 11054 26732 11060 26784
rect 11112 26732 11118 26784
rect 11624 26772 11652 26812
rect 12176 26772 12204 26880
rect 12434 26868 12440 26880
rect 12492 26908 12498 26920
rect 14047 26911 14105 26917
rect 14047 26908 14059 26911
rect 12492 26880 14059 26908
rect 12492 26868 12498 26880
rect 14047 26877 14059 26880
rect 14093 26908 14105 26911
rect 14093 26880 14686 26908
rect 14093 26877 14105 26880
rect 14047 26871 14105 26877
rect 12250 26800 12256 26852
rect 12308 26840 12314 26852
rect 12308 26812 13584 26840
rect 12308 26800 12314 26812
rect 11624 26744 12204 26772
rect 12342 26732 12348 26784
rect 12400 26772 12406 26784
rect 12529 26775 12587 26781
rect 12529 26772 12541 26775
rect 12400 26744 12541 26772
rect 12400 26732 12406 26744
rect 12529 26741 12541 26744
rect 12575 26741 12587 26775
rect 13556 26772 13584 26812
rect 13630 26800 13636 26852
rect 13688 26800 13694 26852
rect 14550 26772 14556 26784
rect 13556 26744 14556 26772
rect 12529 26735 12587 26741
rect 14550 26732 14556 26744
rect 14608 26732 14614 26784
rect 14658 26772 14686 26880
rect 16942 26868 16948 26920
rect 17000 26868 17006 26920
rect 18504 26840 18532 26948
rect 19061 26945 19073 26948
rect 19107 26945 19119 26979
rect 19061 26939 19119 26945
rect 19337 26979 19395 26985
rect 19337 26945 19349 26979
rect 19383 26945 19395 26979
rect 19337 26939 19395 26945
rect 19613 26979 19671 26985
rect 19613 26945 19625 26979
rect 19659 26945 19671 26979
rect 19613 26939 19671 26945
rect 18598 26868 18604 26920
rect 18656 26868 18662 26920
rect 18782 26868 18788 26920
rect 18840 26908 18846 26920
rect 19352 26908 19380 26939
rect 18840 26880 19380 26908
rect 18840 26868 18846 26880
rect 17604 26812 18532 26840
rect 15286 26772 15292 26784
rect 14658 26744 15292 26772
rect 15286 26732 15292 26744
rect 15344 26732 15350 26784
rect 16485 26775 16543 26781
rect 16485 26741 16497 26775
rect 16531 26772 16543 26775
rect 17034 26772 17040 26784
rect 16531 26744 17040 26772
rect 16531 26741 16543 26744
rect 16485 26735 16543 26741
rect 17034 26732 17040 26744
rect 17092 26732 17098 26784
rect 17310 26732 17316 26784
rect 17368 26772 17374 26784
rect 17604 26772 17632 26812
rect 19058 26800 19064 26852
rect 19116 26840 19122 26852
rect 19628 26840 19656 26939
rect 21542 26868 21548 26920
rect 21600 26908 21606 26920
rect 21910 26908 21916 26920
rect 21600 26880 21916 26908
rect 21600 26868 21606 26880
rect 21910 26868 21916 26880
rect 21968 26868 21974 26920
rect 19116 26812 19656 26840
rect 19116 26800 19122 26812
rect 17368 26744 17632 26772
rect 17368 26732 17374 26744
rect 17678 26732 17684 26784
rect 17736 26772 17742 26784
rect 17862 26772 17868 26784
rect 17736 26744 17868 26772
rect 17736 26732 17742 26744
rect 17862 26732 17868 26744
rect 17920 26772 17926 26784
rect 17957 26775 18015 26781
rect 17957 26772 17969 26775
rect 17920 26744 17969 26772
rect 17920 26732 17926 26744
rect 17957 26741 17969 26744
rect 18003 26741 18015 26775
rect 17957 26735 18015 26741
rect 18509 26775 18567 26781
rect 18509 26741 18521 26775
rect 18555 26772 18567 26775
rect 19702 26772 19708 26784
rect 18555 26744 19708 26772
rect 18555 26741 18567 26744
rect 18509 26735 18567 26741
rect 19702 26732 19708 26744
rect 19760 26732 19766 26784
rect 19886 26732 19892 26784
rect 19944 26732 19950 26784
rect 20441 26775 20499 26781
rect 20441 26741 20453 26775
rect 20487 26772 20499 26775
rect 20622 26772 20628 26784
rect 20487 26744 20628 26772
rect 20487 26741 20499 26744
rect 20441 26735 20499 26741
rect 20622 26732 20628 26744
rect 20680 26732 20686 26784
rect 1104 26682 20884 26704
rect 1104 26630 3422 26682
rect 3474 26630 3486 26682
rect 3538 26630 3550 26682
rect 3602 26630 3614 26682
rect 3666 26630 3678 26682
rect 3730 26630 8367 26682
rect 8419 26630 8431 26682
rect 8483 26630 8495 26682
rect 8547 26630 8559 26682
rect 8611 26630 8623 26682
rect 8675 26630 13312 26682
rect 13364 26630 13376 26682
rect 13428 26630 13440 26682
rect 13492 26630 13504 26682
rect 13556 26630 13568 26682
rect 13620 26630 18257 26682
rect 18309 26630 18321 26682
rect 18373 26630 18385 26682
rect 18437 26630 18449 26682
rect 18501 26630 18513 26682
rect 18565 26630 20884 26682
rect 1104 26608 20884 26630
rect 1302 26528 1308 26580
rect 1360 26568 1366 26580
rect 3234 26568 3240 26580
rect 1360 26540 3240 26568
rect 1360 26528 1366 26540
rect 3234 26528 3240 26540
rect 3292 26528 3298 26580
rect 3421 26571 3479 26577
rect 3421 26537 3433 26571
rect 3467 26568 3479 26571
rect 4798 26568 4804 26580
rect 3467 26540 4804 26568
rect 3467 26537 3479 26540
rect 3421 26531 3479 26537
rect 4798 26528 4804 26540
rect 4856 26528 4862 26580
rect 4890 26528 4896 26580
rect 4948 26568 4954 26580
rect 5537 26571 5595 26577
rect 5537 26568 5549 26571
rect 4948 26540 5549 26568
rect 4948 26528 4954 26540
rect 5537 26537 5549 26540
rect 5583 26537 5595 26571
rect 5537 26531 5595 26537
rect 7098 26528 7104 26580
rect 7156 26568 7162 26580
rect 7282 26568 7288 26580
rect 7156 26540 7288 26568
rect 7156 26528 7162 26540
rect 7282 26528 7288 26540
rect 7340 26528 7346 26580
rect 7558 26528 7564 26580
rect 7616 26568 7622 26580
rect 8205 26571 8263 26577
rect 8205 26568 8217 26571
rect 7616 26540 8217 26568
rect 7616 26528 7622 26540
rect 8205 26537 8217 26540
rect 8251 26537 8263 26571
rect 8205 26531 8263 26537
rect 9122 26528 9128 26580
rect 9180 26568 9186 26580
rect 10134 26568 10140 26580
rect 9180 26540 10140 26568
rect 9180 26528 9186 26540
rect 10134 26528 10140 26540
rect 10192 26528 10198 26580
rect 13630 26528 13636 26580
rect 13688 26528 13694 26580
rect 14826 26528 14832 26580
rect 14884 26568 14890 26580
rect 17310 26568 17316 26580
rect 14884 26540 17316 26568
rect 14884 26528 14890 26540
rect 17310 26528 17316 26540
rect 17368 26528 17374 26580
rect 17862 26528 17868 26580
rect 17920 26568 17926 26580
rect 18046 26568 18052 26580
rect 17920 26540 18052 26568
rect 17920 26528 17926 26540
rect 18046 26528 18052 26540
rect 18104 26528 18110 26580
rect 18598 26568 18604 26580
rect 18248 26540 18604 26568
rect 3050 26460 3056 26512
rect 3108 26460 3114 26512
rect 3329 26503 3387 26509
rect 3329 26469 3341 26503
rect 3375 26500 3387 26503
rect 3970 26500 3976 26512
rect 3375 26472 3976 26500
rect 3375 26469 3387 26472
rect 3329 26463 3387 26469
rect 3970 26460 3976 26472
rect 4028 26460 4034 26512
rect 5442 26460 5448 26512
rect 5500 26500 5506 26512
rect 7006 26500 7012 26512
rect 5500 26472 7012 26500
rect 5500 26460 5506 26472
rect 7006 26460 7012 26472
rect 7064 26460 7070 26512
rect 11974 26460 11980 26512
rect 12032 26460 12038 26512
rect 3528 26404 4476 26432
rect 1302 26324 1308 26376
rect 1360 26364 1366 26376
rect 1489 26367 1547 26373
rect 1489 26364 1501 26367
rect 1360 26336 1501 26364
rect 1360 26324 1366 26336
rect 1489 26333 1501 26336
rect 1535 26333 1547 26367
rect 1762 26364 1768 26376
rect 1723 26336 1768 26364
rect 1489 26327 1547 26333
rect 1762 26324 1768 26336
rect 1820 26324 1826 26376
rect 2869 26367 2927 26373
rect 2869 26333 2881 26367
rect 2915 26364 2927 26367
rect 3050 26364 3056 26376
rect 2915 26336 3056 26364
rect 2915 26333 2927 26336
rect 2869 26327 2927 26333
rect 3050 26324 3056 26336
rect 3108 26324 3114 26376
rect 3142 26324 3148 26376
rect 3200 26324 3206 26376
rect 3528 26296 3556 26404
rect 3605 26367 3663 26373
rect 3605 26333 3617 26367
rect 3651 26333 3663 26367
rect 3605 26327 3663 26333
rect 1596 26268 3556 26296
rect 1596 26240 1624 26268
rect 3620 26240 3648 26327
rect 4448 26296 4476 26404
rect 6822 26392 6828 26444
rect 6880 26432 6886 26444
rect 7193 26435 7251 26441
rect 7193 26432 7205 26435
rect 6880 26404 7205 26432
rect 6880 26392 6886 26404
rect 7193 26401 7205 26404
rect 7239 26401 7251 26435
rect 7193 26395 7251 26401
rect 11054 26392 11060 26444
rect 11112 26392 11118 26444
rect 16206 26392 16212 26444
rect 16264 26432 16270 26444
rect 16574 26432 16580 26444
rect 16264 26404 16580 26432
rect 16264 26392 16270 26404
rect 16574 26392 16580 26404
rect 16632 26392 16638 26444
rect 16684 26404 18184 26432
rect 4522 26324 4528 26376
rect 4580 26324 4586 26376
rect 4706 26324 4712 26376
rect 4764 26364 4770 26376
rect 4799 26367 4857 26373
rect 4799 26364 4811 26367
rect 4764 26336 4811 26364
rect 4764 26324 4770 26336
rect 4799 26333 4811 26336
rect 4845 26364 4857 26367
rect 7467 26367 7525 26373
rect 7467 26364 7479 26367
rect 4845 26336 7479 26364
rect 4845 26333 4857 26336
rect 4799 26327 4857 26333
rect 7467 26333 7479 26336
rect 7513 26364 7525 26367
rect 7513 26336 8064 26364
rect 7513 26333 7525 26336
rect 7467 26327 7525 26333
rect 8036 26308 8064 26336
rect 8662 26324 8668 26376
rect 8720 26364 8726 26376
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 8720 26336 9137 26364
rect 8720 26324 8726 26336
rect 9125 26333 9137 26336
rect 9171 26333 9183 26367
rect 9367 26367 9425 26373
rect 9367 26364 9379 26367
rect 9125 26327 9183 26333
rect 9214 26336 9379 26364
rect 7558 26296 7564 26308
rect 4448 26268 7564 26296
rect 7558 26256 7564 26268
rect 7616 26256 7622 26308
rect 8018 26256 8024 26308
rect 8076 26256 8082 26308
rect 8110 26256 8116 26308
rect 8168 26296 8174 26308
rect 9214 26296 9242 26336
rect 9367 26333 9379 26336
rect 9413 26333 9425 26367
rect 9367 26327 9425 26333
rect 10962 26324 10968 26376
rect 11020 26324 11026 26376
rect 11790 26364 11796 26376
rect 11072 26336 11796 26364
rect 8168 26268 9242 26296
rect 8168 26256 8174 26268
rect 10318 26256 10324 26308
rect 10376 26296 10382 26308
rect 10594 26296 10600 26308
rect 10376 26268 10600 26296
rect 10376 26256 10382 26268
rect 10594 26256 10600 26268
rect 10652 26256 10658 26308
rect 11072 26305 11100 26336
rect 11790 26324 11796 26336
rect 11848 26324 11854 26376
rect 12526 26324 12532 26376
rect 12584 26364 12590 26376
rect 12621 26367 12679 26373
rect 12621 26364 12633 26367
rect 12584 26336 12633 26364
rect 12584 26324 12590 26336
rect 12621 26333 12633 26336
rect 12667 26364 12679 26367
rect 12894 26364 12900 26376
rect 12667 26336 12756 26364
rect 12855 26336 12900 26364
rect 12667 26333 12679 26336
rect 12621 26327 12679 26333
rect 10689 26299 10747 26305
rect 10689 26265 10701 26299
rect 10735 26296 10747 26299
rect 11057 26299 11115 26305
rect 10735 26268 11008 26296
rect 10735 26265 10747 26268
rect 10689 26259 10747 26265
rect 1578 26188 1584 26240
rect 1636 26188 1642 26240
rect 2038 26188 2044 26240
rect 2096 26228 2102 26240
rect 2222 26228 2228 26240
rect 2096 26200 2228 26228
rect 2096 26188 2102 26200
rect 2222 26188 2228 26200
rect 2280 26188 2286 26240
rect 2498 26188 2504 26240
rect 2556 26188 2562 26240
rect 2590 26188 2596 26240
rect 2648 26228 2654 26240
rect 3510 26228 3516 26240
rect 2648 26200 3516 26228
rect 2648 26188 2654 26200
rect 3510 26188 3516 26200
rect 3568 26188 3574 26240
rect 3602 26188 3608 26240
rect 3660 26188 3666 26240
rect 4982 26188 4988 26240
rect 5040 26228 5046 26240
rect 5626 26228 5632 26240
rect 5040 26200 5632 26228
rect 5040 26188 5046 26200
rect 5626 26188 5632 26200
rect 5684 26188 5690 26240
rect 7006 26188 7012 26240
rect 7064 26228 7070 26240
rect 9398 26228 9404 26240
rect 7064 26200 9404 26228
rect 7064 26188 7070 26200
rect 9398 26188 9404 26200
rect 9456 26188 9462 26240
rect 10042 26188 10048 26240
rect 10100 26228 10106 26240
rect 10137 26231 10195 26237
rect 10137 26228 10149 26231
rect 10100 26200 10149 26228
rect 10100 26188 10106 26200
rect 10137 26197 10149 26200
rect 10183 26197 10195 26231
rect 10980 26228 11008 26268
rect 11057 26265 11069 26299
rect 11103 26265 11115 26299
rect 11057 26259 11115 26265
rect 11425 26299 11483 26305
rect 11425 26265 11437 26299
rect 11471 26296 11483 26299
rect 11698 26296 11704 26308
rect 11471 26268 11704 26296
rect 11471 26265 11483 26268
rect 11425 26259 11483 26265
rect 11698 26256 11704 26268
rect 11756 26296 11762 26308
rect 11756 26268 12020 26296
rect 11756 26256 11762 26268
rect 11992 26240 12020 26268
rect 12728 26240 12756 26336
rect 12894 26324 12900 26336
rect 12952 26324 12958 26376
rect 14550 26324 14556 26376
rect 14608 26324 14614 26376
rect 15105 26367 15163 26373
rect 15105 26333 15117 26367
rect 15151 26364 15163 26367
rect 15194 26364 15200 26376
rect 15151 26336 15200 26364
rect 15151 26333 15163 26336
rect 15105 26327 15163 26333
rect 15194 26324 15200 26336
rect 15252 26364 15258 26376
rect 16684 26364 16712 26404
rect 18156 26376 18184 26404
rect 15252 26336 16712 26364
rect 15252 26324 15258 26336
rect 16758 26324 16764 26376
rect 16816 26324 16822 26376
rect 16942 26324 16948 26376
rect 17000 26324 17006 26376
rect 17034 26324 17040 26376
rect 17092 26364 17098 26376
rect 17497 26367 17555 26373
rect 17497 26364 17509 26367
rect 17092 26336 17509 26364
rect 17092 26324 17098 26336
rect 17497 26333 17509 26336
rect 17543 26333 17555 26367
rect 17497 26327 17555 26333
rect 17678 26324 17684 26376
rect 17736 26324 17742 26376
rect 17865 26367 17923 26373
rect 17865 26333 17877 26367
rect 17911 26333 17923 26367
rect 17865 26327 17923 26333
rect 13078 26256 13084 26308
rect 13136 26296 13142 26308
rect 14366 26296 14372 26308
rect 13136 26268 14372 26296
rect 13136 26256 13142 26268
rect 14366 26256 14372 26268
rect 14424 26256 14430 26308
rect 14568 26296 14596 26324
rect 15010 26296 15016 26308
rect 14568 26268 15016 26296
rect 15010 26256 15016 26268
rect 15068 26296 15074 26308
rect 15350 26299 15408 26305
rect 15350 26296 15362 26299
rect 15068 26268 15362 26296
rect 15068 26256 15074 26268
rect 15350 26265 15362 26268
rect 15396 26265 15408 26299
rect 15350 26259 15408 26265
rect 16390 26256 16396 26308
rect 16448 26296 16454 26308
rect 16853 26299 16911 26305
rect 16853 26296 16865 26299
rect 16448 26268 16865 26296
rect 16448 26256 16454 26268
rect 16853 26265 16865 26268
rect 16899 26265 16911 26299
rect 17880 26296 17908 26327
rect 18138 26324 18144 26376
rect 18196 26324 18202 26376
rect 18248 26296 18276 26540
rect 18598 26528 18604 26540
rect 18656 26528 18662 26580
rect 18693 26571 18751 26577
rect 18693 26537 18705 26571
rect 18739 26568 18751 26571
rect 18739 26540 20576 26568
rect 18739 26537 18751 26540
rect 18693 26531 18751 26537
rect 18325 26503 18383 26509
rect 18325 26469 18337 26503
rect 18371 26500 18383 26503
rect 18782 26500 18788 26512
rect 18371 26472 18788 26500
rect 18371 26469 18383 26472
rect 18325 26463 18383 26469
rect 18782 26460 18788 26472
rect 18840 26460 18846 26512
rect 18877 26503 18935 26509
rect 18877 26469 18889 26503
rect 18923 26469 18935 26503
rect 18877 26463 18935 26469
rect 18892 26432 18920 26463
rect 19334 26460 19340 26512
rect 19392 26500 19398 26512
rect 19392 26472 19564 26500
rect 19392 26460 19398 26472
rect 19536 26441 19564 26472
rect 20070 26460 20076 26512
rect 20128 26460 20134 26512
rect 20254 26460 20260 26512
rect 20312 26500 20318 26512
rect 20312 26472 20392 26500
rect 20312 26460 20318 26472
rect 19521 26435 19579 26441
rect 18892 26404 19472 26432
rect 18506 26324 18512 26376
rect 18564 26324 18570 26376
rect 18601 26367 18659 26373
rect 18601 26333 18613 26367
rect 18647 26333 18659 26367
rect 18601 26327 18659 26333
rect 16853 26259 16911 26265
rect 17328 26268 17908 26296
rect 17972 26268 18276 26296
rect 18616 26296 18644 26327
rect 18782 26324 18788 26376
rect 18840 26324 18846 26376
rect 18874 26324 18880 26376
rect 18932 26364 18938 26376
rect 19444 26373 19472 26404
rect 19521 26401 19533 26435
rect 19567 26401 19579 26435
rect 20088 26432 20116 26460
rect 20364 26441 20392 26472
rect 20548 26441 20576 26540
rect 19904 26404 20116 26432
rect 20349 26435 20407 26441
rect 19904 26402 19932 26404
rect 19521 26395 19579 26401
rect 19812 26374 19932 26402
rect 20349 26401 20361 26435
rect 20395 26401 20407 26435
rect 20349 26395 20407 26401
rect 20533 26435 20591 26441
rect 20533 26401 20545 26435
rect 20579 26401 20591 26435
rect 20533 26395 20591 26401
rect 19812 26373 19840 26374
rect 19061 26367 19119 26373
rect 19061 26364 19073 26367
rect 18932 26336 19073 26364
rect 18932 26324 18938 26336
rect 19061 26333 19073 26336
rect 19107 26333 19119 26367
rect 19061 26327 19119 26333
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26333 19487 26367
rect 19429 26327 19487 26333
rect 19779 26367 19840 26373
rect 19779 26333 19791 26367
rect 19825 26336 19840 26367
rect 20254 26364 20260 26376
rect 19996 26336 20260 26364
rect 19825 26333 19837 26336
rect 19779 26327 19837 26333
rect 18616 26268 19334 26296
rect 11606 26228 11612 26240
rect 10980 26200 11612 26228
rect 10137 26191 10195 26197
rect 11606 26188 11612 26200
rect 11664 26188 11670 26240
rect 11793 26231 11851 26237
rect 11793 26197 11805 26231
rect 11839 26228 11851 26231
rect 11882 26228 11888 26240
rect 11839 26200 11888 26228
rect 11839 26197 11851 26200
rect 11793 26191 11851 26197
rect 11882 26188 11888 26200
rect 11940 26188 11946 26240
rect 11974 26188 11980 26240
rect 12032 26188 12038 26240
rect 12710 26188 12716 26240
rect 12768 26188 12774 26240
rect 13170 26188 13176 26240
rect 13228 26228 13234 26240
rect 15654 26228 15660 26240
rect 13228 26200 15660 26228
rect 13228 26188 13234 26200
rect 15654 26188 15660 26200
rect 15712 26188 15718 26240
rect 16482 26188 16488 26240
rect 16540 26188 16546 26240
rect 17328 26237 17356 26268
rect 17313 26231 17371 26237
rect 17313 26197 17325 26231
rect 17359 26197 17371 26231
rect 17313 26191 17371 26197
rect 17865 26231 17923 26237
rect 17865 26197 17877 26231
rect 17911 26228 17923 26231
rect 17972 26228 18000 26268
rect 17911 26200 18000 26228
rect 19306 26228 19334 26268
rect 19996 26228 20024 26336
rect 20254 26324 20260 26336
rect 20312 26324 20318 26376
rect 21266 26364 21272 26376
rect 20456 26336 21272 26364
rect 20165 26299 20223 26305
rect 20165 26265 20177 26299
rect 20211 26296 20223 26299
rect 20456 26296 20484 26336
rect 21266 26324 21272 26336
rect 21324 26324 21330 26376
rect 20211 26268 20484 26296
rect 20211 26265 20223 26268
rect 20165 26259 20223 26265
rect 19306 26200 20024 26228
rect 17911 26197 17923 26200
rect 17865 26191 17923 26197
rect 20070 26188 20076 26240
rect 20128 26228 20134 26240
rect 20438 26228 20444 26240
rect 20128 26200 20444 26228
rect 20128 26188 20134 26200
rect 20438 26188 20444 26200
rect 20496 26188 20502 26240
rect 20530 26188 20536 26240
rect 20588 26188 20594 26240
rect 20714 26188 20720 26240
rect 20772 26228 20778 26240
rect 21910 26228 21916 26240
rect 20772 26200 21916 26228
rect 20772 26188 20778 26200
rect 21910 26188 21916 26200
rect 21968 26188 21974 26240
rect 382 26120 388 26172
rect 440 26160 446 26172
rect 842 26160 848 26172
rect 440 26132 848 26160
rect 440 26120 446 26132
rect 842 26120 848 26132
rect 900 26120 906 26172
rect 1104 26138 21043 26160
rect 1104 26086 5894 26138
rect 5946 26086 5958 26138
rect 6010 26086 6022 26138
rect 6074 26086 6086 26138
rect 6138 26086 6150 26138
rect 6202 26086 10839 26138
rect 10891 26086 10903 26138
rect 10955 26086 10967 26138
rect 11019 26086 11031 26138
rect 11083 26086 11095 26138
rect 11147 26086 15784 26138
rect 15836 26086 15848 26138
rect 15900 26086 15912 26138
rect 15964 26086 15976 26138
rect 16028 26086 16040 26138
rect 16092 26086 20729 26138
rect 20781 26086 20793 26138
rect 20845 26086 20857 26138
rect 20909 26086 20921 26138
rect 20973 26086 20985 26138
rect 21037 26086 21043 26138
rect 1104 26064 21043 26086
rect 1581 26027 1639 26033
rect 1581 25993 1593 26027
rect 1627 26024 1639 26027
rect 1670 26024 1676 26036
rect 1627 25996 1676 26024
rect 1627 25993 1639 25996
rect 1581 25987 1639 25993
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 1857 26027 1915 26033
rect 1857 25993 1869 26027
rect 1903 26024 1915 26027
rect 2314 26024 2320 26036
rect 1903 25996 2320 26024
rect 1903 25993 1915 25996
rect 1857 25987 1915 25993
rect 2314 25984 2320 25996
rect 2372 25984 2378 26036
rect 2590 25984 2596 26036
rect 2648 26024 2654 26036
rect 5166 26024 5172 26036
rect 2648 25996 5172 26024
rect 2648 25984 2654 25996
rect 5166 25984 5172 25996
rect 5224 25984 5230 26036
rect 5258 25984 5264 26036
rect 5316 26024 5322 26036
rect 5534 26024 5540 26036
rect 5316 25996 5540 26024
rect 5316 25984 5322 25996
rect 5534 25984 5540 25996
rect 5592 25984 5598 26036
rect 5626 25984 5632 26036
rect 5684 26024 5690 26036
rect 5810 26024 5816 26036
rect 5684 25996 5816 26024
rect 5684 25984 5690 25996
rect 5810 25984 5816 25996
rect 5868 25984 5874 26036
rect 6270 25984 6276 26036
rect 6328 25984 6334 26036
rect 7834 26024 7840 26036
rect 7208 25996 7840 26024
rect 1946 25916 1952 25968
rect 2004 25956 2010 25968
rect 2133 25959 2191 25965
rect 2133 25956 2145 25959
rect 2004 25928 2145 25956
rect 2004 25916 2010 25928
rect 2133 25925 2145 25928
rect 2179 25925 2191 25959
rect 2133 25919 2191 25925
rect 2222 25916 2228 25968
rect 2280 25916 2286 25968
rect 2866 25916 2872 25968
rect 2924 25916 2930 25968
rect 2961 25959 3019 25965
rect 2961 25925 2973 25959
rect 3007 25925 3019 25959
rect 2961 25919 3019 25925
rect 3528 25928 4108 25956
rect 750 25848 756 25900
rect 808 25888 814 25900
rect 1397 25891 1455 25897
rect 1397 25888 1409 25891
rect 808 25860 1409 25888
rect 808 25848 814 25860
rect 1397 25857 1409 25860
rect 1443 25857 1455 25891
rect 1397 25851 1455 25857
rect 2498 25848 2504 25900
rect 2556 25848 2562 25900
rect 2593 25891 2651 25897
rect 2593 25857 2605 25891
rect 2639 25888 2651 25891
rect 2884 25888 2912 25916
rect 2639 25860 2912 25888
rect 2639 25857 2651 25860
rect 2593 25851 2651 25857
rect 2516 25806 2544 25848
rect 2990 25820 3018 25919
rect 3234 25848 3240 25900
rect 3292 25888 3298 25900
rect 3528 25897 3556 25928
rect 3513 25891 3571 25897
rect 3513 25888 3525 25891
rect 3292 25860 3525 25888
rect 3292 25848 3298 25860
rect 3513 25857 3525 25860
rect 3559 25857 3571 25891
rect 3513 25851 3571 25857
rect 3694 25848 3700 25900
rect 3752 25888 3758 25900
rect 3787 25891 3845 25897
rect 3787 25888 3799 25891
rect 3752 25860 3799 25888
rect 3752 25848 3758 25860
rect 3787 25857 3799 25860
rect 3833 25857 3845 25891
rect 4080 25888 4108 25928
rect 4154 25916 4160 25968
rect 4212 25956 4218 25968
rect 6288 25956 6316 25984
rect 7098 25956 7104 25968
rect 4212 25928 6316 25956
rect 6840 25928 7104 25956
rect 4212 25916 4218 25928
rect 4522 25888 4528 25900
rect 4080 25860 4528 25888
rect 3787 25851 3845 25857
rect 4522 25848 4528 25860
rect 4580 25848 4586 25900
rect 5166 25888 5172 25900
rect 5127 25860 5172 25888
rect 5166 25848 5172 25860
rect 5224 25848 5230 25900
rect 6840 25897 6868 25928
rect 7098 25916 7104 25928
rect 7156 25916 7162 25968
rect 7208 25897 7236 25996
rect 7834 25984 7840 25996
rect 7892 26024 7898 26036
rect 8481 26027 8539 26033
rect 8481 26024 8493 26027
rect 7892 25996 8493 26024
rect 7892 25984 7898 25996
rect 8481 25993 8493 25996
rect 8527 25993 8539 26027
rect 8481 25987 8539 25993
rect 9214 25984 9220 26036
rect 9272 26024 9278 26036
rect 9398 26024 9404 26036
rect 9272 25996 9404 26024
rect 9272 25984 9278 25996
rect 9398 25984 9404 25996
rect 9456 25984 9462 26036
rect 10042 26024 10048 26036
rect 9784 25996 10048 26024
rect 7926 25956 7932 25968
rect 7482 25928 7932 25956
rect 6825 25891 6883 25897
rect 6825 25857 6837 25891
rect 6871 25857 6883 25891
rect 6825 25851 6883 25857
rect 6917 25891 6975 25897
rect 6917 25857 6929 25891
rect 6963 25857 6975 25891
rect 6917 25851 6975 25857
rect 7193 25891 7251 25897
rect 7193 25857 7205 25891
rect 7239 25857 7251 25891
rect 7193 25851 7251 25857
rect 7377 25891 7435 25897
rect 7377 25857 7389 25891
rect 7423 25888 7435 25891
rect 7482 25888 7510 25928
rect 7926 25916 7932 25928
rect 7984 25916 7990 25968
rect 8294 25916 8300 25968
rect 8352 25956 8358 25968
rect 9784 25965 9812 25996
rect 10042 25984 10048 25996
rect 10100 25984 10106 26036
rect 11514 26024 11520 26036
rect 10152 25996 11520 26024
rect 10152 25968 10180 25996
rect 11514 25984 11520 25996
rect 11572 25984 11578 26036
rect 12342 26024 12348 26036
rect 12084 25996 12348 26024
rect 9769 25959 9827 25965
rect 8352 25928 9260 25956
rect 8352 25916 8358 25928
rect 7742 25897 7748 25900
rect 7423 25860 7510 25888
rect 7711 25891 7748 25897
rect 7423 25857 7435 25860
rect 7377 25851 7435 25857
rect 7711 25857 7723 25891
rect 7800 25888 7806 25900
rect 7800 25860 9168 25888
rect 7711 25851 7748 25857
rect 2990 25792 3262 25820
rect 3142 25644 3148 25696
rect 3200 25644 3206 25696
rect 3234 25684 3262 25792
rect 4798 25780 4804 25832
rect 4856 25820 4862 25832
rect 4893 25823 4951 25829
rect 4893 25820 4905 25823
rect 4856 25792 4905 25820
rect 4856 25780 4862 25792
rect 4893 25789 4905 25792
rect 4939 25789 4951 25823
rect 6932 25820 6960 25851
rect 7742 25848 7748 25851
rect 7800 25848 7806 25860
rect 4893 25783 4951 25789
rect 6656 25792 6960 25820
rect 6656 25761 6684 25792
rect 7006 25780 7012 25832
rect 7064 25820 7070 25832
rect 7282 25820 7288 25832
rect 7064 25792 7288 25820
rect 7064 25780 7070 25792
rect 7282 25780 7288 25792
rect 7340 25820 7346 25832
rect 7469 25823 7527 25829
rect 7469 25820 7481 25823
rect 7340 25792 7481 25820
rect 7340 25780 7346 25792
rect 7469 25789 7481 25792
rect 7515 25789 7527 25823
rect 7469 25783 7527 25789
rect 6641 25755 6699 25761
rect 4172 25724 4660 25752
rect 4172 25684 4200 25724
rect 3234 25656 4200 25684
rect 4522 25644 4528 25696
rect 4580 25644 4586 25696
rect 4632 25684 4660 25724
rect 6641 25721 6653 25755
rect 6687 25721 6699 25755
rect 6641 25715 6699 25721
rect 5166 25684 5172 25696
rect 4632 25656 5172 25684
rect 5166 25644 5172 25656
rect 5224 25644 5230 25696
rect 5810 25644 5816 25696
rect 5868 25684 5874 25696
rect 5905 25687 5963 25693
rect 5905 25684 5917 25687
rect 5868 25656 5917 25684
rect 5868 25644 5874 25656
rect 5905 25653 5917 25656
rect 5951 25653 5963 25687
rect 5905 25647 5963 25653
rect 7006 25644 7012 25696
rect 7064 25644 7070 25696
rect 7285 25687 7343 25693
rect 7285 25653 7297 25687
rect 7331 25684 7343 25687
rect 8202 25684 8208 25696
rect 7331 25656 8208 25684
rect 7331 25653 7343 25656
rect 7285 25647 7343 25653
rect 8202 25644 8208 25656
rect 8260 25644 8266 25696
rect 9140 25684 9168 25860
rect 9232 25806 9260 25928
rect 9769 25925 9781 25959
rect 9815 25925 9827 25959
rect 9769 25919 9827 25925
rect 10134 25916 10140 25968
rect 10192 25916 10198 25968
rect 11238 25956 11244 25968
rect 10428 25928 11244 25956
rect 9677 25891 9735 25897
rect 9677 25857 9689 25891
rect 9723 25888 9735 25891
rect 10428 25888 10456 25928
rect 11238 25916 11244 25928
rect 11296 25956 11302 25968
rect 12084 25956 12112 25996
rect 12342 25984 12348 25996
rect 12400 25984 12406 26036
rect 12894 25984 12900 26036
rect 12952 26024 12958 26036
rect 14734 26024 14740 26036
rect 12952 25996 14740 26024
rect 12952 25984 12958 25996
rect 11296 25928 12112 25956
rect 11296 25916 11302 25928
rect 12158 25916 12164 25968
rect 12216 25956 12222 25968
rect 13541 25959 13599 25965
rect 12216 25928 13400 25956
rect 12216 25916 12222 25928
rect 9723 25860 10456 25888
rect 10519 25891 10577 25897
rect 9723 25857 9735 25860
rect 9677 25851 9735 25857
rect 10519 25857 10531 25891
rect 10565 25888 10577 25891
rect 10686 25888 10692 25900
rect 10565 25860 10692 25888
rect 10565 25857 10577 25860
rect 10519 25851 10577 25857
rect 10612 25696 10640 25860
rect 10686 25848 10692 25860
rect 10744 25848 10750 25900
rect 11943 25891 12001 25897
rect 11943 25857 11955 25891
rect 11989 25888 12001 25891
rect 12176 25888 12204 25916
rect 11989 25860 12204 25888
rect 11989 25857 12001 25860
rect 11943 25851 12001 25857
rect 12526 25848 12532 25900
rect 12584 25888 12590 25900
rect 13265 25891 13323 25897
rect 13265 25888 13277 25891
rect 12584 25860 13277 25888
rect 12584 25848 12590 25860
rect 13265 25857 13277 25860
rect 13311 25857 13323 25891
rect 13265 25851 13323 25857
rect 13372 25832 13400 25928
rect 13541 25925 13553 25959
rect 13587 25956 13599 25959
rect 13722 25956 13728 25968
rect 13587 25928 13728 25956
rect 13587 25925 13599 25928
rect 13541 25919 13599 25925
rect 13722 25916 13728 25928
rect 13780 25916 13786 25968
rect 13998 25927 14026 25996
rect 14734 25984 14740 25996
rect 14792 25984 14798 26036
rect 15010 25984 15016 26036
rect 15068 25984 15074 26036
rect 15657 26027 15715 26033
rect 15657 25993 15669 26027
rect 15703 25993 15715 26027
rect 15657 25987 15715 25993
rect 13983 25921 14041 25927
rect 13633 25891 13691 25897
rect 13633 25857 13645 25891
rect 13679 25857 13691 25891
rect 13983 25887 13995 25921
rect 14029 25887 14041 25921
rect 13983 25881 14041 25887
rect 15028 25888 15056 25984
rect 15102 25916 15108 25968
rect 15160 25956 15166 25968
rect 15470 25956 15476 25968
rect 15160 25928 15476 25956
rect 15160 25916 15166 25928
rect 15470 25916 15476 25928
rect 15528 25916 15534 25968
rect 15672 25956 15700 25987
rect 16206 25984 16212 26036
rect 16264 26024 16270 26036
rect 16485 26027 16543 26033
rect 16485 26024 16497 26027
rect 16264 25996 16497 26024
rect 16264 25984 16270 25996
rect 16485 25993 16497 25996
rect 16531 25993 16543 26027
rect 16485 25987 16543 25993
rect 16758 25984 16764 26036
rect 16816 26024 16822 26036
rect 17681 26027 17739 26033
rect 17681 26024 17693 26027
rect 16816 25996 17693 26024
rect 16816 25984 16822 25996
rect 17681 25993 17693 25996
rect 17727 25993 17739 26027
rect 17681 25987 17739 25993
rect 18141 26027 18199 26033
rect 18141 25993 18153 26027
rect 18187 26024 18199 26027
rect 18782 26024 18788 26036
rect 18187 25996 18788 26024
rect 18187 25993 18199 25996
rect 18141 25987 18199 25993
rect 18782 25984 18788 25996
rect 18840 25984 18846 26036
rect 19797 26027 19855 26033
rect 19797 25993 19809 26027
rect 19843 25993 19855 26027
rect 19797 25987 19855 25993
rect 15672 25928 15976 25956
rect 15948 25897 15976 25928
rect 15841 25891 15899 25897
rect 15841 25888 15853 25891
rect 15028 25860 15853 25888
rect 13633 25851 13691 25857
rect 15841 25857 15853 25860
rect 15887 25857 15899 25891
rect 15841 25851 15899 25857
rect 15933 25891 15991 25897
rect 15933 25857 15945 25891
rect 15979 25857 15991 25891
rect 15933 25851 15991 25857
rect 16209 25891 16267 25897
rect 16209 25857 16221 25891
rect 16255 25888 16267 25891
rect 16776 25888 16804 25984
rect 19812 25956 19840 25987
rect 18340 25928 19840 25956
rect 16911 25904 16969 25907
rect 16255 25860 16804 25888
rect 16255 25857 16267 25860
rect 16209 25851 16267 25857
rect 16850 25852 16856 25904
rect 16908 25901 16969 25904
rect 16908 25867 16923 25901
rect 16957 25867 16969 25901
rect 18340 25897 18368 25928
rect 18690 25897 18696 25900
rect 16908 25861 16969 25867
rect 18325 25891 18383 25897
rect 16908 25860 16968 25861
rect 16908 25852 16914 25860
rect 18325 25857 18337 25891
rect 18371 25857 18383 25891
rect 18684 25888 18696 25897
rect 18651 25860 18696 25888
rect 18325 25851 18383 25857
rect 18684 25851 18696 25860
rect 11701 25823 11759 25829
rect 11701 25789 11713 25823
rect 11747 25789 11759 25823
rect 11701 25783 11759 25789
rect 13081 25823 13139 25829
rect 13081 25789 13093 25823
rect 13127 25789 13139 25823
rect 13081 25783 13139 25789
rect 11716 25752 11744 25783
rect 11716 25724 11836 25752
rect 11808 25696 11836 25724
rect 12710 25712 12716 25764
rect 12768 25752 12774 25764
rect 13096 25752 13124 25783
rect 13354 25780 13360 25832
rect 13412 25780 13418 25832
rect 12768 25724 13124 25752
rect 12768 25712 12774 25724
rect 9214 25684 9220 25696
rect 9140 25656 9220 25684
rect 9214 25644 9220 25656
rect 9272 25644 9278 25696
rect 10594 25644 10600 25696
rect 10652 25644 10658 25696
rect 10686 25644 10692 25696
rect 10744 25644 10750 25696
rect 11790 25644 11796 25696
rect 11848 25644 11854 25696
rect 12158 25644 12164 25696
rect 12216 25684 12222 25696
rect 13648 25684 13676 25851
rect 18690 25848 18696 25851
rect 18748 25848 18754 25900
rect 20165 25891 20223 25897
rect 20165 25888 20177 25891
rect 19444 25860 20177 25888
rect 13722 25780 13728 25832
rect 13780 25780 13786 25832
rect 14642 25780 14648 25832
rect 14700 25820 14706 25832
rect 15102 25820 15108 25832
rect 14700 25792 15108 25820
rect 14700 25780 14706 25792
rect 15102 25780 15108 25792
rect 15160 25780 15166 25832
rect 15286 25780 15292 25832
rect 15344 25820 15350 25832
rect 15562 25820 15568 25832
rect 15344 25792 15568 25820
rect 15344 25780 15350 25792
rect 15562 25780 15568 25792
rect 15620 25780 15626 25832
rect 16390 25780 16396 25832
rect 16448 25820 16454 25832
rect 16485 25823 16543 25829
rect 16485 25820 16497 25823
rect 16448 25792 16497 25820
rect 16448 25780 16454 25792
rect 16485 25789 16497 25792
rect 16531 25789 16543 25823
rect 16485 25783 16543 25789
rect 16669 25823 16727 25829
rect 16669 25789 16681 25823
rect 16715 25789 16727 25823
rect 16669 25783 16727 25789
rect 15304 25752 15332 25780
rect 14382 25724 15332 25752
rect 16684 25752 16712 25783
rect 18138 25780 18144 25832
rect 18196 25820 18202 25832
rect 18417 25823 18475 25829
rect 18417 25820 18429 25823
rect 18196 25792 18429 25820
rect 18196 25780 18202 25792
rect 18417 25789 18429 25792
rect 18463 25789 18475 25823
rect 18417 25783 18475 25789
rect 16684 25724 16804 25752
rect 12216 25656 13676 25684
rect 12216 25644 12222 25656
rect 13722 25644 13728 25696
rect 13780 25684 13786 25696
rect 14382 25684 14410 25724
rect 16776 25696 16804 25724
rect 17770 25712 17776 25764
rect 17828 25712 17834 25764
rect 13780 25656 14410 25684
rect 13780 25644 13786 25656
rect 14734 25644 14740 25696
rect 14792 25644 14798 25696
rect 16025 25687 16083 25693
rect 16025 25653 16037 25687
rect 16071 25684 16083 25687
rect 16301 25687 16359 25693
rect 16301 25684 16313 25687
rect 16071 25656 16313 25684
rect 16071 25653 16083 25656
rect 16025 25647 16083 25653
rect 16301 25653 16313 25656
rect 16347 25653 16359 25687
rect 16301 25647 16359 25653
rect 16758 25644 16764 25696
rect 16816 25644 16822 25696
rect 17788 25684 17816 25712
rect 19444 25684 19472 25860
rect 20165 25857 20177 25860
rect 20211 25857 20223 25891
rect 20165 25851 20223 25857
rect 17788 25656 19472 25684
rect 20438 25644 20444 25696
rect 20496 25644 20502 25696
rect 1104 25594 20884 25616
rect 1104 25542 3422 25594
rect 3474 25542 3486 25594
rect 3538 25542 3550 25594
rect 3602 25542 3614 25594
rect 3666 25542 3678 25594
rect 3730 25542 8367 25594
rect 8419 25542 8431 25594
rect 8483 25542 8495 25594
rect 8547 25542 8559 25594
rect 8611 25542 8623 25594
rect 8675 25542 13312 25594
rect 13364 25542 13376 25594
rect 13428 25542 13440 25594
rect 13492 25542 13504 25594
rect 13556 25542 13568 25594
rect 13620 25542 18257 25594
rect 18309 25542 18321 25594
rect 18373 25542 18385 25594
rect 18437 25542 18449 25594
rect 18501 25542 18513 25594
rect 18565 25542 20884 25594
rect 1104 25520 20884 25542
rect 2222 25440 2228 25492
rect 2280 25480 2286 25492
rect 2777 25483 2835 25489
rect 2777 25480 2789 25483
rect 2280 25452 2789 25480
rect 2280 25440 2286 25452
rect 2777 25449 2789 25452
rect 2823 25449 2835 25483
rect 2777 25443 2835 25449
rect 5810 25440 5816 25492
rect 5868 25480 5874 25492
rect 6914 25480 6920 25492
rect 5868 25452 6224 25480
rect 5868 25440 5874 25452
rect 2498 25372 2504 25424
rect 2556 25412 2562 25424
rect 3234 25412 3240 25424
rect 2556 25384 3240 25412
rect 2556 25372 2562 25384
rect 3234 25372 3240 25384
rect 3292 25372 3298 25424
rect 3976 25356 4028 25362
rect 1302 25304 1308 25356
rect 1360 25344 1366 25356
rect 1360 25316 1808 25344
rect 1360 25304 1366 25316
rect 1780 25288 1808 25316
rect 6196 25344 6224 25452
rect 6405 25452 6920 25480
rect 6273 25347 6331 25353
rect 6273 25344 6285 25347
rect 6196 25316 6285 25344
rect 6273 25313 6285 25316
rect 6319 25313 6331 25347
rect 6405 25344 6433 25452
rect 6914 25440 6920 25452
rect 6972 25440 6978 25492
rect 7006 25440 7012 25492
rect 7064 25480 7070 25492
rect 7064 25452 8064 25480
rect 7064 25440 7070 25452
rect 7282 25372 7288 25424
rect 7340 25372 7346 25424
rect 7374 25372 7380 25424
rect 7432 25372 7438 25424
rect 7834 25412 7840 25424
rect 7760 25384 7840 25412
rect 6549 25347 6607 25353
rect 6549 25344 6561 25347
rect 6405 25316 6561 25344
rect 6273 25307 6331 25313
rect 6549 25313 6561 25316
rect 6595 25313 6607 25347
rect 6549 25307 6607 25313
rect 7006 25304 7012 25356
rect 7064 25344 7070 25356
rect 7300 25344 7328 25372
rect 7064 25316 7328 25344
rect 7064 25304 7070 25316
rect 3976 25298 4028 25304
rect 658 25236 664 25288
rect 716 25276 722 25288
rect 1397 25279 1455 25285
rect 1397 25276 1409 25279
rect 716 25248 1409 25276
rect 716 25236 722 25248
rect 1397 25245 1409 25248
rect 1443 25245 1455 25279
rect 1397 25239 1455 25245
rect 1762 25236 1768 25288
rect 1820 25236 1826 25288
rect 2039 25279 2097 25285
rect 2039 25245 2051 25279
rect 2085 25276 2097 25279
rect 2130 25276 2136 25288
rect 2085 25248 2136 25276
rect 2085 25245 2097 25248
rect 2039 25239 2097 25245
rect 2130 25236 2136 25248
rect 2188 25276 2194 25288
rect 2406 25276 2412 25288
rect 2188 25248 2412 25276
rect 2188 25236 2194 25248
rect 2406 25236 2412 25248
rect 2464 25236 2470 25288
rect 3329 25279 3387 25285
rect 3329 25245 3341 25279
rect 3375 25245 3387 25279
rect 4706 25276 4712 25288
rect 3329 25239 3387 25245
rect 4172 25248 4712 25276
rect 1302 25168 1308 25220
rect 1360 25208 1366 25220
rect 3344 25208 3372 25239
rect 4172 25208 4200 25248
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 5626 25236 5632 25288
rect 5684 25236 5690 25288
rect 5718 25236 5724 25288
rect 5776 25276 5782 25288
rect 6730 25285 6736 25288
rect 5813 25279 5871 25285
rect 5813 25276 5825 25279
rect 5776 25248 5825 25276
rect 5776 25236 5782 25248
rect 5813 25245 5825 25248
rect 5859 25245 5871 25279
rect 5813 25239 5871 25245
rect 6687 25279 6736 25285
rect 6687 25245 6699 25279
rect 6733 25245 6736 25279
rect 6687 25239 6736 25245
rect 6702 25238 6736 25239
rect 6730 25236 6736 25238
rect 6788 25236 6794 25288
rect 6822 25236 6828 25288
rect 6880 25236 6886 25288
rect 1360 25180 3372 25208
rect 3896 25180 4200 25208
rect 1360 25168 1366 25180
rect 1581 25143 1639 25149
rect 1581 25109 1593 25143
rect 1627 25140 1639 25143
rect 2590 25140 2596 25152
rect 1627 25112 2596 25140
rect 1627 25109 1639 25112
rect 1581 25103 1639 25109
rect 2590 25100 2596 25112
rect 2648 25100 2654 25152
rect 3145 25143 3203 25149
rect 3145 25109 3157 25143
rect 3191 25140 3203 25143
rect 3896 25140 3924 25180
rect 4246 25168 4252 25220
rect 4304 25168 4310 25220
rect 4341 25211 4399 25217
rect 4341 25177 4353 25211
rect 4387 25208 4399 25211
rect 4614 25208 4620 25220
rect 4387 25180 4620 25208
rect 4387 25177 4399 25180
rect 4341 25171 4399 25177
rect 4614 25168 4620 25180
rect 4672 25168 4678 25220
rect 4798 25168 4804 25220
rect 4856 25208 4862 25220
rect 7392 25208 7420 25372
rect 7760 25353 7788 25384
rect 7834 25372 7840 25384
rect 7892 25372 7898 25424
rect 7745 25347 7803 25353
rect 7745 25313 7757 25347
rect 7791 25313 7803 25347
rect 7745 25307 7803 25313
rect 8036 25285 8064 25452
rect 8202 25440 8208 25492
rect 8260 25440 8266 25492
rect 9030 25440 9036 25492
rect 9088 25480 9094 25492
rect 9088 25452 11542 25480
rect 9088 25440 9094 25452
rect 8021 25279 8079 25285
rect 8021 25245 8033 25279
rect 8067 25245 8079 25279
rect 8220 25276 8248 25440
rect 10042 25304 10048 25356
rect 10100 25344 10106 25356
rect 11422 25344 11428 25356
rect 10100 25316 11428 25344
rect 10100 25304 10106 25316
rect 11422 25304 11428 25316
rect 11480 25304 11486 25356
rect 8481 25279 8539 25285
rect 8481 25276 8493 25279
rect 8220 25248 8493 25276
rect 8021 25239 8079 25245
rect 8481 25245 8493 25248
rect 8527 25245 8539 25279
rect 8481 25239 8539 25245
rect 8570 25236 8576 25288
rect 8628 25276 8634 25288
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8628 25248 8953 25276
rect 8628 25236 8634 25248
rect 8941 25245 8953 25248
rect 8987 25276 8999 25279
rect 8987 25248 9076 25276
rect 9214 25255 9220 25288
rect 8987 25245 8999 25248
rect 8941 25239 8999 25245
rect 8202 25208 8208 25220
rect 4856 25180 5488 25208
rect 7392 25180 8208 25208
rect 4856 25168 4862 25180
rect 5460 25152 5488 25180
rect 8202 25168 8208 25180
rect 8260 25168 8266 25220
rect 8754 25168 8760 25220
rect 8812 25168 8818 25220
rect 9048 25152 9076 25248
rect 9199 25249 9220 25255
rect 9199 25215 9211 25249
rect 9272 25236 9278 25288
rect 10778 25276 10784 25288
rect 9324 25248 10784 25276
rect 9245 25215 9257 25236
rect 9199 25209 9257 25215
rect 3191 25112 3924 25140
rect 3973 25143 4031 25149
rect 3191 25109 3203 25112
rect 3145 25103 3203 25109
rect 3973 25109 3985 25143
rect 4019 25140 4031 25143
rect 4062 25140 4068 25152
rect 4019 25112 4068 25140
rect 4019 25109 4031 25112
rect 3973 25103 4031 25109
rect 4062 25100 4068 25112
rect 4120 25100 4126 25152
rect 5074 25100 5080 25152
rect 5132 25100 5138 25152
rect 5258 25100 5264 25152
rect 5316 25100 5322 25152
rect 5442 25100 5448 25152
rect 5500 25100 5506 25152
rect 7466 25100 7472 25152
rect 7524 25100 7530 25152
rect 9030 25100 9036 25152
rect 9088 25100 9094 25152
rect 9214 25100 9220 25152
rect 9272 25140 9278 25152
rect 9324 25140 9352 25248
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 11238 25208 11244 25220
rect 9416 25180 11244 25208
rect 9416 25152 9444 25180
rect 11238 25168 11244 25180
rect 11296 25168 11302 25220
rect 11514 25208 11542 25452
rect 12158 25440 12164 25492
rect 12216 25440 12222 25492
rect 12437 25483 12495 25489
rect 12437 25449 12449 25483
rect 12483 25480 12495 25483
rect 12526 25480 12532 25492
rect 12483 25452 12532 25480
rect 12483 25449 12495 25452
rect 12437 25443 12495 25449
rect 12526 25440 12532 25452
rect 12584 25440 12590 25492
rect 13354 25480 13360 25492
rect 12728 25452 13360 25480
rect 12728 25412 12756 25452
rect 13354 25440 13360 25452
rect 13412 25440 13418 25492
rect 13906 25440 13912 25492
rect 13964 25480 13970 25492
rect 16390 25480 16396 25492
rect 13964 25452 16396 25480
rect 13964 25440 13970 25452
rect 16390 25440 16396 25452
rect 16448 25440 16454 25492
rect 16853 25483 16911 25489
rect 16853 25449 16865 25483
rect 16899 25480 16911 25483
rect 16942 25480 16948 25492
rect 16899 25452 16948 25480
rect 16899 25449 16911 25452
rect 16853 25443 16911 25449
rect 16942 25440 16948 25452
rect 17000 25440 17006 25492
rect 17218 25440 17224 25492
rect 17276 25480 17282 25492
rect 19058 25480 19064 25492
rect 17276 25452 19064 25480
rect 17276 25440 17282 25452
rect 19058 25440 19064 25452
rect 19116 25440 19122 25492
rect 20254 25440 20260 25492
rect 20312 25440 20318 25492
rect 12636 25384 12756 25412
rect 12636 25344 12664 25384
rect 14090 25372 14096 25424
rect 14148 25372 14154 25424
rect 16206 25372 16212 25424
rect 16264 25412 16270 25424
rect 17034 25412 17040 25424
rect 16264 25384 17040 25412
rect 16264 25372 16270 25384
rect 17034 25372 17040 25384
rect 17092 25372 17098 25424
rect 18966 25372 18972 25424
rect 19024 25372 19030 25424
rect 14108 25344 14136 25372
rect 12544 25316 12664 25344
rect 13280 25316 14136 25344
rect 12066 25236 12072 25288
rect 12124 25236 12130 25288
rect 12250 25236 12256 25288
rect 12308 25236 12314 25288
rect 12345 25279 12403 25285
rect 12345 25245 12357 25279
rect 12391 25276 12403 25279
rect 12544 25276 12572 25316
rect 13280 25288 13308 25316
rect 15286 25304 15292 25356
rect 15344 25344 15350 25356
rect 15473 25347 15531 25353
rect 15473 25344 15485 25347
rect 15344 25316 15485 25344
rect 15344 25304 15350 25316
rect 15473 25313 15485 25316
rect 15519 25313 15531 25347
rect 16574 25344 16580 25356
rect 15473 25307 15531 25313
rect 16408 25316 16580 25344
rect 12391 25248 12572 25276
rect 12391 25245 12403 25248
rect 12345 25239 12403 25245
rect 12618 25236 12624 25288
rect 12676 25236 12682 25288
rect 12895 25279 12953 25285
rect 12895 25245 12907 25279
rect 12941 25276 12953 25279
rect 13262 25276 13268 25288
rect 12941 25248 13268 25276
rect 12941 25245 12953 25248
rect 12895 25239 12953 25245
rect 13262 25236 13268 25248
rect 13320 25236 13326 25288
rect 13722 25236 13728 25288
rect 13780 25276 13786 25288
rect 13906 25276 13912 25288
rect 13780 25248 13912 25276
rect 13780 25236 13786 25248
rect 13906 25236 13912 25248
rect 13964 25276 13970 25288
rect 14093 25279 14151 25285
rect 14093 25276 14105 25279
rect 13964 25248 14105 25276
rect 13964 25236 13970 25248
rect 14093 25245 14105 25248
rect 14139 25245 14151 25279
rect 14335 25269 14393 25275
rect 14335 25252 14347 25269
rect 14093 25239 14151 25245
rect 14200 25235 14347 25252
rect 14381 25235 14393 25269
rect 15731 25249 15789 25255
rect 15731 25246 15743 25249
rect 14200 25229 14393 25235
rect 14200 25224 14378 25229
rect 14200 25208 14228 25224
rect 15730 25215 15743 25246
rect 15777 25215 15789 25249
rect 15730 25209 15789 25215
rect 15730 25208 15758 25209
rect 11514 25180 14228 25208
rect 15580 25180 15758 25208
rect 16408 25208 16436 25316
rect 16574 25304 16580 25316
rect 16632 25304 16638 25356
rect 16850 25304 16856 25356
rect 16908 25344 16914 25356
rect 17126 25344 17132 25356
rect 16908 25316 17132 25344
rect 16908 25304 16914 25316
rect 17126 25304 17132 25316
rect 17184 25344 17190 25356
rect 18984 25344 19012 25372
rect 17184 25316 19288 25344
rect 17184 25304 17190 25316
rect 16482 25236 16488 25288
rect 16540 25276 16546 25288
rect 19260 25285 19288 25316
rect 17037 25279 17095 25285
rect 17037 25276 17049 25279
rect 16540 25248 17049 25276
rect 16540 25236 16546 25248
rect 17037 25245 17049 25248
rect 17083 25245 17095 25279
rect 18969 25279 19027 25285
rect 18969 25276 18981 25279
rect 17037 25239 17095 25245
rect 17926 25248 18981 25276
rect 17126 25208 17132 25220
rect 16408 25180 17132 25208
rect 15580 25152 15608 25180
rect 17126 25168 17132 25180
rect 17184 25168 17190 25220
rect 17926 25152 17954 25248
rect 18969 25245 18981 25248
rect 19015 25245 19027 25279
rect 18969 25239 19027 25245
rect 19245 25279 19303 25285
rect 19245 25245 19257 25279
rect 19291 25245 19303 25279
rect 19245 25239 19303 25245
rect 19518 25236 19524 25288
rect 19576 25236 19582 25288
rect 9272 25112 9352 25140
rect 9272 25100 9278 25112
rect 9398 25100 9404 25152
rect 9456 25100 9462 25152
rect 9950 25100 9956 25152
rect 10008 25100 10014 25152
rect 10134 25100 10140 25152
rect 10192 25140 10198 25152
rect 10594 25140 10600 25152
rect 10192 25112 10600 25140
rect 10192 25100 10198 25112
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 13633 25143 13691 25149
rect 13633 25109 13645 25143
rect 13679 25140 13691 25143
rect 14090 25140 14096 25152
rect 13679 25112 14096 25140
rect 13679 25109 13691 25112
rect 13633 25103 13691 25109
rect 14090 25100 14096 25112
rect 14148 25100 14154 25152
rect 14274 25100 14280 25152
rect 14332 25140 14338 25152
rect 14826 25140 14832 25152
rect 14332 25112 14832 25140
rect 14332 25100 14338 25112
rect 14826 25100 14832 25112
rect 14884 25100 14890 25152
rect 15105 25143 15163 25149
rect 15105 25109 15117 25143
rect 15151 25140 15163 25143
rect 15286 25140 15292 25152
rect 15151 25112 15292 25140
rect 15151 25109 15163 25112
rect 15105 25103 15163 25109
rect 15286 25100 15292 25112
rect 15344 25100 15350 25152
rect 15562 25100 15568 25152
rect 15620 25100 15626 25152
rect 16485 25143 16543 25149
rect 16485 25109 16497 25143
rect 16531 25140 16543 25143
rect 16574 25140 16580 25152
rect 16531 25112 16580 25140
rect 16531 25109 16543 25112
rect 16485 25103 16543 25109
rect 16574 25100 16580 25112
rect 16632 25100 16638 25152
rect 17862 25100 17868 25152
rect 17920 25112 17954 25152
rect 18785 25143 18843 25149
rect 17920 25100 17926 25112
rect 18785 25109 18797 25143
rect 18831 25140 18843 25143
rect 19334 25140 19340 25152
rect 18831 25112 19340 25140
rect 18831 25109 18843 25112
rect 18785 25103 18843 25109
rect 19334 25100 19340 25112
rect 19392 25100 19398 25152
rect 1104 25050 21043 25072
rect 1104 24998 5894 25050
rect 5946 24998 5958 25050
rect 6010 24998 6022 25050
rect 6074 24998 6086 25050
rect 6138 24998 6150 25050
rect 6202 24998 10839 25050
rect 10891 24998 10903 25050
rect 10955 24998 10967 25050
rect 11019 24998 11031 25050
rect 11083 24998 11095 25050
rect 11147 24998 15784 25050
rect 15836 24998 15848 25050
rect 15900 24998 15912 25050
rect 15964 24998 15976 25050
rect 16028 24998 16040 25050
rect 16092 24998 20729 25050
rect 20781 24998 20793 25050
rect 20845 24998 20857 25050
rect 20909 24998 20921 25050
rect 20973 24998 20985 25050
rect 21037 24998 21043 25050
rect 1104 24976 21043 24998
rect 1762 24896 1768 24948
rect 1820 24936 1826 24948
rect 1820 24908 2820 24936
rect 1820 24896 1826 24908
rect 2682 24828 2688 24880
rect 2740 24828 2746 24880
rect 2792 24868 2820 24908
rect 3970 24896 3976 24948
rect 4028 24896 4034 24948
rect 4154 24896 4160 24948
rect 4212 24936 4218 24948
rect 4525 24939 4583 24945
rect 4525 24936 4537 24939
rect 4212 24908 4537 24936
rect 4212 24896 4218 24908
rect 4525 24905 4537 24908
rect 4571 24905 4583 24939
rect 4525 24899 4583 24905
rect 4706 24896 4712 24948
rect 4764 24936 4770 24948
rect 5629 24939 5687 24945
rect 5629 24936 5641 24939
rect 4764 24908 5641 24936
rect 4764 24896 4770 24908
rect 5629 24905 5641 24908
rect 5675 24905 5687 24939
rect 5629 24899 5687 24905
rect 6178 24896 6184 24948
rect 6236 24936 6242 24948
rect 6362 24936 6368 24948
rect 6236 24908 6368 24936
rect 6236 24896 6242 24908
rect 6362 24896 6368 24908
rect 6420 24896 6426 24948
rect 7377 24939 7435 24945
rect 7377 24936 7389 24939
rect 6840 24908 7389 24936
rect 6840 24880 6868 24908
rect 7377 24905 7389 24908
rect 7423 24905 7435 24939
rect 7377 24899 7435 24905
rect 7466 24896 7472 24948
rect 7524 24896 7530 24948
rect 7926 24896 7932 24948
rect 7984 24896 7990 24948
rect 9217 24939 9275 24945
rect 9217 24905 9229 24939
rect 9263 24905 9275 24939
rect 9217 24899 9275 24905
rect 2792 24840 5488 24868
rect 1210 24760 1216 24812
rect 1268 24800 1274 24812
rect 2317 24803 2375 24809
rect 2317 24800 2329 24803
rect 1268 24772 2329 24800
rect 1268 24760 1274 24772
rect 2317 24769 2329 24772
rect 2363 24769 2375 24803
rect 2317 24763 2375 24769
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24769 2651 24803
rect 2700 24800 2728 24828
rect 5460 24812 5488 24840
rect 6822 24828 6828 24880
rect 6880 24828 6886 24880
rect 3234 24809 3240 24812
rect 3203 24803 3240 24809
rect 3203 24800 3215 24803
rect 2700 24772 3215 24800
rect 2593 24763 2651 24769
rect 3203 24769 3215 24772
rect 3203 24763 3240 24769
rect 1394 24692 1400 24744
rect 1452 24692 1458 24744
rect 2608 24732 2636 24763
rect 3234 24760 3240 24763
rect 3292 24760 3298 24812
rect 4154 24760 4160 24812
rect 4212 24800 4218 24812
rect 4448 24800 4660 24810
rect 4706 24800 4712 24812
rect 4212 24782 4712 24800
rect 4212 24772 4476 24782
rect 4632 24772 4712 24782
rect 4212 24760 4218 24772
rect 4706 24760 4712 24772
rect 4764 24760 4770 24812
rect 4798 24760 4804 24812
rect 4856 24760 4862 24812
rect 4890 24760 4896 24812
rect 4948 24760 4954 24812
rect 5258 24760 5264 24812
rect 5316 24760 5322 24812
rect 5442 24760 5448 24812
rect 5500 24800 5506 24812
rect 5500 24772 5672 24800
rect 5500 24760 5506 24772
rect 4528 24744 4580 24750
rect 2332 24704 2636 24732
rect 1302 24624 1308 24676
rect 1360 24664 1366 24676
rect 2332 24664 2360 24704
rect 2866 24692 2872 24744
rect 2924 24732 2930 24744
rect 2961 24735 3019 24741
rect 2961 24732 2973 24735
rect 2924 24704 2973 24732
rect 2924 24692 2930 24704
rect 2961 24701 2973 24704
rect 3007 24701 3019 24735
rect 2961 24695 3019 24701
rect 5644 24732 5672 24772
rect 5902 24760 5908 24812
rect 5960 24800 5966 24812
rect 6639 24803 6697 24809
rect 6639 24800 6651 24803
rect 5960 24772 6651 24800
rect 5960 24760 5966 24772
rect 6639 24769 6651 24772
rect 6685 24800 6697 24803
rect 6730 24800 6736 24812
rect 6685 24772 6736 24800
rect 6685 24769 6697 24772
rect 6639 24763 6697 24769
rect 6730 24760 6736 24772
rect 6788 24760 6794 24812
rect 7484 24800 7512 24896
rect 8938 24868 8944 24880
rect 8220 24840 8944 24868
rect 8220 24809 8248 24840
rect 8938 24828 8944 24840
rect 8996 24828 9002 24880
rect 9232 24868 9260 24899
rect 9398 24896 9404 24948
rect 9456 24936 9462 24948
rect 9674 24936 9680 24948
rect 9456 24908 9680 24936
rect 9456 24896 9462 24908
rect 9674 24896 9680 24908
rect 9732 24896 9738 24948
rect 10410 24896 10416 24948
rect 10468 24936 10474 24948
rect 10594 24936 10600 24948
rect 10468 24908 10600 24936
rect 10468 24896 10474 24908
rect 10594 24896 10600 24908
rect 10652 24896 10658 24948
rect 11422 24896 11428 24948
rect 11480 24936 11486 24948
rect 11480 24908 12204 24936
rect 11480 24896 11486 24908
rect 10502 24868 10508 24880
rect 9232 24840 10508 24868
rect 10502 24828 10508 24840
rect 10560 24828 10566 24880
rect 11882 24828 11888 24880
rect 11940 24828 11946 24880
rect 12176 24868 12204 24908
rect 12250 24896 12256 24948
rect 12308 24936 12314 24948
rect 13449 24939 13507 24945
rect 13449 24936 13461 24939
rect 12308 24908 13461 24936
rect 12308 24896 12314 24908
rect 13449 24905 13461 24908
rect 13495 24905 13507 24939
rect 17862 24936 17868 24948
rect 13449 24899 13507 24905
rect 13832 24908 17868 24936
rect 12176 24840 13768 24868
rect 8113 24803 8171 24809
rect 8113 24800 8125 24803
rect 7484 24772 8125 24800
rect 8113 24769 8125 24772
rect 8159 24769 8171 24803
rect 8113 24763 8171 24769
rect 8205 24803 8263 24809
rect 8205 24769 8217 24803
rect 8251 24769 8263 24803
rect 8205 24763 8263 24769
rect 8478 24760 8484 24812
rect 8536 24800 8542 24812
rect 8536 24772 8579 24800
rect 8536 24760 8542 24772
rect 9398 24760 9404 24812
rect 9456 24800 9462 24812
rect 9827 24803 9885 24809
rect 9827 24800 9839 24803
rect 9456 24772 9839 24800
rect 9456 24760 9462 24772
rect 9827 24769 9839 24772
rect 9873 24769 9885 24803
rect 9827 24763 9885 24769
rect 10318 24760 10324 24812
rect 10376 24800 10382 24812
rect 10778 24800 10784 24812
rect 10376 24772 10784 24800
rect 10376 24760 10382 24772
rect 10778 24760 10784 24772
rect 10836 24760 10842 24812
rect 11900 24800 11928 24828
rect 13740 24812 13768 24840
rect 12035 24803 12093 24809
rect 12035 24800 12047 24803
rect 11900 24772 12047 24800
rect 12035 24769 12047 24772
rect 12081 24800 12093 24803
rect 12894 24800 12900 24812
rect 12081 24772 12900 24800
rect 12081 24769 12093 24772
rect 12035 24763 12093 24769
rect 12894 24760 12900 24772
rect 12952 24760 12958 24812
rect 13170 24760 13176 24812
rect 13228 24800 13234 24812
rect 13357 24803 13415 24809
rect 13357 24800 13369 24803
rect 13228 24772 13369 24800
rect 13228 24760 13234 24772
rect 13357 24769 13369 24772
rect 13403 24769 13415 24803
rect 13357 24763 13415 24769
rect 13630 24760 13636 24812
rect 13688 24760 13694 24812
rect 13722 24760 13728 24812
rect 13780 24760 13786 24812
rect 5994 24732 6000 24744
rect 5644 24704 6000 24732
rect 5994 24692 6000 24704
rect 6052 24732 6058 24744
rect 6365 24735 6423 24741
rect 6365 24732 6377 24735
rect 6052 24704 6377 24732
rect 6052 24692 6058 24704
rect 6365 24701 6377 24704
rect 6411 24701 6423 24735
rect 6365 24695 6423 24701
rect 9140 24704 9352 24732
rect 4528 24686 4580 24692
rect 1360 24636 2360 24664
rect 1360 24624 1366 24636
rect 2498 24624 2504 24676
rect 2556 24624 2562 24676
rect 1627 24599 1685 24605
rect 1627 24565 1639 24599
rect 1673 24596 1685 24599
rect 2682 24596 2688 24608
rect 1673 24568 2688 24596
rect 1673 24565 1685 24568
rect 1627 24559 1685 24565
rect 2682 24556 2688 24568
rect 2740 24556 2746 24608
rect 2777 24599 2835 24605
rect 2777 24565 2789 24599
rect 2823 24596 2835 24599
rect 3970 24596 3976 24608
rect 2823 24568 3976 24596
rect 2823 24565 2835 24568
rect 2777 24559 2835 24565
rect 3970 24556 3976 24568
rect 4028 24556 4034 24608
rect 5813 24599 5871 24605
rect 5813 24565 5825 24599
rect 5859 24596 5871 24599
rect 9140 24596 9168 24704
rect 5859 24568 9168 24596
rect 9324 24596 9352 24704
rect 9490 24692 9496 24744
rect 9548 24732 9554 24744
rect 9585 24735 9643 24741
rect 9585 24732 9597 24735
rect 9548 24704 9597 24732
rect 9548 24692 9554 24704
rect 9585 24701 9597 24704
rect 9631 24701 9643 24735
rect 9585 24695 9643 24701
rect 10244 24704 10732 24732
rect 10244 24596 10272 24704
rect 10318 24624 10324 24676
rect 10376 24664 10382 24676
rect 10376 24636 10640 24664
rect 10376 24624 10382 24636
rect 10612 24605 10640 24636
rect 9324 24568 10272 24596
rect 10597 24599 10655 24605
rect 5859 24565 5871 24568
rect 5813 24559 5871 24565
rect 10597 24565 10609 24599
rect 10643 24565 10655 24599
rect 10704 24596 10732 24704
rect 11790 24692 11796 24744
rect 11848 24692 11854 24744
rect 13832 24732 13860 24908
rect 17862 24896 17868 24908
rect 17920 24936 17926 24948
rect 17920 24896 17954 24936
rect 17926 24868 17954 24896
rect 18478 24871 18536 24877
rect 18478 24868 18490 24871
rect 17926 24840 18490 24868
rect 18478 24837 18490 24840
rect 18524 24837 18536 24871
rect 18478 24831 18536 24837
rect 18598 24828 18604 24880
rect 18656 24828 18662 24880
rect 14826 24809 14832 24812
rect 14783 24803 14832 24809
rect 14783 24769 14795 24803
rect 14829 24769 14832 24803
rect 14783 24763 14832 24769
rect 14826 24760 14832 24763
rect 14884 24760 14890 24812
rect 16574 24760 16580 24812
rect 16632 24760 16638 24812
rect 17095 24803 17153 24809
rect 17095 24800 17107 24803
rect 16684 24772 17107 24800
rect 12452 24704 13860 24732
rect 13909 24735 13967 24741
rect 12452 24596 12480 24704
rect 13909 24701 13921 24735
rect 13955 24701 13967 24735
rect 13909 24695 13967 24701
rect 13173 24667 13231 24673
rect 13173 24633 13185 24667
rect 13219 24664 13231 24667
rect 13354 24664 13360 24676
rect 13219 24636 13360 24664
rect 13219 24633 13231 24636
rect 13173 24627 13231 24633
rect 13354 24624 13360 24636
rect 13412 24624 13418 24676
rect 13924 24608 13952 24695
rect 14274 24692 14280 24744
rect 14332 24732 14338 24744
rect 14645 24735 14703 24741
rect 14645 24732 14657 24735
rect 14332 24704 14657 24732
rect 14332 24692 14338 24704
rect 14645 24701 14657 24704
rect 14691 24701 14703 24735
rect 14645 24695 14703 24701
rect 14921 24735 14979 24741
rect 14921 24701 14933 24735
rect 14967 24732 14979 24735
rect 16592 24732 16620 24760
rect 14967 24704 16620 24732
rect 14967 24701 14979 24704
rect 14921 24695 14979 24701
rect 14369 24667 14427 24673
rect 14369 24633 14381 24667
rect 14415 24633 14427 24667
rect 14369 24627 14427 24633
rect 10704 24568 12480 24596
rect 10597 24559 10655 24565
rect 12802 24556 12808 24608
rect 12860 24556 12866 24608
rect 12986 24556 12992 24608
rect 13044 24596 13050 24608
rect 13906 24596 13912 24608
rect 13044 24568 13912 24596
rect 13044 24556 13050 24568
rect 13906 24556 13912 24568
rect 13964 24556 13970 24608
rect 14384 24596 14412 24627
rect 16114 24624 16120 24676
rect 16172 24664 16178 24676
rect 16684 24664 16712 24772
rect 17095 24769 17107 24772
rect 17141 24769 17153 24803
rect 18616 24800 18644 24828
rect 19981 24803 20039 24809
rect 18616 24772 19656 24800
rect 17095 24763 17153 24769
rect 19628 24744 19656 24772
rect 19981 24769 19993 24803
rect 20027 24769 20039 24803
rect 19981 24763 20039 24769
rect 16850 24692 16856 24744
rect 16908 24692 16914 24744
rect 17678 24692 17684 24744
rect 17736 24732 17742 24744
rect 18138 24732 18144 24744
rect 17736 24704 18144 24732
rect 17736 24692 17742 24704
rect 18138 24692 18144 24704
rect 18196 24732 18202 24744
rect 18233 24735 18291 24741
rect 18233 24732 18245 24735
rect 18196 24704 18245 24732
rect 18196 24692 18202 24704
rect 18233 24701 18245 24704
rect 18279 24701 18291 24735
rect 18233 24695 18291 24701
rect 19610 24692 19616 24744
rect 19668 24692 19674 24744
rect 19996 24664 20024 24763
rect 16172 24636 16712 24664
rect 19306 24636 20024 24664
rect 16172 24624 16178 24636
rect 15286 24596 15292 24608
rect 14384 24568 15292 24596
rect 15286 24556 15292 24568
rect 15344 24556 15350 24608
rect 15562 24556 15568 24608
rect 15620 24556 15626 24608
rect 17862 24556 17868 24608
rect 17920 24556 17926 24608
rect 18598 24556 18604 24608
rect 18656 24596 18662 24608
rect 19306 24596 19334 24636
rect 18656 24568 19334 24596
rect 18656 24556 18662 24568
rect 19426 24556 19432 24608
rect 19484 24596 19490 24608
rect 19613 24599 19671 24605
rect 19613 24596 19625 24599
rect 19484 24568 19625 24596
rect 19484 24556 19490 24568
rect 19613 24565 19625 24568
rect 19659 24565 19671 24599
rect 19613 24559 19671 24565
rect 20254 24556 20260 24608
rect 20312 24556 20318 24608
rect 1104 24506 20884 24528
rect 1104 24454 3422 24506
rect 3474 24454 3486 24506
rect 3538 24454 3550 24506
rect 3602 24454 3614 24506
rect 3666 24454 3678 24506
rect 3730 24454 8367 24506
rect 8419 24454 8431 24506
rect 8483 24454 8495 24506
rect 8547 24454 8559 24506
rect 8611 24454 8623 24506
rect 8675 24454 13312 24506
rect 13364 24454 13376 24506
rect 13428 24454 13440 24506
rect 13492 24454 13504 24506
rect 13556 24454 13568 24506
rect 13620 24454 18257 24506
rect 18309 24454 18321 24506
rect 18373 24454 18385 24506
rect 18437 24454 18449 24506
rect 18501 24454 18513 24506
rect 18565 24454 20884 24506
rect 1104 24432 20884 24454
rect 4062 24352 4068 24404
rect 4120 24392 4126 24404
rect 4120 24364 4568 24392
rect 4120 24352 4126 24364
rect 842 24216 848 24268
rect 900 24256 906 24268
rect 1486 24256 1492 24268
rect 900 24228 1492 24256
rect 900 24216 906 24228
rect 1486 24216 1492 24228
rect 1544 24216 1550 24268
rect 2958 24216 2964 24268
rect 3016 24256 3022 24268
rect 3789 24259 3847 24265
rect 3789 24256 3801 24259
rect 3016 24228 3801 24256
rect 3016 24216 3022 24228
rect 3789 24225 3801 24228
rect 3835 24225 3847 24259
rect 4540 24256 4568 24364
rect 4614 24352 4620 24404
rect 4672 24392 4678 24404
rect 4801 24395 4859 24401
rect 4801 24392 4813 24395
rect 4672 24364 4813 24392
rect 4672 24352 4678 24364
rect 4801 24361 4813 24364
rect 4847 24361 4859 24395
rect 4801 24355 4859 24361
rect 4890 24352 4896 24404
rect 4948 24392 4954 24404
rect 5718 24392 5724 24404
rect 4948 24364 5724 24392
rect 4948 24352 4954 24364
rect 5718 24352 5724 24364
rect 5776 24352 5782 24404
rect 5810 24352 5816 24404
rect 5868 24352 5874 24404
rect 5994 24352 6000 24404
rect 6052 24392 6058 24404
rect 6052 24364 6868 24392
rect 6052 24352 6058 24364
rect 4706 24284 4712 24336
rect 4764 24324 4770 24336
rect 5828 24324 5856 24352
rect 5905 24327 5963 24333
rect 5905 24324 5917 24327
rect 4764 24296 5396 24324
rect 5828 24296 5917 24324
rect 4764 24284 4770 24296
rect 5258 24256 5264 24268
rect 4540 24228 5264 24256
rect 3789 24219 3847 24225
rect 5258 24216 5264 24228
rect 5316 24216 5322 24268
rect 5368 24256 5396 24296
rect 5905 24293 5917 24296
rect 5951 24293 5963 24327
rect 6840 24324 6868 24364
rect 7098 24352 7104 24404
rect 7156 24352 7162 24404
rect 7190 24352 7196 24404
rect 7248 24392 7254 24404
rect 8754 24392 8760 24404
rect 7248 24364 8760 24392
rect 7248 24352 7254 24364
rect 8754 24352 8760 24364
rect 8812 24352 8818 24404
rect 8938 24352 8944 24404
rect 8996 24392 9002 24404
rect 9490 24392 9496 24404
rect 8996 24364 9496 24392
rect 8996 24352 9002 24364
rect 9490 24352 9496 24364
rect 9548 24352 9554 24404
rect 10778 24352 10784 24404
rect 10836 24352 10842 24404
rect 13265 24395 13323 24401
rect 12176 24364 13032 24392
rect 7006 24324 7012 24336
rect 6840 24296 7012 24324
rect 5905 24287 5963 24293
rect 7006 24284 7012 24296
rect 7064 24324 7070 24336
rect 12176 24324 12204 24364
rect 7064 24296 7236 24324
rect 7064 24284 7070 24296
rect 6298 24259 6356 24265
rect 6298 24256 6310 24259
rect 5368 24228 6310 24256
rect 6298 24225 6310 24228
rect 6344 24225 6356 24259
rect 6298 24219 6356 24225
rect 6457 24259 6515 24265
rect 6457 24225 6469 24259
rect 6503 24256 6515 24259
rect 6822 24256 6828 24268
rect 6503 24228 6828 24256
rect 6503 24225 6515 24228
rect 6457 24219 6515 24225
rect 6822 24216 6828 24228
rect 6880 24216 6886 24268
rect 1763 24191 1821 24197
rect 1763 24157 1775 24191
rect 1809 24188 1821 24191
rect 2222 24188 2228 24200
rect 1809 24160 2228 24188
rect 1809 24157 1821 24160
rect 1763 24151 1821 24157
rect 2222 24148 2228 24160
rect 2280 24148 2286 24200
rect 2869 24191 2927 24197
rect 2869 24188 2881 24191
rect 2746 24160 2881 24188
rect 1302 24080 1308 24132
rect 1360 24120 1366 24132
rect 2746 24120 2774 24160
rect 2869 24157 2881 24160
rect 2915 24157 2927 24191
rect 3694 24188 3700 24200
rect 2869 24151 2927 24157
rect 2976 24160 3700 24188
rect 1360 24092 2774 24120
rect 1360 24080 1366 24092
rect 2976 24064 3004 24160
rect 3694 24148 3700 24160
rect 3752 24148 3758 24200
rect 4063 24191 4121 24197
rect 4063 24157 4075 24191
rect 4109 24188 4121 24191
rect 4614 24188 4620 24200
rect 4109 24160 4620 24188
rect 4109 24157 4121 24160
rect 4063 24151 4121 24157
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 5074 24148 5080 24200
rect 5132 24188 5138 24200
rect 5442 24188 5448 24200
rect 5132 24160 5448 24188
rect 5132 24148 5138 24160
rect 5442 24148 5448 24160
rect 5500 24148 5506 24200
rect 6178 24148 6184 24200
rect 6236 24148 6242 24200
rect 7208 24197 7236 24296
rect 10980 24296 12204 24324
rect 10508 24268 10560 24274
rect 10778 24256 10784 24268
rect 10508 24210 10560 24216
rect 10704 24228 10784 24256
rect 7193 24191 7251 24197
rect 7193 24157 7205 24191
rect 7239 24157 7251 24191
rect 7193 24151 7251 24157
rect 7467 24191 7525 24197
rect 7467 24157 7479 24191
rect 7513 24188 7525 24191
rect 8202 24188 8208 24200
rect 7513 24160 8208 24188
rect 7513 24157 7525 24160
rect 7467 24151 7525 24157
rect 3234 24080 3240 24132
rect 3292 24120 3298 24132
rect 4154 24120 4160 24132
rect 3292 24092 4160 24120
rect 3292 24080 3298 24092
rect 4154 24080 4160 24092
rect 4212 24080 4218 24132
rect 7208 24120 7236 24151
rect 8202 24148 8208 24160
rect 8260 24148 8266 24200
rect 8294 24148 8300 24200
rect 8352 24148 8358 24200
rect 9766 24148 9772 24200
rect 9824 24148 9830 24200
rect 9861 24191 9919 24197
rect 9861 24157 9873 24191
rect 9907 24188 9919 24191
rect 10318 24188 10324 24200
rect 9907 24160 10324 24188
rect 9907 24157 9919 24160
rect 9861 24151 9919 24157
rect 10318 24148 10324 24160
rect 10376 24148 10382 24200
rect 7834 24120 7840 24132
rect 7208 24092 7840 24120
rect 2406 24012 2412 24064
rect 2464 24052 2470 24064
rect 2501 24055 2559 24061
rect 2501 24052 2513 24055
rect 2464 24024 2513 24052
rect 2464 24012 2470 24024
rect 2501 24021 2513 24024
rect 2547 24021 2559 24055
rect 2501 24015 2559 24021
rect 2958 24012 2964 24064
rect 3016 24012 3022 24064
rect 3053 24055 3111 24061
rect 3053 24021 3065 24055
rect 3099 24052 3111 24055
rect 4062 24052 4068 24064
rect 3099 24024 4068 24052
rect 3099 24021 3111 24024
rect 3053 24015 3111 24021
rect 4062 24012 4068 24024
rect 4120 24012 4126 24064
rect 5074 24012 5080 24064
rect 5132 24052 5138 24064
rect 7208 24052 7236 24092
rect 7834 24080 7840 24092
rect 7892 24080 7898 24132
rect 8312 24120 8340 24148
rect 9950 24120 9956 24132
rect 8312 24092 9956 24120
rect 9950 24080 9956 24092
rect 10008 24080 10014 24132
rect 10134 24080 10140 24132
rect 10192 24120 10198 24132
rect 10229 24123 10287 24129
rect 10229 24120 10241 24123
rect 10192 24092 10241 24120
rect 10192 24080 10198 24092
rect 10229 24089 10241 24092
rect 10275 24120 10287 24123
rect 10502 24120 10508 24132
rect 10275 24092 10508 24120
rect 10275 24089 10287 24092
rect 10229 24083 10287 24089
rect 10502 24080 10508 24092
rect 10560 24080 10566 24132
rect 10597 24123 10655 24129
rect 10597 24089 10609 24123
rect 10643 24120 10655 24123
rect 10704 24120 10732 24228
rect 10778 24216 10784 24228
rect 10836 24216 10842 24268
rect 10980 24120 11008 24296
rect 11422 24216 11428 24268
rect 11480 24216 11486 24268
rect 12066 24216 12072 24268
rect 12124 24216 12130 24268
rect 12176 24256 12204 24296
rect 12462 24259 12520 24265
rect 12462 24256 12474 24259
rect 12176 24228 12474 24256
rect 12462 24225 12474 24228
rect 12508 24225 12520 24259
rect 12462 24219 12520 24225
rect 12621 24259 12679 24265
rect 12621 24225 12633 24259
rect 12667 24256 12679 24259
rect 12802 24256 12808 24268
rect 12667 24228 12808 24256
rect 12667 24225 12679 24228
rect 12621 24219 12679 24225
rect 12802 24216 12808 24228
rect 12860 24216 12866 24268
rect 13004 24256 13032 24364
rect 13265 24361 13277 24395
rect 13311 24392 13323 24395
rect 13538 24392 13544 24404
rect 13311 24364 13544 24392
rect 13311 24361 13323 24364
rect 13265 24355 13323 24361
rect 13538 24352 13544 24364
rect 13596 24352 13602 24404
rect 15562 24352 15568 24404
rect 15620 24352 15626 24404
rect 17678 24392 17684 24404
rect 16408 24364 17684 24392
rect 14096 24268 14148 24274
rect 13004 24228 13676 24256
rect 13648 24200 13676 24228
rect 13740 24228 14044 24256
rect 13740 24200 13768 24228
rect 11609 24191 11667 24197
rect 11609 24157 11621 24191
rect 11655 24157 11667 24191
rect 11609 24151 11667 24157
rect 10643 24092 10732 24120
rect 10796 24092 11008 24120
rect 10643 24089 10655 24092
rect 10597 24083 10655 24089
rect 5132 24024 7236 24052
rect 5132 24012 5138 24024
rect 7558 24012 7564 24064
rect 7616 24052 7622 24064
rect 8205 24055 8263 24061
rect 8205 24052 8217 24055
rect 7616 24024 8217 24052
rect 7616 24012 7622 24024
rect 8205 24021 8217 24024
rect 8251 24021 8263 24055
rect 8205 24015 8263 24021
rect 9490 24012 9496 24064
rect 9548 24052 9554 24064
rect 10796 24052 10824 24092
rect 9548 24024 10824 24052
rect 9548 24012 9554 24024
rect 10870 24012 10876 24064
rect 10928 24052 10934 24064
rect 11422 24052 11428 24064
rect 10928 24024 11428 24052
rect 10928 24012 10934 24024
rect 11422 24012 11428 24024
rect 11480 24012 11486 24064
rect 11624 24052 11652 24151
rect 12342 24148 12348 24200
rect 12400 24148 12406 24200
rect 13630 24148 13636 24200
rect 13688 24148 13694 24200
rect 13722 24148 13728 24200
rect 13780 24148 13786 24200
rect 13906 24148 13912 24200
rect 13964 24148 13970 24200
rect 14016 24178 14044 24228
rect 14096 24210 14148 24216
rect 14200 24178 14486 24188
rect 14016 24160 14486 24178
rect 14016 24150 14228 24160
rect 13924 24120 13952 24148
rect 14458 24120 14486 24160
rect 14550 24148 14556 24200
rect 14608 24148 14614 24200
rect 14645 24191 14703 24197
rect 14645 24157 14657 24191
rect 14691 24188 14703 24191
rect 14734 24188 14740 24200
rect 14691 24160 14740 24188
rect 14691 24157 14703 24160
rect 14645 24151 14703 24157
rect 14734 24148 14740 24160
rect 14792 24148 14798 24200
rect 15580 24188 15608 24352
rect 16408 24265 16436 24364
rect 17678 24352 17684 24364
rect 17736 24352 17742 24404
rect 18049 24395 18107 24401
rect 18049 24361 18061 24395
rect 18095 24392 18107 24395
rect 18230 24392 18236 24404
rect 18095 24364 18236 24392
rect 18095 24361 18107 24364
rect 18049 24355 18107 24361
rect 18230 24352 18236 24364
rect 18288 24352 18294 24404
rect 18877 24395 18935 24401
rect 18877 24392 18889 24395
rect 18432 24364 18889 24392
rect 17957 24327 18015 24333
rect 17957 24293 17969 24327
rect 18003 24324 18015 24327
rect 18325 24327 18383 24333
rect 18325 24324 18337 24327
rect 18003 24296 18337 24324
rect 18003 24293 18015 24296
rect 17957 24287 18015 24293
rect 18325 24293 18337 24296
rect 18371 24293 18383 24327
rect 18325 24287 18383 24293
rect 16393 24259 16451 24265
rect 16393 24225 16405 24259
rect 16439 24225 16451 24259
rect 18141 24264 18199 24265
rect 18141 24259 18276 24264
rect 16393 24219 16451 24225
rect 17420 24228 18000 24256
rect 16301 24191 16359 24197
rect 16301 24188 16313 24191
rect 15580 24160 16313 24188
rect 16301 24157 16313 24160
rect 16347 24188 16359 24191
rect 16649 24191 16707 24197
rect 16649 24188 16661 24191
rect 16347 24160 16661 24188
rect 16347 24157 16359 24160
rect 16301 24151 16359 24157
rect 16649 24157 16661 24160
rect 16695 24157 16707 24191
rect 16649 24151 16707 24157
rect 15013 24123 15071 24129
rect 15013 24120 15025 24123
rect 13924 24092 14394 24120
rect 14458 24092 15025 24120
rect 13906 24052 13912 24064
rect 11624 24024 13912 24052
rect 13906 24012 13912 24024
rect 13964 24012 13970 24064
rect 14090 24012 14096 24064
rect 14148 24052 14154 24064
rect 14277 24055 14335 24061
rect 14277 24052 14289 24055
rect 14148 24024 14289 24052
rect 14148 24012 14154 24024
rect 14277 24021 14289 24024
rect 14323 24021 14335 24055
rect 14366 24052 14394 24092
rect 15013 24089 15025 24092
rect 15059 24089 15071 24123
rect 17420 24120 17448 24228
rect 17862 24148 17868 24200
rect 17920 24148 17926 24200
rect 17972 24188 18000 24228
rect 18141 24225 18153 24259
rect 18187 24256 18276 24259
rect 18432 24256 18460 24364
rect 18877 24361 18889 24364
rect 18923 24361 18935 24395
rect 18877 24355 18935 24361
rect 18509 24327 18567 24333
rect 18509 24293 18521 24327
rect 18555 24324 18567 24327
rect 18555 24296 18920 24324
rect 18555 24293 18567 24296
rect 18509 24287 18567 24293
rect 18187 24236 18460 24256
rect 18187 24225 18199 24236
rect 18248 24228 18460 24236
rect 18616 24228 18828 24256
rect 18141 24219 18199 24225
rect 18233 24191 18291 24197
rect 18233 24188 18245 24191
rect 17972 24160 18245 24188
rect 18233 24157 18245 24160
rect 18279 24157 18291 24191
rect 18616 24188 18644 24228
rect 18800 24197 18828 24228
rect 18233 24151 18291 24157
rect 18340 24160 18644 24188
rect 18693 24191 18751 24197
rect 15013 24083 15071 24089
rect 16132 24092 17448 24120
rect 17880 24120 17908 24148
rect 18340 24120 18368 24160
rect 18693 24157 18705 24191
rect 18739 24157 18751 24191
rect 18693 24151 18751 24157
rect 18785 24191 18843 24197
rect 18785 24157 18797 24191
rect 18831 24157 18843 24191
rect 18892 24188 18920 24296
rect 18966 24284 18972 24336
rect 19024 24284 19030 24336
rect 18984 24256 19012 24284
rect 19245 24259 19303 24265
rect 19245 24256 19257 24259
rect 18984 24228 19257 24256
rect 19245 24225 19257 24228
rect 19291 24225 19303 24259
rect 19245 24219 19303 24225
rect 18969 24191 19027 24197
rect 18969 24188 18981 24191
rect 18892 24160 18981 24188
rect 18785 24151 18843 24157
rect 18969 24157 18981 24160
rect 19015 24157 19027 24191
rect 18969 24151 19027 24157
rect 19503 24161 19561 24167
rect 18708 24120 18736 24151
rect 19503 24127 19515 24161
rect 19549 24158 19561 24161
rect 19549 24127 19562 24158
rect 20346 24148 20352 24200
rect 20404 24188 20410 24200
rect 20622 24188 20628 24200
rect 20404 24160 20628 24188
rect 20404 24148 20410 24160
rect 20622 24148 20628 24160
rect 20680 24148 20686 24200
rect 19503 24121 19562 24127
rect 17880 24092 18368 24120
rect 18524 24092 18736 24120
rect 19534 24120 19562 24121
rect 19610 24120 19616 24132
rect 19534 24092 19616 24120
rect 15381 24055 15439 24061
rect 15381 24052 15393 24055
rect 14366 24024 15393 24052
rect 14277 24015 14335 24021
rect 15381 24021 15393 24024
rect 15427 24021 15439 24055
rect 15381 24015 15439 24021
rect 15565 24055 15623 24061
rect 15565 24021 15577 24055
rect 15611 24052 15623 24055
rect 15654 24052 15660 24064
rect 15611 24024 15660 24052
rect 15611 24021 15623 24024
rect 15565 24015 15623 24021
rect 15654 24012 15660 24024
rect 15712 24012 15718 24064
rect 16132 24061 16160 24092
rect 16117 24055 16175 24061
rect 16117 24021 16129 24055
rect 16163 24021 16175 24055
rect 16117 24015 16175 24021
rect 17773 24055 17831 24061
rect 17773 24021 17785 24055
rect 17819 24052 17831 24055
rect 18524 24052 18552 24092
rect 19610 24080 19616 24092
rect 19668 24080 19674 24132
rect 17819 24024 18552 24052
rect 17819 24021 17831 24024
rect 17773 24015 17831 24021
rect 18598 24012 18604 24064
rect 18656 24052 18662 24064
rect 20254 24052 20260 24064
rect 18656 24024 20260 24052
rect 18656 24012 18662 24024
rect 20254 24012 20260 24024
rect 20312 24012 20318 24064
rect 1104 23962 21043 23984
rect 1104 23910 5894 23962
rect 5946 23910 5958 23962
rect 6010 23910 6022 23962
rect 6074 23910 6086 23962
rect 6138 23910 6150 23962
rect 6202 23910 10839 23962
rect 10891 23910 10903 23962
rect 10955 23910 10967 23962
rect 11019 23910 11031 23962
rect 11083 23910 11095 23962
rect 11147 23910 15784 23962
rect 15836 23910 15848 23962
rect 15900 23910 15912 23962
rect 15964 23910 15976 23962
rect 16028 23910 16040 23962
rect 16092 23910 20729 23962
rect 20781 23910 20793 23962
rect 20845 23910 20857 23962
rect 20909 23910 20921 23962
rect 20973 23910 20985 23962
rect 21037 23910 21043 23962
rect 1104 23888 21043 23910
rect 1581 23851 1639 23857
rect 1581 23817 1593 23851
rect 1627 23848 1639 23851
rect 2958 23848 2964 23860
rect 1627 23820 2964 23848
rect 1627 23817 1639 23820
rect 1581 23811 1639 23817
rect 2958 23808 2964 23820
rect 3016 23808 3022 23860
rect 3234 23808 3240 23860
rect 3292 23808 3298 23860
rect 3694 23808 3700 23860
rect 3752 23848 3758 23860
rect 3752 23820 8064 23848
rect 3752 23808 3758 23820
rect 2130 23740 2136 23792
rect 2188 23740 2194 23792
rect 2409 23783 2467 23789
rect 2409 23749 2421 23783
rect 2455 23780 2467 23783
rect 8036 23780 8064 23820
rect 9490 23808 9496 23860
rect 9548 23808 9554 23860
rect 11238 23848 11244 23860
rect 10244 23820 11244 23848
rect 9766 23789 9772 23792
rect 9765 23780 9772 23789
rect 2455 23752 5580 23780
rect 8036 23752 8294 23780
rect 9727 23752 9772 23780
rect 2455 23749 2467 23752
rect 2409 23743 2467 23749
rect 750 23672 756 23724
rect 808 23712 814 23724
rect 1397 23715 1455 23721
rect 1397 23712 1409 23715
rect 808 23684 1409 23712
rect 808 23672 814 23684
rect 1397 23681 1409 23684
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 1670 23672 1676 23724
rect 1728 23672 1734 23724
rect 2501 23715 2559 23721
rect 2501 23681 2513 23715
rect 2547 23712 2559 23715
rect 2682 23712 2688 23724
rect 2547 23684 2688 23712
rect 2547 23681 2559 23684
rect 2501 23675 2559 23681
rect 2682 23672 2688 23684
rect 2740 23672 2746 23724
rect 2774 23672 2780 23724
rect 2832 23712 2838 23724
rect 2869 23715 2927 23721
rect 2869 23712 2881 23715
rect 2832 23684 2881 23712
rect 2832 23672 2838 23684
rect 2869 23681 2881 23684
rect 2915 23681 2927 23715
rect 2869 23675 2927 23681
rect 4893 23715 4951 23721
rect 4893 23681 4905 23715
rect 4939 23712 4951 23715
rect 5074 23712 5080 23724
rect 4939 23684 5080 23712
rect 4939 23681 4951 23684
rect 4893 23675 4951 23681
rect 5074 23672 5080 23684
rect 5132 23672 5138 23724
rect 5166 23672 5172 23724
rect 5224 23672 5230 23724
rect 2406 23604 2412 23656
rect 2464 23604 2470 23656
rect 3786 23604 3792 23656
rect 3844 23604 3850 23656
rect 1854 23536 1860 23588
rect 1912 23536 1918 23588
rect 3421 23579 3479 23585
rect 3421 23545 3433 23579
rect 3467 23576 3479 23579
rect 3804 23576 3832 23604
rect 3467 23548 3832 23576
rect 3467 23545 3479 23548
rect 3421 23539 3479 23545
rect 3878 23468 3884 23520
rect 3936 23508 3942 23520
rect 5166 23508 5172 23520
rect 3936 23480 5172 23508
rect 3936 23468 3942 23480
rect 5166 23468 5172 23480
rect 5224 23468 5230 23520
rect 5552 23508 5580 23752
rect 6270 23672 6276 23724
rect 6328 23712 6334 23724
rect 6365 23715 6423 23721
rect 6365 23712 6377 23715
rect 6328 23684 6377 23712
rect 6328 23672 6334 23684
rect 6365 23681 6377 23684
rect 6411 23681 6423 23715
rect 6365 23675 6423 23681
rect 7558 23672 7564 23724
rect 7616 23672 7622 23724
rect 8266 23712 8294 23752
rect 9765 23743 9772 23752
rect 9766 23740 9772 23743
rect 9824 23740 9830 23792
rect 9861 23783 9919 23789
rect 9861 23749 9873 23783
rect 9907 23780 9919 23783
rect 9950 23780 9956 23792
rect 9907 23752 9956 23780
rect 9907 23749 9919 23752
rect 9861 23743 9919 23749
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 10244 23789 10272 23820
rect 11238 23808 11244 23820
rect 11296 23808 11302 23860
rect 12986 23848 12992 23860
rect 11532 23820 12992 23848
rect 10229 23783 10287 23789
rect 10229 23749 10241 23783
rect 10275 23749 10287 23783
rect 10229 23743 10287 23749
rect 10597 23783 10655 23789
rect 10597 23749 10609 23783
rect 10643 23780 10655 23783
rect 11422 23780 11428 23792
rect 10643 23752 11428 23780
rect 10643 23749 10655 23752
rect 10597 23743 10655 23749
rect 11422 23740 11428 23752
rect 11480 23740 11486 23792
rect 11532 23721 11560 23820
rect 12986 23808 12992 23820
rect 13044 23808 13050 23860
rect 13170 23808 13176 23860
rect 13228 23848 13234 23860
rect 13357 23851 13415 23857
rect 13357 23848 13369 23851
rect 13228 23820 13369 23848
rect 13228 23808 13234 23820
rect 13357 23817 13369 23820
rect 13403 23817 13415 23851
rect 13357 23811 13415 23817
rect 14182 23808 14188 23860
rect 14240 23848 14246 23860
rect 14550 23848 14556 23860
rect 14240 23820 14556 23848
rect 14240 23808 14246 23820
rect 14550 23808 14556 23820
rect 14608 23808 14614 23860
rect 15010 23808 15016 23860
rect 15068 23848 15074 23860
rect 16114 23848 16120 23860
rect 15068 23820 16120 23848
rect 15068 23808 15074 23820
rect 16114 23808 16120 23820
rect 16172 23808 16178 23860
rect 17862 23848 17868 23860
rect 16684 23820 17868 23848
rect 16684 23780 16712 23820
rect 17862 23808 17868 23820
rect 17920 23808 17926 23860
rect 19426 23808 19432 23860
rect 19484 23808 19490 23860
rect 20254 23848 20260 23860
rect 19720 23820 20260 23848
rect 14200 23752 16712 23780
rect 11517 23715 11575 23721
rect 11517 23712 11529 23715
rect 8266 23684 11529 23712
rect 11517 23681 11529 23684
rect 11563 23681 11575 23715
rect 11517 23675 11575 23681
rect 13814 23672 13820 23724
rect 13872 23712 13878 23724
rect 14200 23721 14228 23752
rect 14185 23715 14243 23721
rect 14185 23712 14197 23715
rect 13872 23684 14197 23712
rect 13872 23672 13878 23684
rect 14185 23681 14197 23684
rect 14231 23681 14243 23715
rect 14185 23675 14243 23681
rect 14459 23715 14517 23721
rect 14459 23681 14471 23715
rect 14505 23712 14517 23715
rect 14826 23712 14832 23724
rect 14505 23684 14832 23712
rect 14505 23681 14517 23684
rect 14459 23675 14517 23681
rect 14826 23672 14832 23684
rect 14884 23672 14890 23724
rect 16684 23721 16712 23752
rect 17126 23740 17132 23792
rect 17184 23740 17190 23792
rect 19444 23780 19472 23808
rect 19260 23752 19472 23780
rect 16943 23725 17001 23731
rect 16669 23715 16727 23721
rect 16669 23681 16681 23715
rect 16715 23681 16727 23715
rect 16943 23691 16955 23725
rect 16989 23712 17001 23725
rect 17144 23712 17172 23740
rect 19260 23721 19288 23752
rect 16989 23691 17172 23712
rect 16943 23685 17172 23691
rect 16960 23684 17172 23685
rect 19245 23715 19303 23721
rect 16669 23675 16727 23681
rect 19245 23681 19257 23715
rect 19291 23681 19303 23715
rect 19245 23675 19303 23681
rect 19334 23672 19340 23724
rect 19392 23672 19398 23724
rect 19720 23721 19748 23820
rect 20254 23808 20260 23820
rect 20312 23808 20318 23860
rect 19981 23783 20039 23789
rect 19981 23749 19993 23783
rect 20027 23780 20039 23783
rect 20165 23783 20223 23789
rect 20165 23780 20177 23783
rect 20027 23752 20177 23780
rect 20027 23749 20039 23752
rect 19981 23743 20039 23749
rect 20165 23749 20177 23752
rect 20211 23749 20223 23783
rect 20165 23743 20223 23749
rect 19705 23715 19763 23721
rect 19705 23681 19717 23715
rect 19751 23681 19763 23715
rect 19705 23675 19763 23681
rect 6454 23604 6460 23656
rect 6512 23644 6518 23656
rect 6549 23647 6607 23653
rect 6549 23644 6561 23647
rect 6512 23616 6561 23644
rect 6512 23604 6518 23616
rect 6549 23613 6561 23616
rect 6595 23644 6607 23647
rect 6638 23644 6644 23656
rect 6595 23616 6644 23644
rect 6595 23613 6607 23616
rect 6549 23607 6607 23613
rect 6638 23604 6644 23616
rect 6696 23604 6702 23656
rect 7098 23604 7104 23656
rect 7156 23644 7162 23656
rect 7466 23653 7472 23656
rect 7285 23647 7343 23653
rect 7285 23644 7297 23647
rect 7156 23616 7297 23644
rect 7156 23604 7162 23616
rect 7285 23613 7297 23616
rect 7331 23613 7343 23647
rect 7285 23607 7343 23613
rect 7423 23647 7472 23653
rect 7423 23613 7435 23647
rect 7469 23613 7472 23647
rect 7423 23607 7472 23613
rect 7466 23604 7472 23607
rect 7524 23604 7530 23656
rect 10042 23604 10048 23656
rect 10100 23604 10106 23656
rect 11422 23604 11428 23656
rect 11480 23644 11486 23656
rect 11701 23647 11759 23653
rect 11701 23644 11713 23647
rect 11480 23616 11713 23644
rect 11480 23604 11486 23616
rect 11701 23613 11713 23616
rect 11747 23613 11759 23647
rect 11701 23607 11759 23613
rect 12434 23604 12440 23656
rect 12492 23604 12498 23656
rect 12526 23604 12532 23656
rect 12584 23653 12590 23656
rect 12584 23647 12612 23653
rect 12600 23613 12612 23647
rect 12584 23607 12612 23613
rect 12723 23647 12781 23653
rect 12723 23613 12735 23647
rect 12769 23644 12781 23647
rect 12769 23616 13216 23644
rect 12769 23613 12781 23616
rect 12723 23607 12781 23613
rect 12584 23604 12590 23607
rect 13188 23588 13216 23616
rect 18690 23604 18696 23656
rect 18748 23644 18754 23656
rect 19981 23647 20039 23653
rect 19981 23644 19993 23647
rect 18748 23616 19993 23644
rect 18748 23604 18754 23616
rect 19981 23613 19993 23616
rect 20027 23613 20039 23647
rect 19981 23607 20039 23613
rect 5905 23579 5963 23585
rect 5905 23545 5917 23579
rect 5951 23576 5963 23579
rect 6822 23576 6828 23588
rect 5951 23548 6828 23576
rect 5951 23545 5963 23548
rect 5905 23539 5963 23545
rect 6822 23536 6828 23548
rect 6880 23576 6886 23588
rect 7009 23579 7067 23585
rect 7009 23576 7021 23579
rect 6880 23548 7021 23576
rect 6880 23536 6886 23548
rect 7009 23545 7021 23548
rect 7055 23545 7067 23579
rect 7009 23539 7067 23545
rect 11238 23536 11244 23588
rect 11296 23576 11302 23588
rect 11882 23576 11888 23588
rect 11296 23548 11888 23576
rect 11296 23536 11302 23548
rect 11882 23536 11888 23548
rect 11940 23536 11946 23588
rect 12161 23579 12219 23585
rect 12161 23545 12173 23579
rect 12207 23545 12219 23579
rect 12161 23539 12219 23545
rect 6362 23508 6368 23520
rect 5552 23480 6368 23508
rect 6362 23468 6368 23480
rect 6420 23468 6426 23520
rect 8202 23468 8208 23520
rect 8260 23468 8266 23520
rect 10778 23468 10784 23520
rect 10836 23468 10842 23520
rect 11146 23468 11152 23520
rect 11204 23508 11210 23520
rect 11790 23508 11796 23520
rect 11204 23480 11796 23508
rect 11204 23468 11210 23480
rect 11790 23468 11796 23480
rect 11848 23468 11854 23520
rect 12066 23468 12072 23520
rect 12124 23508 12130 23520
rect 12176 23508 12204 23539
rect 13170 23536 13176 23588
rect 13228 23536 13234 23588
rect 19334 23536 19340 23588
rect 19392 23576 19398 23588
rect 20070 23576 20076 23588
rect 19392 23548 20076 23576
rect 19392 23536 19398 23548
rect 20070 23536 20076 23548
rect 20128 23536 20134 23588
rect 12124 23480 12204 23508
rect 12124 23468 12130 23480
rect 12434 23468 12440 23520
rect 12492 23508 12498 23520
rect 14274 23508 14280 23520
rect 12492 23480 14280 23508
rect 12492 23468 12498 23480
rect 14274 23468 14280 23480
rect 14332 23468 14338 23520
rect 15194 23468 15200 23520
rect 15252 23468 15258 23520
rect 15654 23468 15660 23520
rect 15712 23508 15718 23520
rect 17681 23511 17739 23517
rect 17681 23508 17693 23511
rect 15712 23480 17693 23508
rect 15712 23468 15718 23480
rect 17681 23477 17693 23480
rect 17727 23477 17739 23511
rect 17681 23471 17739 23477
rect 19058 23468 19064 23520
rect 19116 23468 19122 23520
rect 19429 23511 19487 23517
rect 19429 23477 19441 23511
rect 19475 23508 19487 23511
rect 19797 23511 19855 23517
rect 19797 23508 19809 23511
rect 19475 23480 19809 23508
rect 19475 23477 19487 23480
rect 19429 23471 19487 23477
rect 19797 23477 19809 23480
rect 19843 23477 19855 23511
rect 19797 23471 19855 23477
rect 20438 23468 20444 23520
rect 20496 23468 20502 23520
rect 1104 23418 20884 23440
rect 1104 23366 3422 23418
rect 3474 23366 3486 23418
rect 3538 23366 3550 23418
rect 3602 23366 3614 23418
rect 3666 23366 3678 23418
rect 3730 23366 8367 23418
rect 8419 23366 8431 23418
rect 8483 23366 8495 23418
rect 8547 23366 8559 23418
rect 8611 23366 8623 23418
rect 8675 23366 13312 23418
rect 13364 23366 13376 23418
rect 13428 23366 13440 23418
rect 13492 23366 13504 23418
rect 13556 23366 13568 23418
rect 13620 23366 18257 23418
rect 18309 23366 18321 23418
rect 18373 23366 18385 23418
rect 18437 23366 18449 23418
rect 18501 23366 18513 23418
rect 18565 23366 20884 23418
rect 1104 23344 20884 23366
rect 1857 23307 1915 23313
rect 1857 23273 1869 23307
rect 1903 23304 1915 23307
rect 2314 23304 2320 23316
rect 1903 23276 2320 23304
rect 1903 23273 1915 23276
rect 1857 23267 1915 23273
rect 2314 23264 2320 23276
rect 2372 23264 2378 23316
rect 2682 23264 2688 23316
rect 2740 23304 2746 23316
rect 2961 23307 3019 23313
rect 2961 23304 2973 23307
rect 2740 23276 2973 23304
rect 2740 23264 2746 23276
rect 2961 23273 2973 23276
rect 3007 23273 3019 23307
rect 5350 23304 5356 23316
rect 2961 23267 3019 23273
rect 3804 23276 5356 23304
rect 1581 23239 1639 23245
rect 1581 23205 1593 23239
rect 1627 23236 1639 23239
rect 1946 23236 1952 23248
rect 1627 23208 1952 23236
rect 1627 23205 1639 23208
rect 1581 23199 1639 23205
rect 1946 23196 1952 23208
rect 2004 23196 2010 23248
rect 3694 23128 3700 23180
rect 3752 23168 3758 23180
rect 3804 23177 3832 23276
rect 5350 23264 5356 23276
rect 5408 23264 5414 23316
rect 6380 23276 8156 23304
rect 5258 23196 5264 23248
rect 5316 23236 5322 23248
rect 5994 23236 6000 23248
rect 5316 23208 6000 23236
rect 5316 23196 5322 23208
rect 5994 23196 6000 23208
rect 6052 23196 6058 23248
rect 3789 23171 3847 23177
rect 3789 23168 3801 23171
rect 3752 23140 3801 23168
rect 3752 23128 3758 23140
rect 3789 23137 3801 23140
rect 3835 23137 3847 23171
rect 3789 23131 3847 23137
rect 5350 23128 5356 23180
rect 5408 23168 5414 23180
rect 5626 23168 5632 23180
rect 5408 23140 5632 23168
rect 5408 23128 5414 23140
rect 5626 23128 5632 23140
rect 5684 23128 5690 23180
rect 750 23060 756 23112
rect 808 23100 814 23112
rect 1397 23103 1455 23109
rect 1397 23100 1409 23103
rect 808 23072 1409 23100
rect 808 23060 814 23072
rect 1397 23069 1409 23072
rect 1443 23069 1455 23103
rect 1397 23063 1455 23069
rect 1673 23103 1731 23109
rect 1673 23069 1685 23103
rect 1719 23069 1731 23103
rect 1673 23063 1731 23069
rect 1949 23103 2007 23109
rect 1949 23069 1961 23103
rect 1995 23069 2007 23103
rect 2682 23100 2688 23112
rect 1949 23063 2007 23069
rect 2207 23073 2265 23079
rect 934 22992 940 23044
rect 992 23032 998 23044
rect 1688 23032 1716 23063
rect 992 23004 1716 23032
rect 992 22992 998 23004
rect 1964 22976 1992 23063
rect 2207 23039 2219 23073
rect 2253 23070 2265 23073
rect 2516 23072 2688 23100
rect 2253 23039 2266 23070
rect 2516 23044 2544 23072
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 4062 23100 4068 23112
rect 4023 23072 4068 23100
rect 4062 23060 4068 23072
rect 4120 23060 4126 23112
rect 2207 23033 2266 23039
rect 2238 23032 2266 23033
rect 2498 23032 2504 23044
rect 2238 23004 2504 23032
rect 2498 22992 2504 23004
rect 2556 22992 2562 23044
rect 6380 23032 6408 23276
rect 6822 23196 6828 23248
rect 6880 23236 6886 23248
rect 7101 23239 7159 23245
rect 7101 23236 7113 23239
rect 6880 23208 7113 23236
rect 6880 23196 6886 23208
rect 7101 23205 7113 23208
rect 7147 23205 7159 23239
rect 7101 23199 7159 23205
rect 6454 23128 6460 23180
rect 6512 23168 6518 23180
rect 6730 23168 6736 23180
rect 6512 23140 6736 23168
rect 6512 23128 6518 23140
rect 6730 23128 6736 23140
rect 6788 23128 6794 23180
rect 7206 23168 7234 23276
rect 7377 23171 7435 23177
rect 7377 23168 7389 23171
rect 7206 23140 7389 23168
rect 7377 23137 7389 23140
rect 7423 23137 7435 23171
rect 7377 23131 7435 23137
rect 7466 23128 7472 23180
rect 7524 23177 7530 23180
rect 7524 23171 7552 23177
rect 7540 23137 7552 23171
rect 7524 23131 7552 23137
rect 7524 23128 7530 23131
rect 7650 23128 7656 23180
rect 7708 23128 7714 23180
rect 8128 23168 8156 23276
rect 8202 23264 8208 23316
rect 8260 23304 8266 23316
rect 8260 23276 8616 23304
rect 8260 23264 8266 23276
rect 8202 23168 8208 23180
rect 8128 23140 8208 23168
rect 8202 23128 8208 23140
rect 8260 23128 8266 23180
rect 6546 23060 6552 23112
rect 6604 23100 6610 23112
rect 6641 23103 6699 23109
rect 6641 23100 6653 23103
rect 6604 23072 6653 23100
rect 6604 23060 6610 23072
rect 6641 23069 6653 23072
rect 6687 23100 6699 23103
rect 6822 23100 6828 23112
rect 6687 23072 6828 23100
rect 6687 23069 6699 23072
rect 6641 23063 6699 23069
rect 6822 23060 6828 23072
rect 6880 23060 6886 23112
rect 8588 23109 8616 23276
rect 9030 23264 9036 23316
rect 9088 23304 9094 23316
rect 9490 23304 9496 23316
rect 9088 23276 9496 23304
rect 9088 23264 9094 23276
rect 9490 23264 9496 23276
rect 9548 23264 9554 23316
rect 9950 23264 9956 23316
rect 10008 23304 10014 23316
rect 10597 23307 10655 23313
rect 10597 23304 10609 23307
rect 10008 23276 10609 23304
rect 10008 23264 10014 23276
rect 10597 23273 10609 23276
rect 10643 23273 10655 23307
rect 10597 23267 10655 23273
rect 11514 23264 11520 23316
rect 11572 23304 11578 23316
rect 11572 23276 12020 23304
rect 11572 23264 11578 23276
rect 8662 23196 8668 23248
rect 8720 23236 8726 23248
rect 9214 23236 9220 23248
rect 8720 23208 9220 23236
rect 8720 23196 8726 23208
rect 9214 23196 9220 23208
rect 9272 23196 9278 23248
rect 11992 23168 12020 23276
rect 12066 23264 12072 23316
rect 12124 23304 12130 23316
rect 12253 23307 12311 23313
rect 12253 23304 12265 23307
rect 12124 23276 12265 23304
rect 12124 23264 12130 23276
rect 12253 23273 12265 23276
rect 12299 23273 12311 23307
rect 12253 23267 12311 23273
rect 13906 23264 13912 23316
rect 13964 23264 13970 23316
rect 15194 23304 15200 23316
rect 15120 23276 15200 23304
rect 13722 23196 13728 23248
rect 13780 23236 13786 23248
rect 13924 23236 13952 23264
rect 15120 23245 15148 23276
rect 15194 23264 15200 23276
rect 15252 23264 15258 23316
rect 16114 23264 16120 23316
rect 16172 23304 16178 23316
rect 18046 23304 18052 23316
rect 16172 23276 18052 23304
rect 16172 23264 16178 23276
rect 18046 23264 18052 23276
rect 18104 23264 18110 23316
rect 18601 23307 18659 23313
rect 18601 23273 18613 23307
rect 18647 23304 18659 23307
rect 18690 23304 18696 23316
rect 18647 23276 18696 23304
rect 18647 23273 18659 23276
rect 18601 23267 18659 23273
rect 18690 23264 18696 23276
rect 18748 23264 18754 23316
rect 19058 23264 19064 23316
rect 19116 23264 19122 23316
rect 19886 23304 19892 23316
rect 19168 23276 19892 23304
rect 15111 23239 15169 23245
rect 13780 23208 14780 23236
rect 13780 23196 13786 23208
rect 11992 23140 13492 23168
rect 9125 23119 9183 23125
rect 9125 23116 9137 23119
rect 8573 23103 8631 23109
rect 8573 23069 8585 23103
rect 8619 23069 8631 23103
rect 9048 23100 9137 23116
rect 8573 23063 8631 23069
rect 8772 23088 9137 23100
rect 8772 23072 9076 23088
rect 9125 23085 9137 23088
rect 9171 23085 9183 23119
rect 9125 23079 9183 23085
rect 3988 23004 6408 23032
rect 8297 23035 8355 23041
rect 1578 22924 1584 22976
rect 1636 22964 1642 22976
rect 1946 22964 1952 22976
rect 1636 22936 1952 22964
rect 1636 22924 1642 22936
rect 1946 22924 1952 22936
rect 2004 22924 2010 22976
rect 2314 22924 2320 22976
rect 2372 22964 2378 22976
rect 3988 22964 4016 23004
rect 8297 23001 8309 23035
rect 8343 23032 8355 23035
rect 8772 23032 8800 23072
rect 9490 23060 9496 23112
rect 9548 23100 9554 23112
rect 9585 23103 9643 23109
rect 9585 23100 9597 23103
rect 9548 23072 9597 23100
rect 9548 23060 9554 23072
rect 9585 23069 9597 23072
rect 9631 23069 9643 23103
rect 11241 23103 11299 23109
rect 11241 23100 11253 23103
rect 9843 23073 9901 23079
rect 9843 23070 9855 23073
rect 9585 23063 9643 23069
rect 8343 23004 8800 23032
rect 8343 23001 8355 23004
rect 8297 22995 8355 23001
rect 9030 22992 9036 23044
rect 9088 23032 9094 23044
rect 9784 23042 9855 23070
rect 9784 23032 9812 23042
rect 9843 23039 9855 23042
rect 9889 23039 9901 23073
rect 11164 23072 11253 23100
rect 11164 23044 11192 23072
rect 11241 23069 11253 23072
rect 11287 23069 11299 23103
rect 11241 23063 11299 23069
rect 11515 23103 11573 23109
rect 11515 23069 11527 23103
rect 11561 23100 11573 23103
rect 12894 23100 12900 23112
rect 11561 23072 12900 23100
rect 11561 23069 11573 23072
rect 11515 23063 11573 23069
rect 12894 23060 12900 23072
rect 12952 23100 12958 23112
rect 13078 23100 13084 23112
rect 12952 23072 13084 23100
rect 12952 23060 12958 23072
rect 13078 23060 13084 23072
rect 13136 23060 13142 23112
rect 13464 23100 13492 23140
rect 13906 23128 13912 23180
rect 13964 23168 13970 23180
rect 14645 23171 14703 23177
rect 14645 23168 14657 23171
rect 13964 23140 14657 23168
rect 13964 23128 13970 23140
rect 14645 23137 14657 23140
rect 14691 23137 14703 23171
rect 14752 23168 14780 23208
rect 15111 23205 15123 23239
rect 15157 23205 15169 23239
rect 15111 23199 15169 23205
rect 16206 23196 16212 23248
rect 16264 23236 16270 23248
rect 18874 23236 18880 23248
rect 16264 23208 18880 23236
rect 16264 23196 16270 23208
rect 18874 23196 18880 23208
rect 18932 23196 18938 23248
rect 15194 23168 15200 23180
rect 14752 23140 15200 23168
rect 14645 23131 14703 23137
rect 15166 23129 15200 23140
rect 15194 23128 15200 23129
rect 15252 23128 15258 23180
rect 15378 23128 15384 23180
rect 15436 23128 15442 23180
rect 15488 23140 16252 23168
rect 13814 23100 13820 23112
rect 13464 23072 13820 23100
rect 13814 23060 13820 23072
rect 13872 23100 13878 23112
rect 14461 23103 14519 23109
rect 14461 23100 14473 23103
rect 13872 23072 14473 23100
rect 13872 23060 13878 23072
rect 14461 23069 14473 23072
rect 14507 23069 14519 23103
rect 14826 23100 14832 23112
rect 14461 23063 14519 23069
rect 14566 23072 14832 23100
rect 9843 23033 9901 23039
rect 9088 23004 9812 23032
rect 9088 22992 9094 23004
rect 10502 22992 10508 23044
rect 10560 22992 10566 23044
rect 11146 22992 11152 23044
rect 11204 22992 11210 23044
rect 11882 22992 11888 23044
rect 11940 23032 11946 23044
rect 14566 23032 14594 23072
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 15488 23109 15516 23140
rect 15488 23103 15556 23109
rect 15488 23072 15510 23103
rect 15498 23069 15510 23072
rect 15544 23069 15556 23103
rect 15498 23063 15556 23069
rect 15654 23060 15660 23112
rect 15712 23060 15718 23112
rect 11940 23004 14594 23032
rect 11940 22992 11946 23004
rect 2372 22936 4016 22964
rect 2372 22924 2378 22936
rect 4062 22924 4068 22976
rect 4120 22964 4126 22976
rect 4801 22967 4859 22973
rect 4801 22964 4813 22967
rect 4120 22936 4813 22964
rect 4120 22924 4126 22936
rect 4801 22933 4813 22936
rect 4847 22933 4859 22967
rect 4801 22927 4859 22933
rect 5166 22924 5172 22976
rect 5224 22964 5230 22976
rect 5442 22964 5448 22976
rect 5224 22936 5448 22964
rect 5224 22924 5230 22936
rect 5442 22924 5448 22936
rect 5500 22924 5506 22976
rect 8389 22967 8447 22973
rect 8389 22933 8401 22967
rect 8435 22964 8447 22967
rect 8754 22964 8760 22976
rect 8435 22936 8760 22964
rect 8435 22933 8447 22936
rect 8389 22927 8447 22933
rect 8754 22924 8760 22936
rect 8812 22924 8818 22976
rect 8941 22967 8999 22973
rect 8941 22933 8953 22967
rect 8987 22964 8999 22967
rect 9306 22964 9312 22976
rect 8987 22936 9312 22964
rect 8987 22933 8999 22936
rect 8941 22927 8999 22933
rect 9306 22924 9312 22936
rect 9364 22924 9370 22976
rect 10520 22964 10548 22992
rect 15194 22964 15200 22976
rect 10520 22936 15200 22964
rect 15194 22924 15200 22936
rect 15252 22964 15258 22976
rect 16224 22964 16252 23140
rect 17678 23128 17684 23180
rect 17736 23168 17742 23180
rect 17954 23168 17960 23180
rect 17736 23140 17960 23168
rect 17736 23128 17742 23140
rect 17954 23128 17960 23140
rect 18012 23128 18018 23180
rect 19076 23168 19104 23264
rect 19168 23248 19196 23276
rect 19886 23264 19892 23276
rect 19944 23264 19950 23316
rect 20070 23264 20076 23316
rect 20128 23304 20134 23316
rect 21634 23304 21640 23316
rect 20128 23276 21640 23304
rect 20128 23264 20134 23276
rect 21634 23264 21640 23276
rect 21692 23264 21698 23316
rect 19150 23196 19156 23248
rect 19208 23196 19214 23248
rect 19702 23196 19708 23248
rect 19760 23236 19766 23248
rect 20254 23236 20260 23248
rect 19760 23208 20260 23236
rect 19760 23196 19766 23208
rect 20254 23196 20260 23208
rect 20312 23196 20318 23248
rect 18708 23140 19104 23168
rect 19429 23171 19487 23177
rect 18509 23103 18567 23109
rect 18509 23069 18521 23103
rect 18555 23100 18567 23103
rect 18598 23100 18604 23112
rect 18555 23072 18604 23100
rect 18555 23069 18567 23072
rect 18509 23063 18567 23069
rect 18598 23060 18604 23072
rect 18656 23060 18662 23112
rect 18708 23109 18736 23140
rect 19429 23137 19441 23171
rect 19475 23168 19487 23171
rect 19797 23171 19855 23177
rect 19797 23168 19809 23171
rect 19475 23140 19809 23168
rect 19475 23137 19487 23140
rect 19429 23131 19487 23137
rect 19797 23137 19809 23140
rect 19843 23137 19855 23171
rect 19797 23131 19855 23137
rect 19886 23128 19892 23180
rect 19944 23168 19950 23180
rect 19981 23171 20039 23177
rect 19981 23168 19993 23171
rect 19944 23140 19993 23168
rect 19944 23128 19950 23140
rect 19981 23137 19993 23140
rect 20027 23137 20039 23171
rect 19981 23131 20039 23137
rect 18693 23103 18751 23109
rect 18693 23069 18705 23103
rect 18739 23069 18751 23103
rect 18969 23103 19027 23109
rect 18969 23100 18981 23103
rect 18693 23063 18751 23069
rect 18800 23072 18981 23100
rect 16301 23035 16359 23041
rect 16301 23001 16313 23035
rect 16347 23032 16359 23035
rect 18800 23032 18828 23072
rect 18969 23069 18981 23072
rect 19015 23069 19027 23103
rect 18969 23063 19027 23069
rect 19337 23103 19395 23109
rect 19337 23069 19349 23103
rect 19383 23069 19395 23103
rect 19337 23063 19395 23069
rect 16347 23004 18828 23032
rect 16347 23001 16359 23004
rect 16301 22995 16359 23001
rect 18708 22976 18736 23004
rect 15252 22936 16252 22964
rect 15252 22924 15258 22936
rect 18690 22924 18696 22976
rect 18748 22924 18754 22976
rect 18785 22967 18843 22973
rect 18785 22933 18797 22967
rect 18831 22964 18843 22967
rect 19352 22964 19380 23063
rect 19702 23060 19708 23112
rect 19760 23100 19766 23112
rect 19760 23072 20300 23100
rect 19760 23060 19766 23072
rect 20272 23044 20300 23072
rect 20070 22992 20076 23044
rect 20128 23032 20134 23044
rect 20165 23035 20223 23041
rect 20165 23032 20177 23035
rect 20128 23004 20177 23032
rect 20128 22992 20134 23004
rect 20165 23001 20177 23004
rect 20211 23001 20223 23035
rect 20165 22995 20223 23001
rect 20254 22992 20260 23044
rect 20312 22992 20318 23044
rect 20533 23035 20591 23041
rect 20533 23001 20545 23035
rect 20579 23032 20591 23035
rect 21266 23032 21272 23044
rect 20579 23004 21272 23032
rect 20579 23001 20591 23004
rect 20533 22995 20591 23001
rect 21266 22992 21272 23004
rect 21324 22992 21330 23044
rect 18831 22936 19380 22964
rect 19981 22967 20039 22973
rect 18831 22933 18843 22936
rect 18785 22927 18843 22933
rect 19981 22933 19993 22967
rect 20027 22964 20039 22967
rect 20438 22964 20444 22976
rect 20027 22936 20444 22964
rect 20027 22933 20039 22936
rect 19981 22927 20039 22933
rect 20438 22924 20444 22936
rect 20496 22924 20502 22976
rect 1104 22874 21043 22896
rect 1104 22822 5894 22874
rect 5946 22822 5958 22874
rect 6010 22822 6022 22874
rect 6074 22822 6086 22874
rect 6138 22822 6150 22874
rect 6202 22822 10839 22874
rect 10891 22822 10903 22874
rect 10955 22822 10967 22874
rect 11019 22822 11031 22874
rect 11083 22822 11095 22874
rect 11147 22822 15784 22874
rect 15836 22822 15848 22874
rect 15900 22822 15912 22874
rect 15964 22822 15976 22874
rect 16028 22822 16040 22874
rect 16092 22822 20729 22874
rect 20781 22822 20793 22874
rect 20845 22822 20857 22874
rect 20909 22822 20921 22874
rect 20973 22822 20985 22874
rect 21037 22822 21043 22874
rect 1104 22800 21043 22822
rect 1026 22720 1032 22772
rect 1084 22760 1090 22772
rect 1670 22760 1676 22772
rect 1084 22732 1676 22760
rect 1084 22720 1090 22732
rect 1670 22720 1676 22732
rect 1728 22720 1734 22772
rect 2041 22763 2099 22769
rect 2041 22729 2053 22763
rect 2087 22760 2099 22763
rect 2087 22732 3294 22760
rect 2087 22729 2099 22732
rect 2041 22723 2099 22729
rect 106 22652 112 22704
rect 164 22692 170 22704
rect 1302 22692 1308 22704
rect 164 22664 1308 22692
rect 164 22652 170 22664
rect 1302 22652 1308 22664
rect 1360 22652 1366 22704
rect 2314 22652 2320 22704
rect 2372 22652 2378 22704
rect 3142 22652 3148 22704
rect 3200 22652 3206 22704
rect 3266 22692 3294 22732
rect 3326 22720 3332 22772
rect 3384 22720 3390 22772
rect 3697 22763 3755 22769
rect 3697 22729 3709 22763
rect 3743 22760 3755 22763
rect 3970 22760 3976 22772
rect 3743 22732 3976 22760
rect 3743 22729 3755 22732
rect 3697 22723 3755 22729
rect 3970 22720 3976 22732
rect 4028 22720 4034 22772
rect 4338 22720 4344 22772
rect 4396 22760 4402 22772
rect 4614 22760 4620 22772
rect 4396 22732 4620 22760
rect 4396 22720 4402 22732
rect 4614 22720 4620 22732
rect 4672 22760 4678 22772
rect 4985 22763 5043 22769
rect 4985 22760 4997 22763
rect 4672 22732 4997 22760
rect 4672 22720 4678 22732
rect 4985 22729 4997 22732
rect 5031 22729 5043 22763
rect 4985 22723 5043 22729
rect 7558 22720 7564 22772
rect 7616 22760 7622 22772
rect 8846 22760 8852 22772
rect 7616 22732 8852 22760
rect 7616 22720 7622 22732
rect 8846 22720 8852 22732
rect 8904 22720 8910 22772
rect 9030 22720 9036 22772
rect 9088 22760 9094 22772
rect 9214 22760 9220 22772
rect 9088 22732 9220 22760
rect 9088 22720 9094 22732
rect 9214 22720 9220 22732
rect 9272 22720 9278 22772
rect 9398 22720 9404 22772
rect 9456 22720 9462 22772
rect 9582 22720 9588 22772
rect 9640 22760 9646 22772
rect 9766 22760 9772 22772
rect 9640 22732 9772 22760
rect 9640 22720 9646 22732
rect 9766 22720 9772 22732
rect 9824 22720 9830 22772
rect 10226 22720 10232 22772
rect 10284 22760 10290 22772
rect 10502 22760 10508 22772
rect 10284 22732 10508 22760
rect 10284 22720 10290 22732
rect 10502 22720 10508 22732
rect 10560 22720 10566 22772
rect 13814 22720 13820 22772
rect 13872 22760 13878 22772
rect 15562 22760 15568 22772
rect 13872 22732 15568 22760
rect 13872 22720 13878 22732
rect 15562 22720 15568 22732
rect 15620 22720 15626 22772
rect 19702 22760 19708 22772
rect 18156 22732 19708 22760
rect 4430 22692 4436 22704
rect 3266 22664 4436 22692
rect 4430 22652 4436 22664
rect 4488 22652 4494 22704
rect 4801 22695 4859 22701
rect 4801 22661 4813 22695
rect 4847 22692 4859 22695
rect 5166 22692 5172 22704
rect 4847 22664 5172 22692
rect 4847 22661 4859 22664
rect 4801 22655 4859 22661
rect 5166 22652 5172 22664
rect 5224 22652 5230 22704
rect 750 22584 756 22636
rect 808 22624 814 22636
rect 1397 22627 1455 22633
rect 1397 22624 1409 22627
rect 808 22596 1409 22624
rect 808 22584 814 22596
rect 1397 22593 1409 22596
rect 1443 22593 1455 22627
rect 1397 22587 1455 22593
rect 2406 22584 2412 22636
rect 2464 22584 2470 22636
rect 2774 22584 2780 22636
rect 2832 22624 2838 22636
rect 3602 22624 3608 22636
rect 2832 22596 3608 22624
rect 2832 22584 2838 22596
rect 3602 22584 3608 22596
rect 3660 22584 3666 22636
rect 3970 22584 3976 22636
rect 4028 22584 4034 22636
rect 4062 22584 4068 22636
rect 4120 22584 4126 22636
rect 4982 22584 4988 22636
rect 5040 22624 5046 22636
rect 5902 22624 5908 22636
rect 5040 22596 5908 22624
rect 5040 22584 5046 22596
rect 5902 22584 5908 22596
rect 5960 22584 5966 22636
rect 5994 22584 6000 22636
rect 6052 22624 6058 22636
rect 6822 22624 6828 22636
rect 6052 22596 6828 22624
rect 6052 22584 6058 22596
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 8295 22627 8353 22633
rect 8295 22593 8307 22627
rect 8341 22624 8353 22627
rect 9416 22624 9444 22720
rect 10134 22692 10140 22704
rect 9968 22664 10140 22692
rect 8341 22596 9444 22624
rect 8341 22593 8353 22596
rect 8295 22587 8353 22593
rect 9582 22584 9588 22636
rect 9640 22584 9646 22636
rect 9968 22633 9996 22664
rect 10134 22652 10140 22664
rect 10192 22652 10198 22704
rect 16758 22692 16764 22704
rect 10244 22664 10456 22692
rect 9953 22627 10011 22633
rect 9953 22593 9965 22627
rect 9999 22593 10011 22627
rect 10244 22624 10272 22664
rect 9953 22587 10011 22593
rect 10060 22596 10272 22624
rect 2498 22516 2504 22568
rect 2556 22516 2562 22568
rect 3878 22516 3884 22568
rect 3936 22516 3942 22568
rect 4798 22516 4804 22568
rect 4856 22556 4862 22568
rect 5169 22559 5227 22565
rect 5169 22556 5181 22559
rect 4856 22528 5181 22556
rect 4856 22516 4862 22528
rect 5169 22525 5181 22528
rect 5215 22525 5227 22559
rect 5169 22519 5227 22525
rect 5445 22559 5503 22565
rect 5445 22525 5457 22559
rect 5491 22556 5503 22559
rect 7190 22556 7196 22568
rect 5491 22528 7196 22556
rect 5491 22525 5503 22528
rect 5445 22519 5503 22525
rect 7190 22516 7196 22528
rect 7248 22516 7254 22568
rect 7834 22516 7840 22568
rect 7892 22556 7898 22568
rect 8021 22559 8079 22565
rect 8021 22556 8033 22559
rect 7892 22528 8033 22556
rect 7892 22516 7898 22528
rect 8021 22525 8033 22528
rect 8067 22525 8079 22559
rect 8021 22519 8079 22525
rect 9401 22559 9459 22565
rect 9401 22525 9413 22559
rect 9447 22525 9459 22559
rect 9401 22519 9459 22525
rect 8036 22432 8064 22519
rect 9033 22491 9091 22497
rect 9033 22457 9045 22491
rect 9079 22488 9091 22491
rect 9214 22488 9220 22500
rect 9079 22460 9220 22488
rect 9079 22457 9091 22460
rect 9033 22451 9091 22457
rect 9214 22448 9220 22460
rect 9272 22488 9278 22500
rect 9416 22488 9444 22519
rect 9490 22516 9496 22568
rect 9548 22556 9554 22568
rect 10060 22565 10088 22596
rect 10318 22584 10324 22636
rect 10376 22584 10382 22636
rect 10428 22624 10456 22664
rect 16316 22664 16764 22692
rect 11775 22657 11833 22663
rect 10428 22596 10644 22624
rect 10045 22559 10103 22565
rect 10045 22556 10057 22559
rect 9548 22528 10057 22556
rect 9548 22516 9554 22528
rect 9272 22460 9444 22488
rect 9272 22448 9278 22460
rect 1578 22380 1584 22432
rect 1636 22380 1642 22432
rect 5074 22380 5080 22432
rect 5132 22420 5138 22432
rect 6549 22423 6607 22429
rect 6549 22420 6561 22423
rect 5132 22392 6561 22420
rect 5132 22380 5138 22392
rect 6549 22389 6561 22392
rect 6595 22389 6607 22423
rect 6549 22383 6607 22389
rect 6914 22380 6920 22432
rect 6972 22420 6978 22432
rect 7190 22420 7196 22432
rect 6972 22392 7196 22420
rect 6972 22380 6978 22392
rect 7190 22380 7196 22392
rect 7248 22380 7254 22432
rect 8018 22380 8024 22432
rect 8076 22380 8082 22432
rect 8846 22380 8852 22432
rect 8904 22420 8910 22432
rect 9600 22420 9628 22528
rect 10045 22525 10057 22528
rect 10091 22525 10103 22559
rect 10616 22556 10644 22596
rect 11330 22584 11336 22636
rect 11388 22624 11394 22636
rect 11775 22624 11787 22657
rect 11388 22623 11787 22624
rect 11821 22623 11833 22657
rect 11388 22617 11833 22623
rect 11388 22596 11818 22617
rect 11388 22584 11394 22596
rect 12250 22584 12256 22636
rect 12308 22624 12314 22636
rect 13078 22624 13084 22636
rect 12308 22596 13084 22624
rect 12308 22584 12314 22596
rect 13078 22584 13084 22596
rect 13136 22584 13142 22636
rect 13906 22584 13912 22636
rect 13964 22624 13970 22636
rect 16316 22633 16344 22664
rect 16758 22652 16764 22664
rect 16816 22652 16822 22704
rect 17218 22652 17224 22704
rect 17276 22652 17282 22704
rect 14461 22627 14519 22633
rect 14461 22624 14473 22627
rect 13964 22596 14473 22624
rect 13964 22584 13970 22596
rect 14461 22593 14473 22596
rect 14507 22593 14519 22627
rect 14461 22587 14519 22593
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22593 16359 22627
rect 16301 22587 16359 22593
rect 16482 22584 16488 22636
rect 16540 22624 16546 22636
rect 16669 22627 16727 22633
rect 16669 22624 16681 22627
rect 16540 22596 16681 22624
rect 16540 22584 16546 22596
rect 16669 22593 16681 22596
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 16943 22627 17001 22633
rect 16943 22593 16955 22627
rect 16989 22624 17001 22627
rect 17236 22624 17264 22652
rect 18156 22633 18184 22732
rect 19702 22720 19708 22732
rect 19760 22720 19766 22772
rect 19886 22720 19892 22772
rect 19944 22720 19950 22772
rect 18690 22701 18696 22704
rect 18233 22695 18291 22701
rect 18233 22661 18245 22695
rect 18279 22692 18291 22695
rect 18279 22664 18644 22692
rect 18279 22661 18291 22664
rect 18233 22655 18291 22661
rect 16989 22596 17264 22624
rect 18141 22627 18199 22633
rect 16989 22593 17001 22596
rect 16943 22587 17001 22593
rect 18141 22593 18153 22627
rect 18187 22593 18199 22627
rect 18141 22587 18199 22593
rect 18325 22627 18383 22633
rect 18325 22593 18337 22627
rect 18371 22624 18383 22627
rect 18506 22624 18512 22636
rect 18371 22596 18512 22624
rect 18371 22593 18383 22596
rect 18325 22587 18383 22593
rect 18506 22584 18512 22596
rect 18564 22584 18570 22636
rect 18616 22624 18644 22664
rect 18684 22655 18696 22701
rect 18748 22692 18754 22704
rect 18748 22664 18784 22692
rect 18690 22652 18696 22655
rect 18748 22652 18754 22664
rect 19904 22624 19932 22720
rect 20165 22695 20223 22701
rect 20165 22661 20177 22695
rect 20211 22692 20223 22695
rect 20438 22692 20444 22704
rect 20211 22664 20444 22692
rect 20211 22661 20223 22664
rect 20165 22655 20223 22661
rect 20438 22652 20444 22664
rect 20496 22652 20502 22704
rect 18616 22596 19932 22624
rect 11146 22556 11152 22568
rect 10616 22528 11152 22556
rect 10045 22519 10103 22525
rect 11146 22516 11152 22528
rect 11204 22556 11210 22568
rect 15562 22565 15568 22568
rect 11517 22559 11575 22565
rect 11517 22556 11529 22559
rect 11204 22528 11529 22556
rect 11204 22516 11210 22528
rect 11517 22525 11529 22528
rect 11563 22525 11575 22559
rect 14645 22559 14703 22565
rect 14645 22556 14657 22559
rect 11517 22519 11575 22525
rect 14200 22528 14657 22556
rect 12250 22448 12256 22500
rect 12308 22488 12314 22500
rect 12529 22491 12587 22497
rect 12529 22488 12541 22491
rect 12308 22460 12541 22488
rect 12308 22448 12314 22460
rect 12529 22457 12541 22460
rect 12575 22457 12587 22491
rect 12529 22451 12587 22457
rect 14200 22432 14228 22528
rect 14645 22525 14657 22528
rect 14691 22525 14703 22559
rect 15381 22559 15439 22565
rect 15381 22556 15393 22559
rect 14645 22519 14703 22525
rect 15212 22528 15393 22556
rect 15102 22448 15108 22500
rect 15160 22448 15166 22500
rect 8904 22392 9628 22420
rect 9861 22423 9919 22429
rect 8904 22380 8910 22392
rect 9861 22389 9873 22423
rect 9907 22420 9919 22423
rect 10502 22420 10508 22432
rect 9907 22392 10508 22420
rect 9907 22389 9919 22392
rect 9861 22383 9919 22389
rect 10502 22380 10508 22392
rect 10560 22380 10566 22432
rect 11054 22380 11060 22432
rect 11112 22380 11118 22432
rect 11422 22380 11428 22432
rect 11480 22420 11486 22432
rect 14182 22420 14188 22432
rect 11480 22392 14188 22420
rect 11480 22380 11486 22392
rect 14182 22380 14188 22392
rect 14240 22380 14246 22432
rect 14642 22380 14648 22432
rect 14700 22420 14706 22432
rect 15212 22420 15240 22528
rect 15381 22525 15393 22528
rect 15427 22525 15439 22559
rect 15381 22519 15439 22525
rect 15519 22559 15568 22565
rect 15519 22525 15531 22559
rect 15565 22525 15568 22559
rect 15519 22519 15568 22525
rect 15562 22516 15568 22519
rect 15620 22516 15626 22568
rect 15657 22559 15715 22565
rect 15657 22525 15669 22559
rect 15703 22556 15715 22559
rect 18417 22559 18475 22565
rect 15703 22528 16712 22556
rect 15703 22525 15715 22528
rect 15657 22519 15715 22525
rect 14700 22392 15240 22420
rect 16684 22420 16712 22528
rect 18417 22525 18429 22559
rect 18463 22525 18475 22559
rect 18417 22519 18475 22525
rect 18138 22448 18144 22500
rect 18196 22488 18202 22500
rect 18432 22488 18460 22519
rect 18196 22460 18460 22488
rect 18196 22448 18202 22460
rect 17681 22423 17739 22429
rect 17681 22420 17693 22423
rect 16684 22392 17693 22420
rect 14700 22380 14706 22392
rect 17681 22389 17693 22392
rect 17727 22389 17739 22423
rect 17681 22383 17739 22389
rect 19058 22380 19064 22432
rect 19116 22420 19122 22432
rect 19797 22423 19855 22429
rect 19797 22420 19809 22423
rect 19116 22392 19809 22420
rect 19116 22380 19122 22392
rect 19797 22389 19809 22392
rect 19843 22389 19855 22423
rect 19797 22383 19855 22389
rect 20438 22380 20444 22432
rect 20496 22380 20502 22432
rect 1104 22330 20884 22352
rect 1104 22278 3422 22330
rect 3474 22278 3486 22330
rect 3538 22278 3550 22330
rect 3602 22278 3614 22330
rect 3666 22278 3678 22330
rect 3730 22278 8367 22330
rect 8419 22278 8431 22330
rect 8483 22278 8495 22330
rect 8547 22278 8559 22330
rect 8611 22278 8623 22330
rect 8675 22278 13312 22330
rect 13364 22278 13376 22330
rect 13428 22278 13440 22330
rect 13492 22278 13504 22330
rect 13556 22278 13568 22330
rect 13620 22278 18257 22330
rect 18309 22278 18321 22330
rect 18373 22278 18385 22330
rect 18437 22278 18449 22330
rect 18501 22278 18513 22330
rect 18565 22278 20884 22330
rect 1104 22256 20884 22278
rect 1857 22219 1915 22225
rect 1857 22185 1869 22219
rect 1903 22216 1915 22219
rect 2774 22216 2780 22228
rect 1903 22188 2780 22216
rect 1903 22185 1915 22188
rect 1857 22179 1915 22185
rect 2774 22176 2780 22188
rect 2832 22176 2838 22228
rect 3970 22176 3976 22228
rect 4028 22216 4034 22228
rect 4433 22219 4491 22225
rect 4433 22216 4445 22219
rect 4028 22188 4445 22216
rect 4028 22176 4034 22188
rect 4433 22185 4445 22188
rect 4479 22185 4491 22219
rect 4433 22179 4491 22185
rect 6362 22176 6368 22228
rect 6420 22216 6426 22228
rect 7834 22216 7840 22228
rect 6420 22188 7840 22216
rect 6420 22176 6426 22188
rect 7834 22176 7840 22188
rect 7892 22176 7898 22228
rect 9033 22219 9091 22225
rect 9033 22185 9045 22219
rect 9079 22216 9091 22219
rect 9582 22216 9588 22228
rect 9079 22188 9588 22216
rect 9079 22185 9091 22188
rect 9033 22179 9091 22185
rect 9582 22176 9588 22188
rect 9640 22176 9646 22228
rect 14734 22216 14740 22228
rect 11624 22188 14740 22216
rect 4154 22148 4160 22160
rect 3160 22120 4160 22148
rect 1946 22040 1952 22092
rect 2004 22040 2010 22092
rect 2774 22040 2780 22092
rect 2832 22080 2838 22092
rect 3160 22080 3188 22120
rect 4154 22108 4160 22120
rect 4212 22108 4218 22160
rect 5994 22108 6000 22160
rect 6052 22108 6058 22160
rect 11624 22157 11652 22188
rect 14734 22176 14740 22188
rect 14792 22176 14798 22228
rect 15102 22176 15108 22228
rect 15160 22216 15166 22228
rect 15381 22219 15439 22225
rect 15381 22216 15393 22219
rect 15160 22188 15393 22216
rect 15160 22176 15166 22188
rect 15381 22185 15393 22188
rect 15427 22185 15439 22219
rect 16942 22216 16948 22228
rect 15381 22179 15439 22185
rect 16592 22188 16948 22216
rect 11609 22151 11667 22157
rect 11609 22117 11621 22151
rect 11655 22117 11667 22151
rect 11609 22111 11667 22117
rect 12250 22108 12256 22160
rect 12308 22108 12314 22160
rect 13262 22108 13268 22160
rect 13320 22148 13326 22160
rect 13357 22151 13415 22157
rect 13357 22148 13369 22151
rect 13320 22120 13369 22148
rect 13320 22108 13326 22120
rect 13357 22117 13369 22120
rect 13403 22117 13415 22151
rect 13357 22111 13415 22117
rect 2832 22052 3188 22080
rect 3234 22052 4016 22080
rect 2832 22040 2838 22052
rect 842 21972 848 22024
rect 900 22012 906 22024
rect 1673 22015 1731 22021
rect 1673 22012 1685 22015
rect 900 21984 1685 22012
rect 900 21972 906 21984
rect 1673 21981 1685 21984
rect 1719 21981 1731 22015
rect 1964 22012 1992 22040
rect 2041 22015 2099 22021
rect 2041 22012 2053 22015
rect 1964 21984 2053 22012
rect 1673 21975 1731 21981
rect 2041 21981 2053 21984
rect 2087 21981 2099 22015
rect 2315 22015 2373 22021
rect 2315 22012 2327 22015
rect 2041 21975 2099 21981
rect 2148 21984 2327 22012
rect 1026 21836 1032 21888
rect 1084 21876 1090 21888
rect 2148 21876 2176 21984
rect 2315 21981 2327 21984
rect 2361 22012 2373 22015
rect 3234 22012 3262 22052
rect 3988 22024 4016 22052
rect 5534 22040 5540 22092
rect 5592 22040 5598 22092
rect 5902 22040 5908 22092
rect 5960 22080 5966 22092
rect 6733 22083 6791 22089
rect 6733 22080 6745 22083
rect 5960 22052 6745 22080
rect 5960 22040 5966 22052
rect 6733 22049 6745 22052
rect 6779 22049 6791 22083
rect 6733 22043 6791 22049
rect 9306 22040 9312 22092
rect 9364 22080 9370 22092
rect 12268 22080 12296 22108
rect 9364 22052 9444 22080
rect 11362 22052 12296 22080
rect 9364 22040 9370 22052
rect 2361 21984 3262 22012
rect 2361 21981 2373 21984
rect 2315 21975 2373 21981
rect 3418 21972 3424 22024
rect 3476 21972 3482 22024
rect 3970 21972 3976 22024
rect 4028 21972 4034 22024
rect 4430 21972 4436 22024
rect 4488 21972 4494 22024
rect 4982 21972 4988 22024
rect 5040 21972 5046 22024
rect 5077 22015 5135 22021
rect 5077 21981 5089 22015
rect 5123 22012 5135 22015
rect 6178 22012 6184 22024
rect 5123 21984 6184 22012
rect 5123 21981 5135 21984
rect 5077 21975 5135 21981
rect 6178 21972 6184 21984
rect 6236 21972 6242 22024
rect 6362 21972 6368 22024
rect 6420 22012 6426 22024
rect 7007 22015 7065 22021
rect 7007 22012 7019 22015
rect 6420 22008 6684 22012
rect 6840 22008 7019 22012
rect 6420 21984 7019 22008
rect 6420 21972 6426 21984
rect 6656 21980 6868 21984
rect 4448 21944 4476 21972
rect 5445 21947 5503 21953
rect 5445 21944 5457 21947
rect 4448 21916 5457 21944
rect 5445 21913 5457 21916
rect 5491 21913 5503 21947
rect 6932 21944 6960 21984
rect 7007 21981 7019 21984
rect 7053 21981 7065 22015
rect 7007 21975 7065 21981
rect 8754 21972 8760 22024
rect 8812 22012 8818 22024
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8812 21984 8953 22012
rect 8812 21972 8818 21984
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 9214 21972 9220 22024
rect 9272 21972 9278 22024
rect 9416 22021 9444 22052
rect 9401 22015 9459 22021
rect 9401 21981 9413 22015
rect 9447 21981 9459 22015
rect 9401 21975 9459 21981
rect 9766 21972 9772 22024
rect 9824 22012 9830 22024
rect 10502 22012 10508 22024
rect 9824 21984 10508 22012
rect 9824 21972 9830 21984
rect 10502 21972 10508 21984
rect 10560 22012 10566 22024
rect 10597 22015 10655 22021
rect 10597 22012 10609 22015
rect 10560 21984 10609 22012
rect 10560 21972 10566 21984
rect 10597 21981 10609 21984
rect 10643 21981 10655 22015
rect 10597 21975 10655 21981
rect 10689 22015 10747 22021
rect 10689 21981 10701 22015
rect 10735 22012 10747 22015
rect 11146 22012 11152 22024
rect 10735 21984 11152 22012
rect 10735 21981 10747 21984
rect 10689 21975 10747 21981
rect 11146 21972 11152 21984
rect 11204 21972 11210 22024
rect 11422 21972 11428 22024
rect 11480 22021 11486 22024
rect 11480 22015 11497 22021
rect 11485 21981 11497 22015
rect 11480 21975 11497 21981
rect 11480 21972 11486 21975
rect 12066 21972 12072 22024
rect 12124 21972 12130 22024
rect 12250 21972 12256 22024
rect 12308 22012 12314 22024
rect 12345 22015 12403 22021
rect 12345 22012 12357 22015
rect 12308 21984 12357 22012
rect 12308 21972 12314 21984
rect 12345 21981 12357 21984
rect 12391 21981 12403 22015
rect 12345 21975 12403 21981
rect 12619 22015 12677 22021
rect 12619 21981 12631 22015
rect 12665 22012 12677 22015
rect 13906 22012 13912 22024
rect 12665 21984 13912 22012
rect 12665 21981 12677 21984
rect 12619 21975 12677 21981
rect 9309 21947 9367 21953
rect 6932 21916 7880 21944
rect 5445 21907 5503 21913
rect 1084 21848 2176 21876
rect 1084 21836 1090 21848
rect 2406 21836 2412 21888
rect 2464 21876 2470 21888
rect 3053 21879 3111 21885
rect 3053 21876 3065 21879
rect 2464 21848 3065 21876
rect 2464 21836 2470 21848
rect 3053 21845 3065 21848
rect 3099 21845 3111 21879
rect 3053 21839 3111 21845
rect 3602 21836 3608 21888
rect 3660 21836 3666 21888
rect 4706 21836 4712 21888
rect 4764 21836 4770 21888
rect 4982 21836 4988 21888
rect 5040 21876 5046 21888
rect 5626 21876 5632 21888
rect 5040 21848 5632 21876
rect 5040 21836 5046 21848
rect 5626 21836 5632 21848
rect 5684 21876 5690 21888
rect 5813 21879 5871 21885
rect 5813 21876 5825 21879
rect 5684 21848 5825 21876
rect 5684 21836 5690 21848
rect 5813 21845 5825 21848
rect 5859 21845 5871 21879
rect 5813 21839 5871 21845
rect 6178 21836 6184 21888
rect 6236 21876 6242 21888
rect 7745 21879 7803 21885
rect 7745 21876 7757 21879
rect 6236 21848 7757 21876
rect 6236 21836 6242 21848
rect 7745 21845 7757 21848
rect 7791 21845 7803 21879
rect 7852 21876 7880 21916
rect 9309 21913 9321 21947
rect 9355 21944 9367 21947
rect 10134 21944 10140 21956
rect 9355 21916 10140 21944
rect 9355 21913 9367 21916
rect 9309 21907 9367 21913
rect 10134 21904 10140 21916
rect 10192 21904 10198 21956
rect 10226 21904 10232 21956
rect 10284 21944 10290 21956
rect 10321 21947 10379 21953
rect 10321 21944 10333 21947
rect 10284 21916 10333 21944
rect 10284 21904 10290 21916
rect 10321 21913 10333 21916
rect 10367 21913 10379 21947
rect 10321 21907 10379 21913
rect 11057 21947 11115 21953
rect 11057 21913 11069 21947
rect 11103 21944 11115 21947
rect 12084 21944 12112 21972
rect 11103 21916 12112 21944
rect 12360 21944 12388 21975
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14369 22015 14427 22021
rect 14369 21981 14381 22015
rect 14415 21981 14427 22015
rect 14369 21975 14427 21981
rect 14643 22015 14701 22021
rect 14643 21981 14655 22015
rect 14689 22012 14701 22015
rect 15010 22012 15016 22024
rect 14689 21984 15016 22012
rect 14689 21981 14701 21984
rect 14643 21975 14701 21981
rect 12526 21944 12532 21956
rect 12360 21916 12532 21944
rect 11103 21913 11115 21916
rect 11057 21907 11115 21913
rect 12526 21904 12532 21916
rect 12584 21944 12590 21956
rect 14384 21944 14412 21975
rect 15010 21972 15016 21984
rect 15068 21972 15074 22024
rect 16592 22012 16620 22188
rect 16942 22176 16948 22188
rect 17000 22176 17006 22228
rect 18598 22176 18604 22228
rect 18656 22216 18662 22228
rect 18877 22219 18935 22225
rect 18877 22216 18889 22219
rect 18656 22188 18889 22216
rect 18656 22176 18662 22188
rect 18877 22185 18889 22188
rect 18923 22185 18935 22219
rect 18877 22179 18935 22185
rect 20254 22176 20260 22228
rect 20312 22176 20318 22228
rect 18141 22151 18199 22157
rect 18141 22117 18153 22151
rect 18187 22148 18199 22151
rect 18414 22148 18420 22160
rect 18187 22120 18420 22148
rect 18187 22117 18199 22120
rect 18141 22111 18199 22117
rect 18414 22108 18420 22120
rect 18472 22108 18478 22160
rect 18690 22108 18696 22160
rect 18748 22148 18754 22160
rect 19150 22148 19156 22160
rect 18748 22120 19156 22148
rect 18748 22108 18754 22120
rect 19150 22108 19156 22120
rect 19208 22108 19214 22160
rect 18322 22040 18328 22092
rect 18380 22080 18386 22092
rect 18966 22080 18972 22092
rect 18380 22052 18972 22080
rect 18380 22040 18386 22052
rect 18966 22040 18972 22052
rect 19024 22080 19030 22092
rect 19245 22083 19303 22089
rect 19245 22080 19257 22083
rect 19024 22052 19257 22080
rect 19024 22040 19030 22052
rect 19245 22049 19257 22052
rect 19291 22049 19303 22083
rect 19245 22043 19303 22049
rect 16669 22015 16727 22021
rect 16669 22012 16681 22015
rect 16592 21984 16681 22012
rect 16669 21981 16681 21984
rect 16715 21981 16727 22015
rect 16669 21975 16727 21981
rect 16390 21944 16396 21956
rect 12584 21916 16396 21944
rect 12584 21904 12590 21916
rect 16390 21904 16396 21916
rect 16448 21904 16454 21956
rect 16684 21944 16712 21975
rect 16758 21972 16764 22024
rect 16816 22012 16822 22024
rect 18138 22012 18144 22024
rect 16816 21984 18144 22012
rect 16816 21972 16822 21984
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 18233 22015 18291 22021
rect 18233 21981 18245 22015
rect 18279 21981 18291 22015
rect 18233 21975 18291 21981
rect 17006 21947 17064 21953
rect 17006 21944 17018 21947
rect 16684 21916 17018 21944
rect 17006 21913 17018 21916
rect 17052 21913 17064 21947
rect 17006 21907 17064 21913
rect 14826 21876 14832 21888
rect 7852 21848 14832 21876
rect 7745 21839 7803 21845
rect 14826 21836 14832 21848
rect 14884 21836 14890 21888
rect 15286 21836 15292 21888
rect 15344 21876 15350 21888
rect 16298 21876 16304 21888
rect 15344 21848 16304 21876
rect 15344 21836 15350 21848
rect 16298 21836 16304 21848
rect 16356 21836 16362 21888
rect 16485 21879 16543 21885
rect 16485 21845 16497 21879
rect 16531 21876 16543 21879
rect 18248 21876 18276 21975
rect 18414 21972 18420 22024
rect 18472 22012 18478 22024
rect 18693 22015 18751 22021
rect 18693 22012 18705 22015
rect 18472 21984 18705 22012
rect 18472 21972 18478 21984
rect 18693 21981 18705 21984
rect 18739 21981 18751 22015
rect 18693 21975 18751 21981
rect 19058 21972 19064 22024
rect 19116 21972 19122 22024
rect 19519 22015 19577 22021
rect 19519 21981 19531 22015
rect 19565 22012 19577 22015
rect 21542 22012 21548 22024
rect 19565 21984 21548 22012
rect 19565 21981 19577 21984
rect 19519 21975 19577 21981
rect 21542 21972 21548 21984
rect 21600 21972 21606 22024
rect 18966 21904 18972 21956
rect 19024 21944 19030 21956
rect 19702 21944 19708 21956
rect 19024 21916 19708 21944
rect 19024 21904 19030 21916
rect 19702 21904 19708 21916
rect 19760 21904 19766 21956
rect 16531 21848 18276 21876
rect 16531 21845 16543 21848
rect 16485 21839 16543 21845
rect 18322 21836 18328 21888
rect 18380 21836 18386 21888
rect 18509 21879 18567 21885
rect 18509 21845 18521 21879
rect 18555 21876 18567 21879
rect 19242 21876 19248 21888
rect 18555 21848 19248 21876
rect 18555 21845 18567 21848
rect 18509 21839 18567 21845
rect 19242 21836 19248 21848
rect 19300 21836 19306 21888
rect 1104 21786 21043 21808
rect 1104 21734 5894 21786
rect 5946 21734 5958 21786
rect 6010 21734 6022 21786
rect 6074 21734 6086 21786
rect 6138 21734 6150 21786
rect 6202 21734 10839 21786
rect 10891 21734 10903 21786
rect 10955 21734 10967 21786
rect 11019 21734 11031 21786
rect 11083 21734 11095 21786
rect 11147 21734 15784 21786
rect 15836 21734 15848 21786
rect 15900 21734 15912 21786
rect 15964 21734 15976 21786
rect 16028 21734 16040 21786
rect 16092 21734 20729 21786
rect 20781 21734 20793 21786
rect 20845 21734 20857 21786
rect 20909 21734 20921 21786
rect 20973 21734 20985 21786
rect 21037 21734 21043 21786
rect 1104 21712 21043 21734
rect 1578 21632 1584 21684
rect 1636 21672 1642 21684
rect 2038 21672 2044 21684
rect 1636 21644 2044 21672
rect 1636 21632 1642 21644
rect 2038 21632 2044 21644
rect 2096 21632 2102 21684
rect 2498 21632 2504 21684
rect 2556 21632 2562 21684
rect 4065 21675 4123 21681
rect 4065 21641 4077 21675
rect 4111 21641 4123 21675
rect 4065 21635 4123 21641
rect 1946 21604 1952 21616
rect 1504 21576 1952 21604
rect 1504 21545 1532 21576
rect 1946 21564 1952 21576
rect 2004 21564 2010 21616
rect 3068 21576 3832 21604
rect 1489 21539 1547 21545
rect 1489 21505 1501 21539
rect 1535 21505 1547 21539
rect 1489 21499 1547 21505
rect 1670 21496 1676 21548
rect 1728 21536 1734 21548
rect 1763 21539 1821 21545
rect 1763 21536 1775 21539
rect 1728 21508 1775 21536
rect 1728 21496 1734 21508
rect 1763 21505 1775 21508
rect 1809 21536 1821 21539
rect 2406 21536 2412 21548
rect 1809 21508 2412 21536
rect 1809 21505 1821 21508
rect 1763 21499 1821 21505
rect 2406 21496 2412 21508
rect 2464 21496 2470 21548
rect 3068 21545 3096 21576
rect 3804 21548 3832 21576
rect 3878 21564 3884 21616
rect 3936 21604 3942 21616
rect 4080 21604 4108 21635
rect 4890 21632 4896 21684
rect 4948 21632 4954 21684
rect 5534 21632 5540 21684
rect 5592 21672 5598 21684
rect 5629 21675 5687 21681
rect 5629 21672 5641 21675
rect 5592 21644 5641 21672
rect 5592 21632 5598 21644
rect 5629 21641 5641 21644
rect 5675 21641 5687 21675
rect 5629 21635 5687 21641
rect 7650 21632 7656 21684
rect 7708 21672 7714 21684
rect 8021 21675 8079 21681
rect 8021 21672 8033 21675
rect 7708 21644 8033 21672
rect 7708 21632 7714 21644
rect 8021 21641 8033 21644
rect 8067 21641 8079 21675
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 8021 21635 8079 21641
rect 8128 21644 9137 21672
rect 4908 21604 4936 21632
rect 5074 21604 5080 21616
rect 3936 21576 4108 21604
rect 4632 21576 5080 21604
rect 3936 21564 3942 21576
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21505 3111 21539
rect 3053 21499 3111 21505
rect 3234 21496 3240 21548
rect 3292 21536 3298 21548
rect 3327 21539 3385 21545
rect 3327 21536 3339 21539
rect 3292 21508 3339 21536
rect 3292 21496 3298 21508
rect 3327 21505 3339 21508
rect 3373 21505 3385 21539
rect 3327 21499 3385 21505
rect 3786 21496 3792 21548
rect 3844 21536 3850 21548
rect 4154 21536 4160 21548
rect 3844 21508 4160 21536
rect 3844 21496 3850 21508
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4430 21496 4436 21548
rect 4488 21536 4494 21548
rect 4632 21545 4660 21576
rect 5074 21564 5080 21576
rect 5132 21564 5138 21616
rect 7742 21604 7748 21616
rect 6654 21576 7748 21604
rect 6654 21575 6682 21576
rect 6623 21569 6682 21575
rect 4617 21539 4675 21545
rect 4617 21536 4629 21539
rect 4488 21508 4629 21536
rect 4488 21496 4494 21508
rect 4617 21505 4629 21508
rect 4663 21505 4675 21539
rect 4617 21499 4675 21505
rect 4891 21539 4949 21545
rect 4891 21505 4903 21539
rect 4937 21536 4949 21539
rect 5442 21536 5448 21548
rect 4937 21508 5448 21536
rect 4937 21505 4949 21508
rect 4891 21499 4949 21505
rect 5442 21496 5448 21508
rect 5500 21496 5506 21548
rect 6623 21535 6635 21569
rect 6669 21538 6682 21569
rect 7742 21564 7748 21576
rect 7800 21564 7806 21616
rect 8128 21604 8156 21644
rect 9125 21641 9137 21644
rect 9171 21641 9183 21675
rect 9125 21635 9183 21641
rect 10410 21632 10416 21684
rect 10468 21672 10474 21684
rect 11422 21672 11428 21684
rect 10468 21644 11428 21672
rect 10468 21632 10474 21644
rect 11422 21632 11428 21644
rect 11480 21632 11486 21684
rect 12986 21672 12992 21684
rect 12268 21644 12992 21672
rect 7852 21576 8156 21604
rect 6669 21535 6681 21538
rect 6623 21529 6681 21535
rect 6730 21496 6736 21548
rect 6788 21536 6794 21548
rect 7852 21536 7880 21576
rect 8202 21564 8208 21616
rect 8260 21604 8266 21616
rect 8297 21607 8355 21613
rect 8297 21604 8309 21607
rect 8260 21576 8309 21604
rect 8260 21564 8266 21576
rect 8297 21573 8309 21576
rect 8343 21573 8355 21607
rect 8297 21567 8355 21573
rect 8389 21607 8447 21613
rect 8389 21573 8401 21607
rect 8435 21604 8447 21607
rect 9030 21604 9036 21616
rect 8435 21576 9036 21604
rect 8435 21573 8447 21576
rect 8389 21567 8447 21573
rect 9030 21564 9036 21576
rect 9088 21564 9094 21616
rect 12268 21604 12296 21644
rect 12986 21632 12992 21644
rect 13044 21632 13050 21684
rect 13814 21632 13820 21684
rect 13872 21632 13878 21684
rect 16758 21632 16764 21684
rect 16816 21672 16822 21684
rect 17218 21672 17224 21684
rect 16816 21644 17224 21672
rect 16816 21632 16822 21644
rect 17218 21632 17224 21644
rect 17276 21632 17282 21684
rect 18322 21632 18328 21684
rect 18380 21632 18386 21684
rect 20441 21675 20499 21681
rect 20441 21641 20453 21675
rect 20487 21672 20499 21675
rect 21266 21672 21272 21684
rect 20487 21644 21272 21672
rect 20487 21641 20499 21644
rect 20441 21635 20499 21641
rect 21266 21632 21272 21644
rect 21324 21632 21330 21684
rect 10302 21576 12296 21604
rect 6788 21508 7880 21536
rect 8757 21539 8815 21545
rect 6788 21496 6794 21508
rect 8757 21505 8769 21539
rect 8803 21536 8815 21539
rect 8846 21536 8852 21548
rect 8803 21508 8852 21536
rect 8803 21505 8815 21508
rect 8757 21499 8815 21505
rect 8846 21496 8852 21508
rect 8904 21496 8910 21548
rect 9490 21496 9496 21548
rect 9548 21536 9554 21548
rect 10302 21545 10330 21576
rect 10287 21539 10345 21545
rect 10287 21536 10299 21539
rect 9548 21508 10299 21536
rect 9548 21496 9554 21508
rect 10287 21505 10299 21508
rect 10333 21505 10345 21539
rect 10287 21499 10345 21505
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 13078 21496 13084 21548
rect 13136 21545 13142 21548
rect 13136 21539 13164 21545
rect 13152 21505 13164 21539
rect 13136 21499 13164 21505
rect 13136 21496 13142 21499
rect 13262 21496 13268 21548
rect 13320 21496 13326 21548
rect 13832 21536 13860 21632
rect 18340 21604 18368 21632
rect 18340 21576 18828 21604
rect 14001 21539 14059 21545
rect 14001 21536 14013 21539
rect 13832 21508 14013 21536
rect 14001 21505 14013 21508
rect 14047 21505 14059 21539
rect 14001 21499 14059 21505
rect 14182 21496 14188 21548
rect 14240 21496 14246 21548
rect 15010 21496 15016 21548
rect 15068 21545 15074 21548
rect 18800 21545 18828 21576
rect 18874 21564 18880 21616
rect 18932 21604 18938 21616
rect 18932 21576 19564 21604
rect 18932 21564 18938 21576
rect 15068 21539 15096 21545
rect 15084 21505 15096 21539
rect 15068 21499 15096 21505
rect 15841 21539 15899 21545
rect 15841 21505 15853 21539
rect 15887 21536 15899 21539
rect 16117 21539 16175 21545
rect 16117 21536 16129 21539
rect 15887 21508 16129 21536
rect 15887 21505 15899 21508
rect 15841 21499 15899 21505
rect 16117 21505 16129 21508
rect 16163 21505 16175 21539
rect 17555 21539 17613 21545
rect 17555 21536 17567 21539
rect 16117 21499 16175 21505
rect 16224 21508 17567 21536
rect 15068 21496 15074 21499
rect 2314 21428 2320 21480
rect 2372 21468 2378 21480
rect 2498 21468 2504 21480
rect 2372 21440 2504 21468
rect 2372 21428 2378 21440
rect 2498 21428 2504 21440
rect 2556 21428 2562 21480
rect 6365 21471 6423 21477
rect 6365 21437 6377 21471
rect 6411 21437 6423 21471
rect 6365 21431 6423 21437
rect 14 21360 20 21412
rect 72 21400 78 21412
rect 1210 21400 1216 21412
rect 72 21372 1216 21400
rect 72 21360 78 21372
rect 1210 21360 1216 21372
rect 1268 21360 1274 21412
rect 382 21292 388 21344
rect 440 21332 446 21344
rect 1026 21332 1032 21344
rect 440 21304 1032 21332
rect 440 21292 446 21304
rect 1026 21292 1032 21304
rect 1084 21292 1090 21344
rect 1946 21292 1952 21344
rect 2004 21332 2010 21344
rect 3326 21332 3332 21344
rect 2004 21304 3332 21332
rect 2004 21292 2010 21304
rect 3326 21292 3332 21304
rect 3384 21292 3390 21344
rect 4614 21292 4620 21344
rect 4672 21332 4678 21344
rect 6380 21332 6408 21431
rect 8202 21428 8208 21480
rect 8260 21428 8266 21480
rect 9398 21428 9404 21480
rect 9456 21468 9462 21480
rect 9950 21468 9956 21480
rect 9456 21440 9956 21468
rect 9456 21428 9462 21440
rect 9950 21428 9956 21440
rect 10008 21428 10014 21480
rect 10042 21428 10048 21480
rect 10100 21428 10106 21480
rect 11974 21468 11980 21480
rect 10702 21440 11980 21468
rect 9306 21360 9312 21412
rect 9364 21360 9370 21412
rect 7282 21332 7288 21344
rect 4672 21304 7288 21332
rect 4672 21292 4678 21304
rect 7282 21292 7288 21304
rect 7340 21292 7346 21344
rect 7374 21292 7380 21344
rect 7432 21292 7438 21344
rect 9950 21292 9956 21344
rect 10008 21332 10014 21344
rect 10702 21332 10730 21440
rect 11974 21428 11980 21440
rect 12032 21468 12038 21480
rect 12253 21471 12311 21477
rect 12253 21468 12265 21471
rect 12032 21440 12265 21468
rect 12032 21428 12038 21440
rect 12253 21437 12265 21440
rect 12299 21437 12311 21471
rect 12253 21431 12311 21437
rect 12986 21428 12992 21480
rect 13044 21428 13050 21480
rect 14921 21471 14979 21477
rect 14921 21468 14933 21471
rect 13648 21440 14933 21468
rect 11057 21403 11115 21409
rect 11057 21369 11069 21403
rect 11103 21400 11115 21403
rect 12066 21400 12072 21412
rect 11103 21372 12072 21400
rect 11103 21369 11115 21372
rect 11057 21363 11115 21369
rect 12066 21360 12072 21372
rect 12124 21360 12130 21412
rect 12710 21360 12716 21412
rect 12768 21360 12774 21412
rect 10008 21304 10730 21332
rect 10008 21292 10014 21304
rect 11790 21292 11796 21344
rect 11848 21332 11854 21344
rect 11977 21335 12035 21341
rect 11977 21332 11989 21335
rect 11848 21304 11989 21332
rect 11848 21292 11854 21304
rect 11977 21301 11989 21304
rect 12023 21301 12035 21335
rect 11977 21295 12035 21301
rect 12434 21292 12440 21344
rect 12492 21332 12498 21344
rect 13648 21332 13676 21440
rect 14921 21437 14933 21440
rect 14967 21437 14979 21471
rect 14921 21431 14979 21437
rect 15197 21471 15255 21477
rect 15197 21437 15209 21471
rect 15243 21468 15255 21471
rect 15378 21468 15384 21480
rect 15243 21440 15384 21468
rect 15243 21437 15255 21440
rect 15197 21431 15255 21437
rect 15378 21428 15384 21440
rect 15436 21428 15442 21480
rect 16224 21468 16252 21508
rect 17555 21505 17567 21508
rect 17601 21505 17613 21539
rect 18693 21539 18751 21545
rect 18693 21536 18705 21539
rect 17555 21499 17613 21505
rect 18340 21508 18705 21536
rect 15856 21440 16252 21468
rect 17313 21471 17371 21477
rect 14645 21403 14703 21409
rect 14645 21369 14657 21403
rect 14691 21369 14703 21403
rect 14645 21363 14703 21369
rect 12492 21304 13676 21332
rect 12492 21292 12498 21304
rect 13722 21292 13728 21344
rect 13780 21332 13786 21344
rect 13909 21335 13967 21341
rect 13909 21332 13921 21335
rect 13780 21304 13921 21332
rect 13780 21292 13786 21304
rect 13909 21301 13921 21304
rect 13955 21301 13967 21335
rect 13909 21295 13967 21301
rect 14458 21292 14464 21344
rect 14516 21332 14522 21344
rect 14660 21332 14688 21363
rect 14516 21304 14688 21332
rect 14516 21292 14522 21304
rect 14918 21292 14924 21344
rect 14976 21332 14982 21344
rect 15856 21332 15884 21440
rect 17313 21437 17325 21471
rect 17359 21437 17371 21471
rect 17313 21431 17371 21437
rect 14976 21304 15884 21332
rect 14976 21292 14982 21304
rect 15930 21292 15936 21344
rect 15988 21292 15994 21344
rect 17328 21332 17356 21431
rect 18340 21409 18368 21508
rect 18693 21505 18705 21508
rect 18739 21505 18751 21539
rect 18693 21499 18751 21505
rect 18785 21539 18843 21545
rect 18785 21505 18797 21539
rect 18831 21505 18843 21539
rect 19061 21539 19119 21545
rect 19061 21536 19073 21539
rect 18785 21499 18843 21505
rect 18892 21508 19073 21536
rect 18708 21468 18736 21499
rect 18892 21468 18920 21508
rect 19061 21505 19073 21508
rect 19107 21505 19119 21539
rect 19061 21499 19119 21505
rect 19242 21496 19248 21548
rect 19300 21496 19306 21548
rect 19536 21545 19564 21576
rect 20162 21564 20168 21616
rect 20220 21564 20226 21616
rect 19521 21539 19579 21545
rect 19521 21505 19533 21539
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 19705 21539 19763 21545
rect 19705 21505 19717 21539
rect 19751 21536 19763 21539
rect 20530 21536 20536 21548
rect 19751 21508 20536 21536
rect 19751 21505 19763 21508
rect 19705 21499 19763 21505
rect 20530 21496 20536 21508
rect 20588 21496 20594 21548
rect 18708 21440 18920 21468
rect 18969 21471 19027 21477
rect 18969 21437 18981 21471
rect 19015 21468 19027 21471
rect 19153 21471 19211 21477
rect 19153 21468 19165 21471
rect 19015 21440 19165 21468
rect 19015 21437 19027 21440
rect 18969 21431 19027 21437
rect 19153 21437 19165 21440
rect 19199 21437 19211 21471
rect 19153 21431 19211 21437
rect 19334 21428 19340 21480
rect 19392 21468 19398 21480
rect 20438 21468 20444 21480
rect 19392 21440 20444 21468
rect 19392 21428 19398 21440
rect 20438 21428 20444 21440
rect 20496 21428 20502 21480
rect 18325 21403 18383 21409
rect 18325 21369 18337 21403
rect 18371 21369 18383 21403
rect 18325 21363 18383 21369
rect 18138 21332 18144 21344
rect 17328 21304 18144 21332
rect 18138 21292 18144 21304
rect 18196 21292 18202 21344
rect 18877 21335 18935 21341
rect 18877 21301 18889 21335
rect 18923 21332 18935 21335
rect 19242 21332 19248 21344
rect 18923 21304 19248 21332
rect 18923 21301 18935 21304
rect 18877 21295 18935 21301
rect 19242 21292 19248 21304
rect 19300 21292 19306 21344
rect 19334 21292 19340 21344
rect 19392 21292 19398 21344
rect 19886 21292 19892 21344
rect 19944 21292 19950 21344
rect 1104 21242 20884 21264
rect 1104 21190 3422 21242
rect 3474 21190 3486 21242
rect 3538 21190 3550 21242
rect 3602 21190 3614 21242
rect 3666 21190 3678 21242
rect 3730 21190 8367 21242
rect 8419 21190 8431 21242
rect 8483 21190 8495 21242
rect 8547 21190 8559 21242
rect 8611 21190 8623 21242
rect 8675 21190 13312 21242
rect 13364 21190 13376 21242
rect 13428 21190 13440 21242
rect 13492 21190 13504 21242
rect 13556 21190 13568 21242
rect 13620 21190 18257 21242
rect 18309 21190 18321 21242
rect 18373 21190 18385 21242
rect 18437 21190 18449 21242
rect 18501 21190 18513 21242
rect 18565 21190 20884 21242
rect 1104 21168 20884 21190
rect 3804 21100 4844 21128
rect 3145 21063 3203 21069
rect 3145 21029 3157 21063
rect 3191 21060 3203 21063
rect 3694 21060 3700 21072
rect 3191 21032 3700 21060
rect 3191 21029 3203 21032
rect 3145 21023 3203 21029
rect 3694 21020 3700 21032
rect 3752 21020 3758 21072
rect 3804 20992 3832 21100
rect 4816 21069 4844 21100
rect 7374 21088 7380 21140
rect 7432 21088 7438 21140
rect 8202 21088 8208 21140
rect 8260 21128 8266 21140
rect 8481 21131 8539 21137
rect 8481 21128 8493 21131
rect 8260 21100 8493 21128
rect 8260 21088 8266 21100
rect 8481 21097 8493 21100
rect 8527 21097 8539 21131
rect 8481 21091 8539 21097
rect 9030 21088 9036 21140
rect 9088 21128 9094 21140
rect 9953 21131 10011 21137
rect 9953 21128 9965 21131
rect 9088 21100 9965 21128
rect 9088 21088 9094 21100
rect 9953 21097 9965 21100
rect 9999 21097 10011 21131
rect 9953 21091 10011 21097
rect 11330 21088 11336 21140
rect 11388 21128 11394 21140
rect 12434 21128 12440 21140
rect 11388 21100 12440 21128
rect 11388 21088 11394 21100
rect 12434 21088 12440 21100
rect 12492 21088 12498 21140
rect 12986 21088 12992 21140
rect 13044 21128 13050 21140
rect 13173 21131 13231 21137
rect 13173 21128 13185 21131
rect 13044 21100 13185 21128
rect 13044 21088 13050 21100
rect 13173 21097 13185 21100
rect 13219 21097 13231 21131
rect 13173 21091 13231 21097
rect 15930 21088 15936 21140
rect 15988 21088 15994 21140
rect 17034 21088 17040 21140
rect 17092 21128 17098 21140
rect 17092 21100 18368 21128
rect 17092 21088 17098 21100
rect 4801 21063 4859 21069
rect 4801 21029 4813 21063
rect 4847 21029 4859 21063
rect 4801 21023 4859 21029
rect 2898 20964 3832 20992
rect 5828 20936 5856 20978
rect 1581 20927 1639 20933
rect 1581 20893 1593 20927
rect 1627 20924 1639 20927
rect 2133 20927 2191 20933
rect 2133 20924 2145 20927
rect 1627 20896 2145 20924
rect 1627 20893 1639 20896
rect 1581 20887 1639 20893
rect 2133 20893 2145 20896
rect 2179 20893 2191 20927
rect 2133 20887 2191 20893
rect 3329 20927 3387 20933
rect 3329 20893 3341 20927
rect 3375 20924 3387 20927
rect 3418 20924 3424 20936
rect 3375 20896 3424 20924
rect 3375 20893 3387 20896
rect 3329 20887 3387 20893
rect 3418 20884 3424 20896
rect 3476 20884 3482 20936
rect 3602 20884 3608 20936
rect 3660 20924 3666 20936
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 3660 20896 3801 20924
rect 3660 20884 3666 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 4031 20927 4089 20933
rect 4031 20924 4043 20927
rect 3789 20887 3847 20893
rect 3896 20896 4043 20924
rect 290 20816 296 20868
rect 348 20856 354 20868
rect 1118 20856 1124 20868
rect 348 20828 1124 20856
rect 348 20816 354 20828
rect 1118 20816 1124 20828
rect 1176 20856 1182 20868
rect 1857 20859 1915 20865
rect 1857 20856 1869 20859
rect 1176 20828 1869 20856
rect 1176 20816 1182 20828
rect 1857 20825 1869 20828
rect 1903 20825 1915 20859
rect 1857 20819 1915 20825
rect 2222 20816 2228 20868
rect 2280 20816 2286 20868
rect 2498 20816 2504 20868
rect 2556 20856 2562 20868
rect 2593 20859 2651 20865
rect 2593 20856 2605 20859
rect 2556 20828 2605 20856
rect 2556 20816 2562 20828
rect 2593 20825 2605 20828
rect 2639 20825 2651 20859
rect 2593 20819 2651 20825
rect 2961 20859 3019 20865
rect 2961 20825 2973 20859
rect 3007 20856 3019 20859
rect 3050 20856 3056 20868
rect 3007 20828 3056 20856
rect 3007 20825 3019 20828
rect 2961 20819 3019 20825
rect 3050 20816 3056 20828
rect 3108 20816 3114 20868
rect 3896 20856 3924 20896
rect 4031 20893 4043 20896
rect 4077 20893 4089 20927
rect 4031 20887 4089 20893
rect 4890 20884 4896 20936
rect 4948 20924 4954 20936
rect 5166 20924 5172 20936
rect 4948 20896 5172 20924
rect 4948 20884 4954 20896
rect 5166 20884 5172 20896
rect 5224 20884 5230 20936
rect 5810 20884 5816 20936
rect 5868 20884 5874 20936
rect 5902 20884 5908 20936
rect 5960 20924 5966 20936
rect 5997 20927 6055 20933
rect 5997 20924 6009 20927
rect 5960 20896 6009 20924
rect 5960 20884 5966 20896
rect 5997 20893 6009 20896
rect 6043 20893 6055 20927
rect 5997 20887 6055 20893
rect 6089 20927 6147 20933
rect 6089 20893 6101 20927
rect 6135 20924 6147 20927
rect 7392 20924 7420 21088
rect 10502 21020 10508 21072
rect 10560 21060 10566 21072
rect 10560 21032 11652 21060
rect 10560 21020 10566 21032
rect 10594 20952 10600 21004
rect 10652 20992 10658 21004
rect 10873 20995 10931 21001
rect 10873 20992 10885 20995
rect 10652 20964 10885 20992
rect 10652 20952 10658 20964
rect 10873 20961 10885 20964
rect 10919 20961 10931 20995
rect 11422 20992 11428 21004
rect 10873 20955 10931 20961
rect 11072 20964 11428 20992
rect 11072 20936 11100 20964
rect 11422 20952 11428 20964
rect 11480 20952 11486 21004
rect 11514 20952 11520 21004
rect 11572 20952 11578 21004
rect 11624 20992 11652 21032
rect 13538 21020 13544 21072
rect 13596 21060 13602 21072
rect 13596 21032 14320 21060
rect 13596 21020 13602 21032
rect 14292 21001 14320 21032
rect 14642 21020 14648 21072
rect 14700 21060 14706 21072
rect 14700 21032 14872 21060
rect 14700 21020 14706 21032
rect 11910 20995 11968 21001
rect 11910 20992 11922 20995
rect 11624 20964 11922 20992
rect 11910 20961 11922 20964
rect 11956 20992 11968 20995
rect 14277 20995 14335 21001
rect 11956 20964 14044 20992
rect 11956 20961 11968 20964
rect 11910 20955 11968 20961
rect 6135 20896 7420 20924
rect 7469 20927 7527 20933
rect 6135 20893 6147 20896
rect 6089 20887 6147 20893
rect 7469 20893 7481 20927
rect 7515 20893 7527 20927
rect 7469 20887 7527 20893
rect 7743 20927 7801 20933
rect 7743 20893 7755 20927
rect 7789 20924 7801 20927
rect 8662 20924 8668 20936
rect 7789 20896 8668 20924
rect 7789 20893 7801 20896
rect 7743 20887 7801 20893
rect 3436 20828 3924 20856
rect 2866 20748 2872 20800
rect 2924 20788 2930 20800
rect 3436 20788 3464 20828
rect 4246 20816 4252 20868
rect 4304 20816 4310 20868
rect 4982 20816 4988 20868
rect 5040 20856 5046 20868
rect 5040 20828 5854 20856
rect 5040 20816 5046 20828
rect 2924 20760 3464 20788
rect 3513 20791 3571 20797
rect 2924 20748 2930 20760
rect 3513 20757 3525 20791
rect 3559 20788 3571 20791
rect 4062 20788 4068 20800
rect 3559 20760 4068 20788
rect 3559 20757 3571 20760
rect 3513 20751 3571 20757
rect 4062 20748 4068 20760
rect 4120 20748 4126 20800
rect 4264 20788 4292 20816
rect 5721 20791 5779 20797
rect 5721 20788 5733 20791
rect 4264 20760 5733 20788
rect 5721 20757 5733 20760
rect 5767 20757 5779 20791
rect 5826 20788 5854 20828
rect 6362 20816 6368 20868
rect 6420 20856 6426 20868
rect 6457 20859 6515 20865
rect 6457 20856 6469 20859
rect 6420 20828 6469 20856
rect 6420 20816 6426 20828
rect 6457 20825 6469 20828
rect 6503 20825 6515 20859
rect 6457 20819 6515 20825
rect 7282 20816 7288 20868
rect 7340 20856 7346 20868
rect 7484 20856 7512 20887
rect 8662 20884 8668 20896
rect 8720 20884 8726 20936
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20924 8999 20927
rect 9215 20927 9273 20933
rect 8987 20896 9076 20924
rect 8987 20893 8999 20896
rect 8941 20887 8999 20893
rect 9048 20868 9076 20896
rect 9215 20893 9227 20927
rect 9261 20924 9273 20927
rect 9261 20896 11008 20924
rect 9261 20893 9273 20896
rect 9215 20887 9273 20893
rect 8754 20856 8760 20868
rect 7340 20828 8760 20856
rect 7340 20816 7346 20828
rect 8754 20816 8760 20828
rect 8812 20856 8818 20868
rect 9030 20856 9036 20868
rect 8812 20828 9036 20856
rect 8812 20816 8818 20828
rect 9030 20816 9036 20828
rect 9088 20816 9094 20868
rect 10980 20856 11008 20896
rect 11054 20884 11060 20936
rect 11112 20884 11118 20936
rect 11790 20884 11796 20936
rect 11848 20933 11854 20936
rect 11848 20927 11869 20933
rect 11857 20893 11869 20927
rect 11848 20887 11869 20893
rect 11848 20884 11854 20887
rect 12066 20884 12072 20936
rect 12124 20884 12130 20936
rect 12713 20927 12771 20933
rect 12713 20893 12725 20927
rect 12759 20924 12771 20927
rect 13538 20924 13544 20936
rect 12759 20896 13544 20924
rect 12759 20893 12771 20896
rect 12713 20887 12771 20893
rect 13538 20884 13544 20896
rect 13596 20884 13602 20936
rect 10980 20828 11098 20856
rect 6825 20791 6883 20797
rect 6825 20788 6837 20791
rect 5826 20760 6837 20788
rect 5721 20751 5779 20757
rect 6825 20757 6837 20760
rect 6871 20757 6883 20791
rect 6825 20751 6883 20757
rect 7009 20791 7067 20797
rect 7009 20757 7021 20791
rect 7055 20788 7067 20791
rect 8018 20788 8024 20800
rect 7055 20760 8024 20788
rect 7055 20757 7067 20760
rect 7009 20751 7067 20757
rect 8018 20748 8024 20760
rect 8076 20748 8082 20800
rect 8202 20748 8208 20800
rect 8260 20788 8266 20800
rect 10962 20788 10968 20800
rect 8260 20760 10968 20788
rect 8260 20748 8266 20760
rect 10962 20748 10968 20760
rect 11020 20748 11026 20800
rect 11070 20788 11098 20828
rect 12158 20788 12164 20800
rect 11070 20760 12164 20788
rect 12158 20748 12164 20760
rect 12216 20788 12222 20800
rect 12618 20788 12624 20800
rect 12216 20760 12624 20788
rect 12216 20748 12222 20760
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 13078 20748 13084 20800
rect 13136 20788 13142 20800
rect 13814 20788 13820 20800
rect 13136 20760 13820 20788
rect 13136 20748 13142 20760
rect 13814 20748 13820 20760
rect 13872 20748 13878 20800
rect 14016 20788 14044 20964
rect 14277 20961 14289 20995
rect 14323 20961 14335 20995
rect 14737 20995 14795 21001
rect 14737 20992 14749 20995
rect 14277 20955 14335 20961
rect 14476 20964 14749 20992
rect 14090 20884 14096 20936
rect 14148 20884 14154 20936
rect 14182 20816 14188 20868
rect 14240 20856 14246 20868
rect 14292 20856 14320 20955
rect 14476 20936 14504 20964
rect 14737 20961 14749 20964
rect 14783 20961 14795 20995
rect 14844 20992 14872 21032
rect 15130 20995 15188 21001
rect 15130 20992 15142 20995
rect 14844 20964 15142 20992
rect 14737 20955 14795 20961
rect 15130 20961 15142 20964
rect 15176 20961 15188 20995
rect 15948 20992 15976 21088
rect 18340 21060 18368 21100
rect 18414 21088 18420 21140
rect 18472 21128 18478 21140
rect 19702 21128 19708 21140
rect 18472 21100 19708 21128
rect 18472 21088 18478 21100
rect 19702 21088 19708 21100
rect 19760 21088 19766 21140
rect 19886 21060 19892 21072
rect 18340 21032 19892 21060
rect 19886 21020 19892 21032
rect 19944 21020 19950 21072
rect 19334 20992 19340 21004
rect 15948 20964 16712 20992
rect 15130 20955 15188 20961
rect 14458 20884 14464 20936
rect 14516 20884 14522 20936
rect 15010 20884 15016 20936
rect 15068 20884 15074 20936
rect 15286 20884 15292 20936
rect 15344 20884 15350 20936
rect 16209 20927 16267 20933
rect 16209 20893 16221 20927
rect 16255 20893 16267 20927
rect 16209 20887 16267 20893
rect 14240 20828 14320 20856
rect 14240 20816 14246 20828
rect 15010 20788 15016 20800
rect 14016 20760 15016 20788
rect 15010 20748 15016 20760
rect 15068 20748 15074 20800
rect 15933 20791 15991 20797
rect 15933 20757 15945 20791
rect 15979 20788 15991 20791
rect 16114 20788 16120 20800
rect 15979 20760 16120 20788
rect 15979 20757 15991 20760
rect 15933 20751 15991 20757
rect 16114 20748 16120 20760
rect 16172 20748 16178 20800
rect 16224 20788 16252 20887
rect 16390 20884 16396 20936
rect 16448 20884 16454 20936
rect 16684 20933 16712 20964
rect 18616 20964 19340 20992
rect 18616 20933 18644 20964
rect 19334 20952 19340 20964
rect 19392 20952 19398 21004
rect 20346 20952 20352 21004
rect 20404 20992 20410 21004
rect 21726 20992 21732 21004
rect 20404 20964 21732 20992
rect 20404 20952 20410 20964
rect 21726 20952 21732 20964
rect 21784 20952 21790 21004
rect 16669 20927 16727 20933
rect 16669 20893 16681 20927
rect 16715 20893 16727 20927
rect 16669 20887 16727 20893
rect 18601 20927 18659 20933
rect 18601 20893 18613 20927
rect 18647 20893 18659 20927
rect 18601 20887 18659 20893
rect 18874 20884 18880 20936
rect 18932 20884 18938 20936
rect 18966 20884 18972 20936
rect 19024 20924 19030 20936
rect 19061 20927 19119 20933
rect 19061 20924 19073 20927
rect 19024 20896 19073 20924
rect 19024 20884 19030 20896
rect 19061 20893 19073 20896
rect 19107 20893 19119 20927
rect 19061 20887 19119 20893
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 19978 20884 19984 20936
rect 20036 20884 20042 20936
rect 16482 20816 16488 20868
rect 16540 20816 16546 20868
rect 16574 20816 16580 20868
rect 16632 20816 16638 20868
rect 18693 20859 18751 20865
rect 18693 20825 18705 20859
rect 18739 20856 18751 20859
rect 19334 20856 19340 20868
rect 18739 20828 19340 20856
rect 18739 20825 18751 20828
rect 18693 20819 18751 20825
rect 19334 20816 19340 20828
rect 19392 20816 19398 20868
rect 19797 20859 19855 20865
rect 19797 20825 19809 20859
rect 19843 20856 19855 20859
rect 21266 20856 21272 20868
rect 19843 20828 21272 20856
rect 19843 20825 19855 20828
rect 19797 20819 19855 20825
rect 21266 20816 21272 20828
rect 21324 20816 21330 20868
rect 16761 20791 16819 20797
rect 16761 20788 16773 20791
rect 16224 20760 16773 20788
rect 16761 20757 16773 20760
rect 16807 20757 16819 20791
rect 16761 20751 16819 20757
rect 17126 20748 17132 20800
rect 17184 20788 17190 20800
rect 17494 20788 17500 20800
rect 17184 20760 17500 20788
rect 17184 20748 17190 20760
rect 17494 20748 17500 20760
rect 17552 20748 17558 20800
rect 19061 20791 19119 20797
rect 19061 20757 19073 20791
rect 19107 20788 19119 20791
rect 19702 20788 19708 20800
rect 19107 20760 19708 20788
rect 19107 20757 19119 20760
rect 19061 20751 19119 20757
rect 19702 20748 19708 20760
rect 19760 20748 19766 20800
rect 20257 20791 20315 20797
rect 20257 20757 20269 20791
rect 20303 20788 20315 20791
rect 21542 20788 21548 20800
rect 20303 20760 21548 20788
rect 20303 20757 20315 20760
rect 20257 20751 20315 20757
rect 21542 20748 21548 20760
rect 21600 20748 21606 20800
rect 1104 20698 21043 20720
rect 1104 20646 5894 20698
rect 5946 20646 5958 20698
rect 6010 20646 6022 20698
rect 6074 20646 6086 20698
rect 6138 20646 6150 20698
rect 6202 20646 10839 20698
rect 10891 20646 10903 20698
rect 10955 20646 10967 20698
rect 11019 20646 11031 20698
rect 11083 20646 11095 20698
rect 11147 20646 15784 20698
rect 15836 20646 15848 20698
rect 15900 20646 15912 20698
rect 15964 20646 15976 20698
rect 16028 20646 16040 20698
rect 16092 20646 20729 20698
rect 20781 20646 20793 20698
rect 20845 20646 20857 20698
rect 20909 20646 20921 20698
rect 20973 20646 20985 20698
rect 21037 20646 21043 20698
rect 1104 20624 21043 20646
rect 1578 20544 1584 20596
rect 1636 20584 1642 20596
rect 1854 20584 1860 20596
rect 1636 20556 1860 20584
rect 1636 20544 1642 20556
rect 1854 20544 1860 20556
rect 1912 20544 1918 20596
rect 2222 20544 2228 20596
rect 2280 20584 2286 20596
rect 2593 20587 2651 20593
rect 2593 20584 2605 20587
rect 2280 20556 2605 20584
rect 2280 20544 2286 20556
rect 2593 20553 2605 20556
rect 2639 20553 2651 20587
rect 3602 20584 3608 20596
rect 2593 20547 2651 20553
rect 2700 20556 3608 20584
rect 2700 20516 2728 20556
rect 3602 20544 3608 20556
rect 3660 20584 3666 20596
rect 3660 20556 5654 20584
rect 3660 20544 3666 20556
rect 3878 20516 3884 20528
rect 1596 20488 2728 20516
rect 3434 20488 3884 20516
rect 1596 20457 1624 20488
rect 1581 20451 1639 20457
rect 1581 20417 1593 20451
rect 1627 20417 1639 20451
rect 1854 20448 1860 20460
rect 1815 20420 1860 20448
rect 1581 20411 1639 20417
rect 1854 20408 1860 20420
rect 1912 20408 1918 20460
rect 3434 20457 3462 20488
rect 3878 20476 3884 20488
rect 3936 20516 3942 20528
rect 4614 20516 4620 20528
rect 3936 20488 4620 20516
rect 3936 20476 3942 20488
rect 4614 20476 4620 20488
rect 4672 20476 4678 20528
rect 5626 20516 5654 20556
rect 6730 20544 6736 20596
rect 6788 20584 6794 20596
rect 8294 20584 8300 20596
rect 6788 20556 8300 20584
rect 6788 20544 6794 20556
rect 8294 20544 8300 20556
rect 8352 20584 8358 20596
rect 11606 20584 11612 20596
rect 8352 20556 11612 20584
rect 8352 20544 8358 20556
rect 11606 20544 11612 20556
rect 11664 20584 11670 20596
rect 11664 20556 11986 20584
rect 11664 20544 11670 20556
rect 5182 20488 5598 20516
rect 5626 20488 7512 20516
rect 3419 20451 3477 20457
rect 3419 20417 3431 20451
rect 3465 20417 3477 20451
rect 3419 20411 3477 20417
rect 3510 20408 3516 20460
rect 3568 20448 3574 20460
rect 4525 20451 4583 20457
rect 4525 20448 4537 20451
rect 3568 20420 4537 20448
rect 3568 20408 3574 20420
rect 4525 20417 4537 20420
rect 4571 20417 4583 20451
rect 4525 20411 4583 20417
rect 4706 20408 4712 20460
rect 4764 20448 4770 20460
rect 5182 20457 5210 20488
rect 4893 20451 4951 20457
rect 4893 20448 4905 20451
rect 4764 20420 4905 20448
rect 4764 20408 4770 20420
rect 4893 20417 4905 20420
rect 4939 20417 4951 20451
rect 4893 20411 4951 20417
rect 5167 20451 5225 20457
rect 5167 20417 5179 20451
rect 5213 20417 5225 20451
rect 5167 20411 5225 20417
rect 3145 20383 3203 20389
rect 3145 20349 3157 20383
rect 3191 20349 3203 20383
rect 5570 20380 5598 20488
rect 7116 20457 7144 20488
rect 7484 20460 7512 20488
rect 8938 20476 8944 20528
rect 8996 20516 9002 20528
rect 10870 20516 10876 20528
rect 8996 20488 10876 20516
rect 8996 20476 9002 20488
rect 10870 20476 10876 20488
rect 10928 20476 10934 20528
rect 11790 20476 11796 20528
rect 11848 20476 11854 20528
rect 11958 20487 11986 20556
rect 12710 20544 12716 20596
rect 12768 20544 12774 20596
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 14277 20587 14335 20593
rect 13136 20556 13676 20584
rect 13136 20544 13142 20556
rect 13648 20516 13676 20556
rect 14277 20553 14289 20587
rect 14323 20584 14335 20587
rect 14458 20584 14464 20596
rect 14323 20556 14464 20584
rect 14323 20553 14335 20556
rect 14277 20547 14335 20553
rect 14458 20544 14464 20556
rect 14516 20544 14522 20596
rect 15286 20544 15292 20596
rect 15344 20584 15350 20596
rect 15657 20587 15715 20593
rect 15657 20584 15669 20587
rect 15344 20556 15669 20584
rect 15344 20544 15350 20556
rect 15657 20553 15669 20556
rect 15703 20553 15715 20587
rect 15657 20547 15715 20553
rect 16114 20544 16120 20596
rect 16172 20544 16178 20596
rect 16390 20544 16396 20596
rect 16448 20544 16454 20596
rect 16485 20587 16543 20593
rect 16485 20553 16497 20587
rect 16531 20584 16543 20587
rect 16574 20584 16580 20596
rect 16531 20556 16580 20584
rect 16531 20553 16543 20556
rect 16485 20547 16543 20553
rect 16574 20544 16580 20556
rect 16632 20544 16638 20596
rect 16850 20544 16856 20596
rect 16908 20544 16914 20596
rect 17770 20544 17776 20596
rect 17828 20584 17834 20596
rect 18049 20587 18107 20593
rect 18049 20584 18061 20587
rect 17828 20556 18061 20584
rect 17828 20544 17834 20556
rect 18049 20553 18061 20556
rect 18095 20553 18107 20587
rect 18049 20547 18107 20553
rect 18782 20544 18788 20596
rect 18840 20584 18846 20596
rect 18840 20556 18920 20584
rect 18840 20544 18846 20556
rect 16022 20516 16028 20528
rect 13648 20488 16028 20516
rect 11958 20481 12017 20487
rect 7101 20451 7159 20457
rect 7101 20417 7113 20451
rect 7147 20417 7159 20451
rect 7374 20448 7380 20460
rect 7335 20420 7380 20448
rect 7101 20411 7159 20417
rect 7374 20408 7380 20420
rect 7432 20408 7438 20460
rect 7466 20408 7472 20460
rect 7524 20408 7530 20460
rect 7834 20408 7840 20460
rect 7892 20448 7898 20460
rect 8754 20448 8760 20460
rect 7892 20420 8760 20448
rect 7892 20408 7898 20420
rect 8754 20408 8760 20420
rect 8812 20408 8818 20460
rect 9215 20451 9273 20457
rect 9215 20417 9227 20451
rect 9261 20448 9273 20451
rect 10778 20448 10784 20460
rect 9261 20420 10784 20448
rect 9261 20417 9273 20420
rect 9215 20411 9273 20417
rect 10778 20408 10784 20420
rect 10836 20448 10842 20460
rect 11808 20448 11836 20476
rect 11958 20450 11971 20481
rect 10836 20420 11836 20448
rect 11959 20447 11971 20450
rect 12005 20447 12017 20481
rect 13523 20481 13581 20487
rect 13523 20478 13535 20481
rect 11959 20441 12017 20447
rect 10836 20408 10842 20420
rect 12066 20408 12072 20460
rect 12124 20448 12130 20460
rect 13522 20448 13535 20478
rect 12124 20447 13535 20448
rect 13569 20448 13581 20481
rect 16022 20476 16028 20488
rect 16080 20476 16086 20528
rect 13569 20447 14044 20448
rect 12124 20420 14044 20447
rect 12124 20408 12130 20420
rect 6730 20380 6736 20392
rect 5570 20352 6736 20380
rect 3145 20343 3203 20349
rect 2314 20204 2320 20256
rect 2372 20244 2378 20256
rect 3160 20244 3188 20343
rect 6730 20340 6736 20352
rect 6788 20340 6794 20392
rect 8202 20380 8208 20392
rect 8036 20352 8208 20380
rect 4430 20312 4436 20324
rect 3802 20284 4436 20312
rect 3802 20244 3830 20284
rect 4430 20272 4436 20284
rect 4488 20272 4494 20324
rect 5810 20272 5816 20324
rect 5868 20312 5874 20324
rect 5905 20315 5963 20321
rect 5905 20312 5917 20315
rect 5868 20284 5917 20312
rect 5868 20272 5874 20284
rect 5905 20281 5917 20284
rect 5951 20281 5963 20315
rect 5905 20275 5963 20281
rect 2372 20216 3830 20244
rect 2372 20204 2378 20216
rect 4062 20204 4068 20256
rect 4120 20244 4126 20256
rect 4157 20247 4215 20253
rect 4157 20244 4169 20247
rect 4120 20216 4169 20244
rect 4120 20204 4126 20216
rect 4157 20213 4169 20216
rect 4203 20213 4215 20247
rect 4157 20207 4215 20213
rect 4709 20247 4767 20253
rect 4709 20213 4721 20247
rect 4755 20244 4767 20247
rect 8036 20244 8064 20352
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 8941 20383 8999 20389
rect 8941 20380 8953 20383
rect 8680 20352 8953 20380
rect 8680 20256 8708 20352
rect 8941 20349 8953 20352
rect 8987 20349 8999 20383
rect 8941 20343 8999 20349
rect 10594 20340 10600 20392
rect 10652 20380 10658 20392
rect 11701 20383 11759 20389
rect 11701 20380 11713 20383
rect 10652 20352 11713 20380
rect 10652 20340 10658 20352
rect 11701 20349 11713 20352
rect 11747 20349 11759 20383
rect 11701 20343 11759 20349
rect 4755 20216 8064 20244
rect 8113 20247 8171 20253
rect 4755 20213 4767 20216
rect 4709 20207 4767 20213
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 8202 20244 8208 20256
rect 8159 20216 8208 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 8202 20204 8208 20216
rect 8260 20204 8266 20256
rect 8662 20204 8668 20256
rect 8720 20204 8726 20256
rect 8846 20204 8852 20256
rect 8904 20204 8910 20256
rect 9950 20204 9956 20256
rect 10008 20204 10014 20256
rect 11716 20244 11744 20343
rect 13170 20340 13176 20392
rect 13228 20380 13234 20392
rect 13265 20383 13323 20389
rect 13265 20380 13277 20383
rect 13228 20352 13277 20380
rect 13228 20340 13234 20352
rect 13265 20349 13277 20352
rect 13311 20349 13323 20383
rect 13265 20343 13323 20349
rect 12158 20244 12164 20256
rect 11716 20216 12164 20244
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12526 20204 12532 20256
rect 12584 20244 12590 20256
rect 13078 20244 13084 20256
rect 12584 20216 13084 20244
rect 12584 20204 12590 20216
rect 13078 20204 13084 20216
rect 13136 20204 13142 20256
rect 14016 20244 14044 20420
rect 14090 20408 14096 20460
rect 14148 20448 14154 20460
rect 14458 20448 14464 20460
rect 14148 20420 14464 20448
rect 14148 20408 14154 20420
rect 14458 20408 14464 20420
rect 14516 20408 14522 20460
rect 14918 20448 14924 20460
rect 14879 20420 14924 20448
rect 14918 20408 14924 20420
rect 14976 20408 14982 20460
rect 16132 20448 16160 20544
rect 16209 20451 16267 20457
rect 16209 20448 16221 20451
rect 16132 20420 16221 20448
rect 16209 20417 16221 20420
rect 16255 20417 16267 20451
rect 16209 20411 16267 20417
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20448 16359 20451
rect 16408 20448 16436 20544
rect 16347 20420 16436 20448
rect 16485 20451 16543 20457
rect 16347 20417 16359 20420
rect 16301 20411 16359 20417
rect 16485 20417 16497 20451
rect 16531 20417 16543 20451
rect 16868 20448 16896 20544
rect 18892 20525 18920 20556
rect 18868 20519 18926 20525
rect 18868 20485 18880 20519
rect 18914 20485 18926 20519
rect 18868 20479 18926 20485
rect 19352 20488 20208 20516
rect 19352 20460 19380 20488
rect 16925 20451 16983 20457
rect 16925 20448 16937 20451
rect 16868 20420 16937 20448
rect 16485 20411 16543 20417
rect 16925 20417 16937 20420
rect 16971 20417 16983 20451
rect 16925 20411 16983 20417
rect 14645 20383 14703 20389
rect 14645 20380 14657 20383
rect 14108 20352 14657 20380
rect 14108 20324 14136 20352
rect 14645 20349 14657 20352
rect 14691 20349 14703 20383
rect 16500 20380 16528 20411
rect 17494 20408 17500 20460
rect 17552 20448 17558 20460
rect 18414 20448 18420 20460
rect 17552 20420 18420 20448
rect 17552 20408 17558 20420
rect 18414 20408 18420 20420
rect 18472 20408 18478 20460
rect 19334 20408 19340 20460
rect 19392 20408 19398 20460
rect 20070 20448 20076 20460
rect 19628 20420 20076 20448
rect 14645 20343 14703 20349
rect 16040 20352 16528 20380
rect 14090 20272 14096 20324
rect 14148 20272 14154 20324
rect 16040 20321 16068 20352
rect 16666 20340 16672 20392
rect 16724 20340 16730 20392
rect 18601 20383 18659 20389
rect 18601 20349 18613 20383
rect 18647 20349 18659 20383
rect 18601 20343 18659 20349
rect 16025 20315 16083 20321
rect 16025 20281 16037 20315
rect 16071 20281 16083 20315
rect 16025 20275 16083 20281
rect 16574 20244 16580 20256
rect 14016 20216 16580 20244
rect 16574 20204 16580 20216
rect 16632 20204 16638 20256
rect 16684 20244 16712 20340
rect 17954 20244 17960 20256
rect 16684 20216 17960 20244
rect 17954 20204 17960 20216
rect 18012 20244 18018 20256
rect 18616 20244 18644 20343
rect 18012 20216 18644 20244
rect 18012 20204 18018 20216
rect 18874 20204 18880 20256
rect 18932 20244 18938 20256
rect 19628 20244 19656 20420
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20180 20457 20208 20488
rect 20165 20451 20223 20457
rect 20165 20417 20177 20451
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 19702 20340 19708 20392
rect 19760 20380 19766 20392
rect 20349 20383 20407 20389
rect 20349 20380 20361 20383
rect 19760 20352 20361 20380
rect 19760 20340 19766 20352
rect 20349 20349 20361 20352
rect 20395 20349 20407 20383
rect 20349 20343 20407 20349
rect 18932 20216 19656 20244
rect 18932 20204 18938 20216
rect 19978 20204 19984 20256
rect 20036 20204 20042 20256
rect 20254 20204 20260 20256
rect 20312 20204 20318 20256
rect 1104 20154 20884 20176
rect 198 20068 204 20120
rect 256 20068 262 20120
rect 1104 20102 3422 20154
rect 3474 20102 3486 20154
rect 3538 20102 3550 20154
rect 3602 20102 3614 20154
rect 3666 20102 3678 20154
rect 3730 20102 8367 20154
rect 8419 20102 8431 20154
rect 8483 20102 8495 20154
rect 8547 20102 8559 20154
rect 8611 20102 8623 20154
rect 8675 20102 13312 20154
rect 13364 20102 13376 20154
rect 13428 20102 13440 20154
rect 13492 20102 13504 20154
rect 13556 20102 13568 20154
rect 13620 20102 18257 20154
rect 18309 20102 18321 20154
rect 18373 20102 18385 20154
rect 18437 20102 18449 20154
rect 18501 20102 18513 20154
rect 18565 20102 20884 20154
rect 1104 20080 20884 20102
rect 216 20040 244 20068
rect 3694 20040 3700 20052
rect 216 20012 3700 20040
rect 3694 20000 3700 20012
rect 3752 20000 3758 20052
rect 5552 20012 6776 20040
rect 4068 19916 4120 19922
rect 1394 19864 1400 19916
rect 1452 19864 1458 19916
rect 1670 19864 1676 19916
rect 1728 19864 1734 19916
rect 2314 19864 2320 19916
rect 2372 19864 2378 19916
rect 5166 19864 5172 19916
rect 5224 19904 5230 19916
rect 5552 19913 5580 20012
rect 6748 19984 6776 20012
rect 7466 20000 7472 20052
rect 7524 20040 7530 20052
rect 7524 20012 8156 20040
rect 7524 20000 7530 20012
rect 6730 19932 6736 19984
rect 6788 19932 6794 19984
rect 7484 19913 7512 20000
rect 5537 19907 5595 19913
rect 5537 19904 5549 19907
rect 5224 19876 5549 19904
rect 5224 19864 5230 19876
rect 5537 19873 5549 19876
rect 5583 19873 5595 19907
rect 5537 19867 5595 19873
rect 7469 19907 7527 19913
rect 7469 19873 7481 19907
rect 7515 19873 7527 19907
rect 7469 19867 7527 19873
rect 4068 19858 4120 19864
rect 2591 19839 2649 19845
rect 2591 19805 2603 19839
rect 2637 19836 2649 19839
rect 2682 19836 2688 19848
rect 2637 19808 2688 19836
rect 2637 19805 2649 19808
rect 2591 19799 2649 19805
rect 2682 19796 2688 19808
rect 2740 19796 2746 19848
rect 4341 19839 4399 19845
rect 4341 19836 4353 19839
rect 4172 19808 4353 19836
rect 3234 19728 3240 19780
rect 3292 19768 3298 19780
rect 4065 19771 4123 19777
rect 4065 19768 4077 19771
rect 3292 19740 4077 19768
rect 3292 19728 3298 19740
rect 4065 19737 4077 19740
rect 4111 19737 4123 19771
rect 4065 19731 4123 19737
rect 3326 19660 3332 19712
rect 3384 19660 3390 19712
rect 3694 19660 3700 19712
rect 3752 19700 3758 19712
rect 3878 19700 3884 19712
rect 3752 19672 3884 19700
rect 3752 19660 3758 19672
rect 3878 19660 3884 19672
rect 3936 19700 3942 19712
rect 4172 19700 4200 19808
rect 4341 19805 4353 19808
rect 4387 19805 4399 19839
rect 4341 19799 4399 19805
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19836 4491 19839
rect 4479 19808 5488 19836
rect 4479 19805 4491 19808
rect 4433 19799 4491 19805
rect 4246 19728 4252 19780
rect 4304 19768 4310 19780
rect 4801 19771 4859 19777
rect 4801 19768 4813 19771
rect 4304 19740 4813 19768
rect 4304 19728 4310 19740
rect 4801 19737 4813 19740
rect 4847 19737 4859 19771
rect 5460 19768 5488 19808
rect 5718 19796 5724 19848
rect 5776 19836 5782 19848
rect 5811 19839 5869 19845
rect 5811 19836 5823 19839
rect 5776 19808 5823 19836
rect 5776 19796 5782 19808
rect 5811 19805 5823 19808
rect 5857 19805 5869 19839
rect 5811 19799 5869 19805
rect 6362 19796 6368 19848
rect 6420 19836 6426 19848
rect 7711 19839 7769 19845
rect 7711 19836 7723 19839
rect 6420 19808 7723 19836
rect 6420 19796 6426 19808
rect 7711 19805 7723 19808
rect 7757 19805 7769 19839
rect 7711 19799 7769 19805
rect 8128 19768 8156 20012
rect 9232 20012 11284 20040
rect 8570 19932 8576 19984
rect 8628 19972 8634 19984
rect 8846 19972 8852 19984
rect 8628 19944 8852 19972
rect 8628 19932 8634 19944
rect 8846 19932 8852 19944
rect 8904 19932 8910 19984
rect 8662 19904 8668 19916
rect 8220 19876 8668 19904
rect 8220 19848 8248 19876
rect 8662 19864 8668 19876
rect 8720 19904 8726 19916
rect 9232 19913 9260 20012
rect 9217 19907 9275 19913
rect 9217 19904 9229 19907
rect 8720 19876 9229 19904
rect 8720 19864 8726 19876
rect 9217 19873 9229 19876
rect 9263 19873 9275 19907
rect 11256 19904 11284 20012
rect 11514 20000 11520 20052
rect 11572 20040 11578 20052
rect 11609 20043 11667 20049
rect 11609 20040 11621 20043
rect 11572 20012 11621 20040
rect 11572 20000 11578 20012
rect 11609 20009 11621 20012
rect 11655 20009 11667 20043
rect 11609 20003 11667 20009
rect 12250 20000 12256 20052
rect 12308 20040 12314 20052
rect 13170 20040 13176 20052
rect 12308 20012 13176 20040
rect 12308 20000 12314 20012
rect 13170 20000 13176 20012
rect 13228 20040 13234 20052
rect 14090 20040 14096 20052
rect 13228 20012 14096 20040
rect 13228 20000 13234 20012
rect 14090 20000 14096 20012
rect 14148 20040 14154 20052
rect 14148 20012 15516 20040
rect 14148 20000 14154 20012
rect 11514 19904 11520 19916
rect 11256 19876 11520 19904
rect 9217 19867 9275 19873
rect 11514 19864 11520 19876
rect 11572 19904 11578 19916
rect 11977 19907 12035 19913
rect 11977 19904 11989 19907
rect 11572 19876 11989 19904
rect 11572 19864 11578 19876
rect 11977 19873 11989 19876
rect 12023 19873 12035 19907
rect 11977 19867 12035 19873
rect 15378 19864 15384 19916
rect 15436 19864 15442 19916
rect 15488 19913 15516 20012
rect 16390 20000 16396 20052
rect 16448 20040 16454 20052
rect 16485 20043 16543 20049
rect 16485 20040 16497 20043
rect 16448 20012 16497 20040
rect 16448 20000 16454 20012
rect 16485 20009 16497 20012
rect 16531 20009 16543 20043
rect 16485 20003 16543 20009
rect 16850 20000 16856 20052
rect 16908 20000 16914 20052
rect 17770 20000 17776 20052
rect 17828 20000 17834 20052
rect 18877 20043 18935 20049
rect 18877 20009 18889 20043
rect 18923 20040 18935 20043
rect 18966 20040 18972 20052
rect 18923 20012 18972 20040
rect 18923 20009 18935 20012
rect 18877 20003 18935 20009
rect 18966 20000 18972 20012
rect 19024 20000 19030 20052
rect 19978 20040 19984 20052
rect 19076 20012 19984 20040
rect 15473 19907 15531 19913
rect 15473 19873 15485 19907
rect 15519 19873 15531 19907
rect 15473 19867 15531 19873
rect 16390 19864 16396 19916
rect 16448 19904 16454 19916
rect 16758 19904 16764 19916
rect 16448 19876 16764 19904
rect 16448 19864 16454 19876
rect 16758 19864 16764 19876
rect 16816 19864 16822 19916
rect 8202 19796 8208 19848
rect 8260 19796 8266 19848
rect 8310 19808 9076 19836
rect 8310 19768 8338 19808
rect 5460 19740 6592 19768
rect 8128 19740 8338 19768
rect 4801 19731 4859 19737
rect 3936 19672 4200 19700
rect 3936 19660 3942 19672
rect 4614 19660 4620 19712
rect 4672 19700 4678 19712
rect 4890 19700 4896 19712
rect 4672 19672 4896 19700
rect 4672 19660 4678 19672
rect 4890 19660 4896 19672
rect 4948 19700 4954 19712
rect 5169 19703 5227 19709
rect 5169 19700 5181 19703
rect 4948 19672 5181 19700
rect 4948 19660 4954 19672
rect 5169 19669 5181 19672
rect 5215 19669 5227 19703
rect 5169 19663 5227 19669
rect 5353 19703 5411 19709
rect 5353 19669 5365 19703
rect 5399 19700 5411 19703
rect 5626 19700 5632 19712
rect 5399 19672 5632 19700
rect 5399 19669 5411 19672
rect 5353 19663 5411 19669
rect 5626 19660 5632 19672
rect 5684 19660 5690 19712
rect 6564 19709 6592 19740
rect 6549 19703 6607 19709
rect 6549 19669 6561 19703
rect 6595 19669 6607 19703
rect 6549 19663 6607 19669
rect 8481 19703 8539 19709
rect 8481 19669 8493 19703
rect 8527 19700 8539 19703
rect 8846 19700 8852 19712
rect 8527 19672 8852 19700
rect 8527 19669 8539 19672
rect 8481 19663 8539 19669
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9048 19700 9076 19808
rect 9122 19796 9128 19848
rect 9180 19796 9186 19848
rect 9490 19836 9496 19848
rect 9451 19808 9496 19836
rect 9490 19796 9496 19808
rect 9548 19796 9554 19848
rect 10042 19796 10048 19848
rect 10100 19836 10106 19848
rect 10594 19836 10600 19848
rect 10100 19808 10600 19836
rect 10100 19796 10106 19808
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 10778 19796 10784 19848
rect 10836 19836 10842 19848
rect 10871 19839 10929 19845
rect 10871 19836 10883 19839
rect 10836 19808 10883 19836
rect 10836 19796 10842 19808
rect 10871 19805 10883 19808
rect 10917 19805 10929 19839
rect 12219 19839 12277 19845
rect 12219 19836 12231 19839
rect 10871 19799 10929 19805
rect 11992 19808 12231 19836
rect 9508 19768 9536 19796
rect 9508 19740 10640 19768
rect 10612 19712 10640 19740
rect 11992 19712 12020 19808
rect 12219 19805 12231 19808
rect 12265 19805 12277 19839
rect 12219 19799 12277 19805
rect 13538 19796 13544 19848
rect 13596 19796 13602 19848
rect 13909 19839 13967 19845
rect 13909 19805 13921 19839
rect 13955 19805 13967 19839
rect 13909 19799 13967 19805
rect 13924 19768 13952 19799
rect 14090 19796 14096 19848
rect 14148 19796 14154 19848
rect 14366 19836 14372 19848
rect 14327 19808 14372 19836
rect 14366 19796 14372 19808
rect 14424 19836 14430 19848
rect 15396 19836 15424 19864
rect 15715 19839 15773 19845
rect 15715 19836 15727 19839
rect 14424 19808 15727 19836
rect 14424 19796 14430 19808
rect 15715 19805 15727 19808
rect 15761 19805 15773 19839
rect 16868 19836 16896 20000
rect 17129 19839 17187 19845
rect 17129 19836 17141 19839
rect 16868 19808 17141 19836
rect 15715 19799 15773 19805
rect 17129 19805 17141 19808
rect 17175 19805 17187 19839
rect 17129 19799 17187 19805
rect 17497 19839 17555 19845
rect 17497 19805 17509 19839
rect 17543 19805 17555 19839
rect 17788 19836 17816 20000
rect 18138 19864 18144 19916
rect 18196 19864 18202 19916
rect 18049 19839 18107 19845
rect 18049 19836 18061 19839
rect 17788 19808 18061 19836
rect 17497 19799 17555 19805
rect 18049 19805 18061 19808
rect 18095 19805 18107 19839
rect 18049 19799 18107 19805
rect 14826 19768 14832 19780
rect 12176 19740 13860 19768
rect 13924 19740 14832 19768
rect 12176 19712 12204 19740
rect 10042 19700 10048 19712
rect 9048 19672 10048 19700
rect 10042 19660 10048 19672
rect 10100 19660 10106 19712
rect 10226 19660 10232 19712
rect 10284 19660 10290 19712
rect 10594 19660 10600 19712
rect 10652 19660 10658 19712
rect 11974 19660 11980 19712
rect 12032 19660 12038 19712
rect 12158 19660 12164 19712
rect 12216 19660 12222 19712
rect 12986 19660 12992 19712
rect 13044 19660 13050 19712
rect 13832 19700 13860 19740
rect 14826 19728 14832 19740
rect 14884 19728 14890 19780
rect 17512 19768 17540 19799
rect 16960 19740 17540 19768
rect 18156 19768 18184 19864
rect 19076 19845 19104 20012
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 20070 20000 20076 20052
rect 20128 20040 20134 20052
rect 20257 20043 20315 20049
rect 20257 20040 20269 20043
rect 20128 20012 20269 20040
rect 20128 20000 20134 20012
rect 20257 20009 20269 20012
rect 20303 20009 20315 20043
rect 20257 20003 20315 20009
rect 19061 19839 19119 19845
rect 19061 19805 19073 19839
rect 19107 19805 19119 19839
rect 19061 19799 19119 19805
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19487 19839 19545 19845
rect 19487 19805 19499 19839
rect 19533 19805 19545 19839
rect 19487 19799 19545 19805
rect 19260 19768 19288 19799
rect 18156 19740 19288 19768
rect 14366 19700 14372 19712
rect 13832 19672 14372 19700
rect 14366 19660 14372 19672
rect 14424 19660 14430 19712
rect 14642 19660 14648 19712
rect 14700 19700 14706 19712
rect 15105 19703 15163 19709
rect 15105 19700 15117 19703
rect 14700 19672 15117 19700
rect 14700 19660 14706 19672
rect 15105 19669 15117 19672
rect 15151 19669 15163 19703
rect 15105 19663 15163 19669
rect 15654 19660 15660 19712
rect 15712 19700 15718 19712
rect 16206 19700 16212 19712
rect 15712 19672 16212 19700
rect 15712 19660 15718 19672
rect 16206 19660 16212 19672
rect 16264 19660 16270 19712
rect 16960 19709 16988 19740
rect 19076 19712 19104 19740
rect 19334 19728 19340 19780
rect 19392 19768 19398 19780
rect 19502 19768 19530 19799
rect 19392 19740 19530 19768
rect 19392 19728 19398 19740
rect 16945 19703 17003 19709
rect 16945 19669 16957 19703
rect 16991 19669 17003 19703
rect 16945 19663 17003 19669
rect 17586 19660 17592 19712
rect 17644 19660 17650 19712
rect 17865 19703 17923 19709
rect 17865 19669 17877 19703
rect 17911 19700 17923 19703
rect 18414 19700 18420 19712
rect 17911 19672 18420 19700
rect 17911 19669 17923 19672
rect 17865 19663 17923 19669
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 19058 19660 19064 19712
rect 19116 19660 19122 19712
rect 19518 19660 19524 19712
rect 19576 19700 19582 19712
rect 20990 19700 20996 19712
rect 19576 19672 20996 19700
rect 19576 19660 19582 19672
rect 20990 19660 20996 19672
rect 21048 19660 21054 19712
rect 1104 19610 21043 19632
rect 1104 19558 5894 19610
rect 5946 19558 5958 19610
rect 6010 19558 6022 19610
rect 6074 19558 6086 19610
rect 6138 19558 6150 19610
rect 6202 19558 10839 19610
rect 10891 19558 10903 19610
rect 10955 19558 10967 19610
rect 11019 19558 11031 19610
rect 11083 19558 11095 19610
rect 11147 19558 15784 19610
rect 15836 19558 15848 19610
rect 15900 19558 15912 19610
rect 15964 19558 15976 19610
rect 16028 19558 16040 19610
rect 16092 19558 20729 19610
rect 20781 19558 20793 19610
rect 20845 19558 20857 19610
rect 20909 19558 20921 19610
rect 20973 19558 20985 19610
rect 21037 19558 21043 19610
rect 1104 19536 21043 19558
rect 3234 19456 3240 19508
rect 3292 19456 3298 19508
rect 3326 19456 3332 19508
rect 3384 19496 3390 19508
rect 3384 19468 3648 19496
rect 3384 19456 3390 19468
rect 750 19388 756 19440
rect 808 19428 814 19440
rect 1489 19431 1547 19437
rect 1489 19428 1501 19431
rect 808 19400 1501 19428
rect 808 19388 814 19400
rect 1489 19397 1501 19400
rect 1535 19397 1547 19431
rect 1489 19391 1547 19397
rect 2130 19388 2136 19440
rect 2188 19388 2194 19440
rect 3252 19428 3280 19456
rect 3513 19431 3571 19437
rect 3513 19428 3525 19431
rect 3252 19400 3525 19428
rect 3513 19397 3525 19400
rect 3559 19397 3571 19431
rect 3513 19391 3571 19397
rect 2148 19360 2176 19388
rect 2223 19363 2281 19369
rect 2223 19360 2235 19363
rect 2148 19332 2235 19360
rect 2223 19329 2235 19332
rect 2269 19329 2281 19363
rect 3620 19360 3648 19468
rect 4338 19456 4344 19508
rect 4396 19496 4402 19508
rect 7282 19496 7288 19508
rect 4396 19468 7288 19496
rect 4396 19456 4402 19468
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 8938 19496 8944 19508
rect 7852 19468 8944 19496
rect 3694 19388 3700 19440
rect 3752 19428 3758 19440
rect 3789 19431 3847 19437
rect 3789 19428 3801 19431
rect 3752 19400 3801 19428
rect 3752 19388 3758 19400
rect 3789 19397 3801 19400
rect 3835 19397 3847 19431
rect 3789 19391 3847 19397
rect 4614 19388 4620 19440
rect 4672 19388 4678 19440
rect 5258 19388 5264 19440
rect 5316 19428 5322 19440
rect 7852 19428 7880 19468
rect 8938 19456 8944 19468
rect 8996 19456 9002 19508
rect 9122 19456 9128 19508
rect 9180 19496 9186 19508
rect 9180 19468 10088 19496
rect 9180 19456 9186 19468
rect 5316 19400 7880 19428
rect 5316 19388 5322 19400
rect 3881 19363 3939 19369
rect 3881 19360 3893 19363
rect 3620 19332 3893 19360
rect 2223 19323 2281 19329
rect 3881 19329 3893 19332
rect 3927 19329 3939 19363
rect 3881 19323 3939 19329
rect 4246 19320 4252 19372
rect 4304 19320 4310 19372
rect 4706 19320 4712 19372
rect 4764 19360 4770 19372
rect 5626 19360 5632 19372
rect 4764 19332 5632 19360
rect 4764 19320 4770 19332
rect 5626 19320 5632 19332
rect 5684 19320 5690 19372
rect 7650 19320 7656 19372
rect 7708 19320 7714 19372
rect 7852 19369 7880 19400
rect 9674 19388 9680 19440
rect 9732 19428 9738 19440
rect 10060 19437 10088 19468
rect 10226 19456 10232 19508
rect 10284 19456 10290 19508
rect 11882 19456 11888 19508
rect 11940 19496 11946 19508
rect 12161 19499 12219 19505
rect 12161 19496 12173 19499
rect 11940 19468 12173 19496
rect 11940 19456 11946 19468
rect 12161 19465 12173 19468
rect 12207 19465 12219 19499
rect 13538 19496 13544 19508
rect 12161 19459 12219 19465
rect 12452 19468 13544 19496
rect 9769 19431 9827 19437
rect 9769 19428 9781 19431
rect 9732 19400 9781 19428
rect 9732 19388 9738 19400
rect 9769 19397 9781 19400
rect 9815 19397 9827 19431
rect 9769 19391 9827 19397
rect 10045 19431 10103 19437
rect 10045 19397 10057 19431
rect 10091 19397 10103 19431
rect 10045 19391 10103 19397
rect 10137 19431 10195 19437
rect 10137 19397 10149 19431
rect 10183 19428 10195 19431
rect 10244 19428 10272 19456
rect 12452 19437 12480 19468
rect 13538 19456 13544 19468
rect 13596 19456 13602 19508
rect 14366 19456 14372 19508
rect 14424 19496 14430 19508
rect 15102 19496 15108 19508
rect 14424 19468 15108 19496
rect 14424 19456 14430 19468
rect 15102 19456 15108 19468
rect 15160 19456 15166 19508
rect 15654 19456 15660 19508
rect 15712 19496 15718 19508
rect 17862 19496 17868 19508
rect 15712 19468 17868 19496
rect 15712 19456 15718 19468
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 17957 19499 18015 19505
rect 17957 19465 17969 19499
rect 18003 19465 18015 19499
rect 17957 19459 18015 19465
rect 10183 19400 10272 19428
rect 10873 19431 10931 19437
rect 10183 19397 10195 19400
rect 10137 19391 10195 19397
rect 10873 19397 10885 19431
rect 10919 19428 10931 19431
rect 12437 19431 12495 19437
rect 10919 19400 11192 19428
rect 10919 19397 10931 19400
rect 10873 19391 10931 19397
rect 11164 19372 11192 19400
rect 12437 19397 12449 19431
rect 12483 19397 12495 19431
rect 12437 19391 12495 19397
rect 13078 19388 13084 19440
rect 13136 19428 13142 19440
rect 13265 19431 13323 19437
rect 13265 19428 13277 19431
rect 13136 19400 13277 19428
rect 13136 19388 13142 19400
rect 13265 19397 13277 19400
rect 13311 19397 13323 19431
rect 13265 19391 13323 19397
rect 13354 19388 13360 19440
rect 13412 19428 13418 19440
rect 13412 19400 14136 19428
rect 13412 19388 13418 19400
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19329 7895 19363
rect 7837 19323 7895 19329
rect 8570 19320 8576 19372
rect 8628 19320 8634 19372
rect 8662 19320 8668 19372
rect 8720 19369 8726 19372
rect 8720 19363 8748 19369
rect 8736 19329 8748 19363
rect 8720 19323 8748 19329
rect 8720 19320 8726 19323
rect 8846 19320 8852 19372
rect 8904 19320 8910 19372
rect 10502 19320 10508 19372
rect 10560 19320 10566 19372
rect 11146 19320 11152 19372
rect 11204 19320 11210 19372
rect 12526 19320 12532 19372
rect 12584 19320 12590 19372
rect 12897 19363 12955 19369
rect 12897 19329 12909 19363
rect 12943 19360 12955 19363
rect 13909 19363 13967 19369
rect 13909 19360 13921 19363
rect 12943 19332 13921 19360
rect 12943 19329 12955 19332
rect 12897 19323 12955 19329
rect 13909 19329 13921 19332
rect 13955 19360 13967 19363
rect 13998 19360 14004 19372
rect 13955 19332 14004 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 13998 19320 14004 19332
rect 14056 19320 14062 19372
rect 14108 19369 14136 19400
rect 14093 19363 14151 19369
rect 14093 19329 14105 19363
rect 14139 19329 14151 19363
rect 14093 19323 14151 19329
rect 14826 19320 14832 19372
rect 14884 19320 14890 19372
rect 17218 19320 17224 19372
rect 17276 19320 17282 19372
rect 17586 19320 17592 19372
rect 17644 19320 17650 19372
rect 17972 19360 18000 19459
rect 18414 19456 18420 19508
rect 18472 19456 18478 19508
rect 20254 19496 20260 19508
rect 19812 19468 20260 19496
rect 18432 19428 18460 19456
rect 19812 19437 19840 19468
rect 20254 19456 20260 19468
rect 20312 19456 20318 19508
rect 19797 19431 19855 19437
rect 18432 19400 18920 19428
rect 18892 19369 18920 19400
rect 19797 19397 19809 19431
rect 19843 19397 19855 19431
rect 19797 19391 19855 19397
rect 19978 19388 19984 19440
rect 20036 19428 20042 19440
rect 20533 19431 20591 19437
rect 20533 19428 20545 19431
rect 20036 19400 20545 19428
rect 20036 19388 20042 19400
rect 20533 19397 20545 19400
rect 20579 19397 20591 19431
rect 20533 19391 20591 19397
rect 18325 19363 18383 19369
rect 18325 19360 18337 19363
rect 17972 19332 18337 19360
rect 18325 19329 18337 19332
rect 18371 19360 18383 19363
rect 18693 19363 18751 19369
rect 18693 19360 18705 19363
rect 18371 19332 18705 19360
rect 18371 19329 18383 19332
rect 18325 19323 18383 19329
rect 18693 19329 18705 19332
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19329 18935 19363
rect 18877 19323 18935 19329
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 20254 19320 20260 19372
rect 20312 19320 20318 19372
rect 1949 19295 2007 19301
rect 1949 19261 1961 19295
rect 1995 19261 2007 19295
rect 1949 19255 2007 19261
rect 2976 19264 3358 19292
rect 1302 19116 1308 19168
rect 1360 19156 1366 19168
rect 1581 19159 1639 19165
rect 1581 19156 1593 19159
rect 1360 19128 1593 19156
rect 1360 19116 1366 19128
rect 1581 19125 1593 19128
rect 1627 19125 1639 19159
rect 1964 19156 1992 19255
rect 2976 19233 3004 19264
rect 8294 19252 8300 19304
rect 8352 19252 8358 19304
rect 9950 19252 9956 19304
rect 10008 19252 10014 19304
rect 12986 19252 12992 19304
rect 13044 19252 13050 19304
rect 14553 19295 14611 19301
rect 14553 19261 14565 19295
rect 14599 19292 14611 19295
rect 14642 19292 14648 19304
rect 14599 19264 14648 19292
rect 14599 19261 14611 19264
rect 14553 19255 14611 19261
rect 14642 19252 14648 19264
rect 14700 19252 14706 19304
rect 15010 19301 15016 19304
rect 14967 19295 15016 19301
rect 14967 19261 14979 19295
rect 15013 19261 15016 19295
rect 14967 19255 15016 19261
rect 15010 19252 15016 19255
rect 15068 19252 15074 19304
rect 15102 19252 15108 19304
rect 15160 19252 15166 19304
rect 16945 19295 17003 19301
rect 16945 19261 16957 19295
rect 16991 19261 17003 19295
rect 17604 19292 17632 19320
rect 18417 19295 18475 19301
rect 18417 19292 18429 19295
rect 17604 19264 18429 19292
rect 16945 19255 17003 19261
rect 18417 19261 18429 19264
rect 18463 19261 18475 19295
rect 18417 19255 18475 19261
rect 18601 19295 18659 19301
rect 18601 19261 18613 19295
rect 18647 19292 18659 19295
rect 18785 19295 18843 19301
rect 18785 19292 18797 19295
rect 18647 19264 18797 19292
rect 18647 19261 18659 19264
rect 18601 19255 18659 19261
rect 18785 19261 18797 19264
rect 18831 19261 18843 19295
rect 18785 19255 18843 19261
rect 2961 19227 3019 19233
rect 2961 19193 2973 19227
rect 3007 19193 3019 19227
rect 2961 19187 3019 19193
rect 4798 19184 4804 19236
rect 4856 19184 4862 19236
rect 4890 19184 4896 19236
rect 4948 19224 4954 19236
rect 4948 19196 5396 19224
rect 4948 19184 4954 19196
rect 2038 19156 2044 19168
rect 1964 19128 2044 19156
rect 1581 19119 1639 19125
rect 2038 19116 2044 19128
rect 2096 19156 2102 19168
rect 2314 19156 2320 19168
rect 2096 19128 2320 19156
rect 2096 19116 2102 19128
rect 2314 19116 2320 19128
rect 2372 19116 2378 19168
rect 2774 19116 2780 19168
rect 2832 19156 2838 19168
rect 3418 19156 3424 19168
rect 2832 19128 3424 19156
rect 2832 19116 2838 19128
rect 3418 19116 3424 19128
rect 3476 19116 3482 19168
rect 4816 19156 4844 19184
rect 5258 19156 5264 19168
rect 4816 19128 5264 19156
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 5368 19156 5396 19196
rect 6822 19184 6828 19236
rect 6880 19224 6886 19236
rect 8110 19224 8116 19236
rect 6880 19196 8116 19224
rect 6880 19184 6886 19196
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 11054 19184 11060 19236
rect 11112 19184 11118 19236
rect 15749 19227 15807 19233
rect 15749 19193 15761 19227
rect 15795 19224 15807 19227
rect 16114 19224 16120 19236
rect 15795 19196 16120 19224
rect 15795 19193 15807 19196
rect 15749 19187 15807 19193
rect 16114 19184 16120 19196
rect 16172 19184 16178 19236
rect 7558 19156 7564 19168
rect 5368 19128 7564 19156
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 7926 19116 7932 19168
rect 7984 19156 7990 19168
rect 9398 19156 9404 19168
rect 7984 19128 9404 19156
rect 7984 19116 7990 19128
rect 9398 19116 9404 19128
rect 9456 19116 9462 19168
rect 9490 19116 9496 19168
rect 9548 19116 9554 19168
rect 13449 19159 13507 19165
rect 13449 19125 13461 19159
rect 13495 19156 13507 19159
rect 15010 19156 15016 19168
rect 13495 19128 15016 19156
rect 13495 19125 13507 19128
rect 13449 19119 13507 19125
rect 15010 19116 15016 19128
rect 15068 19156 15074 19168
rect 15470 19156 15476 19168
rect 15068 19128 15476 19156
rect 15068 19116 15074 19128
rect 15470 19116 15476 19128
rect 15528 19116 15534 19168
rect 15838 19116 15844 19168
rect 15896 19156 15902 19168
rect 16025 19159 16083 19165
rect 16025 19156 16037 19159
rect 15896 19128 16037 19156
rect 15896 19116 15902 19128
rect 16025 19125 16037 19128
rect 16071 19125 16083 19159
rect 16960 19156 16988 19255
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 20346 19292 20352 19304
rect 19392 19264 20352 19292
rect 19392 19252 19398 19264
rect 20346 19252 20352 19264
rect 20404 19252 20410 19304
rect 20530 19252 20536 19304
rect 20588 19252 20594 19304
rect 18138 19184 18144 19236
rect 18196 19184 18202 19236
rect 18156 19156 18184 19184
rect 16960 19128 18184 19156
rect 18509 19159 18567 19165
rect 16025 19119 16083 19125
rect 18509 19125 18521 19159
rect 18555 19156 18567 19159
rect 19150 19156 19156 19168
rect 18555 19128 19156 19156
rect 18555 19125 18567 19128
rect 18509 19119 18567 19125
rect 19150 19116 19156 19128
rect 19208 19116 19214 19168
rect 19242 19116 19248 19168
rect 19300 19156 19306 19168
rect 19429 19159 19487 19165
rect 19429 19156 19441 19159
rect 19300 19128 19441 19156
rect 19300 19116 19306 19128
rect 19429 19125 19441 19128
rect 19475 19125 19487 19159
rect 19429 19119 19487 19125
rect 20070 19116 20076 19168
rect 20128 19116 20134 19168
rect 20346 19116 20352 19168
rect 20404 19116 20410 19168
rect 1104 19066 20884 19088
rect 1104 19014 3422 19066
rect 3474 19014 3486 19066
rect 3538 19014 3550 19066
rect 3602 19014 3614 19066
rect 3666 19014 3678 19066
rect 3730 19014 8367 19066
rect 8419 19014 8431 19066
rect 8483 19014 8495 19066
rect 8547 19014 8559 19066
rect 8611 19014 8623 19066
rect 8675 19014 13312 19066
rect 13364 19014 13376 19066
rect 13428 19014 13440 19066
rect 13492 19014 13504 19066
rect 13556 19014 13568 19066
rect 13620 19014 18257 19066
rect 18309 19014 18321 19066
rect 18373 19014 18385 19066
rect 18437 19014 18449 19066
rect 18501 19014 18513 19066
rect 18565 19014 20884 19066
rect 1104 18992 20884 19014
rect 3050 18912 3056 18964
rect 3108 18952 3114 18964
rect 3145 18955 3203 18961
rect 3145 18952 3157 18955
rect 3108 18924 3157 18952
rect 3108 18912 3114 18924
rect 3145 18921 3157 18924
rect 3191 18921 3203 18955
rect 3145 18915 3203 18921
rect 3421 18955 3479 18961
rect 3421 18921 3433 18955
rect 3467 18952 3479 18955
rect 4338 18952 4344 18964
rect 3467 18924 4344 18952
rect 3467 18921 3479 18924
rect 3421 18915 3479 18921
rect 4338 18912 4344 18924
rect 4396 18912 4402 18964
rect 5166 18912 5172 18964
rect 5224 18952 5230 18964
rect 6546 18952 6552 18964
rect 5224 18924 6552 18952
rect 5224 18912 5230 18924
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 6730 18912 6736 18964
rect 6788 18952 6794 18964
rect 7558 18952 7564 18964
rect 6788 18924 7564 18952
rect 6788 18912 6794 18924
rect 7558 18912 7564 18924
rect 7616 18952 7622 18964
rect 8294 18952 8300 18964
rect 7616 18924 8300 18952
rect 7616 18912 7622 18924
rect 8294 18912 8300 18924
rect 8352 18912 8358 18964
rect 12526 18912 12532 18964
rect 12584 18952 12590 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 12584 18924 13277 18952
rect 12584 18912 12590 18924
rect 13265 18921 13277 18924
rect 13311 18921 13323 18955
rect 17865 18955 17923 18961
rect 17865 18952 17877 18955
rect 13265 18915 13323 18921
rect 16868 18924 17877 18952
rect 1578 18844 1584 18896
rect 1636 18884 1642 18896
rect 1762 18884 1768 18896
rect 1636 18856 1768 18884
rect 1636 18844 1642 18856
rect 1762 18844 1768 18856
rect 1820 18844 1826 18896
rect 5077 18887 5135 18893
rect 5077 18853 5089 18887
rect 5123 18884 5135 18887
rect 6089 18887 6147 18893
rect 6089 18884 6101 18887
rect 5123 18856 6101 18884
rect 5123 18853 5135 18856
rect 5077 18847 5135 18853
rect 6089 18853 6101 18856
rect 6135 18853 6147 18887
rect 6089 18847 6147 18853
rect 12910 18856 15700 18884
rect 1210 18776 1216 18828
rect 1268 18816 1274 18828
rect 1268 18788 2912 18816
rect 1268 18776 1274 18788
rect 750 18708 756 18760
rect 808 18748 814 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 808 18720 1409 18748
rect 808 18708 814 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 2317 18751 2375 18757
rect 2317 18748 2329 18751
rect 1397 18711 1455 18717
rect 1504 18720 2329 18748
rect 1210 18640 1216 18692
rect 1268 18680 1274 18692
rect 1504 18680 1532 18720
rect 2317 18717 2329 18720
rect 2363 18717 2375 18751
rect 2317 18711 2375 18717
rect 2682 18708 2688 18760
rect 2740 18708 2746 18760
rect 2884 18744 2912 18788
rect 3694 18776 3700 18828
rect 3752 18816 3758 18828
rect 4065 18819 4123 18825
rect 4065 18816 4077 18819
rect 3752 18788 4077 18816
rect 3752 18776 3758 18788
rect 4065 18785 4077 18788
rect 4111 18785 4123 18819
rect 4065 18779 4123 18785
rect 4890 18776 4896 18828
rect 4948 18816 4954 18828
rect 5629 18819 5687 18825
rect 5629 18816 5641 18819
rect 4948 18788 5641 18816
rect 4948 18776 4954 18788
rect 5629 18785 5641 18788
rect 5675 18785 5687 18819
rect 5629 18779 5687 18785
rect 6365 18819 6423 18825
rect 6365 18785 6377 18819
rect 6411 18816 6423 18819
rect 6411 18788 7328 18816
rect 6411 18785 6423 18788
rect 6365 18779 6423 18785
rect 7300 18760 7328 18788
rect 9674 18776 9680 18828
rect 9732 18816 9738 18828
rect 9732 18788 9890 18816
rect 9732 18776 9738 18788
rect 11514 18776 11520 18828
rect 11572 18816 11578 18828
rect 12253 18819 12311 18825
rect 12253 18816 12265 18819
rect 11572 18788 12265 18816
rect 11572 18776 11578 18788
rect 12253 18785 12265 18788
rect 12299 18785 12311 18819
rect 12253 18779 12311 18785
rect 2961 18751 3019 18757
rect 2961 18744 2973 18751
rect 2884 18717 2973 18744
rect 3007 18717 3019 18751
rect 2884 18716 3019 18717
rect 2961 18711 3019 18716
rect 3050 18708 3056 18760
rect 3108 18748 3114 18760
rect 3237 18751 3295 18757
rect 3237 18748 3249 18751
rect 3108 18720 3249 18748
rect 3108 18708 3114 18720
rect 3237 18717 3249 18720
rect 3283 18717 3295 18751
rect 3237 18711 3295 18717
rect 3326 18708 3332 18760
rect 3384 18748 3390 18760
rect 4307 18751 4365 18757
rect 4307 18748 4319 18751
rect 3384 18720 4319 18748
rect 3384 18708 3390 18720
rect 4307 18717 4319 18720
rect 4353 18717 4365 18751
rect 4307 18711 4365 18717
rect 4430 18708 4436 18760
rect 4488 18748 4494 18760
rect 5445 18751 5503 18757
rect 5445 18748 5457 18751
rect 4488 18720 5457 18748
rect 4488 18708 4494 18720
rect 5445 18717 5457 18720
rect 5491 18717 5503 18751
rect 5445 18711 5503 18717
rect 6454 18708 6460 18760
rect 6512 18757 6518 18760
rect 6512 18751 6561 18757
rect 6512 18717 6515 18751
rect 6549 18717 6561 18751
rect 6512 18711 6561 18717
rect 6512 18708 6518 18711
rect 6638 18708 6644 18760
rect 6696 18708 6702 18760
rect 7282 18708 7288 18760
rect 7340 18708 7346 18760
rect 7374 18708 7380 18760
rect 7432 18748 7438 18760
rect 7469 18751 7527 18757
rect 7469 18748 7481 18751
rect 7432 18720 7481 18748
rect 7432 18708 7438 18720
rect 7469 18717 7481 18720
rect 7515 18748 7527 18751
rect 7743 18751 7801 18757
rect 7515 18720 7696 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 1268 18652 1532 18680
rect 1268 18640 1274 18652
rect 1854 18640 1860 18692
rect 1912 18640 1918 18692
rect 2038 18640 2044 18692
rect 2096 18640 2102 18692
rect 5166 18680 5172 18692
rect 2424 18652 5172 18680
rect 1581 18615 1639 18621
rect 1581 18581 1593 18615
rect 1627 18612 1639 18615
rect 2424 18612 2452 18652
rect 5166 18640 5172 18652
rect 5224 18640 5230 18692
rect 7668 18624 7696 18720
rect 7743 18717 7755 18751
rect 7789 18748 7801 18751
rect 12066 18748 12072 18760
rect 7789 18720 12072 18748
rect 7789 18717 7801 18720
rect 7743 18711 7801 18717
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12526 18748 12532 18760
rect 12487 18720 12532 18748
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 9766 18640 9772 18692
rect 9824 18680 9830 18692
rect 10042 18680 10048 18692
rect 9824 18652 10048 18680
rect 9824 18640 9830 18652
rect 10042 18640 10048 18652
rect 10100 18640 10106 18692
rect 10226 18640 10232 18692
rect 10284 18680 10290 18692
rect 10321 18683 10379 18689
rect 10321 18680 10333 18683
rect 10284 18652 10333 18680
rect 10284 18640 10290 18652
rect 10321 18649 10333 18652
rect 10367 18649 10379 18683
rect 10321 18643 10379 18649
rect 10410 18640 10416 18692
rect 10468 18640 10474 18692
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 10781 18683 10839 18689
rect 10781 18680 10793 18683
rect 10560 18652 10793 18680
rect 10560 18640 10566 18652
rect 10781 18649 10793 18652
rect 10827 18649 10839 18683
rect 10781 18643 10839 18649
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 12910 18680 12938 18856
rect 14274 18776 14280 18828
rect 14332 18776 14338 18828
rect 14918 18776 14924 18828
rect 14976 18776 14982 18828
rect 15562 18776 15568 18828
rect 15620 18776 15626 18828
rect 15672 18816 15700 18856
rect 15958 18819 16016 18825
rect 15958 18816 15970 18819
rect 15672 18788 15970 18816
rect 15958 18785 15970 18788
rect 16004 18785 16016 18819
rect 15958 18779 16016 18785
rect 16117 18819 16175 18825
rect 16117 18785 16129 18819
rect 16163 18816 16175 18819
rect 16868 18816 16896 18924
rect 17865 18921 17877 18924
rect 17911 18921 17923 18955
rect 17865 18915 17923 18921
rect 19337 18955 19395 18961
rect 19337 18921 19349 18955
rect 19383 18952 19395 18955
rect 20346 18952 20352 18964
rect 19383 18924 20352 18952
rect 19383 18921 19395 18924
rect 19337 18915 19395 18921
rect 20346 18912 20352 18924
rect 20404 18912 20410 18964
rect 20441 18887 20499 18893
rect 20441 18853 20453 18887
rect 20487 18884 20499 18887
rect 21542 18884 21548 18896
rect 20487 18856 21548 18884
rect 20487 18853 20499 18856
rect 20441 18847 20499 18853
rect 21542 18844 21548 18856
rect 21600 18844 21606 18896
rect 16163 18788 16896 18816
rect 19889 18819 19947 18825
rect 16163 18785 16175 18788
rect 16117 18779 16175 18785
rect 19889 18785 19901 18819
rect 19935 18816 19947 18819
rect 21266 18816 21272 18828
rect 19935 18788 21272 18816
rect 19935 18785 19947 18788
rect 19889 18779 19947 18785
rect 21266 18776 21272 18788
rect 21324 18776 21330 18828
rect 13814 18708 13820 18760
rect 13872 18708 13878 18760
rect 14292 18748 14320 18776
rect 15105 18751 15163 18757
rect 15105 18748 15117 18751
rect 14292 18720 15117 18748
rect 15105 18717 15117 18720
rect 15151 18717 15163 18751
rect 15105 18711 15163 18717
rect 15838 18708 15844 18760
rect 15896 18708 15902 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16684 18720 16865 18748
rect 11112 18652 12938 18680
rect 13832 18680 13860 18708
rect 14918 18680 14924 18692
rect 13832 18652 14924 18680
rect 11112 18640 11118 18652
rect 14918 18640 14924 18652
rect 14976 18640 14982 18692
rect 1627 18584 2452 18612
rect 2501 18615 2559 18621
rect 1627 18581 1639 18584
rect 1581 18575 1639 18581
rect 2501 18581 2513 18615
rect 2547 18612 2559 18615
rect 2774 18612 2780 18624
rect 2547 18584 2780 18612
rect 2547 18581 2559 18584
rect 2501 18575 2559 18581
rect 2774 18572 2780 18584
rect 2832 18572 2838 18624
rect 2869 18615 2927 18621
rect 2869 18581 2881 18615
rect 2915 18612 2927 18615
rect 3142 18612 3148 18624
rect 2915 18584 3148 18612
rect 2915 18581 2927 18584
rect 2869 18575 2927 18581
rect 3142 18572 3148 18584
rect 3200 18572 3206 18624
rect 5442 18572 5448 18624
rect 5500 18612 5506 18624
rect 7285 18615 7343 18621
rect 7285 18612 7297 18615
rect 5500 18584 7297 18612
rect 5500 18572 5506 18584
rect 7285 18581 7297 18584
rect 7331 18581 7343 18615
rect 7285 18575 7343 18581
rect 7650 18572 7656 18624
rect 7708 18612 7714 18624
rect 8202 18612 8208 18624
rect 7708 18584 8208 18612
rect 7708 18572 7714 18584
rect 8202 18572 8208 18584
rect 8260 18572 8266 18624
rect 8481 18615 8539 18621
rect 8481 18581 8493 18615
rect 8527 18612 8539 18615
rect 9214 18612 9220 18624
rect 8527 18584 9220 18612
rect 8527 18581 8539 18584
rect 8481 18575 8539 18581
rect 9214 18572 9220 18584
rect 9272 18572 9278 18624
rect 11146 18572 11152 18624
rect 11204 18572 11210 18624
rect 11330 18572 11336 18624
rect 11388 18572 11394 18624
rect 12066 18572 12072 18624
rect 12124 18612 12130 18624
rect 12894 18612 12900 18624
rect 12124 18584 12900 18612
rect 12124 18572 12130 18584
rect 12894 18572 12900 18584
rect 12952 18572 12958 18624
rect 14090 18572 14096 18624
rect 14148 18612 14154 18624
rect 16684 18612 16712 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 19061 18751 19119 18757
rect 19061 18748 19073 18751
rect 16853 18711 16911 18717
rect 16960 18747 17138 18748
rect 16960 18741 17153 18747
rect 16960 18720 17107 18741
rect 16960 18692 16988 18720
rect 17095 18707 17107 18720
rect 17141 18707 17153 18741
rect 17095 18701 17153 18707
rect 18708 18720 19073 18748
rect 16942 18640 16948 18692
rect 17000 18640 17006 18692
rect 18708 18624 18736 18720
rect 19061 18717 19073 18720
rect 19107 18717 19119 18751
rect 19061 18711 19119 18717
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19260 18680 19288 18711
rect 18892 18652 19288 18680
rect 19628 18680 19656 18711
rect 20162 18708 20168 18760
rect 20220 18708 20226 18760
rect 21634 18680 21640 18692
rect 19628 18652 21640 18680
rect 14148 18584 16712 18612
rect 14148 18572 14154 18584
rect 16758 18572 16764 18624
rect 16816 18572 16822 18624
rect 18690 18572 18696 18624
rect 18748 18572 18754 18624
rect 18892 18621 18920 18652
rect 21634 18640 21640 18652
rect 21692 18640 21698 18692
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18581 18935 18615
rect 18877 18575 18935 18581
rect 1104 18522 21043 18544
rect 1104 18470 5894 18522
rect 5946 18470 5958 18522
rect 6010 18470 6022 18522
rect 6074 18470 6086 18522
rect 6138 18470 6150 18522
rect 6202 18470 10839 18522
rect 10891 18470 10903 18522
rect 10955 18470 10967 18522
rect 11019 18470 11031 18522
rect 11083 18470 11095 18522
rect 11147 18470 15784 18522
rect 15836 18470 15848 18522
rect 15900 18470 15912 18522
rect 15964 18470 15976 18522
rect 16028 18470 16040 18522
rect 16092 18470 20729 18522
rect 20781 18470 20793 18522
rect 20845 18470 20857 18522
rect 20909 18470 20921 18522
rect 20973 18470 20985 18522
rect 21037 18470 21043 18522
rect 1104 18448 21043 18470
rect 1302 18368 1308 18420
rect 1360 18408 1366 18420
rect 1360 18380 3096 18408
rect 1360 18368 1366 18380
rect 3068 18352 3096 18380
rect 3142 18368 3148 18420
rect 3200 18408 3206 18420
rect 4338 18408 4344 18420
rect 3200 18380 4344 18408
rect 3200 18368 3206 18380
rect 4338 18368 4344 18380
rect 4396 18408 4402 18420
rect 4801 18411 4859 18417
rect 4801 18408 4813 18411
rect 4396 18380 4813 18408
rect 4396 18368 4402 18380
rect 4801 18377 4813 18380
rect 4847 18377 4859 18411
rect 4801 18371 4859 18377
rect 5074 18368 5080 18420
rect 5132 18408 5138 18420
rect 7834 18408 7840 18420
rect 5132 18380 7840 18408
rect 5132 18368 5138 18380
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 9490 18368 9496 18420
rect 9548 18408 9554 18420
rect 9548 18380 9628 18408
rect 9548 18368 9554 18380
rect 750 18300 756 18352
rect 808 18340 814 18352
rect 1489 18343 1547 18349
rect 1489 18340 1501 18343
rect 808 18312 1501 18340
rect 808 18300 814 18312
rect 1489 18309 1501 18312
rect 1535 18309 1547 18343
rect 1489 18303 1547 18309
rect 1673 18343 1731 18349
rect 1673 18309 1685 18343
rect 1719 18340 1731 18343
rect 1946 18340 1952 18352
rect 1719 18312 1952 18340
rect 1719 18309 1731 18312
rect 1673 18303 1731 18309
rect 1946 18300 1952 18312
rect 2004 18300 2010 18352
rect 3050 18300 3056 18352
rect 3108 18300 3114 18352
rect 3234 18300 3240 18352
rect 3292 18340 3298 18352
rect 3513 18343 3571 18349
rect 3513 18340 3525 18343
rect 3292 18312 3525 18340
rect 3292 18300 3298 18312
rect 3513 18309 3525 18312
rect 3559 18340 3571 18343
rect 3970 18340 3976 18352
rect 3559 18312 3976 18340
rect 3559 18309 3571 18312
rect 3513 18303 3571 18309
rect 3970 18300 3976 18312
rect 4028 18300 4034 18352
rect 4614 18300 4620 18352
rect 4672 18340 4678 18352
rect 9600 18340 9628 18380
rect 9674 18368 9680 18420
rect 9732 18368 9738 18420
rect 10410 18368 10416 18420
rect 10468 18408 10474 18420
rect 11057 18411 11115 18417
rect 11057 18408 11069 18411
rect 10468 18380 11069 18408
rect 10468 18368 10474 18380
rect 11057 18377 11069 18380
rect 11103 18377 11115 18411
rect 11057 18371 11115 18377
rect 11164 18380 15056 18408
rect 11164 18340 11192 18380
rect 4672 18312 5120 18340
rect 4672 18300 4678 18312
rect 5092 18284 5120 18312
rect 8680 18312 9410 18340
rect 9600 18312 11192 18340
rect 2131 18275 2189 18281
rect 2131 18241 2143 18275
rect 2177 18272 2189 18275
rect 3602 18272 3608 18284
rect 2177 18244 3608 18272
rect 2177 18241 2189 18244
rect 2131 18235 2189 18241
rect 3602 18232 3608 18244
rect 3660 18232 3666 18284
rect 3786 18232 3792 18284
rect 3844 18232 3850 18284
rect 3878 18232 3884 18284
rect 3936 18232 3942 18284
rect 4246 18232 4252 18284
rect 4304 18272 4310 18284
rect 4890 18272 4896 18284
rect 4304 18244 4896 18272
rect 4304 18232 4310 18244
rect 4890 18232 4896 18244
rect 4948 18232 4954 18284
rect 5074 18232 5080 18284
rect 5132 18232 5138 18284
rect 7466 18232 7472 18284
rect 7524 18272 7530 18284
rect 7559 18275 7617 18281
rect 7559 18272 7571 18275
rect 7524 18244 7571 18272
rect 7524 18232 7530 18244
rect 7559 18241 7571 18244
rect 7605 18241 7617 18275
rect 7559 18235 7617 18241
rect 8294 18232 8300 18284
rect 8352 18272 8358 18284
rect 8680 18281 8708 18312
rect 8665 18275 8723 18281
rect 8665 18272 8677 18275
rect 8352 18244 8677 18272
rect 8352 18232 8358 18244
rect 8665 18241 8677 18244
rect 8711 18241 8723 18275
rect 8665 18235 8723 18241
rect 8939 18275 8997 18281
rect 8939 18241 8951 18275
rect 8985 18272 8997 18275
rect 8985 18244 9352 18272
rect 8985 18241 8997 18244
rect 8939 18235 8997 18241
rect 1857 18207 1915 18213
rect 1857 18173 1869 18207
rect 1903 18173 1915 18207
rect 7285 18207 7343 18213
rect 1857 18167 1915 18173
rect 1872 18136 1900 18167
rect 2869 18139 2927 18145
rect 1872 18108 1992 18136
rect 1964 18080 1992 18108
rect 2869 18105 2881 18139
rect 2915 18136 2927 18139
rect 3344 18136 3372 18190
rect 7285 18173 7297 18207
rect 7331 18173 7343 18207
rect 7285 18167 7343 18173
rect 2915 18108 3372 18136
rect 2915 18105 2927 18108
rect 2869 18099 2927 18105
rect 1946 18028 1952 18080
rect 2004 18028 2010 18080
rect 2314 18028 2320 18080
rect 2372 18068 2378 18080
rect 2682 18068 2688 18080
rect 2372 18040 2688 18068
rect 2372 18028 2378 18040
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 7300 18068 7328 18167
rect 9324 18136 9352 18244
rect 9382 18204 9410 18312
rect 11790 18300 11796 18352
rect 11848 18300 11854 18352
rect 12066 18300 12072 18352
rect 12124 18340 12130 18352
rect 12434 18340 12440 18352
rect 12124 18312 12440 18340
rect 12124 18300 12130 18312
rect 12434 18300 12440 18312
rect 12492 18300 12498 18352
rect 12894 18300 12900 18352
rect 12952 18340 12958 18352
rect 13814 18340 13820 18352
rect 12952 18312 13820 18340
rect 12952 18300 12958 18312
rect 13814 18300 13820 18312
rect 13872 18300 13878 18352
rect 14274 18300 14280 18352
rect 14332 18300 14338 18352
rect 15028 18340 15056 18380
rect 15102 18368 15108 18420
rect 15160 18408 15166 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 15160 18380 15209 18408
rect 15160 18368 15166 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 15378 18368 15384 18420
rect 15436 18408 15442 18420
rect 16850 18408 16856 18420
rect 15436 18380 16856 18408
rect 15436 18368 15442 18380
rect 16850 18368 16856 18380
rect 16908 18368 16914 18420
rect 19610 18368 19616 18420
rect 19668 18408 19674 18420
rect 19797 18411 19855 18417
rect 19797 18408 19809 18411
rect 19668 18380 19809 18408
rect 19668 18368 19674 18380
rect 19797 18377 19809 18380
rect 19843 18377 19855 18411
rect 19797 18371 19855 18377
rect 18690 18349 18696 18352
rect 18662 18343 18696 18349
rect 18662 18340 18674 18343
rect 15028 18312 18674 18340
rect 18662 18309 18674 18312
rect 18662 18303 18696 18309
rect 18690 18300 18696 18303
rect 18748 18300 18754 18352
rect 19150 18300 19156 18352
rect 19208 18340 19214 18352
rect 20165 18343 20223 18349
rect 20165 18340 20177 18343
rect 19208 18312 20177 18340
rect 19208 18300 19214 18312
rect 20165 18309 20177 18312
rect 20211 18309 20223 18343
rect 20165 18303 20223 18309
rect 9582 18232 9588 18284
rect 9640 18272 9646 18284
rect 10287 18275 10345 18281
rect 10287 18272 10299 18275
rect 9640 18244 10299 18272
rect 9640 18232 9646 18244
rect 10287 18241 10299 18244
rect 10333 18272 10345 18275
rect 11808 18272 11836 18300
rect 11943 18275 12001 18281
rect 11943 18272 11955 18275
rect 10333 18244 11482 18272
rect 11808 18244 11955 18272
rect 10333 18241 10345 18244
rect 10287 18235 10345 18241
rect 9950 18204 9956 18216
rect 9382 18176 9956 18204
rect 9950 18164 9956 18176
rect 10008 18204 10014 18216
rect 10045 18207 10103 18213
rect 10045 18204 10057 18207
rect 10008 18176 10057 18204
rect 10008 18164 10014 18176
rect 10045 18173 10057 18176
rect 10091 18173 10103 18207
rect 10045 18167 10103 18173
rect 9490 18136 9496 18148
rect 9324 18108 9496 18136
rect 9490 18096 9496 18108
rect 9548 18096 9554 18148
rect 7650 18068 7656 18080
rect 7300 18040 7656 18068
rect 7650 18028 7656 18040
rect 7708 18028 7714 18080
rect 8297 18071 8355 18077
rect 8297 18037 8309 18071
rect 8343 18068 8355 18071
rect 9950 18068 9956 18080
rect 8343 18040 9956 18068
rect 8343 18037 8355 18040
rect 8297 18031 8355 18037
rect 9950 18028 9956 18040
rect 10008 18028 10014 18080
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 10778 18068 10784 18080
rect 10560 18040 10784 18068
rect 10560 18028 10566 18040
rect 10778 18028 10784 18040
rect 10836 18028 10842 18080
rect 11454 18068 11482 18244
rect 11943 18241 11955 18244
rect 11989 18241 12001 18275
rect 14292 18272 14320 18300
rect 14427 18275 14485 18281
rect 14427 18272 14439 18275
rect 11943 18235 12001 18241
rect 12452 18244 14439 18272
rect 12452 18216 12480 18244
rect 14427 18241 14439 18244
rect 14473 18241 14485 18275
rect 14427 18235 14485 18241
rect 15378 18232 15384 18284
rect 15436 18272 15442 18284
rect 16206 18272 16212 18284
rect 15436 18244 16212 18272
rect 15436 18232 15442 18244
rect 16206 18232 16212 18244
rect 16264 18232 16270 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18417 18275 18475 18281
rect 18417 18272 18429 18275
rect 18012 18244 18429 18272
rect 18012 18232 18018 18244
rect 18417 18241 18429 18244
rect 18463 18241 18475 18275
rect 18417 18235 18475 18241
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 11701 18207 11759 18213
rect 11701 18204 11713 18207
rect 11572 18176 11713 18204
rect 11572 18164 11578 18176
rect 11701 18173 11713 18176
rect 11747 18173 11759 18207
rect 11701 18167 11759 18173
rect 12434 18164 12440 18216
rect 12492 18164 12498 18216
rect 12894 18164 12900 18216
rect 12952 18204 12958 18216
rect 13538 18204 13544 18216
rect 12952 18176 13544 18204
rect 12952 18164 12958 18176
rect 13538 18164 13544 18176
rect 13596 18164 13602 18216
rect 14090 18164 14096 18216
rect 14148 18204 14154 18216
rect 14185 18207 14243 18213
rect 14185 18204 14197 18207
rect 14148 18176 14197 18204
rect 14148 18164 14154 18176
rect 14185 18173 14197 18176
rect 14231 18173 14243 18207
rect 14185 18167 14243 18173
rect 15102 18164 15108 18216
rect 15160 18204 15166 18216
rect 17310 18204 17316 18216
rect 15160 18176 17316 18204
rect 15160 18164 15166 18176
rect 17310 18164 17316 18176
rect 17368 18164 17374 18216
rect 12360 18108 12846 18136
rect 12360 18068 12388 18108
rect 11454 18040 12388 18068
rect 12618 18028 12624 18080
rect 12676 18068 12682 18080
rect 12713 18071 12771 18077
rect 12713 18068 12725 18071
rect 12676 18040 12725 18068
rect 12676 18028 12682 18040
rect 12713 18037 12725 18040
rect 12759 18037 12771 18071
rect 12818 18068 12846 18108
rect 16390 18068 16396 18080
rect 12818 18040 16396 18068
rect 12713 18031 12771 18037
rect 16390 18028 16396 18040
rect 16448 18028 16454 18080
rect 20441 18071 20499 18077
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 20990 18068 20996 18080
rect 20487 18040 20996 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 1104 17978 20884 18000
rect 1104 17926 3422 17978
rect 3474 17926 3486 17978
rect 3538 17926 3550 17978
rect 3602 17926 3614 17978
rect 3666 17926 3678 17978
rect 3730 17926 8367 17978
rect 8419 17926 8431 17978
rect 8483 17926 8495 17978
rect 8547 17926 8559 17978
rect 8611 17926 8623 17978
rect 8675 17926 13312 17978
rect 13364 17926 13376 17978
rect 13428 17926 13440 17978
rect 13492 17926 13504 17978
rect 13556 17926 13568 17978
rect 13620 17926 18257 17978
rect 18309 17926 18321 17978
rect 18373 17926 18385 17978
rect 18437 17926 18449 17978
rect 18501 17926 18513 17978
rect 18565 17926 20884 17978
rect 1104 17904 20884 17926
rect 1581 17867 1639 17873
rect 1581 17833 1593 17867
rect 1627 17864 1639 17867
rect 1670 17864 1676 17876
rect 1627 17836 1676 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 1670 17824 1676 17836
rect 1728 17824 1734 17876
rect 2222 17864 2228 17876
rect 1780 17836 2228 17864
rect 1302 17756 1308 17808
rect 1360 17796 1366 17808
rect 1780 17796 1808 17836
rect 2222 17824 2228 17836
rect 2280 17824 2286 17876
rect 2682 17824 2688 17876
rect 2740 17824 2746 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17833 3387 17867
rect 7098 17864 7104 17876
rect 3329 17827 3387 17833
rect 6196 17836 7104 17864
rect 1360 17768 1808 17796
rect 1360 17756 1366 17768
rect 1854 17756 1860 17808
rect 1912 17796 1918 17808
rect 3344 17796 3372 17827
rect 1912 17768 3372 17796
rect 1912 17756 1918 17768
rect 842 17688 848 17740
rect 900 17728 906 17740
rect 1578 17728 1584 17740
rect 900 17700 1584 17728
rect 900 17688 906 17700
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 2222 17688 2228 17740
rect 2280 17728 2286 17740
rect 2406 17728 2412 17740
rect 2280 17700 2412 17728
rect 2280 17688 2286 17700
rect 2406 17688 2412 17700
rect 2464 17688 2470 17740
rect 6196 17737 6224 17836
rect 7098 17824 7104 17836
rect 7156 17864 7162 17876
rect 7466 17864 7472 17876
rect 7156 17836 7472 17864
rect 7156 17824 7162 17836
rect 7466 17824 7472 17836
rect 7524 17824 7530 17876
rect 12268 17836 13676 17864
rect 6181 17731 6239 17737
rect 3344 17700 3818 17728
rect 3344 17672 3372 17700
rect 6181 17697 6193 17731
rect 6227 17697 6239 17731
rect 6181 17691 6239 17697
rect 6822 17688 6828 17740
rect 6880 17688 6886 17740
rect 6914 17688 6920 17740
rect 6972 17728 6978 17740
rect 7218 17731 7276 17737
rect 7218 17728 7230 17731
rect 6972 17700 7230 17728
rect 6972 17688 6978 17700
rect 7218 17697 7230 17700
rect 7264 17697 7276 17731
rect 7218 17691 7276 17697
rect 8846 17688 8852 17740
rect 8904 17728 8910 17740
rect 8904 17700 9982 17728
rect 8904 17688 8910 17700
rect 11514 17688 11520 17740
rect 11572 17728 11578 17740
rect 12268 17737 12296 17836
rect 13648 17796 13676 17836
rect 13722 17824 13728 17876
rect 13780 17864 13786 17876
rect 13780 17836 15516 17864
rect 13780 17824 13786 17836
rect 14550 17796 14556 17808
rect 13648 17768 14556 17796
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 15488 17796 15516 17836
rect 15562 17824 15568 17876
rect 15620 17864 15626 17876
rect 15749 17867 15807 17873
rect 15749 17864 15761 17867
rect 15620 17836 15761 17864
rect 15620 17824 15626 17836
rect 15749 17833 15761 17836
rect 15795 17833 15807 17867
rect 16574 17864 16580 17876
rect 15749 17827 15807 17833
rect 16224 17836 16580 17864
rect 16224 17796 16252 17836
rect 16574 17824 16580 17836
rect 16632 17824 16638 17876
rect 19242 17824 19248 17876
rect 19300 17824 19306 17876
rect 20254 17824 20260 17876
rect 20312 17824 20318 17876
rect 15488 17768 16252 17796
rect 12253 17731 12311 17737
rect 12253 17728 12265 17731
rect 11572 17700 12265 17728
rect 11572 17688 11578 17700
rect 12253 17697 12265 17700
rect 12299 17697 12311 17731
rect 12253 17691 12311 17697
rect 14090 17688 14096 17740
rect 14148 17728 14154 17740
rect 14737 17731 14795 17737
rect 14737 17728 14749 17731
rect 14148 17700 14749 17728
rect 14148 17688 14154 17700
rect 14737 17697 14749 17700
rect 14783 17697 14795 17731
rect 19260 17728 19288 17824
rect 14737 17691 14795 17697
rect 19076 17700 19288 17728
rect 1486 17620 1492 17672
rect 1544 17620 1550 17672
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2087 17632 3096 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2593 17595 2651 17601
rect 2593 17592 2605 17595
rect 1504 17564 2605 17592
rect 1504 17536 1532 17564
rect 2593 17561 2605 17564
rect 2639 17561 2651 17595
rect 2593 17555 2651 17561
rect 1486 17484 1492 17536
rect 1544 17484 1550 17536
rect 2130 17484 2136 17536
rect 2188 17484 2194 17536
rect 3068 17533 3096 17632
rect 3142 17620 3148 17672
rect 3200 17660 3206 17672
rect 3237 17663 3295 17669
rect 3237 17660 3249 17663
rect 3200 17632 3249 17660
rect 3200 17620 3206 17632
rect 3237 17629 3249 17632
rect 3283 17629 3295 17663
rect 3237 17623 3295 17629
rect 3326 17620 3332 17672
rect 3384 17620 3390 17672
rect 3510 17620 3516 17672
rect 3568 17620 3574 17672
rect 4249 17663 4307 17669
rect 4249 17629 4261 17663
rect 4295 17660 4307 17663
rect 4430 17660 4436 17672
rect 4295 17632 4436 17660
rect 4295 17629 4307 17632
rect 4249 17623 4307 17629
rect 4430 17620 4436 17632
rect 4488 17620 4494 17672
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 4890 17660 4896 17672
rect 4755 17632 4896 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 4890 17620 4896 17632
rect 4948 17660 4954 17672
rect 6365 17663 6423 17669
rect 4948 17632 5764 17660
rect 4948 17620 4954 17632
rect 5736 17604 5764 17632
rect 6365 17629 6377 17663
rect 6411 17660 6423 17663
rect 6546 17660 6552 17672
rect 6411 17632 6552 17660
rect 6411 17629 6423 17632
rect 6365 17623 6423 17629
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 7098 17620 7104 17672
rect 7156 17620 7162 17672
rect 7384 17620 7390 17672
rect 7442 17620 7448 17672
rect 9674 17620 9680 17672
rect 9732 17660 9738 17672
rect 10226 17660 10232 17672
rect 9732 17632 10232 17660
rect 9732 17620 9738 17632
rect 10226 17620 10232 17632
rect 10284 17660 10290 17672
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 10284 17632 10425 17660
rect 10284 17620 10290 17632
rect 10413 17629 10425 17632
rect 10459 17660 10471 17663
rect 12066 17660 12072 17672
rect 10459 17632 12072 17660
rect 10459 17629 10471 17632
rect 10413 17623 10471 17629
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 12495 17663 12553 17669
rect 12495 17629 12507 17663
rect 12541 17629 12553 17663
rect 12495 17623 12553 17629
rect 3602 17552 3608 17604
rect 3660 17592 3666 17604
rect 4341 17595 4399 17601
rect 4341 17592 4353 17595
rect 3660 17564 4353 17592
rect 3660 17552 3666 17564
rect 4341 17561 4353 17564
rect 4387 17561 4399 17595
rect 4341 17555 4399 17561
rect 5074 17552 5080 17604
rect 5132 17592 5138 17604
rect 5132 17564 5488 17592
rect 5132 17552 5138 17564
rect 5460 17536 5488 17564
rect 5718 17552 5724 17604
rect 5776 17552 5782 17604
rect 9398 17552 9404 17604
rect 9456 17592 9462 17604
rect 10042 17592 10048 17604
rect 9456 17564 10048 17592
rect 9456 17552 9462 17564
rect 10042 17552 10048 17564
rect 10100 17592 10106 17604
rect 10137 17595 10195 17601
rect 10137 17592 10149 17595
rect 10100 17564 10149 17592
rect 10100 17552 10106 17564
rect 10137 17561 10149 17564
rect 10183 17561 10195 17595
rect 10137 17555 10195 17561
rect 10502 17552 10508 17604
rect 10560 17552 10566 17604
rect 10778 17592 10784 17604
rect 10612 17564 10784 17592
rect 10612 17536 10640 17564
rect 10778 17552 10784 17564
rect 10836 17592 10842 17604
rect 10873 17595 10931 17601
rect 10873 17592 10885 17595
rect 10836 17564 10885 17592
rect 10836 17552 10842 17564
rect 10873 17561 10885 17564
rect 10919 17561 10931 17595
rect 10873 17555 10931 17561
rect 10962 17552 10968 17604
rect 11020 17592 11026 17604
rect 11698 17592 11704 17604
rect 11020 17564 11704 17592
rect 11020 17552 11026 17564
rect 11698 17552 11704 17564
rect 11756 17592 11762 17604
rect 12510 17592 12538 17623
rect 13170 17620 13176 17672
rect 13228 17660 13234 17672
rect 13722 17660 13728 17672
rect 13228 17632 13728 17660
rect 13228 17620 13234 17632
rect 13722 17620 13728 17632
rect 13780 17620 13786 17672
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14366 17660 14372 17672
rect 13872 17632 14372 17660
rect 13872 17620 13878 17632
rect 14366 17620 14372 17632
rect 14424 17660 14430 17672
rect 14979 17663 15037 17669
rect 14979 17660 14991 17663
rect 14424 17632 14991 17660
rect 14424 17620 14430 17632
rect 14979 17629 14991 17632
rect 15025 17629 15037 17663
rect 14979 17623 15037 17629
rect 16117 17663 16175 17669
rect 16117 17629 16129 17663
rect 16163 17629 16175 17663
rect 16390 17660 16396 17672
rect 16351 17632 16396 17660
rect 16117 17623 16175 17629
rect 14458 17592 14464 17604
rect 11756 17564 12538 17592
rect 12887 17564 14464 17592
rect 11756 17552 11762 17564
rect 3053 17527 3111 17533
rect 3053 17493 3065 17527
rect 3099 17493 3111 17527
rect 3053 17487 3111 17493
rect 3970 17484 3976 17536
rect 4028 17484 4034 17536
rect 5166 17484 5172 17536
rect 5224 17524 5230 17536
rect 5261 17527 5319 17533
rect 5261 17524 5273 17527
rect 5224 17496 5273 17524
rect 5224 17484 5230 17496
rect 5261 17493 5273 17496
rect 5307 17524 5319 17527
rect 5350 17524 5356 17536
rect 5307 17496 5356 17524
rect 5307 17493 5319 17496
rect 5261 17487 5319 17493
rect 5350 17484 5356 17496
rect 5408 17484 5414 17536
rect 5442 17484 5448 17536
rect 5500 17484 5506 17536
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 7190 17524 7196 17536
rect 5960 17496 7196 17524
rect 5960 17484 5966 17496
rect 7190 17484 7196 17496
rect 7248 17484 7254 17536
rect 8018 17484 8024 17536
rect 8076 17484 8082 17536
rect 10594 17484 10600 17536
rect 10652 17484 10658 17536
rect 11238 17484 11244 17536
rect 11296 17484 11302 17536
rect 11425 17527 11483 17533
rect 11425 17493 11437 17527
rect 11471 17524 11483 17527
rect 12250 17524 12256 17536
rect 11471 17496 12256 17524
rect 11471 17493 11483 17496
rect 11425 17487 11483 17493
rect 12250 17484 12256 17496
rect 12308 17524 12314 17536
rect 12887 17524 12915 17564
rect 14458 17552 14464 17564
rect 14516 17592 14522 17604
rect 14826 17592 14832 17604
rect 14516 17564 14832 17592
rect 14516 17552 14522 17564
rect 14826 17552 14832 17564
rect 14884 17552 14890 17604
rect 16132 17592 16160 17623
rect 16390 17620 16396 17632
rect 16448 17620 16454 17672
rect 19076 17669 19104 17700
rect 18877 17663 18935 17669
rect 18877 17629 18889 17663
rect 18923 17629 18935 17663
rect 18877 17623 18935 17629
rect 19061 17663 19119 17669
rect 19061 17629 19073 17663
rect 19107 17629 19119 17663
rect 19061 17623 19119 17629
rect 16666 17592 16672 17604
rect 16132 17564 16672 17592
rect 16666 17552 16672 17564
rect 16724 17592 16730 17604
rect 18046 17592 18052 17604
rect 16724 17564 18052 17592
rect 16724 17552 16730 17564
rect 18046 17552 18052 17564
rect 18104 17552 18110 17604
rect 12308 17496 12915 17524
rect 12308 17484 12314 17496
rect 13078 17484 13084 17536
rect 13136 17524 13142 17536
rect 13265 17527 13323 17533
rect 13265 17524 13277 17527
rect 13136 17496 13277 17524
rect 13136 17484 13142 17496
rect 13265 17493 13277 17496
rect 13311 17493 13323 17527
rect 13265 17487 13323 17493
rect 13998 17484 14004 17536
rect 14056 17524 14062 17536
rect 15194 17524 15200 17536
rect 14056 17496 15200 17524
rect 14056 17484 14062 17496
rect 15194 17484 15200 17496
rect 15252 17484 15258 17536
rect 15286 17484 15292 17536
rect 15344 17524 15350 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 15344 17496 17141 17524
rect 15344 17484 15350 17496
rect 17129 17493 17141 17496
rect 17175 17493 17187 17527
rect 18892 17524 18920 17623
rect 19150 17620 19156 17672
rect 19208 17660 19214 17672
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 19208 17632 19257 17660
rect 19208 17620 19214 17632
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 19487 17663 19545 17669
rect 19487 17629 19499 17663
rect 19533 17660 19545 17663
rect 19610 17660 19616 17672
rect 19533 17632 19616 17660
rect 19533 17629 19545 17632
rect 19487 17623 19545 17629
rect 19610 17620 19616 17632
rect 19668 17620 19674 17672
rect 20530 17620 20536 17672
rect 20588 17620 20594 17672
rect 18969 17595 19027 17601
rect 18969 17561 18981 17595
rect 19015 17592 19027 17595
rect 20548 17592 20576 17620
rect 19015 17564 20576 17592
rect 19015 17561 19027 17564
rect 18969 17555 19027 17561
rect 20254 17524 20260 17536
rect 18892 17496 20260 17524
rect 17129 17487 17187 17493
rect 20254 17484 20260 17496
rect 20312 17484 20318 17536
rect 1104 17434 21043 17456
rect 1104 17382 5894 17434
rect 5946 17382 5958 17434
rect 6010 17382 6022 17434
rect 6074 17382 6086 17434
rect 6138 17382 6150 17434
rect 6202 17382 10839 17434
rect 10891 17382 10903 17434
rect 10955 17382 10967 17434
rect 11019 17382 11031 17434
rect 11083 17382 11095 17434
rect 11147 17382 15784 17434
rect 15836 17382 15848 17434
rect 15900 17382 15912 17434
rect 15964 17382 15976 17434
rect 16028 17382 16040 17434
rect 16092 17382 20729 17434
rect 20781 17382 20793 17434
rect 20845 17382 20857 17434
rect 20909 17382 20921 17434
rect 20973 17382 20985 17434
rect 21037 17382 21043 17434
rect 1104 17360 21043 17382
rect 1578 17280 1584 17332
rect 1636 17280 1642 17332
rect 1946 17280 1952 17332
rect 2004 17320 2010 17332
rect 3053 17323 3111 17329
rect 2004 17292 3004 17320
rect 2004 17280 2010 17292
rect 2314 17223 2320 17264
rect 2299 17217 2320 17223
rect 1489 17187 1547 17193
rect 1489 17153 1501 17187
rect 1535 17184 1547 17187
rect 1946 17184 1952 17196
rect 1535 17156 1952 17184
rect 1535 17153 1547 17156
rect 1489 17147 1547 17153
rect 1946 17144 1952 17156
rect 2004 17144 2010 17196
rect 2038 17144 2044 17196
rect 2096 17144 2102 17196
rect 2299 17183 2311 17217
rect 2372 17212 2378 17264
rect 2345 17186 2360 17212
rect 2345 17183 2357 17186
rect 2299 17177 2357 17183
rect 2976 17184 3004 17292
rect 3053 17289 3065 17323
rect 3099 17320 3111 17323
rect 3602 17320 3608 17332
rect 3099 17292 3608 17320
rect 3099 17289 3111 17292
rect 3053 17283 3111 17289
rect 3602 17280 3608 17292
rect 3660 17280 3666 17332
rect 3878 17280 3884 17332
rect 3936 17320 3942 17332
rect 4433 17323 4491 17329
rect 4433 17320 4445 17323
rect 3936 17292 4445 17320
rect 3936 17280 3942 17292
rect 4433 17289 4445 17292
rect 4479 17289 4491 17323
rect 4433 17283 4491 17289
rect 5905 17323 5963 17329
rect 5905 17289 5917 17323
rect 5951 17320 5963 17323
rect 6822 17320 6828 17332
rect 5951 17292 6828 17320
rect 5951 17289 5963 17292
rect 5905 17283 5963 17289
rect 6822 17280 6828 17292
rect 6880 17280 6886 17332
rect 7374 17280 7380 17332
rect 7432 17320 7438 17332
rect 7469 17323 7527 17329
rect 7469 17320 7481 17323
rect 7432 17292 7481 17320
rect 7432 17280 7438 17292
rect 7469 17289 7481 17292
rect 7515 17289 7527 17323
rect 8018 17320 8024 17332
rect 7469 17283 7527 17289
rect 7558 17292 8024 17320
rect 4154 17252 4160 17264
rect 3436 17224 4160 17252
rect 3436 17193 3464 17224
rect 4154 17212 4160 17224
rect 4212 17212 4218 17264
rect 4522 17212 4528 17264
rect 4580 17212 4586 17264
rect 4890 17212 4896 17264
rect 4948 17252 4954 17264
rect 4948 17224 5856 17252
rect 4948 17212 4954 17224
rect 3421 17187 3479 17193
rect 3421 17184 3433 17187
rect 2976 17156 3433 17184
rect 3421 17153 3433 17156
rect 3467 17153 3479 17187
rect 3421 17147 3479 17153
rect 3695 17187 3753 17193
rect 3695 17153 3707 17187
rect 3741 17184 3753 17187
rect 4246 17184 4252 17196
rect 3741 17156 4252 17184
rect 3741 17153 3753 17156
rect 3695 17147 3753 17153
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 4540 17184 4568 17212
rect 5135 17187 5193 17193
rect 5135 17184 5147 17187
rect 4540 17156 5147 17184
rect 5135 17153 5147 17156
rect 5181 17184 5193 17187
rect 5626 17184 5632 17196
rect 5181 17156 5632 17184
rect 5181 17153 5193 17156
rect 5135 17147 5193 17153
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 2866 17076 2872 17128
rect 2924 17116 2930 17128
rect 3050 17116 3056 17128
rect 2924 17088 3056 17116
rect 2924 17076 2930 17088
rect 3050 17076 3056 17088
rect 3108 17076 3114 17128
rect 4522 17076 4528 17128
rect 4580 17116 4586 17128
rect 4890 17116 4896 17128
rect 4580 17088 4896 17116
rect 4580 17076 4586 17088
rect 4890 17076 4896 17088
rect 4948 17076 4954 17128
rect 5828 17116 5856 17224
rect 5994 17212 6000 17264
rect 6052 17252 6058 17264
rect 7558 17252 7586 17292
rect 8018 17280 8024 17292
rect 8076 17280 8082 17332
rect 8846 17280 8852 17332
rect 8904 17280 8910 17332
rect 9398 17280 9404 17332
rect 9456 17280 9462 17332
rect 9766 17280 9772 17332
rect 9824 17280 9830 17332
rect 10410 17280 10416 17332
rect 10468 17320 10474 17332
rect 14458 17320 14464 17332
rect 10468 17292 13768 17320
rect 10468 17280 10474 17292
rect 9784 17252 9812 17280
rect 6052 17224 7586 17252
rect 7622 17224 9812 17252
rect 6052 17212 6058 17224
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 6699 17187 6757 17193
rect 6699 17184 6711 17187
rect 5960 17156 6711 17184
rect 5960 17144 5966 17156
rect 6699 17153 6711 17156
rect 6745 17153 6757 17187
rect 7622 17184 7650 17224
rect 9950 17212 9956 17264
rect 10008 17212 10014 17264
rect 10505 17255 10563 17261
rect 10505 17221 10517 17255
rect 10551 17252 10563 17255
rect 12066 17252 12072 17264
rect 10551 17224 11284 17252
rect 10551 17221 10563 17224
rect 10505 17215 10563 17221
rect 6699 17147 6757 17153
rect 7114 17156 7650 17184
rect 8111 17187 8169 17193
rect 6457 17119 6515 17125
rect 6457 17116 6469 17119
rect 5828 17088 6469 17116
rect 6457 17085 6469 17088
rect 6503 17085 6515 17119
rect 6457 17079 6515 17085
rect 2958 17008 2964 17060
rect 3016 17048 3022 17060
rect 3418 17048 3424 17060
rect 3016 17020 3424 17048
rect 3016 17008 3022 17020
rect 3418 17008 3424 17020
rect 3476 17008 3482 17060
rect 2774 16940 2780 16992
rect 2832 16980 2838 16992
rect 5994 16980 6000 16992
rect 2832 16952 6000 16980
rect 2832 16940 2838 16952
rect 5994 16940 6000 16952
rect 6052 16940 6058 16992
rect 6472 16980 6500 17079
rect 7114 16980 7142 17156
rect 8111 17153 8123 17187
rect 8157 17184 8169 17187
rect 8157 17156 9168 17184
rect 8157 17153 8169 17156
rect 8111 17147 8169 17153
rect 7558 17076 7564 17128
rect 7616 17116 7622 17128
rect 7837 17119 7895 17125
rect 7837 17116 7849 17119
rect 7616 17088 7849 17116
rect 7616 17076 7622 17088
rect 7837 17085 7849 17088
rect 7883 17085 7895 17119
rect 7837 17079 7895 17085
rect 6472 16952 7142 16980
rect 7282 16940 7288 16992
rect 7340 16980 7346 16992
rect 8754 16980 8760 16992
rect 7340 16952 8760 16980
rect 7340 16940 7346 16952
rect 8754 16940 8760 16952
rect 8812 16940 8818 16992
rect 9140 16980 9168 17156
rect 9674 17144 9680 17196
rect 9732 17144 9738 17196
rect 9769 17187 9827 17193
rect 9769 17153 9781 17187
rect 9815 17184 9827 17187
rect 9968 17184 9996 17212
rect 11256 17196 11284 17224
rect 11900 17224 12072 17252
rect 9815 17156 9996 17184
rect 10137 17187 10195 17193
rect 9815 17153 9827 17156
rect 9769 17147 9827 17153
rect 10137 17153 10149 17187
rect 10183 17184 10195 17187
rect 10594 17184 10600 17196
rect 10183 17156 10600 17184
rect 10183 17153 10195 17156
rect 10137 17147 10195 17153
rect 10594 17144 10600 17156
rect 10652 17184 10658 17196
rect 10778 17184 10784 17196
rect 10652 17156 10784 17184
rect 10652 17144 10658 17156
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 11238 17144 11244 17196
rect 11296 17144 11302 17196
rect 11900 17193 11928 17224
rect 12066 17212 12072 17224
rect 12124 17212 12130 17264
rect 13740 17261 13768 17292
rect 14016 17292 14464 17320
rect 13725 17255 13783 17261
rect 13725 17221 13737 17255
rect 13771 17221 13783 17255
rect 13725 17215 13783 17221
rect 11885 17187 11943 17193
rect 11885 17153 11897 17187
rect 11931 17153 11943 17187
rect 11885 17147 11943 17153
rect 13078 17144 13084 17196
rect 13136 17144 13142 17196
rect 13906 17184 13912 17196
rect 13740 17156 13912 17184
rect 9220 17128 9272 17134
rect 10796 17116 10824 17144
rect 12069 17119 12127 17125
rect 12069 17116 12081 17119
rect 10796 17088 12081 17116
rect 12069 17085 12081 17088
rect 12115 17085 12127 17119
rect 12805 17119 12863 17125
rect 12805 17116 12817 17119
rect 12069 17079 12127 17085
rect 12636 17088 12817 17116
rect 9220 17070 9272 17076
rect 12529 17051 12587 17057
rect 12529 17048 12541 17051
rect 12084 17020 12541 17048
rect 12084 16992 12112 17020
rect 12529 17017 12541 17020
rect 12575 17017 12587 17051
rect 12529 17011 12587 17017
rect 9306 16980 9312 16992
rect 9140 16952 9312 16980
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 10594 16940 10600 16992
rect 10652 16980 10658 16992
rect 10689 16983 10747 16989
rect 10689 16980 10701 16983
rect 10652 16952 10701 16980
rect 10652 16940 10658 16952
rect 10689 16949 10701 16952
rect 10735 16949 10747 16983
rect 10689 16943 10747 16949
rect 12066 16940 12072 16992
rect 12124 16940 12130 16992
rect 12636 16980 12664 17088
rect 12805 17085 12817 17088
rect 12851 17085 12863 17119
rect 12805 17079 12863 17085
rect 12943 17119 13001 17125
rect 12943 17085 12955 17119
rect 12989 17116 13001 17119
rect 13740 17116 13768 17156
rect 13906 17144 13912 17156
rect 13964 17144 13970 17196
rect 14016 17193 14044 17292
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 15470 17280 15476 17332
rect 15528 17320 15534 17332
rect 15746 17320 15752 17332
rect 15528 17292 15752 17320
rect 15528 17280 15534 17292
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 17494 17280 17500 17332
rect 17552 17280 17558 17332
rect 19702 17280 19708 17332
rect 19760 17320 19766 17332
rect 20441 17323 20499 17329
rect 19760 17292 20208 17320
rect 19760 17280 19766 17292
rect 15856 17224 16896 17252
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17153 14059 17187
rect 14001 17147 14059 17153
rect 14826 17144 14832 17196
rect 14884 17193 14890 17196
rect 14884 17187 14912 17193
rect 14900 17153 14912 17187
rect 14884 17147 14912 17153
rect 14884 17144 14890 17147
rect 12989 17088 13768 17116
rect 13817 17119 13875 17125
rect 12989 17085 13001 17088
rect 12943 17079 13001 17085
rect 13817 17085 13829 17119
rect 13863 17116 13875 17119
rect 14182 17116 14188 17128
rect 13863 17088 14188 17116
rect 13863 17085 13875 17088
rect 13817 17079 13875 17085
rect 13832 17048 13860 17079
rect 14182 17076 14188 17088
rect 14240 17076 14246 17128
rect 14737 17119 14795 17125
rect 14737 17116 14749 17119
rect 14571 17088 14749 17116
rect 13740 17020 13860 17048
rect 12986 16980 12992 16992
rect 12636 16952 12992 16980
rect 12986 16940 12992 16952
rect 13044 16940 13050 16992
rect 13170 16940 13176 16992
rect 13228 16980 13234 16992
rect 13740 16980 13768 17020
rect 14090 17008 14096 17060
rect 14148 17048 14154 17060
rect 14461 17051 14519 17057
rect 14461 17048 14473 17051
rect 14148 17020 14473 17048
rect 14148 17008 14154 17020
rect 14461 17017 14473 17020
rect 14507 17017 14519 17051
rect 14461 17011 14519 17017
rect 13228 16952 13768 16980
rect 14571 16980 14599 17088
rect 14737 17085 14749 17088
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17116 15071 17119
rect 15194 17116 15200 17128
rect 15059 17088 15200 17116
rect 15059 17085 15071 17088
rect 15013 17079 15071 17085
rect 15194 17076 15200 17088
rect 15252 17076 15258 17128
rect 15378 17076 15384 17128
rect 15436 17116 15442 17128
rect 15856 17116 15884 17224
rect 16868 17184 16896 17224
rect 16943 17187 17001 17193
rect 16943 17184 16955 17187
rect 16868 17156 16955 17184
rect 16943 17153 16955 17156
rect 16989 17184 17001 17187
rect 17512 17184 17540 17280
rect 17770 17212 17776 17264
rect 17828 17252 17834 17264
rect 19610 17252 19616 17264
rect 17828 17224 19616 17252
rect 17828 17212 17834 17224
rect 19610 17212 19616 17224
rect 19668 17212 19674 17264
rect 20180 17261 20208 17292
rect 20441 17289 20453 17323
rect 20487 17320 20499 17323
rect 21266 17320 21272 17332
rect 20487 17292 21272 17320
rect 20487 17289 20499 17292
rect 20441 17283 20499 17289
rect 21266 17280 21272 17292
rect 21324 17280 21330 17332
rect 20165 17255 20223 17261
rect 20165 17221 20177 17255
rect 20211 17221 20223 17255
rect 20165 17215 20223 17221
rect 16989 17156 17540 17184
rect 16989 17153 17001 17156
rect 16943 17147 17001 17153
rect 17954 17144 17960 17196
rect 18012 17144 18018 17196
rect 18046 17144 18052 17196
rect 18104 17184 18110 17196
rect 18489 17187 18547 17193
rect 18489 17184 18501 17187
rect 18104 17156 18501 17184
rect 18104 17144 18110 17156
rect 18489 17153 18501 17156
rect 18535 17184 18547 17187
rect 18782 17184 18788 17196
rect 18535 17156 18788 17184
rect 18535 17153 18547 17156
rect 18489 17147 18547 17153
rect 18782 17144 18788 17156
rect 18840 17144 18846 17196
rect 19705 17187 19763 17193
rect 19705 17153 19717 17187
rect 19751 17184 19763 17187
rect 19978 17184 19984 17196
rect 19751 17156 19984 17184
rect 19751 17153 19763 17156
rect 19705 17147 19763 17153
rect 19978 17144 19984 17156
rect 20036 17144 20042 17196
rect 15436 17088 15884 17116
rect 15436 17076 15442 17088
rect 16666 17076 16672 17128
rect 16724 17076 16730 17128
rect 17972 17116 18000 17144
rect 18233 17119 18291 17125
rect 18233 17116 18245 17119
rect 17972 17088 18245 17116
rect 18233 17085 18245 17088
rect 18279 17085 18291 17119
rect 18233 17079 18291 17085
rect 14826 16980 14832 16992
rect 14571 16952 14832 16980
rect 13228 16940 13234 16952
rect 14826 16940 14832 16952
rect 14884 16980 14890 16992
rect 15102 16980 15108 16992
rect 14884 16952 15108 16980
rect 14884 16940 14890 16952
rect 15102 16940 15108 16952
rect 15160 16940 15166 16992
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15528 16952 15669 16980
rect 15528 16940 15534 16952
rect 15657 16949 15669 16952
rect 15703 16949 15715 16983
rect 15657 16943 15715 16949
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 17681 16983 17739 16989
rect 17681 16980 17693 16983
rect 16264 16952 17693 16980
rect 16264 16940 16270 16952
rect 17681 16949 17693 16952
rect 17727 16949 17739 16983
rect 17681 16943 17739 16949
rect 17862 16940 17868 16992
rect 17920 16980 17926 16992
rect 18046 16980 18052 16992
rect 17920 16952 18052 16980
rect 17920 16940 17926 16952
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 19613 16983 19671 16989
rect 19613 16949 19625 16983
rect 19659 16980 19671 16983
rect 19794 16980 19800 16992
rect 19659 16952 19800 16980
rect 19659 16949 19671 16952
rect 19613 16943 19671 16949
rect 19794 16940 19800 16952
rect 19852 16940 19858 16992
rect 19889 16983 19947 16989
rect 19889 16949 19901 16983
rect 19935 16980 19947 16983
rect 20898 16980 20904 16992
rect 19935 16952 20904 16980
rect 19935 16949 19947 16952
rect 19889 16943 19947 16949
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 1104 16890 20884 16912
rect 1104 16838 3422 16890
rect 3474 16838 3486 16890
rect 3538 16838 3550 16890
rect 3602 16838 3614 16890
rect 3666 16838 3678 16890
rect 3730 16838 8367 16890
rect 8419 16838 8431 16890
rect 8483 16838 8495 16890
rect 8547 16838 8559 16890
rect 8611 16838 8623 16890
rect 8675 16838 13312 16890
rect 13364 16838 13376 16890
rect 13428 16838 13440 16890
rect 13492 16838 13504 16890
rect 13556 16838 13568 16890
rect 13620 16838 18257 16890
rect 18309 16838 18321 16890
rect 18373 16838 18385 16890
rect 18437 16838 18449 16890
rect 18501 16838 18513 16890
rect 18565 16838 20884 16890
rect 1104 16816 20884 16838
rect 1762 16736 1768 16788
rect 1820 16736 1826 16788
rect 2682 16776 2688 16788
rect 1872 16748 2688 16776
rect 1118 16668 1124 16720
rect 1176 16708 1182 16720
rect 1872 16708 1900 16748
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 3326 16736 3332 16788
rect 3384 16736 3390 16788
rect 4264 16748 6592 16776
rect 1176 16680 1900 16708
rect 1176 16668 1182 16680
rect 3050 16668 3056 16720
rect 3108 16708 3114 16720
rect 3789 16711 3847 16717
rect 3789 16708 3801 16711
rect 3108 16680 3801 16708
rect 3108 16668 3114 16680
rect 3789 16677 3801 16680
rect 3835 16677 3847 16711
rect 3789 16671 3847 16677
rect 2038 16600 2044 16652
rect 2096 16640 2102 16652
rect 2317 16643 2375 16649
rect 2317 16640 2329 16643
rect 2096 16612 2329 16640
rect 2096 16600 2102 16612
rect 2317 16609 2329 16612
rect 2363 16609 2375 16643
rect 2317 16603 2375 16609
rect 3804 16612 4154 16640
rect 3804 16584 3832 16612
rect 2591 16575 2649 16581
rect 2591 16541 2603 16575
rect 2637 16572 2649 16575
rect 2958 16572 2964 16584
rect 2637 16544 2964 16572
rect 2637 16541 2649 16544
rect 2591 16535 2649 16541
rect 2958 16532 2964 16544
rect 3016 16572 3022 16584
rect 3016 16544 3372 16572
rect 3016 16532 3022 16544
rect 3344 16516 3372 16544
rect 3786 16532 3792 16584
rect 3844 16532 3850 16584
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 198 16464 204 16516
rect 256 16504 262 16516
rect 658 16504 664 16516
rect 256 16476 664 16504
rect 256 16464 262 16476
rect 658 16464 664 16476
rect 716 16464 722 16516
rect 1673 16507 1731 16513
rect 1673 16473 1685 16507
rect 1719 16504 1731 16507
rect 3050 16504 3056 16516
rect 1719 16476 3056 16504
rect 1719 16473 1731 16476
rect 1673 16467 1731 16473
rect 3050 16464 3056 16476
rect 3108 16464 3114 16516
rect 3326 16464 3332 16516
rect 3384 16464 3390 16516
rect 4126 16504 4154 16612
rect 4264 16581 4292 16748
rect 5350 16668 5356 16720
rect 5408 16668 5414 16720
rect 6564 16708 6592 16748
rect 6638 16736 6644 16788
rect 6696 16776 6702 16788
rect 6733 16779 6791 16785
rect 6733 16776 6745 16779
rect 6696 16748 6745 16776
rect 6696 16736 6702 16748
rect 6733 16745 6745 16748
rect 6779 16745 6791 16779
rect 6733 16739 6791 16745
rect 6822 16736 6828 16788
rect 6880 16776 6886 16788
rect 7006 16776 7012 16788
rect 6880 16748 7012 16776
rect 6880 16736 6886 16748
rect 7006 16736 7012 16748
rect 7064 16736 7070 16788
rect 9950 16776 9956 16788
rect 7576 16748 9956 16776
rect 7576 16708 7604 16748
rect 9950 16736 9956 16748
rect 10008 16736 10014 16788
rect 11330 16736 11336 16788
rect 11388 16776 11394 16788
rect 14090 16776 14096 16788
rect 11388 16748 12664 16776
rect 11388 16736 11394 16748
rect 6564 16680 7604 16708
rect 8481 16711 8539 16717
rect 8481 16677 8493 16711
rect 8527 16677 8539 16711
rect 8481 16671 8539 16677
rect 11241 16711 11299 16717
rect 11241 16677 11253 16711
rect 11287 16708 11299 16711
rect 11287 16680 11468 16708
rect 11287 16677 11299 16680
rect 11241 16671 11299 16677
rect 5721 16643 5779 16649
rect 5721 16640 5733 16643
rect 5000 16612 5733 16640
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4341 16575 4399 16581
rect 4341 16541 4353 16575
rect 4387 16541 4399 16575
rect 4341 16535 4399 16541
rect 4615 16575 4673 16581
rect 4615 16541 4627 16575
rect 4661 16541 4673 16575
rect 4615 16535 4673 16541
rect 4356 16504 4384 16535
rect 3436 16476 3924 16504
rect 4126 16476 4384 16504
rect 4630 16504 4658 16535
rect 4890 16504 4896 16516
rect 4630 16476 4896 16504
rect 2314 16396 2320 16448
rect 2372 16436 2378 16448
rect 3436 16436 3464 16476
rect 2372 16408 3464 16436
rect 3896 16436 3924 16476
rect 4065 16439 4123 16445
rect 4065 16436 4077 16439
rect 3896 16408 4077 16436
rect 2372 16396 2378 16408
rect 4065 16405 4077 16408
rect 4111 16405 4123 16439
rect 4356 16436 4384 16476
rect 4890 16464 4896 16476
rect 4948 16464 4954 16516
rect 5000 16436 5028 16612
rect 5721 16609 5733 16612
rect 5767 16609 5779 16643
rect 5721 16603 5779 16609
rect 7098 16600 7104 16652
rect 7156 16640 7162 16652
rect 7374 16640 7380 16652
rect 7156 16612 7380 16640
rect 7156 16600 7162 16612
rect 7374 16600 7380 16612
rect 7432 16600 7438 16652
rect 8496 16640 8524 16671
rect 8496 16612 9674 16640
rect 5074 16532 5080 16584
rect 5132 16572 5138 16584
rect 5534 16572 5540 16584
rect 5132 16544 5540 16572
rect 5132 16532 5138 16544
rect 5534 16532 5540 16544
rect 5592 16572 5598 16584
rect 5963 16575 6021 16581
rect 5963 16572 5975 16575
rect 5592 16544 5975 16572
rect 5592 16532 5598 16544
rect 5963 16541 5975 16544
rect 6009 16541 6021 16575
rect 5963 16535 6021 16541
rect 7469 16575 7527 16581
rect 7469 16541 7481 16575
rect 7515 16572 7527 16575
rect 7742 16572 7748 16584
rect 7515 16544 7604 16572
rect 7703 16544 7748 16572
rect 7515 16541 7527 16544
rect 7469 16535 7527 16541
rect 7576 16516 7604 16544
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 9646 16572 9674 16612
rect 10134 16600 10140 16652
rect 10192 16600 10198 16652
rect 11330 16600 11336 16652
rect 11388 16600 11394 16652
rect 10321 16575 10379 16581
rect 10321 16572 10333 16575
rect 9646 16544 10333 16572
rect 10321 16541 10333 16544
rect 10367 16541 10379 16575
rect 10321 16535 10379 16541
rect 10410 16532 10416 16584
rect 10468 16572 10474 16584
rect 11348 16572 11376 16600
rect 11440 16584 11468 16680
rect 12636 16640 12664 16748
rect 13004 16748 14096 16776
rect 13004 16717 13032 16748
rect 14090 16736 14096 16748
rect 14148 16736 14154 16788
rect 14182 16736 14188 16788
rect 14240 16736 14246 16788
rect 16206 16776 16212 16788
rect 14844 16748 16212 16776
rect 12989 16711 13047 16717
rect 12989 16677 13001 16711
rect 13035 16677 13047 16711
rect 14200 16708 14228 16736
rect 14844 16717 14872 16748
rect 16206 16736 16212 16748
rect 16264 16736 16270 16788
rect 17494 16776 17500 16788
rect 16408 16748 17500 16776
rect 14829 16711 14887 16717
rect 14200 16680 14318 16708
rect 12989 16671 13047 16677
rect 14185 16643 14243 16649
rect 14185 16640 14197 16643
rect 12636 16612 14197 16640
rect 14185 16609 14197 16612
rect 14231 16609 14243 16643
rect 14290 16640 14318 16680
rect 14829 16677 14841 16711
rect 14875 16677 14887 16711
rect 14829 16671 14887 16677
rect 16301 16711 16359 16717
rect 16301 16677 16313 16711
rect 16347 16677 16359 16711
rect 16301 16671 16359 16677
rect 15222 16643 15280 16649
rect 15222 16640 15234 16643
rect 14290 16612 15234 16640
rect 14185 16603 14243 16609
rect 15222 16609 15234 16612
rect 15268 16609 15280 16643
rect 15746 16640 15752 16652
rect 15222 16603 15280 16609
rect 15329 16612 15752 16640
rect 10468 16544 11376 16572
rect 10468 16532 10474 16544
rect 11422 16532 11428 16584
rect 11480 16532 11486 16584
rect 11790 16532 11796 16584
rect 11848 16572 11854 16584
rect 11977 16575 12035 16581
rect 11977 16572 11989 16575
rect 11848 16544 11989 16572
rect 11848 16532 11854 16544
rect 11977 16541 11989 16544
rect 12023 16541 12035 16575
rect 13170 16572 13176 16584
rect 12251 16565 12309 16571
rect 12251 16562 12263 16565
rect 11977 16535 12035 16541
rect 12250 16531 12263 16562
rect 12297 16531 12309 16565
rect 12250 16525 12309 16531
rect 12452 16544 13176 16572
rect 5350 16464 5356 16516
rect 5408 16504 5414 16516
rect 7006 16504 7012 16516
rect 5408 16476 7012 16504
rect 5408 16464 5414 16476
rect 7006 16464 7012 16476
rect 7064 16464 7070 16516
rect 7558 16464 7564 16516
rect 7616 16504 7622 16516
rect 8938 16504 8944 16516
rect 7616 16476 8944 16504
rect 7616 16464 7622 16476
rect 8938 16464 8944 16476
rect 8996 16464 9002 16516
rect 9858 16464 9864 16516
rect 9916 16464 9922 16516
rect 9953 16507 10011 16513
rect 9953 16473 9965 16507
rect 9999 16504 10011 16507
rect 10042 16504 10048 16516
rect 9999 16476 10048 16504
rect 9999 16473 10011 16476
rect 9953 16467 10011 16473
rect 10042 16464 10048 16476
rect 10100 16464 10106 16516
rect 10226 16464 10232 16516
rect 10284 16464 10290 16516
rect 10689 16507 10747 16513
rect 10689 16473 10701 16507
rect 10735 16504 10747 16507
rect 10778 16504 10784 16516
rect 10735 16476 10784 16504
rect 10735 16473 10747 16476
rect 10689 16467 10747 16473
rect 5810 16436 5816 16448
rect 4356 16408 5816 16436
rect 4065 16399 4123 16405
rect 5810 16396 5816 16408
rect 5868 16396 5874 16448
rect 6178 16396 6184 16448
rect 6236 16436 6242 16448
rect 6362 16436 6368 16448
rect 6236 16408 6368 16436
rect 6236 16396 6242 16408
rect 6362 16396 6368 16408
rect 6420 16396 6426 16448
rect 6546 16396 6552 16448
rect 6604 16436 6610 16448
rect 9766 16436 9772 16448
rect 6604 16408 9772 16436
rect 6604 16396 6610 16408
rect 9766 16396 9772 16408
rect 9824 16396 9830 16448
rect 9876 16436 9904 16464
rect 10704 16436 10732 16467
rect 10778 16464 10784 16476
rect 10836 16464 10842 16516
rect 12158 16504 12164 16516
rect 11348 16476 12164 16504
rect 11348 16448 11376 16476
rect 12158 16464 12164 16476
rect 12216 16504 12222 16516
rect 12250 16504 12278 16525
rect 12216 16476 12278 16504
rect 12216 16464 12222 16476
rect 9876 16408 10732 16436
rect 11057 16439 11115 16445
rect 11057 16405 11069 16439
rect 11103 16436 11115 16439
rect 11238 16436 11244 16448
rect 11103 16408 11244 16436
rect 11103 16405 11115 16408
rect 11057 16399 11115 16405
rect 11238 16396 11244 16408
rect 11296 16396 11302 16448
rect 11330 16396 11336 16448
rect 11388 16396 11394 16448
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 12452 16436 12480 16544
rect 13170 16532 13176 16544
rect 13228 16532 13234 16584
rect 13722 16532 13728 16584
rect 13780 16532 13786 16584
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 12986 16464 12992 16516
rect 13044 16504 13050 16516
rect 13740 16504 13768 16532
rect 13044 16476 13768 16504
rect 13044 16464 13050 16476
rect 11480 16408 12480 16436
rect 14384 16436 14412 16535
rect 15102 16532 15108 16584
rect 15160 16572 15166 16584
rect 15329 16572 15357 16612
rect 15746 16600 15752 16612
rect 15804 16600 15810 16652
rect 16022 16600 16028 16652
rect 16080 16600 16086 16652
rect 15160 16544 15357 16572
rect 15160 16532 15166 16544
rect 15388 16532 15394 16584
rect 15446 16532 15452 16584
rect 16117 16575 16175 16581
rect 16117 16541 16129 16575
rect 16163 16541 16175 16575
rect 16316 16572 16344 16671
rect 16408 16649 16436 16748
rect 17494 16736 17500 16748
rect 17552 16776 17558 16788
rect 17954 16776 17960 16788
rect 17552 16748 17960 16776
rect 17552 16736 17558 16748
rect 17954 16736 17960 16748
rect 18012 16736 18018 16788
rect 18785 16711 18843 16717
rect 18785 16677 18797 16711
rect 18831 16677 18843 16711
rect 18785 16671 18843 16677
rect 16393 16643 16451 16649
rect 16393 16609 16405 16643
rect 16439 16609 16451 16643
rect 16393 16603 16451 16609
rect 17420 16612 17908 16640
rect 17420 16572 17448 16612
rect 17880 16581 17908 16612
rect 17954 16600 17960 16652
rect 18012 16640 18018 16652
rect 18690 16640 18696 16652
rect 18012 16612 18696 16640
rect 18012 16600 18018 16612
rect 18690 16600 18696 16612
rect 18748 16600 18754 16652
rect 18800 16640 18828 16671
rect 19610 16668 19616 16720
rect 19668 16708 19674 16720
rect 19668 16680 20024 16708
rect 19668 16668 19674 16680
rect 19996 16649 20024 16680
rect 19429 16643 19487 16649
rect 18800 16612 19380 16640
rect 16316 16544 17448 16572
rect 17865 16575 17923 16581
rect 16117 16535 16175 16541
rect 17865 16541 17877 16575
rect 17911 16541 17923 16575
rect 18325 16575 18383 16581
rect 18325 16572 18337 16575
rect 17865 16535 17923 16541
rect 18064 16544 18337 16572
rect 16132 16504 16160 16535
rect 16574 16504 16580 16516
rect 16132 16476 16580 16504
rect 16574 16464 16580 16476
rect 16632 16513 16638 16516
rect 16632 16507 16696 16513
rect 16632 16473 16650 16507
rect 16684 16504 16696 16507
rect 18064 16504 18092 16544
rect 18325 16541 18337 16544
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 18414 16532 18420 16584
rect 18472 16532 18478 16584
rect 18601 16575 18659 16581
rect 18601 16541 18613 16575
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 18616 16504 18644 16535
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 19352 16581 19380 16612
rect 19429 16609 19441 16643
rect 19475 16640 19487 16643
rect 19797 16643 19855 16649
rect 19797 16640 19809 16643
rect 19475 16612 19809 16640
rect 19475 16609 19487 16612
rect 19429 16603 19487 16609
rect 19797 16609 19809 16612
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 19981 16643 20039 16649
rect 19981 16609 19993 16643
rect 20027 16609 20039 16643
rect 19981 16603 20039 16609
rect 20438 16600 20444 16652
rect 20496 16600 20502 16652
rect 18969 16575 19027 16581
rect 18969 16572 18981 16575
rect 18840 16544 18981 16572
rect 18840 16532 18846 16544
rect 18969 16541 18981 16544
rect 19015 16541 19027 16575
rect 18969 16535 19027 16541
rect 19337 16575 19395 16581
rect 19337 16541 19349 16575
rect 19383 16541 19395 16575
rect 19337 16535 19395 16541
rect 19702 16532 19708 16584
rect 19760 16532 19766 16584
rect 16684 16476 16725 16504
rect 17788 16476 18092 16504
rect 18156 16476 18644 16504
rect 19981 16507 20039 16513
rect 16684 16473 16696 16476
rect 16632 16467 16696 16473
rect 16632 16464 16638 16467
rect 17678 16436 17684 16448
rect 14384 16408 17684 16436
rect 11480 16396 11486 16408
rect 17678 16396 17684 16408
rect 17736 16396 17742 16448
rect 17788 16445 17816 16476
rect 17773 16439 17831 16445
rect 17773 16405 17785 16439
rect 17819 16405 17831 16439
rect 17773 16399 17831 16405
rect 17957 16439 18015 16445
rect 17957 16405 17969 16439
rect 18003 16436 18015 16439
rect 18046 16436 18052 16448
rect 18003 16408 18052 16436
rect 18003 16405 18015 16408
rect 17957 16399 18015 16405
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 18156 16445 18184 16476
rect 19981 16473 19993 16507
rect 20027 16504 20039 16507
rect 20165 16507 20223 16513
rect 20165 16504 20177 16507
rect 20027 16476 20177 16504
rect 20027 16473 20039 16476
rect 19981 16467 20039 16473
rect 20165 16473 20177 16476
rect 20211 16473 20223 16507
rect 20165 16467 20223 16473
rect 18141 16439 18199 16445
rect 18141 16405 18153 16439
rect 18187 16405 18199 16439
rect 18141 16399 18199 16405
rect 18506 16396 18512 16448
rect 18564 16396 18570 16448
rect 18874 16396 18880 16448
rect 18932 16436 18938 16448
rect 21082 16436 21088 16448
rect 18932 16408 21088 16436
rect 18932 16396 18938 16408
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 1104 16346 21043 16368
rect 1104 16294 5894 16346
rect 5946 16294 5958 16346
rect 6010 16294 6022 16346
rect 6074 16294 6086 16346
rect 6138 16294 6150 16346
rect 6202 16294 10839 16346
rect 10891 16294 10903 16346
rect 10955 16294 10967 16346
rect 11019 16294 11031 16346
rect 11083 16294 11095 16346
rect 11147 16294 15784 16346
rect 15836 16294 15848 16346
rect 15900 16294 15912 16346
rect 15964 16294 15976 16346
rect 16028 16294 16040 16346
rect 16092 16294 20729 16346
rect 20781 16294 20793 16346
rect 20845 16294 20857 16346
rect 20909 16294 20921 16346
rect 20973 16294 20985 16346
rect 21037 16294 21043 16346
rect 1104 16272 21043 16294
rect 1578 16192 1584 16244
rect 1636 16192 1642 16244
rect 1946 16192 1952 16244
rect 2004 16232 2010 16244
rect 2501 16235 2559 16241
rect 2501 16232 2513 16235
rect 2004 16204 2513 16232
rect 2004 16192 2010 16204
rect 2501 16201 2513 16204
rect 2547 16201 2559 16235
rect 2501 16195 2559 16201
rect 3142 16192 3148 16244
rect 3200 16232 3206 16244
rect 6089 16235 6147 16241
rect 6089 16232 6101 16235
rect 3200 16204 4108 16232
rect 3200 16192 3206 16204
rect 1489 16167 1547 16173
rect 1489 16133 1501 16167
rect 1535 16164 1547 16167
rect 1670 16164 1676 16176
rect 1535 16136 1676 16164
rect 1535 16133 1547 16136
rect 1489 16127 1547 16133
rect 1670 16124 1676 16136
rect 1728 16124 1734 16176
rect 2222 16164 2228 16176
rect 1964 16136 2228 16164
rect 1964 16108 1992 16136
rect 2222 16124 2228 16136
rect 2280 16124 2286 16176
rect 3418 16124 3424 16176
rect 3476 16124 3482 16176
rect 3143 16109 3201 16115
rect 3143 16108 3155 16109
rect 3189 16108 3201 16109
rect 1946 16056 1952 16108
rect 2004 16056 2010 16108
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16065 2099 16099
rect 2041 16059 2099 16065
rect 2056 15960 2084 16059
rect 2498 16056 2504 16108
rect 2556 16056 2562 16108
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 2774 16096 2780 16108
rect 2731 16068 2780 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 2774 16056 2780 16068
rect 2832 16056 2838 16108
rect 3142 16056 3148 16108
rect 3200 16056 3206 16108
rect 3436 16096 3464 16124
rect 3436 16068 4016 16096
rect 2516 16028 2544 16056
rect 2869 16031 2927 16037
rect 2869 16028 2881 16031
rect 2516 16000 2881 16028
rect 2869 15997 2881 16000
rect 2915 15997 2927 16031
rect 2869 15991 2927 15997
rect 2056 15932 3004 15960
rect 2130 15852 2136 15904
rect 2188 15852 2194 15904
rect 2976 15892 3004 15932
rect 3786 15892 3792 15904
rect 2976 15864 3792 15892
rect 3786 15852 3792 15864
rect 3844 15852 3850 15904
rect 3878 15852 3884 15904
rect 3936 15852 3942 15904
rect 3988 15892 4016 16068
rect 4080 16028 4108 16204
rect 4172 16204 6101 16232
rect 4172 16028 4200 16204
rect 6089 16201 6101 16204
rect 6135 16201 6147 16235
rect 6089 16195 6147 16201
rect 6454 16192 6460 16244
rect 6512 16232 6518 16244
rect 7374 16232 7380 16244
rect 6512 16204 7380 16232
rect 6512 16192 6518 16204
rect 7374 16192 7380 16204
rect 7432 16192 7438 16244
rect 7650 16192 7656 16244
rect 7708 16232 7714 16244
rect 8110 16232 8116 16244
rect 7708 16204 8116 16232
rect 7708 16192 7714 16204
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 10042 16232 10048 16244
rect 8772 16204 10048 16232
rect 4249 16099 4307 16105
rect 4249 16065 4261 16099
rect 4295 16096 4307 16099
rect 4614 16096 4620 16108
rect 4295 16068 4620 16096
rect 4295 16065 4307 16068
rect 4249 16059 4307 16065
rect 4614 16056 4620 16068
rect 4672 16056 4678 16108
rect 5258 16056 5264 16108
rect 5316 16105 5322 16108
rect 5316 16099 5344 16105
rect 5332 16065 5344 16099
rect 5316 16059 5344 16065
rect 5445 16099 5503 16105
rect 5445 16065 5457 16099
rect 5491 16065 5503 16099
rect 5445 16059 5503 16065
rect 5316 16056 5322 16059
rect 4080 16000 4200 16028
rect 4338 15988 4344 16040
rect 4396 16028 4402 16040
rect 4433 16031 4491 16037
rect 4433 16028 4445 16031
rect 4396 16000 4445 16028
rect 4396 15988 4402 16000
rect 4433 15997 4445 16000
rect 4479 15997 4491 16031
rect 5169 16031 5227 16037
rect 5169 16028 5181 16031
rect 4433 15991 4491 15997
rect 5000 16000 5181 16028
rect 4706 15920 4712 15972
rect 4764 15960 4770 15972
rect 4893 15963 4951 15969
rect 4893 15960 4905 15963
rect 4764 15932 4905 15960
rect 4764 15920 4770 15932
rect 4893 15929 4905 15932
rect 4939 15929 4951 15963
rect 4893 15923 4951 15929
rect 4522 15892 4528 15904
rect 3988 15864 4528 15892
rect 4522 15852 4528 15864
rect 4580 15852 4586 15904
rect 5000 15892 5028 16000
rect 5169 15997 5181 16000
rect 5215 15997 5227 16031
rect 5460 16028 5488 16059
rect 7466 16056 7472 16108
rect 7524 16105 7530 16108
rect 7524 16099 7552 16105
rect 7540 16065 7552 16099
rect 7524 16059 7552 16065
rect 7524 16056 7530 16059
rect 7650 16056 7656 16108
rect 7708 16056 7714 16108
rect 8772 16105 8800 16204
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 13541 16235 13599 16241
rect 13541 16201 13553 16235
rect 13587 16232 13599 16235
rect 13998 16232 14004 16244
rect 13587 16204 14004 16232
rect 13587 16201 13599 16204
rect 13541 16195 13599 16201
rect 13998 16192 14004 16204
rect 14056 16192 14062 16244
rect 14734 16232 14740 16244
rect 14108 16204 14740 16232
rect 11716 16136 13400 16164
rect 11716 16108 11744 16136
rect 8757 16099 8815 16105
rect 8757 16065 8769 16099
rect 8803 16065 8815 16099
rect 8757 16059 8815 16065
rect 9766 16056 9772 16108
rect 9824 16105 9830 16108
rect 9824 16099 9852 16105
rect 9840 16065 9852 16099
rect 9824 16059 9852 16065
rect 9824 16056 9830 16059
rect 11698 16056 11704 16108
rect 11756 16056 11762 16108
rect 12434 16056 12440 16108
rect 12492 16096 12498 16108
rect 12771 16099 12829 16105
rect 12771 16096 12783 16099
rect 12492 16068 12783 16096
rect 12492 16056 12498 16068
rect 12771 16065 12783 16068
rect 12817 16065 12829 16099
rect 12771 16059 12829 16065
rect 5994 16028 6000 16040
rect 5460 16000 6000 16028
rect 5169 15991 5227 15997
rect 5994 15988 6000 16000
rect 6052 15988 6058 16040
rect 6454 15988 6460 16040
rect 6512 15988 6518 16040
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 6641 16031 6699 16037
rect 6641 16028 6653 16031
rect 6604 16000 6653 16028
rect 6604 15988 6610 16000
rect 6641 15997 6653 16000
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 6730 15988 6736 16040
rect 6788 15988 6794 16040
rect 7190 15988 7196 16040
rect 7248 16028 7254 16040
rect 7377 16031 7435 16037
rect 7377 16028 7389 16031
rect 7248 16000 7389 16028
rect 7248 15988 7254 16000
rect 7377 15997 7389 16000
rect 7423 15997 7435 16031
rect 8941 16031 8999 16037
rect 8941 16028 8953 16031
rect 7377 15991 7435 15997
rect 8772 16000 8953 16028
rect 6748 15960 6776 15988
rect 5826 15932 6776 15960
rect 5826 15892 5854 15932
rect 7006 15920 7012 15972
rect 7064 15960 7070 15972
rect 7101 15963 7159 15969
rect 7101 15960 7113 15963
rect 7064 15932 7113 15960
rect 7064 15920 7070 15932
rect 7101 15929 7113 15932
rect 7147 15929 7159 15963
rect 7101 15923 7159 15929
rect 8772 15904 8800 16000
rect 8941 15997 8953 16000
rect 8987 15997 8999 16031
rect 9677 16031 9735 16037
rect 9677 16028 9689 16031
rect 8941 15991 8999 15997
rect 9508 16000 9689 16028
rect 9398 15920 9404 15972
rect 9456 15920 9462 15972
rect 5000 15864 5854 15892
rect 6178 15852 6184 15904
rect 6236 15892 6242 15904
rect 8297 15895 8355 15901
rect 8297 15892 8309 15895
rect 6236 15864 8309 15892
rect 6236 15852 6242 15864
rect 8297 15861 8309 15864
rect 8343 15861 8355 15895
rect 8297 15855 8355 15861
rect 8754 15852 8760 15904
rect 8812 15852 8818 15904
rect 9508 15892 9536 16000
rect 9677 15997 9689 16000
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 9953 16031 10011 16037
rect 9953 15997 9965 16031
rect 9999 16028 10011 16031
rect 10134 16028 10140 16040
rect 9999 16000 10140 16028
rect 9999 15997 10011 16000
rect 9953 15991 10011 15997
rect 10134 15988 10140 16000
rect 10192 15988 10198 16040
rect 10597 16031 10655 16037
rect 10597 16028 10609 16031
rect 10336 16000 10609 16028
rect 9858 15892 9864 15904
rect 9508 15864 9864 15892
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 10042 15852 10048 15904
rect 10100 15892 10106 15904
rect 10336 15892 10364 16000
rect 10597 15997 10609 16000
rect 10643 15997 10655 16031
rect 10597 15991 10655 15997
rect 11790 15988 11796 16040
rect 11848 16028 11854 16040
rect 12529 16031 12587 16037
rect 12529 16028 12541 16031
rect 11848 16000 12541 16028
rect 11848 15988 11854 16000
rect 12529 15997 12541 16000
rect 12575 15997 12587 16031
rect 12529 15991 12587 15997
rect 10100 15864 10364 15892
rect 12544 15892 12572 15991
rect 13372 15960 13400 16136
rect 14108 16105 14136 16204
rect 14734 16192 14740 16204
rect 14792 16192 14798 16244
rect 15194 16192 15200 16244
rect 15252 16232 15258 16244
rect 15933 16235 15991 16241
rect 15933 16232 15945 16235
rect 15252 16204 15945 16232
rect 15252 16192 15258 16204
rect 15933 16201 15945 16204
rect 15979 16201 15991 16235
rect 15933 16195 15991 16201
rect 18046 16192 18052 16244
rect 18104 16192 18110 16244
rect 18414 16192 18420 16244
rect 18472 16192 18478 16244
rect 18506 16192 18512 16244
rect 18564 16192 18570 16244
rect 19702 16192 19708 16244
rect 19760 16192 19766 16244
rect 16942 16164 16948 16176
rect 16592 16136 16948 16164
rect 14093 16099 14151 16105
rect 14093 16065 14105 16099
rect 14139 16065 14151 16099
rect 14093 16059 14151 16065
rect 15010 16056 15016 16108
rect 15068 16056 15074 16108
rect 15286 16056 15292 16108
rect 15344 16056 15350 16108
rect 14274 15988 14280 16040
rect 14332 15988 14338 16040
rect 15130 16031 15188 16037
rect 15130 16028 15142 16031
rect 14366 16000 15142 16028
rect 13372 15932 14044 15960
rect 13814 15892 13820 15904
rect 12544 15864 13820 15892
rect 10100 15852 10106 15864
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 14016 15892 14044 15932
rect 14090 15920 14096 15972
rect 14148 15960 14154 15972
rect 14366 15960 14394 16000
rect 15130 15997 15142 16000
rect 15176 15997 15188 16031
rect 15130 15991 15188 15997
rect 15654 15988 15660 16040
rect 15712 16028 15718 16040
rect 16206 16028 16212 16040
rect 15712 16000 16212 16028
rect 15712 15988 15718 16000
rect 16206 15988 16212 16000
rect 16264 15988 16270 16040
rect 16592 16028 16620 16136
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 18064 16164 18092 16192
rect 18064 16136 18368 16164
rect 16666 16056 16672 16108
rect 16724 16096 16730 16108
rect 18340 16105 18368 16136
rect 17095 16099 17153 16105
rect 17095 16096 17107 16099
rect 16724 16068 17107 16096
rect 16724 16056 16730 16068
rect 17095 16065 17107 16068
rect 17141 16065 17153 16099
rect 17095 16059 17153 16065
rect 18233 16099 18291 16105
rect 18233 16065 18245 16099
rect 18279 16065 18291 16099
rect 18233 16059 18291 16065
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16065 18383 16099
rect 18325 16059 18383 16065
rect 16853 16031 16911 16037
rect 16853 16028 16865 16031
rect 16592 16000 16865 16028
rect 16853 15997 16865 16000
rect 16899 15997 16911 16031
rect 16853 15991 16911 15997
rect 18248 16028 18276 16059
rect 18432 16028 18460 16192
rect 18524 16037 18552 16192
rect 18935 16099 18993 16105
rect 18935 16096 18947 16099
rect 18616 16068 18947 16096
rect 18248 16000 18460 16028
rect 18509 16031 18567 16037
rect 14148 15932 14394 15960
rect 14148 15920 14154 15932
rect 14734 15920 14740 15972
rect 14792 15920 14798 15972
rect 17865 15963 17923 15969
rect 17865 15929 17877 15963
rect 17911 15960 17923 15963
rect 18248 15960 18276 16000
rect 18509 15997 18521 16031
rect 18555 15997 18567 16031
rect 18509 15991 18567 15997
rect 18616 15960 18644 16068
rect 18935 16065 18947 16068
rect 18981 16065 18993 16099
rect 18935 16059 18993 16065
rect 20165 16099 20223 16105
rect 20165 16065 20177 16099
rect 20211 16065 20223 16099
rect 20165 16059 20223 16065
rect 18690 15988 18696 16040
rect 18748 15988 18754 16040
rect 17911 15932 18276 15960
rect 18340 15932 18644 15960
rect 17911 15929 17923 15932
rect 17865 15923 17923 15929
rect 16942 15892 16948 15904
rect 14016 15864 16948 15892
rect 16942 15852 16948 15864
rect 17000 15892 17006 15904
rect 18340 15892 18368 15932
rect 17000 15864 18368 15892
rect 18417 15895 18475 15901
rect 17000 15852 17006 15864
rect 18417 15861 18429 15895
rect 18463 15892 18475 15895
rect 20180 15892 20208 16059
rect 18463 15864 20208 15892
rect 18463 15861 18475 15864
rect 18417 15855 18475 15861
rect 20438 15852 20444 15904
rect 20496 15852 20502 15904
rect 1104 15802 20884 15824
rect 1104 15750 3422 15802
rect 3474 15750 3486 15802
rect 3538 15750 3550 15802
rect 3602 15750 3614 15802
rect 3666 15750 3678 15802
rect 3730 15750 8367 15802
rect 8419 15750 8431 15802
rect 8483 15750 8495 15802
rect 8547 15750 8559 15802
rect 8611 15750 8623 15802
rect 8675 15750 13312 15802
rect 13364 15750 13376 15802
rect 13428 15750 13440 15802
rect 13492 15750 13504 15802
rect 13556 15750 13568 15802
rect 13620 15750 18257 15802
rect 18309 15750 18321 15802
rect 18373 15750 18385 15802
rect 18437 15750 18449 15802
rect 18501 15750 18513 15802
rect 18565 15750 20884 15802
rect 1104 15728 20884 15750
rect 1486 15648 1492 15700
rect 1544 15648 1550 15700
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 1728 15660 3341 15688
rect 1728 15648 1734 15660
rect 3329 15657 3341 15660
rect 3375 15657 3387 15691
rect 6178 15688 6184 15700
rect 3329 15651 3387 15657
rect 4126 15660 6184 15688
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 1765 15487 1823 15493
rect 1765 15453 1777 15487
rect 1811 15453 1823 15487
rect 1765 15447 1823 15453
rect 1688 15348 1716 15447
rect 1780 15416 1808 15447
rect 2038 15444 2044 15496
rect 2096 15444 2102 15496
rect 2130 15444 2136 15496
rect 2188 15444 2194 15496
rect 2774 15444 2780 15496
rect 2832 15484 2838 15496
rect 3142 15484 3148 15496
rect 2832 15456 3148 15484
rect 2832 15444 2838 15456
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15484 4031 15487
rect 4126 15484 4154 15660
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 7101 15691 7159 15697
rect 7101 15657 7113 15691
rect 7147 15688 7159 15691
rect 7558 15688 7564 15700
rect 7147 15660 7564 15688
rect 7147 15657 7159 15660
rect 7101 15651 7159 15657
rect 7558 15648 7564 15660
rect 7616 15648 7622 15700
rect 8481 15691 8539 15697
rect 8481 15657 8493 15691
rect 8527 15688 8539 15691
rect 8527 15660 9720 15688
rect 8527 15657 8539 15660
rect 8481 15651 8539 15657
rect 4522 15580 4528 15632
rect 4580 15580 4586 15632
rect 9692 15620 9720 15660
rect 9950 15648 9956 15700
rect 10008 15688 10014 15700
rect 10045 15691 10103 15697
rect 10045 15688 10057 15691
rect 10008 15660 10057 15688
rect 10008 15648 10014 15660
rect 10045 15657 10057 15660
rect 10091 15657 10103 15691
rect 10045 15651 10103 15657
rect 10134 15648 10140 15700
rect 10192 15648 10198 15700
rect 10502 15648 10508 15700
rect 10560 15688 10566 15700
rect 11425 15691 11483 15697
rect 11425 15688 11437 15691
rect 10560 15660 11437 15688
rect 10560 15648 10566 15660
rect 11425 15657 11437 15660
rect 11471 15657 11483 15691
rect 15194 15688 15200 15700
rect 11425 15651 11483 15657
rect 14476 15660 15200 15688
rect 10152 15620 10180 15648
rect 9692 15592 10180 15620
rect 11790 15580 11796 15632
rect 11848 15580 11854 15632
rect 13906 15580 13912 15632
rect 13964 15620 13970 15632
rect 14476 15620 14504 15660
rect 15194 15648 15200 15660
rect 15252 15648 15258 15700
rect 15378 15648 15384 15700
rect 15436 15688 15442 15700
rect 17037 15691 17095 15697
rect 17037 15688 17049 15691
rect 15436 15660 17049 15688
rect 15436 15648 15442 15660
rect 17037 15657 17049 15660
rect 17083 15657 17095 15691
rect 17037 15651 17095 15657
rect 19610 15648 19616 15700
rect 19668 15648 19674 15700
rect 19702 15648 19708 15700
rect 19760 15648 19766 15700
rect 19794 15648 19800 15700
rect 19852 15648 19858 15700
rect 13964 15592 14504 15620
rect 13964 15580 13970 15592
rect 4540 15552 4568 15580
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 4540 15524 4721 15552
rect 4709 15521 4721 15524
rect 4755 15521 4767 15555
rect 4709 15515 4767 15521
rect 8938 15512 8944 15564
rect 8996 15552 9002 15564
rect 9033 15555 9091 15561
rect 9033 15552 9045 15555
rect 8996 15524 9045 15552
rect 8996 15512 9002 15524
rect 9033 15521 9045 15524
rect 9079 15521 9091 15555
rect 10134 15552 10140 15564
rect 9033 15515 9091 15521
rect 9646 15524 10140 15552
rect 4019 15456 4154 15484
rect 4249 15487 4307 15493
rect 4019 15453 4031 15456
rect 3973 15447 4031 15453
rect 4249 15453 4261 15487
rect 4295 15484 4307 15487
rect 4525 15487 4583 15493
rect 4295 15456 4476 15484
rect 4295 15453 4307 15456
rect 4249 15447 4307 15453
rect 2148 15416 2176 15444
rect 1780 15388 2176 15416
rect 3237 15419 3295 15425
rect 3237 15385 3249 15419
rect 3283 15416 3295 15419
rect 3283 15388 4384 15416
rect 3283 15385 3295 15388
rect 3237 15379 3295 15385
rect 2682 15348 2688 15360
rect 1688 15320 2688 15348
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 2777 15351 2835 15357
rect 2777 15317 2789 15351
rect 2823 15348 2835 15351
rect 2866 15348 2872 15360
rect 2823 15320 2872 15348
rect 2823 15317 2835 15320
rect 2777 15311 2835 15317
rect 2866 15308 2872 15320
rect 2924 15308 2930 15360
rect 3786 15308 3792 15360
rect 3844 15308 3850 15360
rect 3878 15308 3884 15360
rect 3936 15348 3942 15360
rect 4356 15357 4384 15388
rect 4065 15351 4123 15357
rect 4065 15348 4077 15351
rect 3936 15320 4077 15348
rect 3936 15308 3942 15320
rect 4065 15317 4077 15320
rect 4111 15317 4123 15351
rect 4065 15311 4123 15317
rect 4341 15351 4399 15357
rect 4341 15317 4353 15351
rect 4387 15317 4399 15351
rect 4448 15348 4476 15456
rect 4525 15453 4537 15487
rect 4571 15453 4583 15487
rect 4525 15447 4583 15453
rect 4983 15487 5041 15493
rect 4983 15453 4995 15487
rect 5029 15484 5041 15487
rect 5442 15484 5448 15496
rect 5029 15456 5448 15484
rect 5029 15453 5041 15456
rect 4983 15447 5041 15453
rect 4540 15416 4568 15447
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 5810 15444 5816 15496
rect 5868 15484 5874 15496
rect 6089 15487 6147 15493
rect 6089 15484 6101 15487
rect 5868 15456 6101 15484
rect 5868 15444 5874 15456
rect 6089 15453 6101 15456
rect 6135 15453 6147 15487
rect 6089 15447 6147 15453
rect 6270 15444 6276 15496
rect 6328 15484 6334 15496
rect 6363 15487 6421 15493
rect 6363 15484 6375 15487
rect 6328 15456 6375 15484
rect 6328 15444 6334 15456
rect 6363 15453 6375 15456
rect 6409 15453 6421 15487
rect 6363 15447 6421 15453
rect 7466 15444 7472 15496
rect 7524 15444 7530 15496
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 8662 15416 8668 15428
rect 4540 15388 8668 15416
rect 8662 15376 8668 15388
rect 8720 15376 8726 15428
rect 9048 15416 9076 15515
rect 9306 15484 9312 15496
rect 9267 15456 9312 15484
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 9646 15484 9674 15524
rect 10134 15512 10140 15524
rect 10192 15552 10198 15564
rect 10413 15555 10471 15561
rect 10413 15552 10425 15555
rect 10192 15524 10425 15552
rect 10192 15512 10198 15524
rect 10413 15521 10425 15524
rect 10459 15521 10471 15555
rect 11808 15552 11836 15580
rect 10413 15515 10471 15521
rect 11454 15524 11836 15552
rect 10687 15487 10745 15493
rect 9416 15456 9674 15484
rect 10336 15484 10481 15486
rect 10336 15458 10548 15484
rect 9416 15416 9444 15456
rect 9048 15388 9444 15416
rect 9582 15376 9588 15428
rect 9640 15416 9646 15428
rect 10336 15416 10364 15458
rect 10453 15456 10548 15458
rect 9640 15388 10364 15416
rect 10520 15416 10548 15456
rect 10687 15453 10699 15487
rect 10733 15484 10745 15487
rect 11454 15484 11482 15524
rect 13170 15512 13176 15564
rect 13228 15512 13234 15564
rect 14277 15555 14335 15561
rect 14277 15552 14289 15555
rect 13924 15524 14289 15552
rect 10733 15456 11482 15484
rect 10733 15453 10745 15456
rect 10687 15447 10745 15453
rect 11514 15444 11520 15496
rect 11572 15484 11578 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11572 15456 11805 15484
rect 11572 15444 11578 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 11793 15447 11851 15453
rect 12067 15487 12125 15493
rect 12067 15453 12079 15487
rect 12113 15484 12125 15487
rect 12434 15484 12440 15496
rect 12113 15456 12440 15484
rect 12113 15453 12125 15456
rect 12067 15447 12125 15453
rect 12434 15444 12440 15456
rect 12492 15444 12498 15496
rect 13188 15416 13216 15512
rect 13924 15496 13952 15524
rect 14277 15521 14289 15524
rect 14323 15521 14335 15555
rect 14277 15515 14335 15521
rect 14476 15496 14504 15592
rect 14550 15580 14556 15632
rect 14608 15620 14614 15632
rect 14737 15623 14795 15629
rect 14737 15620 14749 15623
rect 14608 15592 14749 15620
rect 14608 15580 14614 15592
rect 14737 15589 14749 15592
rect 14783 15589 14795 15623
rect 14737 15583 14795 15589
rect 18877 15623 18935 15629
rect 18877 15589 18889 15623
rect 18923 15620 18935 15623
rect 19518 15620 19524 15632
rect 18923 15592 19524 15620
rect 18923 15589 18935 15592
rect 18877 15583 18935 15589
rect 19518 15580 19524 15592
rect 19576 15580 19582 15632
rect 15010 15512 15016 15564
rect 15068 15512 15074 15564
rect 15194 15561 15200 15564
rect 15151 15555 15200 15561
rect 15151 15521 15163 15555
rect 15197 15521 15200 15555
rect 15151 15515 15200 15521
rect 15194 15512 15200 15515
rect 15252 15512 15258 15564
rect 15654 15512 15660 15564
rect 15712 15552 15718 15564
rect 15712 15524 16068 15552
rect 15712 15512 15718 15524
rect 13906 15444 13912 15496
rect 13964 15444 13970 15496
rect 14090 15444 14096 15496
rect 14148 15444 14154 15496
rect 14458 15444 14464 15496
rect 14516 15444 14522 15496
rect 15286 15444 15292 15496
rect 15344 15444 15350 15496
rect 16040 15493 16068 15524
rect 17310 15512 17316 15564
rect 17368 15552 17374 15564
rect 19334 15552 19340 15564
rect 17368 15524 19340 15552
rect 17368 15512 17374 15524
rect 19334 15512 19340 15524
rect 19392 15512 19398 15564
rect 19720 15552 19748 15648
rect 19536 15524 19748 15552
rect 19812 15552 19840 15648
rect 19812 15524 20024 15552
rect 16025 15487 16083 15493
rect 16025 15453 16037 15487
rect 16071 15453 16083 15487
rect 16025 15447 16083 15453
rect 14108 15416 14136 15444
rect 10520 15388 12940 15416
rect 13188 15388 14136 15416
rect 15933 15419 15991 15425
rect 9640 15376 9646 15388
rect 5442 15348 5448 15360
rect 4448 15320 5448 15348
rect 4341 15311 4399 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 5721 15351 5779 15357
rect 5721 15317 5733 15351
rect 5767 15348 5779 15351
rect 6638 15348 6644 15360
rect 5767 15320 6644 15348
rect 5767 15317 5779 15320
rect 5721 15311 5779 15317
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 7926 15348 7932 15360
rect 7616 15320 7932 15348
rect 7616 15308 7622 15320
rect 7926 15308 7932 15320
rect 7984 15308 7990 15360
rect 11238 15308 11244 15360
rect 11296 15348 11302 15360
rect 12805 15351 12863 15357
rect 12805 15348 12817 15351
rect 11296 15320 12817 15348
rect 11296 15308 11302 15320
rect 12805 15317 12817 15320
rect 12851 15317 12863 15351
rect 12912 15348 12940 15388
rect 15933 15385 15945 15419
rect 15979 15385 15991 15419
rect 16040 15416 16068 15447
rect 16206 15444 16212 15496
rect 16264 15484 16270 15496
rect 16299 15487 16357 15493
rect 16299 15484 16311 15487
rect 16264 15456 16311 15484
rect 16264 15444 16270 15456
rect 16299 15453 16311 15456
rect 16345 15453 16357 15487
rect 16299 15447 16357 15453
rect 17402 15444 17408 15496
rect 17460 15444 17466 15496
rect 18509 15487 18567 15493
rect 18509 15453 18521 15487
rect 18555 15453 18567 15487
rect 18509 15447 18567 15453
rect 16574 15416 16580 15428
rect 16040 15388 16580 15416
rect 15933 15379 15991 15385
rect 15948 15348 15976 15379
rect 16574 15376 16580 15388
rect 16632 15416 16638 15428
rect 17420 15416 17448 15444
rect 16632 15388 17448 15416
rect 18524 15416 18552 15447
rect 18690 15444 18696 15496
rect 18748 15444 18754 15496
rect 19058 15444 19064 15496
rect 19116 15444 19122 15496
rect 19242 15444 19248 15496
rect 19300 15444 19306 15496
rect 19536 15493 19564 15524
rect 19996 15493 20024 15524
rect 19521 15487 19579 15493
rect 19521 15453 19533 15487
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15484 19763 15487
rect 19981 15487 20039 15493
rect 19751 15456 19840 15484
rect 19751 15453 19763 15456
rect 19705 15447 19763 15453
rect 19150 15416 19156 15428
rect 18524 15388 19156 15416
rect 16632 15376 16638 15388
rect 19150 15376 19156 15388
rect 19208 15376 19214 15428
rect 12912 15320 15976 15348
rect 12805 15311 12863 15317
rect 16942 15308 16948 15360
rect 17000 15348 17006 15360
rect 18598 15348 18604 15360
rect 17000 15320 18604 15348
rect 17000 15308 17006 15320
rect 18598 15308 18604 15320
rect 18656 15308 18662 15360
rect 18693 15351 18751 15357
rect 18693 15317 18705 15351
rect 18739 15348 18751 15351
rect 18782 15348 18788 15360
rect 18739 15320 18788 15348
rect 18739 15317 18751 15320
rect 18693 15311 18751 15317
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 19334 15308 19340 15360
rect 19392 15308 19398 15360
rect 19812 15357 19840 15456
rect 19981 15453 19993 15487
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20165 15419 20223 15425
rect 20165 15385 20177 15419
rect 20211 15385 20223 15419
rect 20165 15379 20223 15385
rect 20533 15419 20591 15425
rect 20533 15385 20545 15419
rect 20579 15416 20591 15419
rect 21266 15416 21272 15428
rect 20579 15388 21272 15416
rect 20579 15385 20591 15388
rect 20533 15379 20591 15385
rect 19797 15351 19855 15357
rect 19797 15317 19809 15351
rect 19843 15317 19855 15351
rect 19797 15311 19855 15317
rect 19978 15308 19984 15360
rect 20036 15348 20042 15360
rect 20180 15348 20208 15379
rect 21266 15376 21272 15388
rect 21324 15376 21330 15428
rect 20036 15320 20208 15348
rect 20036 15308 20042 15320
rect 1104 15258 21043 15280
rect 1104 15206 5894 15258
rect 5946 15206 5958 15258
rect 6010 15206 6022 15258
rect 6074 15206 6086 15258
rect 6138 15206 6150 15258
rect 6202 15206 10839 15258
rect 10891 15206 10903 15258
rect 10955 15206 10967 15258
rect 11019 15206 11031 15258
rect 11083 15206 11095 15258
rect 11147 15206 15784 15258
rect 15836 15206 15848 15258
rect 15900 15206 15912 15258
rect 15964 15206 15976 15258
rect 16028 15206 16040 15258
rect 16092 15206 20729 15258
rect 20781 15206 20793 15258
rect 20845 15206 20857 15258
rect 20909 15206 20921 15258
rect 20973 15206 20985 15258
rect 21037 15206 21043 15258
rect 1104 15184 21043 15206
rect 842 15104 848 15156
rect 900 15144 906 15156
rect 1765 15147 1823 15153
rect 1765 15144 1777 15147
rect 900 15116 1777 15144
rect 900 15104 906 15116
rect 1765 15113 1777 15116
rect 1811 15113 1823 15147
rect 1765 15107 1823 15113
rect 1946 15104 1952 15156
rect 2004 15104 2010 15156
rect 2222 15104 2228 15156
rect 2280 15144 2286 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 2280 15116 8217 15144
rect 2280 15104 2286 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 11330 15144 11336 15156
rect 8205 15107 8263 15113
rect 8922 15116 11336 15144
rect 1670 14968 1676 15020
rect 1728 14968 1734 15020
rect 1964 15008 1992 15104
rect 2682 15076 2688 15088
rect 2422 15048 2688 15076
rect 2422 15047 2450 15048
rect 2391 15041 2450 15047
rect 2038 15008 2044 15020
rect 1964 14980 2044 15008
rect 2038 14968 2044 14980
rect 2096 15008 2102 15020
rect 2133 15011 2191 15017
rect 2133 15008 2145 15011
rect 2096 14980 2145 15008
rect 2096 14968 2102 14980
rect 2133 14977 2145 14980
rect 2179 14977 2191 15011
rect 2391 15007 2403 15041
rect 2437 15010 2450 15041
rect 2682 15036 2688 15048
rect 2740 15036 2746 15088
rect 2958 15036 2964 15088
rect 3016 15076 3022 15088
rect 3878 15076 3884 15088
rect 3016 15048 3884 15076
rect 3016 15036 3022 15048
rect 3878 15036 3884 15048
rect 3936 15036 3942 15088
rect 4062 15036 4068 15088
rect 4120 15076 4126 15088
rect 4120 15036 4154 15076
rect 4246 15036 4252 15088
rect 4304 15076 4310 15088
rect 4304 15048 5120 15076
rect 4304 15036 4310 15048
rect 3787 15011 3845 15017
rect 2437 15007 2449 15010
rect 2391 15001 2449 15007
rect 2133 14971 2191 14977
rect 3787 14977 3799 15011
rect 3833 15008 3845 15011
rect 4126 15008 4154 15036
rect 5092 15020 5120 15048
rect 3833 14980 4292 15008
rect 3833 14977 3845 14980
rect 3787 14971 3845 14977
rect 4264 14952 4292 14980
rect 4522 14968 4528 15020
rect 4580 15008 4586 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4580 14980 4905 15008
rect 4580 14968 4586 14980
rect 4893 14977 4905 14980
rect 4939 14977 4951 15011
rect 4893 14971 4951 14977
rect 5074 14968 5080 15020
rect 5132 15008 5138 15020
rect 5167 15011 5225 15017
rect 5167 15008 5179 15011
rect 5132 14980 5179 15008
rect 5132 14968 5138 14980
rect 5167 14977 5179 14980
rect 5213 14977 5225 15011
rect 5167 14971 5225 14977
rect 7282 14968 7288 15020
rect 7340 14968 7346 15020
rect 8294 14968 8300 15020
rect 8352 15008 8358 15020
rect 8922 15017 8950 15116
rect 11330 15104 11336 15116
rect 11388 15104 11394 15156
rect 11698 15104 11704 15156
rect 11756 15144 11762 15156
rect 12066 15144 12072 15156
rect 11756 15116 12072 15144
rect 11756 15104 11762 15116
rect 12066 15104 12072 15116
rect 12124 15104 12130 15156
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 12618 15144 12624 15156
rect 12308 15116 12624 15144
rect 12308 15104 12314 15116
rect 12618 15104 12624 15116
rect 12676 15104 12682 15156
rect 14734 15104 14740 15156
rect 14792 15144 14798 15156
rect 15013 15147 15071 15153
rect 15013 15144 15025 15147
rect 14792 15116 15025 15144
rect 14792 15104 14798 15116
rect 15013 15113 15025 15116
rect 15059 15113 15071 15147
rect 15013 15107 15071 15113
rect 16114 15104 16120 15156
rect 16172 15104 16178 15156
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 16482 15144 16488 15156
rect 16439 15116 16488 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 16482 15104 16488 15116
rect 16540 15104 16546 15156
rect 16574 15104 16580 15156
rect 16632 15144 16638 15156
rect 20530 15144 20536 15156
rect 16632 15116 20536 15144
rect 16632 15104 16638 15116
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 10962 15076 10968 15088
rect 10060 15048 10968 15076
rect 10060 15017 10088 15048
rect 10962 15036 10968 15048
rect 11020 15036 11026 15088
rect 11054 15036 11060 15088
rect 11112 15076 11118 15088
rect 11514 15076 11520 15088
rect 11112 15048 11520 15076
rect 11112 15036 11118 15048
rect 11514 15036 11520 15048
rect 11572 15036 11578 15088
rect 13814 15036 13820 15088
rect 13872 15076 13878 15088
rect 15654 15076 15660 15088
rect 13872 15048 15660 15076
rect 13872 15036 13878 15048
rect 14016 15020 14044 15048
rect 15654 15036 15660 15048
rect 15712 15036 15718 15088
rect 16132 15076 16160 15104
rect 16914 15079 16972 15085
rect 16914 15076 16926 15079
rect 16132 15048 16926 15076
rect 8907 15011 8965 15017
rect 8907 15008 8919 15011
rect 8352 14980 8919 15008
rect 8352 14968 8358 14980
rect 8907 14977 8919 14980
rect 8953 14977 8965 15011
rect 8907 14971 8965 14977
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 10319 15011 10377 15017
rect 10319 14977 10331 15011
rect 10365 15008 10377 15011
rect 11790 15008 11796 15020
rect 10365 14980 11796 15008
rect 10365 14977 10377 14980
rect 10319 14971 10377 14977
rect 11790 14968 11796 14980
rect 11848 15008 11854 15020
rect 11974 15008 11980 15020
rect 11848 14980 11980 15008
rect 11848 14968 11854 14980
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12069 15011 12127 15017
rect 12069 14977 12081 15011
rect 12115 15008 12127 15011
rect 12158 15008 12164 15020
rect 12115 14980 12164 15008
rect 12115 14977 12127 14980
rect 12069 14971 12127 14977
rect 12158 14968 12164 14980
rect 12216 14968 12222 15020
rect 12986 14968 12992 15020
rect 13044 14968 13050 15020
rect 13998 14968 14004 15020
rect 14056 14968 14062 15020
rect 16132 15017 16160 15048
rect 16914 15045 16926 15048
rect 16960 15045 16972 15079
rect 16914 15039 16972 15045
rect 17678 15036 17684 15088
rect 17736 15076 17742 15088
rect 17736 15048 18368 15076
rect 17736 15036 17742 15048
rect 14275 15011 14333 15017
rect 14275 14977 14287 15011
rect 14321 15008 14333 15011
rect 16117 15011 16175 15017
rect 14321 14980 14872 15008
rect 14321 14977 14333 14980
rect 14275 14971 14333 14977
rect 2958 14900 2964 14952
rect 3016 14940 3022 14952
rect 3513 14943 3571 14949
rect 3513 14940 3525 14943
rect 3016 14912 3525 14940
rect 3016 14900 3022 14912
rect 3513 14909 3525 14912
rect 3559 14909 3571 14943
rect 3513 14903 3571 14909
rect 474 14764 480 14816
rect 532 14804 538 14816
rect 1118 14804 1124 14816
rect 532 14776 1124 14804
rect 532 14764 538 14776
rect 1118 14764 1124 14776
rect 1176 14764 1182 14816
rect 3142 14764 3148 14816
rect 3200 14764 3206 14816
rect 3528 14804 3556 14903
rect 4246 14900 4252 14952
rect 4304 14900 4310 14952
rect 4540 14940 4568 14968
rect 4356 14912 4568 14940
rect 4356 14804 4384 14912
rect 4706 14900 4712 14952
rect 4764 14900 4770 14952
rect 6365 14943 6423 14949
rect 6365 14909 6377 14943
rect 6411 14909 6423 14943
rect 6365 14903 6423 14909
rect 4525 14875 4583 14881
rect 4525 14841 4537 14875
rect 4571 14872 4583 14875
rect 4724 14872 4752 14900
rect 4571 14844 4752 14872
rect 6380 14872 6408 14903
rect 6546 14900 6552 14952
rect 6604 14900 6610 14952
rect 6638 14900 6644 14952
rect 6696 14940 6702 14952
rect 7009 14943 7067 14949
rect 7009 14940 7021 14943
rect 6696 14912 7021 14940
rect 6696 14900 6702 14912
rect 7009 14909 7021 14912
rect 7055 14909 7067 14943
rect 7009 14903 7067 14909
rect 7374 14900 7380 14952
rect 7432 14949 7438 14952
rect 7432 14943 7460 14949
rect 7448 14909 7460 14943
rect 7432 14903 7460 14909
rect 7561 14943 7619 14949
rect 7561 14909 7573 14943
rect 7607 14940 7619 14943
rect 8665 14943 8723 14949
rect 7607 14912 7972 14940
rect 7607 14909 7619 14912
rect 7561 14903 7619 14909
rect 7432 14900 7438 14903
rect 6454 14872 6460 14884
rect 6380 14844 6460 14872
rect 4571 14841 4583 14844
rect 4525 14835 4583 14841
rect 6454 14832 6460 14844
rect 6512 14872 6518 14884
rect 6914 14872 6920 14884
rect 6512 14844 6920 14872
rect 6512 14832 6518 14844
rect 6914 14832 6920 14844
rect 6972 14832 6978 14884
rect 3528 14776 4384 14804
rect 5905 14807 5963 14813
rect 5905 14773 5917 14807
rect 5951 14804 5963 14807
rect 7944 14804 7972 14912
rect 8665 14909 8677 14943
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 8570 14832 8576 14884
rect 8628 14872 8634 14884
rect 8680 14872 8708 14903
rect 10962 14900 10968 14952
rect 11020 14940 11026 14952
rect 11606 14940 11612 14952
rect 11020 14912 11612 14940
rect 11020 14900 11026 14912
rect 11606 14900 11612 14912
rect 11664 14900 11670 14952
rect 12253 14943 12311 14949
rect 11900 14912 12204 14940
rect 9858 14872 9864 14884
rect 8628 14844 8708 14872
rect 9600 14844 9864 14872
rect 8628 14832 8634 14844
rect 5951 14776 7972 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 9122 14764 9128 14816
rect 9180 14804 9186 14816
rect 9600 14804 9628 14844
rect 9858 14832 9864 14844
rect 9916 14832 9922 14884
rect 11057 14875 11115 14881
rect 11057 14841 11069 14875
rect 11103 14872 11115 14875
rect 11900 14872 11928 14912
rect 11103 14844 11928 14872
rect 12176 14872 12204 14912
rect 12253 14909 12265 14943
rect 12299 14940 12311 14943
rect 12434 14940 12440 14952
rect 12299 14912 12440 14940
rect 12299 14909 12311 14912
rect 12253 14903 12311 14909
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 12618 14900 12624 14952
rect 12676 14940 12682 14952
rect 13106 14943 13164 14949
rect 13106 14940 13118 14943
rect 12676 14912 13118 14940
rect 12676 14900 12682 14912
rect 13106 14909 13118 14912
rect 13152 14909 13164 14943
rect 13106 14903 13164 14909
rect 13262 14900 13268 14952
rect 13320 14900 13326 14952
rect 13630 14900 13636 14952
rect 13688 14940 13694 14952
rect 13814 14940 13820 14952
rect 13688 14912 13820 14940
rect 13688 14900 13694 14912
rect 13814 14900 13820 14912
rect 13872 14900 13878 14952
rect 12713 14875 12771 14881
rect 12713 14872 12725 14875
rect 12176 14844 12725 14872
rect 11103 14841 11115 14844
rect 11057 14835 11115 14841
rect 12713 14841 12725 14844
rect 12759 14841 12771 14875
rect 12713 14835 12771 14841
rect 14844 14816 14872 14980
rect 16117 14977 16129 15011
rect 16163 14977 16175 15011
rect 16117 14971 16175 14977
rect 16301 15011 16359 15017
rect 16301 14977 16313 15011
rect 16347 14977 16359 15011
rect 16301 14971 16359 14977
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 17494 15008 17500 15020
rect 16715 14980 17500 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 16316 14940 16344 14971
rect 17494 14968 17500 14980
rect 17552 15008 17558 15020
rect 17552 14980 17998 15008
rect 17552 14968 17558 14980
rect 16132 14912 16344 14940
rect 17970 14940 17998 14980
rect 18138 14968 18144 15020
rect 18196 14968 18202 15020
rect 18340 15017 18368 15048
rect 19426 15036 19432 15088
rect 19484 15076 19490 15088
rect 20165 15079 20223 15085
rect 20165 15076 20177 15079
rect 19484 15048 20177 15076
rect 19484 15036 19490 15048
rect 20165 15045 20177 15048
rect 20211 15045 20223 15079
rect 20165 15039 20223 15045
rect 18325 15011 18383 15017
rect 18325 14977 18337 15011
rect 18371 14977 18383 15011
rect 18325 14971 18383 14977
rect 18506 14968 18512 15020
rect 18564 15008 18570 15020
rect 18690 15017 18696 15020
rect 18673 15011 18696 15017
rect 18673 15008 18685 15011
rect 18564 14980 18685 15008
rect 18564 14968 18570 14980
rect 18673 14977 18685 14980
rect 18673 14971 18696 14977
rect 18690 14968 18696 14971
rect 18748 14968 18754 15020
rect 18417 14943 18475 14949
rect 18417 14940 18429 14943
rect 17970 14912 18429 14940
rect 16132 14816 16160 14912
rect 18417 14909 18429 14912
rect 18463 14909 18475 14943
rect 18417 14903 18475 14909
rect 20070 14872 20076 14884
rect 19628 14844 20076 14872
rect 9180 14776 9628 14804
rect 9677 14807 9735 14813
rect 9180 14764 9186 14776
rect 9677 14773 9689 14807
rect 9723 14804 9735 14807
rect 11606 14804 11612 14816
rect 9723 14776 11612 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 11606 14764 11612 14776
rect 11664 14764 11670 14816
rect 11698 14764 11704 14816
rect 11756 14804 11762 14816
rect 13909 14807 13967 14813
rect 13909 14804 13921 14807
rect 11756 14776 13921 14804
rect 11756 14764 11762 14776
rect 13909 14773 13921 14776
rect 13955 14773 13967 14807
rect 13909 14767 13967 14773
rect 14826 14764 14832 14816
rect 14884 14764 14890 14816
rect 15194 14764 15200 14816
rect 15252 14804 15258 14816
rect 15654 14804 15660 14816
rect 15252 14776 15660 14804
rect 15252 14764 15258 14776
rect 15654 14764 15660 14776
rect 15712 14764 15718 14816
rect 15930 14764 15936 14816
rect 15988 14764 15994 14816
rect 16114 14764 16120 14816
rect 16172 14764 16178 14816
rect 18046 14764 18052 14816
rect 18104 14764 18110 14816
rect 18233 14807 18291 14813
rect 18233 14773 18245 14807
rect 18279 14804 18291 14807
rect 18598 14804 18604 14816
rect 18279 14776 18604 14804
rect 18279 14773 18291 14776
rect 18233 14767 18291 14773
rect 18598 14764 18604 14776
rect 18656 14764 18662 14816
rect 19058 14764 19064 14816
rect 19116 14804 19122 14816
rect 19628 14804 19656 14844
rect 20070 14832 20076 14844
rect 20128 14832 20134 14884
rect 19116 14776 19656 14804
rect 19116 14764 19122 14776
rect 19702 14764 19708 14816
rect 19760 14804 19766 14816
rect 19797 14807 19855 14813
rect 19797 14804 19809 14807
rect 19760 14776 19809 14804
rect 19760 14764 19766 14776
rect 19797 14773 19809 14776
rect 19843 14773 19855 14807
rect 19797 14767 19855 14773
rect 20438 14764 20444 14816
rect 20496 14764 20502 14816
rect 1104 14714 20884 14736
rect 1104 14662 3422 14714
rect 3474 14662 3486 14714
rect 3538 14662 3550 14714
rect 3602 14662 3614 14714
rect 3666 14662 3678 14714
rect 3730 14662 8367 14714
rect 8419 14662 8431 14714
rect 8483 14662 8495 14714
rect 8547 14662 8559 14714
rect 8611 14662 8623 14714
rect 8675 14662 13312 14714
rect 13364 14662 13376 14714
rect 13428 14662 13440 14714
rect 13492 14662 13504 14714
rect 13556 14662 13568 14714
rect 13620 14662 18257 14714
rect 18309 14662 18321 14714
rect 18373 14662 18385 14714
rect 18437 14662 18449 14714
rect 18501 14662 18513 14714
rect 18565 14662 20884 14714
rect 1104 14640 20884 14662
rect 658 14560 664 14612
rect 716 14600 722 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 716 14572 1593 14600
rect 716 14560 722 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 1581 14563 1639 14569
rect 3329 14603 3387 14609
rect 3329 14569 3341 14603
rect 3375 14600 3387 14603
rect 3375 14572 5396 14600
rect 3375 14569 3387 14572
rect 3329 14563 3387 14569
rect 3142 14492 3148 14544
rect 3200 14532 3206 14544
rect 4433 14535 4491 14541
rect 4433 14532 4445 14535
rect 3200 14504 4445 14532
rect 3200 14492 3206 14504
rect 4433 14501 4445 14504
rect 4479 14501 4491 14535
rect 4433 14495 4491 14501
rect 658 14424 664 14476
rect 716 14464 722 14476
rect 1302 14464 1308 14476
rect 716 14436 1308 14464
rect 716 14424 722 14436
rect 1302 14424 1308 14436
rect 1360 14424 1366 14476
rect 2038 14424 2044 14476
rect 2096 14464 2102 14476
rect 2317 14467 2375 14473
rect 2317 14464 2329 14467
rect 2096 14436 2329 14464
rect 2096 14424 2102 14436
rect 2317 14433 2329 14436
rect 2363 14433 2375 14467
rect 2317 14427 2375 14433
rect 3694 14424 3700 14476
rect 3752 14464 3758 14476
rect 4062 14464 4068 14476
rect 3752 14436 4068 14464
rect 3752 14424 3758 14436
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 4706 14424 4712 14476
rect 4764 14424 4770 14476
rect 4798 14424 4804 14476
rect 4856 14473 4862 14476
rect 4856 14467 4884 14473
rect 4872 14433 4884 14467
rect 5368 14464 5396 14572
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 11698 14600 11704 14612
rect 5500 14572 11704 14600
rect 5500 14560 5506 14572
rect 11698 14560 11704 14572
rect 11756 14560 11762 14612
rect 13081 14603 13139 14609
rect 13081 14569 13093 14603
rect 13127 14600 13139 14603
rect 13630 14600 13636 14612
rect 13127 14572 13636 14600
rect 13127 14569 13139 14572
rect 13081 14563 13139 14569
rect 13630 14560 13636 14572
rect 13688 14560 13694 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14976 14572 15117 14600
rect 14976 14560 14982 14572
rect 15105 14569 15117 14572
rect 15151 14569 15163 14603
rect 15105 14563 15163 14569
rect 15930 14560 15936 14612
rect 15988 14600 15994 14612
rect 15988 14572 17816 14600
rect 15988 14560 15994 14572
rect 8481 14535 8539 14541
rect 8481 14501 8493 14535
rect 8527 14532 8539 14535
rect 9398 14532 9404 14544
rect 8527 14504 9404 14532
rect 8527 14501 8539 14504
rect 8481 14495 8539 14501
rect 9398 14492 9404 14504
rect 9456 14492 9462 14544
rect 9858 14492 9864 14544
rect 9916 14532 9922 14544
rect 9916 14504 10088 14532
rect 9916 14492 9922 14504
rect 9953 14467 10011 14473
rect 9953 14464 9965 14467
rect 4856 14427 4884 14433
rect 5000 14436 5396 14464
rect 8588 14436 9965 14464
rect 4856 14424 4862 14427
rect 2222 14356 2228 14408
rect 2280 14356 2286 14408
rect 2590 14396 2596 14408
rect 2551 14368 2596 14396
rect 2590 14356 2596 14368
rect 2648 14396 2654 14408
rect 3142 14396 3148 14408
rect 2648 14368 3148 14396
rect 2648 14356 2654 14368
rect 3142 14356 3148 14368
rect 3200 14356 3206 14408
rect 5000 14405 5028 14436
rect 3789 14399 3847 14405
rect 3789 14365 3801 14399
rect 3835 14365 3847 14399
rect 3789 14359 3847 14365
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14365 4031 14399
rect 3973 14359 4031 14365
rect 4985 14399 5043 14405
rect 4985 14365 4997 14399
rect 5031 14365 5043 14399
rect 4985 14359 5043 14365
rect 1489 14331 1547 14337
rect 1489 14297 1501 14331
rect 1535 14328 1547 14331
rect 3804 14328 3832 14359
rect 1535 14300 2084 14328
rect 1535 14297 1547 14300
rect 1489 14291 1547 14297
rect 2056 14269 2084 14300
rect 2240 14300 3832 14328
rect 2240 14272 2268 14300
rect 2041 14263 2099 14269
rect 2041 14229 2053 14263
rect 2087 14229 2099 14263
rect 2041 14223 2099 14229
rect 2222 14220 2228 14272
rect 2280 14220 2286 14272
rect 2498 14220 2504 14272
rect 2556 14260 2562 14272
rect 3988 14260 4016 14359
rect 5810 14356 5816 14408
rect 5868 14396 5874 14408
rect 6089 14399 6147 14405
rect 6089 14396 6101 14399
rect 5868 14368 6101 14396
rect 5868 14356 5874 14368
rect 6089 14365 6101 14368
rect 6135 14365 6147 14399
rect 6331 14399 6389 14405
rect 6331 14396 6343 14399
rect 6089 14359 6147 14365
rect 6196 14368 6343 14396
rect 6196 14340 6224 14368
rect 6331 14365 6343 14368
rect 6377 14396 6389 14399
rect 6914 14396 6920 14408
rect 6377 14368 6920 14396
rect 6377 14365 6389 14368
rect 6331 14359 6389 14365
rect 6914 14356 6920 14368
rect 6972 14356 6978 14408
rect 7190 14396 7196 14408
rect 7006 14368 7196 14396
rect 6178 14288 6184 14340
rect 6236 14288 6242 14340
rect 4338 14260 4344 14272
rect 2556 14232 4344 14260
rect 2556 14220 2562 14232
rect 4338 14220 4344 14232
rect 4396 14220 4402 14272
rect 4522 14220 4528 14272
rect 4580 14260 4586 14272
rect 5629 14263 5687 14269
rect 5629 14260 5641 14263
rect 4580 14232 5641 14260
rect 4580 14220 4586 14232
rect 5629 14229 5641 14232
rect 5675 14229 5687 14263
rect 5629 14223 5687 14229
rect 6270 14220 6276 14272
rect 6328 14260 6334 14272
rect 7006 14260 7034 14368
rect 7190 14356 7196 14368
rect 7248 14356 7254 14408
rect 7282 14356 7288 14408
rect 7340 14396 7346 14408
rect 7466 14396 7472 14408
rect 7340 14368 7472 14396
rect 7340 14356 7346 14368
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 7742 14356 7748 14408
rect 7800 14356 7806 14408
rect 8588 14328 8616 14436
rect 9953 14433 9965 14436
rect 9999 14433 10011 14467
rect 10060 14464 10088 14504
rect 11612 14476 11664 14482
rect 10229 14467 10287 14473
rect 10229 14464 10241 14467
rect 10060 14436 10241 14464
rect 9953 14427 10011 14433
rect 10229 14433 10241 14436
rect 10275 14433 10287 14467
rect 10229 14427 10287 14433
rect 10318 14424 10324 14476
rect 10376 14473 10382 14476
rect 10376 14467 10404 14473
rect 10392 14433 10404 14467
rect 10376 14427 10404 14433
rect 10376 14424 10382 14427
rect 13998 14424 14004 14476
rect 14056 14464 14062 14476
rect 14093 14467 14151 14473
rect 14093 14464 14105 14467
rect 14056 14436 14105 14464
rect 14056 14424 14062 14436
rect 14093 14433 14105 14436
rect 14139 14433 14151 14467
rect 14093 14427 14151 14433
rect 16850 14424 16856 14476
rect 16908 14424 16914 14476
rect 17788 14464 17816 14572
rect 18598 14560 18604 14612
rect 18656 14560 18662 14612
rect 18877 14603 18935 14609
rect 18877 14569 18889 14603
rect 18923 14600 18935 14603
rect 19242 14600 19248 14612
rect 18923 14572 19248 14600
rect 18923 14569 18935 14572
rect 18877 14563 18935 14569
rect 19242 14560 19248 14572
rect 19300 14560 19306 14612
rect 21910 14600 21916 14612
rect 19352 14572 21916 14600
rect 18509 14467 18567 14473
rect 17788 14436 18460 14464
rect 11612 14418 11664 14424
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 9309 14399 9367 14405
rect 9309 14396 9321 14399
rect 8720 14368 9321 14396
rect 8720 14356 8726 14368
rect 9309 14365 9321 14368
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 9493 14399 9551 14405
rect 9493 14365 9505 14399
rect 9539 14396 9551 14399
rect 9674 14396 9680 14408
rect 9539 14368 9680 14396
rect 9539 14365 9551 14368
rect 9493 14359 9551 14365
rect 9674 14356 9680 14368
rect 9732 14356 9738 14408
rect 10502 14356 10508 14408
rect 10560 14356 10566 14408
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 12066 14356 12072 14408
rect 12124 14356 12130 14408
rect 14366 14396 14372 14408
rect 14327 14368 14372 14396
rect 14366 14356 14372 14368
rect 14424 14356 14430 14408
rect 14734 14356 14740 14408
rect 14792 14396 14798 14408
rect 15010 14396 15016 14408
rect 14792 14368 15016 14396
rect 14792 14356 14798 14368
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15378 14356 15384 14408
rect 15436 14396 15442 14408
rect 15473 14399 15531 14405
rect 15473 14396 15485 14399
rect 15436 14368 15485 14396
rect 15436 14356 15442 14368
rect 15473 14365 15485 14368
rect 15519 14365 15531 14399
rect 15747 14399 15805 14405
rect 15747 14396 15759 14399
rect 15473 14359 15531 14365
rect 15580 14368 15759 14396
rect 7116 14300 8616 14328
rect 11256 14328 11284 14356
rect 12161 14331 12219 14337
rect 12161 14328 12173 14331
rect 11256 14300 12173 14328
rect 7116 14269 7144 14300
rect 12161 14297 12173 14300
rect 12207 14297 12219 14331
rect 12161 14291 12219 14297
rect 12434 14288 12440 14340
rect 12492 14328 12498 14340
rect 12529 14331 12587 14337
rect 12529 14328 12541 14331
rect 12492 14300 12541 14328
rect 12492 14288 12498 14300
rect 12529 14297 12541 14300
rect 12575 14297 12587 14331
rect 12529 14291 12587 14297
rect 12618 14288 12624 14340
rect 12676 14328 12682 14340
rect 15580 14328 15608 14368
rect 15747 14365 15759 14368
rect 15793 14396 15805 14399
rect 16482 14396 16488 14408
rect 15793 14368 16488 14396
rect 15793 14365 15805 14368
rect 15747 14359 15805 14365
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 16868 14396 16896 14424
rect 16868 14368 17080 14396
rect 17144 14375 17724 14396
rect 12676 14300 14412 14328
rect 12676 14288 12682 14300
rect 6328 14232 7034 14260
rect 7101 14263 7159 14269
rect 6328 14220 6334 14232
rect 7101 14229 7113 14263
rect 7147 14229 7159 14263
rect 7101 14223 7159 14229
rect 7466 14220 7472 14272
rect 7524 14260 7530 14272
rect 11149 14263 11207 14269
rect 11149 14260 11161 14263
rect 7524 14232 11161 14260
rect 7524 14220 7530 14232
rect 11149 14229 11161 14232
rect 11195 14229 11207 14263
rect 11149 14223 11207 14229
rect 11793 14263 11851 14269
rect 11793 14229 11805 14263
rect 11839 14260 11851 14263
rect 11974 14260 11980 14272
rect 11839 14232 11980 14260
rect 11839 14229 11851 14232
rect 11793 14223 11851 14229
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12897 14263 12955 14269
rect 12897 14229 12909 14263
rect 12943 14260 12955 14263
rect 12986 14260 12992 14272
rect 12943 14232 12992 14260
rect 12943 14229 12955 14232
rect 12897 14223 12955 14229
rect 12986 14220 12992 14232
rect 13044 14220 13050 14272
rect 14384 14260 14412 14300
rect 14568 14300 15608 14328
rect 14568 14260 14596 14300
rect 16206 14288 16212 14340
rect 16264 14328 16270 14340
rect 16574 14328 16580 14340
rect 16264 14300 16580 14328
rect 16264 14288 16270 14300
rect 16574 14288 16580 14300
rect 16632 14288 16638 14340
rect 14384 14232 14596 14260
rect 14734 14220 14740 14272
rect 14792 14260 14798 14272
rect 16485 14263 16543 14269
rect 16485 14260 16497 14263
rect 14792 14232 16497 14260
rect 14792 14220 14798 14232
rect 16485 14229 16497 14232
rect 16531 14229 16543 14263
rect 17052 14260 17080 14368
rect 17111 14369 17724 14375
rect 17111 14335 17123 14369
rect 17157 14368 17724 14369
rect 17157 14338 17172 14368
rect 17157 14335 17169 14338
rect 17111 14329 17169 14335
rect 17696 14272 17724 14368
rect 18138 14356 18144 14408
rect 18196 14396 18202 14408
rect 18233 14399 18291 14405
rect 18233 14396 18245 14399
rect 18196 14368 18245 14396
rect 18196 14356 18202 14368
rect 18233 14365 18245 14368
rect 18279 14365 18291 14399
rect 18233 14359 18291 14365
rect 18325 14399 18383 14405
rect 18325 14365 18337 14399
rect 18371 14365 18383 14399
rect 18432 14396 18460 14436
rect 18509 14433 18521 14467
rect 18555 14464 18567 14467
rect 18616 14464 18644 14560
rect 18690 14492 18696 14544
rect 18748 14532 18754 14544
rect 19352 14532 19380 14572
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 18748 14504 19380 14532
rect 18748 14492 18754 14504
rect 18555 14436 18644 14464
rect 18555 14433 18567 14436
rect 18509 14427 18567 14433
rect 18782 14424 18788 14476
rect 18840 14424 18846 14476
rect 18966 14424 18972 14476
rect 19024 14464 19030 14476
rect 19242 14464 19248 14476
rect 19024 14436 19248 14464
rect 19024 14424 19030 14436
rect 19242 14424 19248 14436
rect 19300 14424 19306 14476
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18432 14368 18613 14396
rect 18325 14359 18383 14365
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 18800 14396 18828 14424
rect 19061 14399 19119 14405
rect 19061 14396 19073 14399
rect 18800 14368 19073 14396
rect 18601 14359 18659 14365
rect 19061 14365 19073 14368
rect 19107 14365 19119 14399
rect 19061 14359 19119 14365
rect 19503 14369 19561 14375
rect 17402 14260 17408 14272
rect 17052 14232 17408 14260
rect 16485 14223 16543 14229
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 17678 14220 17684 14272
rect 17736 14220 17742 14272
rect 17865 14263 17923 14269
rect 17865 14229 17877 14263
rect 17911 14260 17923 14263
rect 18156 14260 18184 14356
rect 18340 14328 18368 14359
rect 18693 14331 18751 14337
rect 18693 14328 18705 14331
rect 18340 14300 18705 14328
rect 18693 14297 18705 14300
rect 18739 14297 18751 14331
rect 19503 14335 19515 14369
rect 19549 14366 19561 14369
rect 19549 14335 19562 14366
rect 19503 14329 19562 14335
rect 19534 14328 19562 14329
rect 19534 14300 19656 14328
rect 18693 14291 18751 14297
rect 19628 14272 19656 14300
rect 17911 14232 18184 14260
rect 18509 14263 18567 14269
rect 17911 14229 17923 14232
rect 17865 14223 17923 14229
rect 18509 14229 18521 14263
rect 18555 14260 18567 14263
rect 19426 14260 19432 14272
rect 18555 14232 19432 14260
rect 18555 14229 18567 14232
rect 18509 14223 18567 14229
rect 19426 14220 19432 14232
rect 19484 14220 19490 14272
rect 19610 14220 19616 14272
rect 19668 14220 19674 14272
rect 20162 14220 20168 14272
rect 20220 14260 20226 14272
rect 20257 14263 20315 14269
rect 20257 14260 20269 14263
rect 20220 14232 20269 14260
rect 20220 14220 20226 14232
rect 20257 14229 20269 14232
rect 20303 14229 20315 14263
rect 20257 14223 20315 14229
rect 1104 14170 21043 14192
rect 1104 14118 5894 14170
rect 5946 14118 5958 14170
rect 6010 14118 6022 14170
rect 6074 14118 6086 14170
rect 6138 14118 6150 14170
rect 6202 14118 10839 14170
rect 10891 14118 10903 14170
rect 10955 14118 10967 14170
rect 11019 14118 11031 14170
rect 11083 14118 11095 14170
rect 11147 14118 15784 14170
rect 15836 14118 15848 14170
rect 15900 14118 15912 14170
rect 15964 14118 15976 14170
rect 16028 14118 16040 14170
rect 16092 14118 20729 14170
rect 20781 14118 20793 14170
rect 20845 14118 20857 14170
rect 20909 14118 20921 14170
rect 20973 14118 20985 14170
rect 21037 14118 21043 14170
rect 1104 14096 21043 14118
rect 1946 14016 1952 14068
rect 2004 14016 2010 14068
rect 3050 14016 3056 14068
rect 3108 14056 3114 14068
rect 4249 14059 4307 14065
rect 4249 14056 4261 14059
rect 3108 14028 4261 14056
rect 3108 14016 3114 14028
rect 4249 14025 4261 14028
rect 4295 14025 4307 14059
rect 4249 14019 4307 14025
rect 5506 14028 8432 14056
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13988 1731 13991
rect 1762 13988 1768 14000
rect 1719 13960 1768 13988
rect 1719 13957 1731 13960
rect 1673 13951 1731 13957
rect 1762 13948 1768 13960
rect 1820 13948 1826 14000
rect 4062 13948 4068 14000
rect 4120 13988 4126 14000
rect 5506 13988 5534 14028
rect 4120 13960 4568 13988
rect 4120 13948 4126 13960
rect 3326 13880 3332 13932
rect 3384 13929 3390 13932
rect 3384 13923 3412 13929
rect 3400 13889 3412 13923
rect 3384 13883 3412 13889
rect 3384 13880 3390 13883
rect 3510 13880 3516 13932
rect 3568 13880 3574 13932
rect 4154 13880 4160 13932
rect 4212 13880 4218 13932
rect 4430 13880 4436 13932
rect 4488 13880 4494 13932
rect 106 13812 112 13864
rect 164 13852 170 13864
rect 2222 13852 2228 13864
rect 164 13824 2228 13852
rect 164 13812 170 13824
rect 2222 13812 2228 13824
rect 2280 13852 2286 13864
rect 2317 13855 2375 13861
rect 2317 13852 2329 13855
rect 2280 13824 2329 13852
rect 2280 13812 2286 13824
rect 2317 13821 2329 13824
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 2498 13812 2504 13864
rect 2556 13812 2562 13864
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 2961 13855 3019 13861
rect 2961 13852 2973 13855
rect 2924 13824 2973 13852
rect 2924 13812 2930 13824
rect 2961 13821 2973 13824
rect 3007 13821 3019 13855
rect 2961 13815 3019 13821
rect 3237 13855 3295 13861
rect 3237 13821 3249 13855
rect 3283 13852 3295 13855
rect 4172 13852 4200 13880
rect 3283 13824 4200 13852
rect 4540 13852 4568 13960
rect 4724 13960 5534 13988
rect 4724 13929 4752 13960
rect 4709 13923 4767 13929
rect 4709 13889 4721 13923
rect 4755 13889 4767 13923
rect 5074 13920 5080 13932
rect 4709 13883 4767 13889
rect 4816 13892 5080 13920
rect 4816 13852 4844 13892
rect 5074 13880 5080 13892
rect 5132 13929 5138 13932
rect 5132 13923 5193 13929
rect 5132 13889 5147 13923
rect 5181 13889 5193 13923
rect 5132 13883 5193 13889
rect 5132 13880 5138 13883
rect 6546 13880 6552 13932
rect 6604 13880 6610 13932
rect 7282 13880 7288 13932
rect 7340 13880 7346 13932
rect 7374 13880 7380 13932
rect 7432 13929 7438 13932
rect 7432 13923 7460 13929
rect 7448 13889 7460 13923
rect 7432 13883 7460 13889
rect 7432 13880 7438 13883
rect 4540 13824 4844 13852
rect 4893 13855 4951 13861
rect 3283 13821 3295 13824
rect 3237 13815 3295 13821
rect 4062 13784 4068 13796
rect 3896 13756 4068 13784
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 2314 13716 2320 13728
rect 2004 13688 2320 13716
rect 2004 13676 2010 13688
rect 2314 13676 2320 13688
rect 2372 13676 2378 13728
rect 3694 13676 3700 13728
rect 3752 13716 3758 13728
rect 3896 13716 3924 13756
rect 4062 13744 4068 13756
rect 4120 13744 4126 13796
rect 4172 13784 4200 13824
rect 4893 13821 4905 13855
rect 4939 13821 4951 13855
rect 4893 13815 4951 13821
rect 4706 13784 4712 13796
rect 4172 13756 4712 13784
rect 4706 13744 4712 13756
rect 4764 13744 4770 13796
rect 3752 13688 3924 13716
rect 3752 13676 3758 13688
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4157 13719 4215 13725
rect 4157 13716 4169 13719
rect 4028 13688 4169 13716
rect 4028 13676 4034 13688
rect 4157 13685 4169 13688
rect 4203 13685 4215 13719
rect 4157 13679 4215 13685
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 4525 13719 4583 13725
rect 4525 13716 4537 13719
rect 4488 13688 4537 13716
rect 4488 13676 4494 13688
rect 4525 13685 4537 13688
rect 4571 13685 4583 13719
rect 4525 13679 4583 13685
rect 4798 13676 4804 13728
rect 4856 13716 4862 13728
rect 4908 13716 4936 13815
rect 6086 13812 6092 13864
rect 6144 13852 6150 13864
rect 6365 13855 6423 13861
rect 6365 13852 6377 13855
rect 6144 13824 6377 13852
rect 6144 13812 6150 13824
rect 6365 13821 6377 13824
rect 6411 13821 6423 13855
rect 7561 13855 7619 13861
rect 6365 13815 6423 13821
rect 6748 13824 7144 13852
rect 5810 13784 5816 13796
rect 5552 13756 5816 13784
rect 5552 13716 5580 13756
rect 5810 13744 5816 13756
rect 5868 13744 5874 13796
rect 5905 13787 5963 13793
rect 5905 13753 5917 13787
rect 5951 13784 5963 13787
rect 6748 13784 6776 13824
rect 5951 13756 6776 13784
rect 7009 13787 7067 13793
rect 5951 13753 5963 13756
rect 5905 13747 5963 13753
rect 7009 13753 7021 13787
rect 7055 13753 7067 13787
rect 7009 13747 7067 13753
rect 4856 13688 5580 13716
rect 4856 13676 4862 13688
rect 5626 13676 5632 13728
rect 5684 13716 5690 13728
rect 7024 13716 7052 13747
rect 5684 13688 7052 13716
rect 7116 13716 7144 13824
rect 7561 13821 7573 13855
rect 7607 13852 7619 13855
rect 7607 13824 7972 13852
rect 7607 13821 7619 13824
rect 7561 13815 7619 13821
rect 7944 13716 7972 13824
rect 7116 13688 7972 13716
rect 5684 13676 5690 13688
rect 8202 13676 8208 13728
rect 8260 13676 8266 13728
rect 8404 13716 8432 14028
rect 8846 14016 8852 14068
rect 8904 14056 8910 14068
rect 10226 14056 10232 14068
rect 8904 14028 10232 14056
rect 8904 14016 8910 14028
rect 10226 14016 10232 14028
rect 10284 14016 10290 14068
rect 10594 14016 10600 14068
rect 10652 14056 10658 14068
rect 11422 14056 11428 14068
rect 10652 14028 11428 14056
rect 10652 14016 10658 14028
rect 11422 14016 11428 14028
rect 11480 14016 11486 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13357 14059 13415 14065
rect 13357 14056 13369 14059
rect 13228 14028 13369 14056
rect 13228 14016 13234 14028
rect 13357 14025 13369 14028
rect 13403 14025 13415 14059
rect 13357 14019 13415 14025
rect 15654 14016 15660 14068
rect 15712 14016 15718 14068
rect 16301 14059 16359 14065
rect 16301 14025 16313 14059
rect 16347 14056 16359 14059
rect 20162 14056 20168 14068
rect 16347 14028 18184 14056
rect 16347 14025 16359 14028
rect 16301 14019 16359 14025
rect 9030 13948 9036 14000
rect 9088 13988 9094 14000
rect 9490 13988 9496 14000
rect 9088 13960 9496 13988
rect 9088 13948 9094 13960
rect 9490 13948 9496 13960
rect 9548 13948 9554 14000
rect 12526 13948 12532 14000
rect 12584 13988 12590 14000
rect 12894 13988 12900 14000
rect 12584 13960 12900 13988
rect 12584 13948 12590 13960
rect 9048 13892 9352 13920
rect 9048 13864 9076 13892
rect 9030 13812 9036 13864
rect 9088 13812 9094 13864
rect 9324 13852 9352 13892
rect 9858 13880 9864 13932
rect 9916 13880 9922 13932
rect 10594 13929 10600 13932
rect 10551 13923 10600 13929
rect 10551 13889 10563 13923
rect 10597 13889 10600 13923
rect 10551 13883 10600 13889
rect 10594 13880 10600 13883
rect 10652 13880 10658 13932
rect 12634 13929 12662 13960
rect 12894 13948 12900 13960
rect 12952 13948 12958 14000
rect 13814 13948 13820 14000
rect 13872 13948 13878 14000
rect 14182 13948 14188 14000
rect 14240 13988 14246 14000
rect 15672 13988 15700 14016
rect 14240 13960 15700 13988
rect 16132 13960 16528 13988
rect 14240 13948 14246 13960
rect 12619 13923 12677 13929
rect 12619 13889 12631 13923
rect 12665 13889 12677 13923
rect 13832 13920 13860 13948
rect 14275 13923 14333 13929
rect 14275 13920 14287 13923
rect 13832 13892 14287 13920
rect 12619 13883 12677 13889
rect 14275 13889 14287 13892
rect 14321 13920 14333 13923
rect 15194 13920 15200 13932
rect 14321 13892 15200 13920
rect 14321 13889 14333 13892
rect 14275 13883 14333 13889
rect 15194 13880 15200 13892
rect 15252 13880 15258 13932
rect 15654 13880 15660 13932
rect 15712 13920 15718 13932
rect 16132 13920 16160 13960
rect 15712 13892 16160 13920
rect 15712 13880 15718 13892
rect 16206 13880 16212 13932
rect 16264 13880 16270 13932
rect 16500 13929 16528 13960
rect 16684 13960 17540 13988
rect 16684 13929 16712 13960
rect 17512 13932 17540 13960
rect 18046 13948 18052 14000
rect 18104 13948 18110 14000
rect 18156 13988 18184 14028
rect 18892 14028 20168 14056
rect 18690 13988 18696 14000
rect 18156 13960 18696 13988
rect 18690 13948 18696 13960
rect 18748 13948 18754 14000
rect 16485 13923 16543 13929
rect 16485 13889 16497 13923
rect 16531 13889 16543 13923
rect 16485 13883 16543 13889
rect 16669 13923 16727 13929
rect 16669 13889 16681 13923
rect 16715 13889 16727 13923
rect 16925 13923 16983 13929
rect 16925 13920 16937 13923
rect 16669 13883 16727 13889
rect 16776 13892 16937 13920
rect 9493 13855 9551 13861
rect 9493 13852 9505 13855
rect 9324 13824 9505 13852
rect 9493 13821 9505 13824
rect 9539 13821 9551 13855
rect 9493 13815 9551 13821
rect 9677 13855 9735 13861
rect 9677 13821 9689 13855
rect 9723 13821 9735 13855
rect 9876 13852 9904 13880
rect 10413 13855 10471 13861
rect 10413 13852 10425 13855
rect 9876 13824 10425 13852
rect 9677 13815 9735 13821
rect 10413 13821 10425 13824
rect 10459 13821 10471 13855
rect 10413 13815 10471 13821
rect 8662 13744 8668 13796
rect 8720 13784 8726 13796
rect 8846 13784 8852 13796
rect 8720 13756 8852 13784
rect 8720 13744 8726 13756
rect 8846 13744 8852 13756
rect 8904 13744 8910 13796
rect 9122 13744 9128 13796
rect 9180 13784 9186 13796
rect 9398 13784 9404 13796
rect 9180 13756 9404 13784
rect 9180 13744 9186 13756
rect 9398 13744 9404 13756
rect 9456 13784 9462 13796
rect 9692 13784 9720 13815
rect 10686 13812 10692 13864
rect 10744 13812 10750 13864
rect 10870 13812 10876 13864
rect 10928 13852 10934 13864
rect 12250 13852 12256 13864
rect 10928 13824 12256 13852
rect 10928 13812 10934 13824
rect 12250 13812 12256 13824
rect 12308 13812 12314 13864
rect 12345 13855 12403 13861
rect 12345 13821 12357 13855
rect 12391 13821 12403 13855
rect 12345 13815 12403 13821
rect 9456 13756 9720 13784
rect 9456 13744 9462 13756
rect 10134 13744 10140 13796
rect 10192 13744 10198 13796
rect 11333 13719 11391 13725
rect 11333 13716 11345 13719
rect 8404 13688 11345 13716
rect 11333 13685 11345 13688
rect 11379 13685 11391 13719
rect 11333 13679 11391 13685
rect 11422 13676 11428 13728
rect 11480 13716 11486 13728
rect 12360 13716 12388 13815
rect 13998 13812 14004 13864
rect 14056 13812 14062 13864
rect 15286 13812 15292 13864
rect 15344 13812 15350 13864
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 16776 13852 16804 13892
rect 16925 13889 16937 13892
rect 16971 13889 16983 13923
rect 16925 13883 16983 13889
rect 17494 13880 17500 13932
rect 17552 13880 17558 13932
rect 18064 13920 18092 13948
rect 18325 13923 18383 13929
rect 18325 13920 18337 13923
rect 18064 13892 18337 13920
rect 18325 13889 18337 13892
rect 18371 13889 18383 13923
rect 18325 13883 18383 13889
rect 18417 13923 18475 13929
rect 18417 13889 18429 13923
rect 18463 13889 18475 13923
rect 18417 13883 18475 13889
rect 15436 13824 16252 13852
rect 15436 13812 15442 13824
rect 15013 13787 15071 13793
rect 15013 13753 15025 13787
rect 15059 13784 15071 13787
rect 15304 13784 15332 13812
rect 15059 13756 15332 13784
rect 15059 13753 15071 13756
rect 15013 13747 15071 13753
rect 15396 13716 15424 13812
rect 16224 13796 16252 13824
rect 16592 13824 16804 13852
rect 15562 13744 15568 13796
rect 15620 13744 15626 13796
rect 15746 13744 15752 13796
rect 15804 13784 15810 13796
rect 16025 13787 16083 13793
rect 16025 13784 16037 13787
rect 15804 13756 16037 13784
rect 15804 13744 15810 13756
rect 16025 13753 16037 13756
rect 16071 13753 16083 13787
rect 16025 13747 16083 13753
rect 16206 13744 16212 13796
rect 16264 13744 16270 13796
rect 11480 13688 15424 13716
rect 15580 13716 15608 13744
rect 16390 13716 16396 13728
rect 15580 13688 16396 13716
rect 11480 13676 11486 13688
rect 16390 13676 16396 13688
rect 16448 13716 16454 13728
rect 16592 13716 16620 13824
rect 18138 13812 18144 13864
rect 18196 13852 18202 13864
rect 18432 13852 18460 13883
rect 18598 13880 18604 13932
rect 18656 13880 18662 13932
rect 18785 13923 18843 13929
rect 18785 13889 18797 13923
rect 18831 13920 18843 13923
rect 18892 13920 18920 14028
rect 19245 13991 19303 13997
rect 19245 13957 19257 13991
rect 19291 13988 19303 13991
rect 19981 13991 20039 13997
rect 19981 13988 19993 13991
rect 19291 13960 19993 13988
rect 19291 13957 19303 13960
rect 19245 13951 19303 13957
rect 19981 13957 19993 13960
rect 20027 13957 20039 13991
rect 19981 13951 20039 13957
rect 18831 13892 18920 13920
rect 18831 13889 18843 13892
rect 18785 13883 18843 13889
rect 18966 13880 18972 13932
rect 19024 13880 19030 13932
rect 19705 13923 19763 13929
rect 19444 13892 19656 13920
rect 18196 13824 18460 13852
rect 18877 13855 18935 13861
rect 18196 13812 18202 13824
rect 18877 13821 18889 13855
rect 18923 13852 18935 13855
rect 19444 13852 19472 13892
rect 18923 13824 19472 13852
rect 18923 13821 18935 13824
rect 18877 13815 18935 13821
rect 19518 13812 19524 13864
rect 19576 13812 19582 13864
rect 19628 13852 19656 13892
rect 19705 13889 19717 13923
rect 19751 13920 19763 13923
rect 20088 13920 20116 14028
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 20441 14059 20499 14065
rect 20441 14025 20453 14059
rect 20487 14056 20499 14059
rect 21266 14056 21272 14068
rect 20487 14028 21272 14056
rect 20487 14025 20499 14028
rect 20441 14019 20499 14025
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 19751 13892 20116 13920
rect 19751 13889 19763 13892
rect 19705 13883 19763 13889
rect 20162 13880 20168 13932
rect 20220 13880 20226 13932
rect 19981 13855 20039 13861
rect 19981 13852 19993 13855
rect 19628 13824 19993 13852
rect 19981 13821 19993 13824
rect 20027 13821 20039 13855
rect 19981 13815 20039 13821
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13784 18107 13787
rect 19058 13784 19064 13796
rect 18095 13756 19064 13784
rect 18095 13753 18107 13756
rect 18049 13747 18107 13753
rect 19058 13744 19064 13756
rect 19116 13744 19122 13796
rect 19334 13744 19340 13796
rect 19392 13784 19398 13796
rect 19797 13787 19855 13793
rect 19797 13784 19809 13787
rect 19392 13756 19809 13784
rect 19392 13744 19398 13756
rect 19797 13753 19809 13756
rect 19843 13753 19855 13787
rect 19797 13747 19855 13753
rect 16448 13688 16620 13716
rect 16448 13676 16454 13688
rect 17310 13676 17316 13728
rect 17368 13716 17374 13728
rect 17586 13716 17592 13728
rect 17368 13688 17592 13716
rect 17368 13676 17374 13688
rect 17586 13676 17592 13688
rect 17644 13676 17650 13728
rect 18141 13719 18199 13725
rect 18141 13685 18153 13719
rect 18187 13716 18199 13719
rect 18230 13716 18236 13728
rect 18187 13688 18236 13716
rect 18187 13685 18199 13688
rect 18141 13679 18199 13685
rect 18230 13676 18236 13688
rect 18288 13676 18294 13728
rect 18509 13719 18567 13725
rect 18509 13685 18521 13719
rect 18555 13716 18567 13719
rect 18598 13716 18604 13728
rect 18555 13688 18604 13716
rect 18555 13685 18567 13688
rect 18509 13679 18567 13685
rect 18598 13676 18604 13688
rect 18656 13676 18662 13728
rect 1104 13626 20884 13648
rect 1104 13574 3422 13626
rect 3474 13574 3486 13626
rect 3538 13574 3550 13626
rect 3602 13574 3614 13626
rect 3666 13574 3678 13626
rect 3730 13574 8367 13626
rect 8419 13574 8431 13626
rect 8483 13574 8495 13626
rect 8547 13574 8559 13626
rect 8611 13574 8623 13626
rect 8675 13574 13312 13626
rect 13364 13574 13376 13626
rect 13428 13574 13440 13626
rect 13492 13574 13504 13626
rect 13556 13574 13568 13626
rect 13620 13574 18257 13626
rect 18309 13574 18321 13626
rect 18373 13574 18385 13626
rect 18437 13574 18449 13626
rect 18501 13574 18513 13626
rect 18565 13574 20884 13626
rect 1104 13552 20884 13574
rect 1578 13472 1584 13524
rect 1636 13472 1642 13524
rect 3145 13515 3203 13521
rect 2240 13484 3096 13512
rect 2240 13444 2268 13484
rect 1596 13416 2268 13444
rect 3068 13444 3096 13484
rect 3145 13481 3157 13515
rect 3191 13512 3203 13515
rect 3326 13512 3332 13524
rect 3191 13484 3332 13512
rect 3191 13481 3203 13484
rect 3145 13475 3203 13481
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 3970 13472 3976 13524
rect 4028 13472 4034 13524
rect 8202 13512 8208 13524
rect 4126 13484 8208 13512
rect 3694 13444 3700 13456
rect 3068 13416 3700 13444
rect 1596 13320 1624 13416
rect 3694 13404 3700 13416
rect 3752 13404 3758 13456
rect 198 13268 204 13320
rect 256 13268 262 13320
rect 1578 13268 1584 13320
rect 1636 13268 1642 13320
rect 2133 13311 2191 13317
rect 2133 13277 2145 13311
rect 2179 13308 2191 13311
rect 4126 13308 4154 13484
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 9582 13512 9588 13524
rect 9232 13484 9588 13512
rect 9232 13456 9260 13484
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 10410 13512 10416 13524
rect 9968 13484 10416 13512
rect 5629 13447 5687 13453
rect 5629 13413 5641 13447
rect 5675 13444 5687 13447
rect 6454 13444 6460 13456
rect 5675 13416 6460 13444
rect 5675 13413 5687 13416
rect 5629 13407 5687 13413
rect 6454 13404 6460 13416
rect 6512 13404 6518 13456
rect 6638 13404 6644 13456
rect 6696 13404 6702 13456
rect 9214 13404 9220 13456
rect 9272 13404 9278 13456
rect 9398 13404 9404 13456
rect 9456 13444 9462 13456
rect 9968 13444 9996 13484
rect 10410 13472 10416 13484
rect 10468 13512 10474 13524
rect 11606 13512 11612 13524
rect 10468 13484 11612 13512
rect 10468 13472 10474 13484
rect 11606 13472 11612 13484
rect 11664 13472 11670 13524
rect 13357 13515 13415 13521
rect 13357 13481 13369 13515
rect 13403 13512 13415 13515
rect 14090 13512 14096 13524
rect 13403 13484 14096 13512
rect 13403 13481 13415 13484
rect 13357 13475 13415 13481
rect 14090 13472 14096 13484
rect 14148 13512 14154 13524
rect 15286 13512 15292 13524
rect 14148 13484 15292 13512
rect 14148 13472 14154 13484
rect 15286 13472 15292 13484
rect 15344 13472 15350 13524
rect 17037 13515 17095 13521
rect 17037 13512 17049 13515
rect 16040 13484 17049 13512
rect 9456 13416 9996 13444
rect 9456 13404 9462 13416
rect 5997 13379 6055 13385
rect 5997 13376 6009 13379
rect 5506 13348 6009 13376
rect 2179 13280 2268 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 216 13172 244 13268
rect 2240 13252 2268 13280
rect 2391 13281 2449 13287
rect 1489 13243 1547 13249
rect 1489 13209 1501 13243
rect 1535 13240 1547 13243
rect 1854 13240 1860 13252
rect 1535 13212 1860 13240
rect 1535 13209 1547 13212
rect 1489 13203 1547 13209
rect 1854 13200 1860 13212
rect 1912 13200 1918 13252
rect 2222 13200 2228 13252
rect 2280 13200 2286 13252
rect 2391 13247 2403 13281
rect 2437 13278 2449 13281
rect 3160 13280 4154 13308
rect 2437 13247 2450 13278
rect 3160 13252 3188 13280
rect 4522 13268 4528 13320
rect 4580 13268 4586 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 4798 13308 4804 13320
rect 4663 13280 4804 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 4891 13311 4949 13317
rect 4891 13277 4903 13311
rect 4937 13308 4949 13311
rect 4982 13308 4988 13320
rect 4937 13280 4988 13308
rect 4937 13277 4949 13280
rect 4891 13271 4949 13277
rect 4982 13268 4988 13280
rect 5040 13268 5046 13320
rect 5350 13268 5356 13320
rect 5408 13308 5414 13320
rect 5506 13308 5534 13348
rect 5997 13345 6009 13348
rect 6043 13376 6055 13379
rect 6086 13376 6092 13388
rect 6043 13348 6092 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6086 13336 6092 13348
rect 6144 13336 6150 13388
rect 6362 13336 6368 13388
rect 6420 13376 6426 13388
rect 9968 13385 9996 13416
rect 14182 13404 14188 13456
rect 14240 13444 14246 13456
rect 14550 13444 14556 13456
rect 14240 13416 14556 13444
rect 14240 13404 14246 13416
rect 11888 13388 11940 13394
rect 7034 13379 7092 13385
rect 7034 13376 7046 13379
rect 6420 13348 7046 13376
rect 6420 13336 6426 13348
rect 7034 13345 7046 13348
rect 7080 13345 7092 13379
rect 7034 13339 7092 13345
rect 7193 13379 7251 13385
rect 7193 13345 7205 13379
rect 7239 13376 7251 13379
rect 9953 13379 10011 13385
rect 7239 13348 7786 13376
rect 7239 13345 7251 13348
rect 7193 13339 7251 13345
rect 5408 13280 5534 13308
rect 6181 13311 6239 13317
rect 5408 13268 5414 13280
rect 6181 13277 6193 13311
rect 6227 13277 6239 13311
rect 6181 13271 6239 13277
rect 2391 13241 2450 13247
rect 2422 13172 2450 13241
rect 3142 13200 3148 13252
rect 3200 13200 3206 13252
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 4430 13240 4436 13252
rect 3927 13212 4436 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 4430 13200 4436 13212
rect 4488 13200 4494 13252
rect 5092 13212 5534 13240
rect 5092 13184 5120 13212
rect 3602 13172 3608 13184
rect 216 13144 3608 13172
rect 3602 13132 3608 13144
rect 3660 13132 3666 13184
rect 4338 13132 4344 13184
rect 4396 13132 4402 13184
rect 5074 13132 5080 13184
rect 5132 13132 5138 13184
rect 5506 13172 5534 13212
rect 6196 13172 6224 13271
rect 6914 13268 6920 13320
rect 6972 13268 6978 13320
rect 6546 13172 6552 13184
rect 5506 13144 6552 13172
rect 6546 13132 6552 13144
rect 6604 13132 6610 13184
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 7758 13172 7786 13348
rect 9953 13345 9965 13379
rect 9999 13345 10011 13379
rect 10413 13379 10471 13385
rect 10413 13376 10425 13379
rect 9953 13339 10011 13345
rect 10042 13348 10425 13376
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 9122 13308 9128 13320
rect 7892 13280 9128 13308
rect 7892 13268 7898 13280
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9674 13268 9680 13320
rect 9732 13308 9738 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9732 13280 9781 13308
rect 9732 13268 9738 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 10042 13308 10070 13348
rect 10413 13345 10425 13348
rect 10459 13345 10471 13379
rect 11514 13376 11520 13388
rect 10413 13339 10471 13345
rect 10704 13348 11520 13376
rect 10704 13317 10732 13348
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 14290 13385 14318 13416
rect 14550 13404 14556 13416
rect 14608 13404 14614 13456
rect 14734 13404 14740 13456
rect 14792 13404 14798 13456
rect 14277 13379 14335 13385
rect 14277 13345 14289 13379
rect 14323 13345 14335 13379
rect 14277 13339 14335 13345
rect 14642 13336 14648 13388
rect 14700 13376 14706 13388
rect 15130 13379 15188 13385
rect 15130 13376 15142 13379
rect 14700 13348 15142 13376
rect 14700 13336 14706 13348
rect 15130 13345 15142 13348
rect 15176 13345 15188 13379
rect 15130 13339 15188 13345
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 16040 13376 16068 13484
rect 17037 13481 17049 13484
rect 17083 13481 17095 13515
rect 17037 13475 17095 13481
rect 17402 13472 17408 13524
rect 17460 13472 17466 13524
rect 18138 13472 18144 13524
rect 18196 13512 18202 13524
rect 18417 13515 18475 13521
rect 18417 13512 18429 13515
rect 18196 13484 18429 13512
rect 18196 13472 18202 13484
rect 18417 13481 18429 13484
rect 18463 13481 18475 13515
rect 18417 13475 18475 13481
rect 18877 13515 18935 13521
rect 18877 13481 18889 13515
rect 18923 13512 18935 13515
rect 18966 13512 18972 13524
rect 18923 13484 18972 13512
rect 18923 13481 18935 13484
rect 18877 13475 18935 13481
rect 18966 13472 18972 13484
rect 19024 13472 19030 13524
rect 19702 13512 19708 13524
rect 19074 13484 19708 13512
rect 17420 13385 17448 13472
rect 15335 13348 16068 13376
rect 17405 13379 17463 13385
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 17405 13345 17417 13379
rect 17451 13345 17463 13379
rect 17405 13339 17463 13345
rect 11888 13330 11940 13336
rect 19074 13333 19102 13484
rect 19702 13472 19708 13484
rect 19760 13472 19766 13524
rect 19242 13336 19248 13388
rect 19300 13336 19306 13388
rect 19061 13327 19119 13333
rect 9769 13271 9827 13277
rect 9876 13280 10070 13308
rect 10689 13311 10747 13317
rect 9398 13200 9404 13252
rect 9456 13240 9462 13252
rect 9876 13240 9904 13280
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10778 13268 10784 13320
rect 10836 13317 10842 13320
rect 10836 13311 10885 13317
rect 10836 13277 10839 13311
rect 10873 13277 10885 13311
rect 10836 13271 10885 13277
rect 10836 13268 10842 13271
rect 10962 13268 10968 13320
rect 11020 13268 11026 13320
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 12216 13280 12357 13308
rect 12216 13268 12222 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 12526 13268 12532 13320
rect 12584 13308 12590 13320
rect 14093 13311 14151 13317
rect 12584 13280 12848 13308
rect 12584 13268 12590 13280
rect 9456 13212 9904 13240
rect 12437 13243 12495 13249
rect 9456 13200 9462 13212
rect 12437 13209 12449 13243
rect 12483 13240 12495 13243
rect 12710 13240 12716 13252
rect 12483 13212 12716 13240
rect 12483 13209 12495 13212
rect 12437 13203 12495 13209
rect 12710 13200 12716 13212
rect 12768 13200 12774 13252
rect 12820 13249 12848 13280
rect 14093 13277 14105 13311
rect 14139 13308 14151 13311
rect 14182 13308 14188 13320
rect 14139 13280 14188 13308
rect 14139 13277 14151 13280
rect 14093 13271 14151 13277
rect 14182 13268 14188 13280
rect 14240 13268 14246 13320
rect 15010 13268 15016 13320
rect 15068 13268 15074 13320
rect 16025 13311 16083 13317
rect 16025 13277 16037 13311
rect 16071 13308 16083 13311
rect 16206 13308 16212 13320
rect 16071 13280 16212 13308
rect 16071 13277 16083 13280
rect 16025 13271 16083 13277
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16299 13311 16357 13317
rect 16299 13277 16311 13311
rect 16345 13308 16357 13311
rect 16666 13308 16672 13320
rect 16345 13280 16672 13308
rect 16345 13277 16357 13280
rect 16299 13271 16357 13277
rect 16666 13268 16672 13280
rect 16724 13268 16730 13320
rect 19061 13293 19073 13327
rect 19107 13293 19119 13327
rect 19061 13287 19119 13293
rect 19352 13307 19530 13308
rect 19352 13301 19545 13307
rect 17663 13281 17721 13287
rect 17663 13278 17675 13281
rect 12805 13243 12863 13249
rect 12805 13209 12817 13243
rect 12851 13240 12863 13243
rect 13078 13240 13084 13252
rect 12851 13212 13084 13240
rect 12851 13209 12863 13212
rect 12805 13203 12863 13209
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 15930 13200 15936 13252
rect 15988 13200 15994 13252
rect 16482 13200 16488 13252
rect 16540 13240 16546 13252
rect 17034 13240 17040 13252
rect 16540 13212 17040 13240
rect 16540 13200 16546 13212
rect 17034 13200 17040 13212
rect 17092 13240 17098 13252
rect 17662 13247 17675 13278
rect 17709 13247 17721 13281
rect 19352 13280 19499 13301
rect 17662 13241 17721 13247
rect 17662 13240 17690 13241
rect 17092 13212 17690 13240
rect 17092 13200 17098 13212
rect 17862 13200 17868 13252
rect 17920 13240 17926 13252
rect 19352 13240 19380 13280
rect 19487 13267 19499 13280
rect 19533 13267 19545 13301
rect 19487 13261 19545 13267
rect 17920 13212 19380 13240
rect 17920 13200 17926 13212
rect 7064 13144 7786 13172
rect 7064 13132 7070 13144
rect 7834 13132 7840 13184
rect 7892 13132 7898 13184
rect 8202 13132 8208 13184
rect 8260 13172 8266 13184
rect 11609 13175 11667 13181
rect 11609 13172 11621 13175
rect 8260 13144 11621 13172
rect 8260 13132 8266 13144
rect 11609 13141 11621 13144
rect 11655 13141 11667 13175
rect 11609 13135 11667 13141
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 12069 13175 12127 13181
rect 12069 13172 12081 13175
rect 12032 13144 12081 13172
rect 12032 13132 12038 13144
rect 12069 13141 12081 13144
rect 12115 13141 12127 13175
rect 12069 13135 12127 13141
rect 12986 13132 12992 13184
rect 13044 13172 13050 13184
rect 13173 13175 13231 13181
rect 13173 13172 13185 13175
rect 13044 13144 13185 13172
rect 13044 13132 13050 13144
rect 13173 13141 13185 13144
rect 13219 13141 13231 13175
rect 13173 13135 13231 13141
rect 13906 13132 13912 13184
rect 13964 13172 13970 13184
rect 18414 13172 18420 13184
rect 13964 13144 18420 13172
rect 13964 13132 13970 13144
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 18598 13132 18604 13184
rect 18656 13172 18662 13184
rect 20257 13175 20315 13181
rect 20257 13172 20269 13175
rect 18656 13144 20269 13172
rect 18656 13132 18662 13144
rect 20257 13141 20269 13144
rect 20303 13141 20315 13175
rect 20257 13135 20315 13141
rect 1104 13082 21043 13104
rect 1104 13030 5894 13082
rect 5946 13030 5958 13082
rect 6010 13030 6022 13082
rect 6074 13030 6086 13082
rect 6138 13030 6150 13082
rect 6202 13030 10839 13082
rect 10891 13030 10903 13082
rect 10955 13030 10967 13082
rect 11019 13030 11031 13082
rect 11083 13030 11095 13082
rect 11147 13030 15784 13082
rect 15836 13030 15848 13082
rect 15900 13030 15912 13082
rect 15964 13030 15976 13082
rect 16028 13030 16040 13082
rect 16092 13030 20729 13082
rect 20781 13030 20793 13082
rect 20845 13030 20857 13082
rect 20909 13030 20921 13082
rect 20973 13030 20985 13082
rect 21037 13030 21043 13082
rect 1104 13008 21043 13030
rect 1581 12971 1639 12977
rect 1581 12937 1593 12971
rect 1627 12968 1639 12971
rect 1670 12968 1676 12980
rect 1627 12940 1676 12968
rect 1627 12937 1639 12940
rect 1581 12931 1639 12937
rect 1670 12928 1676 12940
rect 1728 12928 1734 12980
rect 4338 12968 4344 12980
rect 1964 12940 4344 12968
rect 1964 12909 1992 12940
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 6641 12971 6699 12977
rect 6641 12968 6653 12971
rect 4448 12940 6653 12968
rect 1949 12903 2007 12909
rect 1949 12869 1961 12903
rect 1995 12869 2007 12903
rect 1949 12863 2007 12869
rect 2501 12903 2559 12909
rect 2501 12869 2513 12903
rect 2547 12900 2559 12903
rect 3786 12900 3792 12912
rect 2547 12872 3792 12900
rect 2547 12869 2559 12872
rect 2501 12863 2559 12869
rect 3786 12860 3792 12872
rect 3844 12860 3850 12912
rect 4448 12900 4476 12940
rect 6641 12937 6653 12940
rect 6687 12937 6699 12971
rect 6641 12931 6699 12937
rect 6730 12928 6736 12980
rect 6788 12968 6794 12980
rect 7558 12968 7564 12980
rect 6788 12940 7564 12968
rect 6788 12928 6794 12940
rect 7558 12928 7564 12940
rect 7616 12928 7622 12980
rect 7834 12928 7840 12980
rect 7892 12928 7898 12980
rect 8294 12928 8300 12980
rect 8352 12928 8358 12980
rect 8662 12928 8668 12980
rect 8720 12968 8726 12980
rect 9677 12971 9735 12977
rect 8720 12940 9444 12968
rect 8720 12928 8726 12940
rect 4126 12872 4476 12900
rect 4617 12903 4675 12909
rect 1765 12835 1823 12841
rect 1765 12801 1777 12835
rect 1811 12832 1823 12835
rect 2866 12832 2872 12844
rect 1811 12804 2872 12832
rect 1811 12801 1823 12804
rect 1765 12795 1823 12801
rect 2866 12792 2872 12804
rect 2924 12792 2930 12844
rect 3234 12832 3240 12844
rect 3195 12804 3240 12832
rect 3234 12792 3240 12804
rect 3292 12792 3298 12844
rect 3602 12792 3608 12844
rect 3660 12792 3666 12844
rect 3694 12792 3700 12844
rect 3752 12832 3758 12844
rect 4126 12832 4154 12872
rect 4617 12869 4629 12903
rect 4663 12900 4675 12903
rect 4982 12900 4988 12912
rect 4663 12872 4988 12900
rect 4663 12869 4675 12872
rect 4617 12863 4675 12869
rect 3752 12804 4154 12832
rect 3752 12792 3758 12804
rect 2314 12724 2320 12776
rect 2372 12764 2378 12776
rect 2958 12764 2964 12776
rect 2372 12736 2964 12764
rect 2372 12724 2378 12736
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3620 12764 3648 12792
rect 4062 12764 4068 12776
rect 3620 12736 4068 12764
rect 4062 12724 4068 12736
rect 4120 12724 4126 12776
rect 4632 12696 4660 12863
rect 4982 12860 4988 12872
rect 5040 12900 5046 12912
rect 7852 12900 7880 12928
rect 9306 12900 9312 12912
rect 5040 12872 5178 12900
rect 5040 12860 5046 12872
rect 5150 12871 5178 12872
rect 6564 12872 7880 12900
rect 8956 12872 9312 12900
rect 5150 12865 5209 12871
rect 5150 12834 5163 12865
rect 5151 12831 5163 12834
rect 5197 12831 5209 12865
rect 6564 12841 6592 12872
rect 8956 12871 8984 12872
rect 8923 12865 8984 12871
rect 5151 12825 5209 12831
rect 6549 12835 6607 12841
rect 6549 12801 6561 12835
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 7466 12832 7472 12844
rect 6871 12804 7472 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 7466 12792 7472 12804
rect 7524 12792 7530 12844
rect 7559 12835 7617 12841
rect 7559 12801 7571 12835
rect 7605 12832 7617 12835
rect 8110 12832 8116 12844
rect 7605 12804 8116 12832
rect 7605 12801 7617 12804
rect 7559 12795 7617 12801
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 8923 12831 8935 12865
rect 8969 12834 8984 12865
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 8969 12831 8981 12834
rect 8923 12825 8981 12831
rect 9416 12832 9444 12940
rect 9677 12937 9689 12971
rect 9723 12968 9735 12971
rect 10502 12968 10508 12980
rect 9723 12940 10508 12968
rect 9723 12937 9735 12940
rect 9677 12931 9735 12937
rect 10502 12928 10508 12940
rect 10560 12928 10566 12980
rect 11057 12971 11115 12977
rect 11057 12937 11069 12971
rect 11103 12968 11115 12971
rect 11882 12968 11888 12980
rect 11103 12940 11888 12968
rect 11103 12937 11115 12940
rect 11057 12931 11115 12937
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 13722 12928 13728 12980
rect 13780 12968 13786 12980
rect 16301 12971 16359 12977
rect 13780 12940 16252 12968
rect 13780 12928 13786 12940
rect 11974 12860 11980 12912
rect 12032 12900 12038 12912
rect 12069 12903 12127 12909
rect 12069 12900 12081 12903
rect 12032 12872 12081 12900
rect 12032 12860 12038 12872
rect 12069 12869 12081 12872
rect 12115 12869 12127 12903
rect 12069 12863 12127 12869
rect 12158 12860 12164 12912
rect 12216 12900 12222 12912
rect 12345 12903 12403 12909
rect 12345 12900 12357 12903
rect 12216 12872 12357 12900
rect 12216 12860 12222 12872
rect 12345 12869 12357 12872
rect 12391 12869 12403 12903
rect 12345 12863 12403 12869
rect 12805 12903 12863 12909
rect 12805 12869 12817 12903
rect 12851 12900 12863 12903
rect 13078 12900 13084 12912
rect 12851 12872 13084 12900
rect 12851 12869 12863 12872
rect 12805 12863 12863 12869
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 13173 12903 13231 12909
rect 13173 12869 13185 12903
rect 13219 12869 13231 12903
rect 13173 12863 13231 12869
rect 10287 12835 10345 12841
rect 10287 12832 10299 12835
rect 9416 12804 10299 12832
rect 10287 12801 10299 12804
rect 10333 12832 10345 12835
rect 11698 12832 11704 12844
rect 10333 12804 11704 12832
rect 10333 12801 10345 12804
rect 10287 12795 10345 12801
rect 11698 12792 11704 12804
rect 11756 12792 11762 12844
rect 12434 12792 12440 12844
rect 12492 12792 12498 12844
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13188 12832 13216 12863
rect 14274 12860 14280 12912
rect 14332 12860 14338 12912
rect 16224 12900 16252 12940
rect 16301 12937 16313 12971
rect 16347 12968 16359 12971
rect 18046 12968 18052 12980
rect 16347 12940 18052 12968
rect 16347 12937 16359 12940
rect 16301 12931 16359 12937
rect 18046 12928 18052 12940
rect 18104 12928 18110 12980
rect 18138 12928 18144 12980
rect 18196 12928 18202 12980
rect 18877 12971 18935 12977
rect 18877 12937 18889 12971
rect 18923 12968 18935 12971
rect 20162 12968 20168 12980
rect 18923 12940 20168 12968
rect 18923 12937 18935 12940
rect 18877 12931 18935 12937
rect 20162 12928 20168 12940
rect 20220 12928 20226 12980
rect 20441 12971 20499 12977
rect 20441 12937 20453 12971
rect 20487 12968 20499 12971
rect 21266 12968 21272 12980
rect 20487 12940 21272 12968
rect 20487 12937 20499 12940
rect 20441 12931 20499 12937
rect 21266 12928 21272 12940
rect 21324 12928 21330 12980
rect 16224 12872 18000 12900
rect 13044 12804 13216 12832
rect 13044 12792 13050 12804
rect 13998 12792 14004 12844
rect 14056 12832 14062 12844
rect 14292 12832 14320 12860
rect 14461 12835 14519 12841
rect 14461 12832 14473 12835
rect 14056 12804 14473 12832
rect 14056 12792 14062 12804
rect 14461 12801 14473 12804
rect 14507 12801 14519 12835
rect 14461 12795 14519 12801
rect 14642 12792 14648 12844
rect 14700 12792 14706 12844
rect 15286 12792 15292 12844
rect 15344 12841 15350 12844
rect 15344 12835 15372 12841
rect 15360 12801 15372 12835
rect 15344 12795 15372 12801
rect 15344 12792 15350 12795
rect 16390 12792 16396 12844
rect 16448 12832 16454 12844
rect 16485 12835 16543 12841
rect 16485 12832 16497 12835
rect 16448 12804 16497 12832
rect 16448 12792 16454 12804
rect 16485 12801 16497 12804
rect 16531 12801 16543 12835
rect 16942 12832 16948 12844
rect 16903 12804 16948 12832
rect 16485 12795 16543 12801
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 4798 12724 4804 12776
rect 4856 12764 4862 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4856 12736 4905 12764
rect 4856 12724 4862 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 7285 12767 7343 12773
rect 7285 12733 7297 12767
rect 7331 12733 7343 12767
rect 7285 12727 7343 12733
rect 3620 12668 4660 12696
rect 2038 12588 2044 12640
rect 2096 12588 2102 12640
rect 2590 12588 2596 12640
rect 2648 12588 2654 12640
rect 2682 12588 2688 12640
rect 2740 12628 2746 12640
rect 3620 12628 3648 12668
rect 5626 12656 5632 12708
rect 5684 12696 5690 12708
rect 5684 12668 5948 12696
rect 5684 12656 5690 12668
rect 2740 12600 3648 12628
rect 3973 12631 4031 12637
rect 2740 12588 2746 12600
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 5810 12628 5816 12640
rect 4019 12600 5816 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 5920 12637 5948 12668
rect 6362 12656 6368 12708
rect 6420 12656 6426 12708
rect 5905 12631 5963 12637
rect 5905 12597 5917 12631
rect 5951 12597 5963 12631
rect 7300 12628 7328 12727
rect 8662 12724 8668 12776
rect 8720 12724 8726 12776
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 7374 12628 7380 12640
rect 7300 12600 7380 12628
rect 5905 12591 5963 12597
rect 7374 12588 7380 12600
rect 7432 12628 7438 12640
rect 8680 12628 8708 12724
rect 10060 12696 10088 12727
rect 12526 12724 12532 12776
rect 12584 12724 12590 12776
rect 13170 12724 13176 12776
rect 13228 12764 13234 12776
rect 14277 12767 14335 12773
rect 14277 12764 14289 12767
rect 13228 12736 14289 12764
rect 13228 12724 13234 12736
rect 14277 12733 14289 12736
rect 14323 12733 14335 12767
rect 14277 12727 14335 12733
rect 13357 12699 13415 12705
rect 10060 12668 10180 12696
rect 10152 12640 10180 12668
rect 13357 12665 13369 12699
rect 13403 12696 13415 12699
rect 14660 12696 14688 12792
rect 15010 12764 15016 12776
rect 13403 12668 14688 12696
rect 14844 12736 15016 12764
rect 13403 12665 13415 12668
rect 13357 12659 13415 12665
rect 7432 12600 8708 12628
rect 7432 12588 7438 12600
rect 10134 12588 10140 12640
rect 10192 12628 10198 12640
rect 11882 12628 11888 12640
rect 10192 12600 11888 12628
rect 10192 12588 10198 12600
rect 11882 12588 11888 12600
rect 11940 12588 11946 12640
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 14844 12628 14872 12736
rect 15010 12724 15016 12736
rect 15068 12764 15074 12776
rect 15197 12767 15255 12773
rect 15197 12764 15209 12767
rect 15068 12736 15209 12764
rect 15068 12724 15074 12736
rect 15197 12733 15209 12736
rect 15243 12733 15255 12767
rect 15197 12727 15255 12733
rect 15473 12767 15531 12773
rect 15473 12733 15485 12767
rect 15519 12764 15531 12767
rect 15519 12736 16068 12764
rect 15519 12733 15531 12736
rect 15473 12727 15531 12733
rect 14921 12699 14979 12705
rect 14921 12665 14933 12699
rect 14967 12665 14979 12699
rect 14921 12659 14979 12665
rect 14700 12600 14872 12628
rect 14936 12628 14964 12659
rect 15562 12628 15568 12640
rect 14936 12600 15568 12628
rect 14700 12588 14706 12600
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 16040 12628 16068 12736
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 16669 12767 16727 12773
rect 16669 12764 16681 12767
rect 16264 12736 16681 12764
rect 16264 12724 16270 12736
rect 16669 12733 16681 12736
rect 16715 12733 16727 12767
rect 17972 12764 18000 12872
rect 18049 12835 18107 12841
rect 18049 12801 18061 12835
rect 18095 12832 18107 12835
rect 18156 12832 18184 12928
rect 19426 12860 19432 12912
rect 19484 12900 19490 12912
rect 19484 12872 20208 12900
rect 19484 12860 19490 12872
rect 18598 12832 18604 12844
rect 18095 12804 18184 12832
rect 18248 12804 18604 12832
rect 18095 12801 18107 12804
rect 18049 12795 18107 12801
rect 18248 12764 18276 12804
rect 18598 12792 18604 12804
rect 18656 12792 18662 12844
rect 18782 12792 18788 12844
rect 18840 12832 18846 12844
rect 20180 12841 20208 12872
rect 19061 12835 19119 12841
rect 19061 12832 19073 12835
rect 18840 12804 19073 12832
rect 18840 12792 18846 12804
rect 19061 12801 19073 12804
rect 19107 12801 19119 12835
rect 19061 12795 19119 12801
rect 19613 12835 19671 12841
rect 19613 12801 19625 12835
rect 19659 12801 19671 12835
rect 19613 12795 19671 12801
rect 20165 12835 20223 12841
rect 20165 12801 20177 12835
rect 20211 12801 20223 12835
rect 20165 12795 20223 12801
rect 17972 12736 18276 12764
rect 16669 12727 16727 12733
rect 18322 12724 18328 12776
rect 18380 12724 18386 12776
rect 18414 12724 18420 12776
rect 18472 12764 18478 12776
rect 18877 12767 18935 12773
rect 18877 12764 18889 12767
rect 18472 12736 18889 12764
rect 18472 12724 18478 12736
rect 18877 12733 18889 12736
rect 18923 12733 18935 12767
rect 19628 12764 19656 12795
rect 21358 12764 21364 12776
rect 19628 12736 21364 12764
rect 18877 12727 18935 12733
rect 21358 12724 21364 12736
rect 21416 12724 21422 12776
rect 16114 12656 16120 12708
rect 16172 12656 16178 12708
rect 19518 12696 19524 12708
rect 18708 12668 19524 12696
rect 17681 12631 17739 12637
rect 17681 12628 17693 12631
rect 16040 12600 17693 12628
rect 17681 12597 17693 12600
rect 17727 12597 17739 12631
rect 17681 12591 17739 12597
rect 18138 12588 18144 12640
rect 18196 12588 18202 12640
rect 18233 12631 18291 12637
rect 18233 12597 18245 12631
rect 18279 12628 18291 12631
rect 18598 12628 18604 12640
rect 18279 12600 18604 12628
rect 18279 12597 18291 12600
rect 18233 12591 18291 12597
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 18708 12637 18736 12668
rect 19518 12656 19524 12668
rect 19576 12656 19582 12708
rect 19978 12656 19984 12708
rect 20036 12696 20042 12708
rect 21266 12696 21272 12708
rect 20036 12668 21272 12696
rect 20036 12656 20042 12668
rect 21266 12656 21272 12668
rect 21324 12656 21330 12708
rect 18693 12631 18751 12637
rect 18693 12597 18705 12631
rect 18739 12597 18751 12631
rect 18693 12591 18751 12597
rect 19334 12588 19340 12640
rect 19392 12588 19398 12640
rect 19886 12588 19892 12640
rect 19944 12588 19950 12640
rect 1104 12538 20884 12560
rect 1104 12486 3422 12538
rect 3474 12486 3486 12538
rect 3538 12486 3550 12538
rect 3602 12486 3614 12538
rect 3666 12486 3678 12538
rect 3730 12486 8367 12538
rect 8419 12486 8431 12538
rect 8483 12486 8495 12538
rect 8547 12486 8559 12538
rect 8611 12486 8623 12538
rect 8675 12486 13312 12538
rect 13364 12486 13376 12538
rect 13428 12486 13440 12538
rect 13492 12486 13504 12538
rect 13556 12486 13568 12538
rect 13620 12486 18257 12538
rect 18309 12486 18321 12538
rect 18373 12486 18385 12538
rect 18437 12486 18449 12538
rect 18501 12486 18513 12538
rect 18565 12486 20884 12538
rect 1104 12464 20884 12486
rect 934 12384 940 12436
rect 992 12424 998 12436
rect 1765 12427 1823 12433
rect 1765 12424 1777 12427
rect 992 12396 1777 12424
rect 992 12384 998 12396
rect 1765 12393 1777 12396
rect 1811 12393 1823 12427
rect 1765 12387 1823 12393
rect 4154 12384 4160 12436
rect 4212 12384 4218 12436
rect 4522 12384 4528 12436
rect 4580 12424 4586 12436
rect 5166 12424 5172 12436
rect 4580 12396 5172 12424
rect 4580 12384 4586 12396
rect 5166 12384 5172 12396
rect 5224 12424 5230 12436
rect 5718 12424 5724 12436
rect 5224 12396 5724 12424
rect 5224 12384 5230 12396
rect 5718 12384 5724 12396
rect 5776 12384 5782 12436
rect 8202 12424 8208 12436
rect 7024 12396 8208 12424
rect 3329 12359 3387 12365
rect 3329 12325 3341 12359
rect 3375 12356 3387 12359
rect 5261 12359 5319 12365
rect 5261 12356 5273 12359
rect 3375 12328 5273 12356
rect 3375 12325 3387 12328
rect 3329 12319 3387 12325
rect 5261 12325 5273 12328
rect 5307 12325 5319 12359
rect 5261 12319 5319 12325
rect 6362 12316 6368 12368
rect 6420 12356 6426 12368
rect 6822 12356 6828 12368
rect 6420 12328 6828 12356
rect 6420 12316 6426 12328
rect 6822 12316 6828 12328
rect 6880 12316 6886 12368
rect 2314 12248 2320 12300
rect 2372 12248 2378 12300
rect 4430 12248 4436 12300
rect 4488 12288 4494 12300
rect 4617 12291 4675 12297
rect 4488 12260 4568 12288
rect 4488 12248 4494 12260
rect 1578 12180 1584 12232
rect 1636 12220 1642 12232
rect 1673 12223 1731 12229
rect 1673 12220 1685 12223
rect 1636 12192 1685 12220
rect 1636 12180 1642 12192
rect 1673 12189 1685 12192
rect 1719 12189 1731 12223
rect 2575 12193 2633 12199
rect 2575 12190 2587 12193
rect 1673 12183 1731 12189
rect 14 12112 20 12164
rect 72 12152 78 12164
rect 2314 12152 2320 12164
rect 72 12124 2320 12152
rect 72 12112 78 12124
rect 2314 12112 2320 12124
rect 2372 12112 2378 12164
rect 2406 12112 2412 12164
rect 2464 12152 2470 12164
rect 2516 12162 2587 12190
rect 2516 12152 2544 12162
rect 2575 12159 2587 12162
rect 2621 12159 2633 12193
rect 3602 12180 3608 12232
rect 3660 12220 3666 12232
rect 3970 12220 3976 12232
rect 3660 12192 3976 12220
rect 3660 12180 3666 12192
rect 3970 12180 3976 12192
rect 4028 12220 4034 12232
rect 4540 12229 4568 12260
rect 4617 12257 4629 12291
rect 4663 12288 4675 12291
rect 5166 12288 5172 12300
rect 4663 12260 5172 12288
rect 4663 12257 4675 12260
rect 4617 12251 4675 12257
rect 5166 12248 5172 12260
rect 5224 12248 5230 12300
rect 5810 12248 5816 12300
rect 5868 12248 5874 12300
rect 4525 12223 4583 12229
rect 4028 12192 4476 12220
rect 4028 12180 4034 12192
rect 2575 12153 2633 12159
rect 3881 12155 3939 12161
rect 2464 12124 2544 12152
rect 2464 12112 2470 12124
rect 2516 12084 2544 12124
rect 3881 12121 3893 12155
rect 3927 12152 3939 12155
rect 4448 12152 4476 12192
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 4801 12223 4859 12229
rect 4801 12189 4813 12223
rect 4847 12189 4859 12223
rect 4801 12183 4859 12189
rect 4816 12152 4844 12183
rect 5534 12180 5540 12232
rect 5592 12180 5598 12232
rect 5718 12229 5724 12232
rect 5675 12223 5724 12229
rect 5675 12220 5687 12223
rect 5669 12216 5687 12220
rect 5644 12189 5687 12216
rect 5721 12189 5724 12223
rect 5644 12182 5724 12189
rect 5718 12180 5724 12182
rect 5776 12180 5782 12232
rect 7024 12229 7052 12396
rect 8202 12384 8208 12396
rect 8260 12384 8266 12436
rect 8481 12427 8539 12433
rect 8481 12393 8493 12427
rect 8527 12424 8539 12427
rect 9398 12424 9404 12436
rect 8527 12396 9404 12424
rect 8527 12393 8539 12396
rect 8481 12387 8539 12393
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9582 12384 9588 12436
rect 9640 12384 9646 12436
rect 11238 12424 11244 12436
rect 9784 12396 11244 12424
rect 8662 12316 8668 12368
rect 8720 12356 8726 12368
rect 9600 12356 9628 12384
rect 8720 12328 9628 12356
rect 8720 12316 8726 12328
rect 7374 12248 7380 12300
rect 7432 12288 7438 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7432 12260 7481 12288
rect 7432 12248 7438 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 8202 12248 8208 12300
rect 8260 12288 8266 12300
rect 9214 12288 9220 12300
rect 8260 12260 9220 12288
rect 8260 12248 8266 12260
rect 9214 12248 9220 12260
rect 9272 12288 9278 12300
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 9272 12260 9597 12288
rect 9272 12248 9278 12260
rect 9585 12257 9597 12260
rect 9631 12288 9643 12291
rect 9784 12288 9812 12396
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 13817 12427 13875 12433
rect 13817 12393 13829 12427
rect 13863 12424 13875 12427
rect 13906 12424 13912 12436
rect 13863 12396 13912 12424
rect 13863 12393 13875 12396
rect 13817 12387 13875 12393
rect 13906 12384 13912 12396
rect 13964 12384 13970 12436
rect 14458 12384 14464 12436
rect 14516 12384 14522 12436
rect 17129 12427 17187 12433
rect 17129 12424 17141 12427
rect 14844 12396 17141 12424
rect 9858 12316 9864 12368
rect 9916 12356 9922 12368
rect 13173 12359 13231 12365
rect 9916 12328 10180 12356
rect 9916 12316 9922 12328
rect 10152 12300 10180 12328
rect 13173 12325 13185 12359
rect 13219 12356 13231 12359
rect 13998 12356 14004 12368
rect 13219 12328 14004 12356
rect 13219 12325 13231 12328
rect 13173 12319 13231 12325
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 14476 12356 14504 12384
rect 14056 12328 14504 12356
rect 14056 12316 14062 12328
rect 14642 12316 14648 12368
rect 14700 12316 14706 12368
rect 14844 12365 14872 12396
rect 17129 12393 17141 12396
rect 17175 12393 17187 12427
rect 17129 12387 17187 12393
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 18417 12427 18475 12433
rect 18417 12424 18429 12427
rect 18196 12396 18429 12424
rect 18196 12384 18202 12396
rect 18417 12393 18429 12396
rect 18463 12393 18475 12427
rect 18417 12387 18475 12393
rect 18969 12427 19027 12433
rect 18969 12393 18981 12427
rect 19015 12424 19027 12427
rect 19058 12424 19064 12436
rect 19015 12396 19064 12424
rect 19015 12393 19027 12396
rect 18969 12387 19027 12393
rect 19058 12384 19064 12396
rect 19116 12384 19122 12436
rect 14829 12359 14887 12365
rect 14829 12325 14841 12359
rect 14875 12325 14887 12359
rect 14829 12319 14887 12325
rect 18230 12316 18236 12368
rect 18288 12356 18294 12368
rect 19150 12356 19156 12368
rect 18288 12328 19156 12356
rect 18288 12316 18294 12328
rect 19150 12316 19156 12328
rect 19208 12316 19214 12368
rect 19242 12316 19248 12368
rect 19300 12356 19306 12368
rect 19978 12356 19984 12368
rect 19300 12328 19984 12356
rect 19300 12316 19306 12328
rect 19978 12316 19984 12328
rect 20036 12316 20042 12368
rect 9631 12260 9812 12288
rect 9631 12257 9643 12260
rect 9585 12251 9643 12257
rect 10042 12248 10048 12300
rect 10100 12248 10106 12300
rect 10134 12248 10140 12300
rect 10192 12288 10198 12300
rect 10321 12291 10379 12297
rect 10321 12288 10333 12291
rect 10192 12260 10333 12288
rect 10192 12248 10198 12260
rect 10321 12257 10333 12260
rect 10367 12257 10379 12291
rect 10321 12251 10379 12257
rect 10410 12248 10416 12300
rect 10468 12297 10474 12300
rect 10468 12291 10496 12297
rect 10484 12257 10496 12291
rect 10468 12251 10496 12257
rect 10468 12248 10474 12251
rect 12618 12248 12624 12300
rect 12676 12248 12682 12300
rect 14090 12288 14096 12300
rect 13924 12260 14096 12288
rect 6733 12223 6791 12229
rect 6733 12189 6745 12223
rect 6779 12189 6791 12223
rect 6733 12183 6791 12189
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12189 7067 12223
rect 7009 12183 7067 12189
rect 7743 12223 7801 12229
rect 7743 12189 7755 12223
rect 7789 12220 7801 12223
rect 8294 12220 8300 12232
rect 7789 12192 8300 12220
rect 7789 12189 7801 12192
rect 7743 12183 7801 12189
rect 3927 12124 4384 12152
rect 4448 12124 4844 12152
rect 6748 12152 6776 12183
rect 8294 12180 8300 12192
rect 8352 12220 8358 12232
rect 8570 12220 8576 12232
rect 8352 12192 8576 12220
rect 8352 12180 8358 12192
rect 8570 12180 8576 12192
rect 8628 12180 8634 12232
rect 8846 12180 8852 12232
rect 8904 12220 8910 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 8904 12192 9413 12220
rect 8904 12180 8910 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9306 12152 9312 12164
rect 6748 12124 9312 12152
rect 3927 12121 3939 12124
rect 3881 12115 3939 12121
rect 2958 12084 2964 12096
rect 2516 12056 2964 12084
rect 2958 12044 2964 12056
rect 3016 12044 3022 12096
rect 4356 12093 4384 12124
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 4341 12087 4399 12093
rect 4341 12053 4353 12087
rect 4387 12053 4399 12087
rect 4341 12047 4399 12053
rect 4430 12044 4436 12096
rect 4488 12084 4494 12096
rect 6457 12087 6515 12093
rect 6457 12084 6469 12087
rect 4488 12056 6469 12084
rect 4488 12044 4494 12056
rect 6457 12053 6469 12056
rect 6503 12053 6515 12087
rect 6457 12047 6515 12053
rect 6546 12044 6552 12096
rect 6604 12044 6610 12096
rect 6822 12044 6828 12096
rect 6880 12044 6886 12096
rect 7098 12044 7104 12096
rect 7156 12084 7162 12096
rect 7374 12084 7380 12096
rect 7156 12056 7380 12084
rect 7156 12044 7162 12056
rect 7374 12044 7380 12056
rect 7432 12044 7438 12096
rect 9416 12084 9444 12183
rect 10594 12180 10600 12232
rect 10652 12180 10658 12232
rect 12158 12180 12164 12232
rect 12216 12180 12222 12232
rect 13078 12180 13084 12232
rect 13136 12180 13142 12232
rect 13722 12180 13728 12232
rect 13780 12180 13786 12232
rect 13924 12229 13952 12260
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14660 12288 14688 12316
rect 15286 12297 15292 12300
rect 15105 12291 15163 12297
rect 15105 12288 15117 12291
rect 14290 12260 15117 12288
rect 13909 12223 13967 12229
rect 13909 12189 13921 12223
rect 13955 12189 13967 12223
rect 13909 12183 13967 12189
rect 14182 12180 14188 12232
rect 14240 12180 14246 12232
rect 11164 12124 12204 12152
rect 9858 12084 9864 12096
rect 9416 12056 9864 12084
rect 9858 12044 9864 12056
rect 9916 12044 9922 12096
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 11164 12084 11192 12124
rect 10468 12056 11192 12084
rect 10468 12044 10474 12056
rect 11238 12044 11244 12096
rect 11296 12044 11302 12096
rect 11885 12087 11943 12093
rect 11885 12053 11897 12087
rect 11931 12084 11943 12087
rect 11974 12084 11980 12096
rect 11931 12056 11980 12084
rect 11931 12053 11943 12056
rect 11885 12047 11943 12053
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12176 12084 12204 12124
rect 12250 12112 12256 12164
rect 12308 12112 12314 12164
rect 12621 12155 12679 12161
rect 12621 12121 12633 12155
rect 12667 12152 12679 12155
rect 13096 12152 13124 12180
rect 12667 12124 13124 12152
rect 12667 12121 12679 12124
rect 12621 12115 12679 12121
rect 12636 12084 12664 12115
rect 13630 12112 13636 12164
rect 13688 12152 13694 12164
rect 14290 12152 14318 12260
rect 15105 12257 15117 12260
rect 15151 12257 15163 12291
rect 15105 12251 15163 12257
rect 15243 12291 15292 12297
rect 15243 12257 15255 12291
rect 15289 12257 15292 12291
rect 15243 12251 15292 12257
rect 15286 12248 15292 12251
rect 15344 12248 15350 12300
rect 15391 12291 15449 12297
rect 15391 12257 15403 12291
rect 15437 12288 15449 12291
rect 15437 12260 16068 12288
rect 15437 12257 15449 12260
rect 15391 12251 15449 12257
rect 16040 12232 16068 12260
rect 17310 12248 17316 12300
rect 17368 12288 17374 12300
rect 20349 12291 20407 12297
rect 20349 12288 20361 12291
rect 17368 12260 20361 12288
rect 17368 12248 17374 12260
rect 20349 12257 20361 12260
rect 20395 12257 20407 12291
rect 20349 12251 20407 12257
rect 14369 12223 14427 12229
rect 14369 12189 14381 12223
rect 14415 12220 14427 12223
rect 14550 12220 14556 12232
rect 14415 12192 14556 12220
rect 14415 12189 14427 12192
rect 14369 12183 14427 12189
rect 14550 12180 14556 12192
rect 14608 12180 14614 12232
rect 16022 12180 16028 12232
rect 16080 12180 16086 12232
rect 16117 12223 16175 12229
rect 16117 12189 16129 12223
rect 16163 12189 16175 12223
rect 16117 12183 16175 12189
rect 16391 12223 16449 12229
rect 16391 12189 16403 12223
rect 16437 12189 16449 12223
rect 16391 12183 16449 12189
rect 13688 12124 14318 12152
rect 13688 12112 13694 12124
rect 15930 12112 15936 12164
rect 15988 12152 15994 12164
rect 16132 12152 16160 12183
rect 15988 12124 16160 12152
rect 16406 12152 16434 12183
rect 16850 12180 16856 12232
rect 16908 12220 16914 12232
rect 17681 12223 17739 12229
rect 17681 12220 17693 12223
rect 16908 12192 17693 12220
rect 16908 12180 16914 12192
rect 17681 12189 17693 12192
rect 17727 12189 17739 12223
rect 17681 12183 17739 12189
rect 17865 12223 17923 12229
rect 17865 12189 17877 12223
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 16758 12152 16764 12164
rect 16406 12124 16764 12152
rect 15988 12112 15994 12124
rect 16758 12112 16764 12124
rect 16816 12152 16822 12164
rect 16942 12152 16948 12164
rect 16816 12124 16948 12152
rect 16816 12112 16822 12124
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 17880 12152 17908 12183
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 18104 12192 18337 12220
rect 18104 12180 18110 12192
rect 18325 12189 18337 12192
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 18598 12180 18604 12232
rect 18656 12220 18662 12232
rect 18693 12223 18751 12229
rect 18693 12220 18705 12223
rect 18656 12192 18705 12220
rect 18656 12180 18662 12192
rect 18693 12189 18705 12192
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 19613 12223 19671 12229
rect 19613 12189 19625 12223
rect 19659 12220 19671 12223
rect 19702 12220 19708 12232
rect 19659 12192 19708 12220
rect 19659 12189 19671 12192
rect 19613 12183 19671 12189
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12189 19855 12223
rect 19797 12183 19855 12189
rect 17512 12124 17908 12152
rect 12176 12056 12664 12084
rect 12986 12044 12992 12096
rect 13044 12044 13050 12096
rect 13078 12044 13084 12096
rect 13136 12084 13142 12096
rect 17512 12093 17540 12124
rect 16025 12087 16083 12093
rect 16025 12084 16037 12087
rect 13136 12056 16037 12084
rect 13136 12044 13142 12056
rect 16025 12053 16037 12056
rect 16071 12053 16083 12087
rect 16025 12047 16083 12053
rect 17497 12087 17555 12093
rect 17497 12053 17509 12087
rect 17543 12053 17555 12087
rect 17497 12047 17555 12053
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12084 18015 12087
rect 18322 12084 18328 12096
rect 18003 12056 18328 12084
rect 18003 12053 18015 12056
rect 17957 12047 18015 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 18506 12044 18512 12096
rect 18564 12084 18570 12096
rect 18874 12084 18880 12096
rect 18564 12056 18880 12084
rect 18564 12044 18570 12056
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 19242 12044 19248 12096
rect 19300 12084 19306 12096
rect 19812 12084 19840 12183
rect 20254 12180 20260 12232
rect 20312 12180 20318 12232
rect 19300 12056 19840 12084
rect 19300 12044 19306 12056
rect 1104 11994 21043 12016
rect 1104 11942 5894 11994
rect 5946 11942 5958 11994
rect 6010 11942 6022 11994
rect 6074 11942 6086 11994
rect 6138 11942 6150 11994
rect 6202 11942 10839 11994
rect 10891 11942 10903 11994
rect 10955 11942 10967 11994
rect 11019 11942 11031 11994
rect 11083 11942 11095 11994
rect 11147 11942 15784 11994
rect 15836 11942 15848 11994
rect 15900 11942 15912 11994
rect 15964 11942 15976 11994
rect 16028 11942 16040 11994
rect 16092 11942 20729 11994
rect 20781 11942 20793 11994
rect 20845 11942 20857 11994
rect 20909 11942 20921 11994
rect 20973 11942 20985 11994
rect 21037 11942 21043 11994
rect 1104 11920 21043 11942
rect 842 11840 848 11892
rect 900 11880 906 11892
rect 1581 11883 1639 11889
rect 1581 11880 1593 11883
rect 900 11852 1593 11880
rect 900 11840 906 11852
rect 1581 11849 1593 11852
rect 1627 11849 1639 11883
rect 1581 11843 1639 11849
rect 3053 11883 3111 11889
rect 3053 11849 3065 11883
rect 3099 11880 3111 11883
rect 3878 11880 3884 11892
rect 3099 11852 3884 11880
rect 3099 11849 3111 11852
rect 3053 11843 3111 11849
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 4948 11852 5210 11880
rect 4948 11840 4954 11852
rect 1026 11772 1032 11824
rect 1084 11812 1090 11824
rect 2590 11812 2596 11824
rect 1084 11784 2596 11812
rect 1084 11772 1090 11784
rect 2590 11772 2596 11784
rect 2648 11772 2654 11824
rect 2866 11772 2872 11824
rect 2924 11812 2930 11824
rect 2924 11784 3556 11812
rect 2924 11772 2930 11784
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1946 11744 1952 11756
rect 1535 11716 1952 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1946 11704 1952 11716
rect 2004 11704 2010 11756
rect 2314 11753 2320 11756
rect 2283 11747 2320 11753
rect 2283 11713 2295 11747
rect 2372 11744 2378 11756
rect 3234 11744 3240 11756
rect 2372 11716 3240 11744
rect 2283 11707 2320 11713
rect 2314 11704 2320 11707
rect 2372 11704 2378 11716
rect 3234 11704 3240 11716
rect 3292 11704 3298 11756
rect 2038 11636 2044 11688
rect 2096 11636 2102 11688
rect 3326 11636 3332 11688
rect 3384 11676 3390 11688
rect 3421 11679 3479 11685
rect 3421 11676 3433 11679
rect 3384 11648 3433 11676
rect 3384 11636 3390 11648
rect 3421 11645 3433 11648
rect 3467 11645 3479 11679
rect 3528 11676 3556 11784
rect 3602 11704 3608 11756
rect 3660 11704 3666 11756
rect 4522 11753 4528 11756
rect 4479 11747 4528 11753
rect 4479 11713 4491 11747
rect 4525 11713 4528 11747
rect 4479 11707 4528 11713
rect 4522 11704 4528 11707
rect 4580 11704 4586 11756
rect 4617 11747 4675 11753
rect 4617 11713 4629 11747
rect 4663 11713 4675 11747
rect 4617 11707 4675 11713
rect 4154 11676 4160 11688
rect 3528 11648 4160 11676
rect 3421 11639 3479 11645
rect 4154 11636 4160 11648
rect 4212 11676 4218 11688
rect 4341 11679 4399 11685
rect 4341 11676 4353 11679
rect 4212 11648 4353 11676
rect 4212 11636 4218 11648
rect 4341 11645 4353 11648
rect 4387 11645 4399 11679
rect 4632 11676 4660 11707
rect 4632 11648 5026 11676
rect 4341 11639 4399 11645
rect 3510 11568 3516 11620
rect 3568 11608 3574 11620
rect 3878 11608 3884 11620
rect 3568 11580 3884 11608
rect 3568 11568 3574 11580
rect 3878 11568 3884 11580
rect 3936 11568 3942 11620
rect 4062 11568 4068 11620
rect 4120 11568 4126 11620
rect 4998 11608 5026 11648
rect 5182 11608 5210 11852
rect 5350 11840 5356 11892
rect 5408 11840 5414 11892
rect 5534 11840 5540 11892
rect 5592 11840 5598 11892
rect 5626 11840 5632 11892
rect 5684 11880 5690 11892
rect 6089 11883 6147 11889
rect 6089 11880 6101 11883
rect 5684 11852 6101 11880
rect 5684 11840 5690 11852
rect 6089 11849 6101 11852
rect 6135 11849 6147 11883
rect 6822 11880 6828 11892
rect 6089 11843 6147 11849
rect 6196 11852 6828 11880
rect 5368 11812 5396 11840
rect 6196 11812 6224 11852
rect 6822 11840 6828 11852
rect 6880 11840 6886 11892
rect 7006 11840 7012 11892
rect 7064 11880 7070 11892
rect 9585 11883 9643 11889
rect 9585 11880 9597 11883
rect 7064 11852 9597 11880
rect 7064 11840 7070 11852
rect 9585 11849 9597 11852
rect 9631 11849 9643 11883
rect 9585 11843 9643 11849
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10226 11880 10232 11892
rect 9815 11852 10232 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10226 11840 10232 11852
rect 10284 11840 10290 11892
rect 10686 11840 10692 11892
rect 10744 11880 10750 11892
rect 10965 11883 11023 11889
rect 10965 11880 10977 11883
rect 10744 11852 10977 11880
rect 10744 11840 10750 11852
rect 10965 11849 10977 11852
rect 11011 11849 11023 11883
rect 10965 11843 11023 11849
rect 12250 11840 12256 11892
rect 12308 11880 12314 11892
rect 14737 11883 14795 11889
rect 14737 11880 14749 11883
rect 12308 11852 14749 11880
rect 12308 11840 12314 11852
rect 14737 11849 14749 11852
rect 14783 11849 14795 11883
rect 14737 11843 14795 11849
rect 15378 11840 15384 11892
rect 15436 11840 15442 11892
rect 15562 11840 15568 11892
rect 15620 11880 15626 11892
rect 16117 11883 16175 11889
rect 16117 11880 16129 11883
rect 15620 11852 16129 11880
rect 15620 11840 15626 11852
rect 16117 11849 16129 11852
rect 16163 11849 16175 11883
rect 18509 11883 18567 11889
rect 16117 11843 16175 11849
rect 16546 11852 18092 11880
rect 5368 11784 6224 11812
rect 8481 11815 8539 11821
rect 8481 11781 8493 11815
rect 8527 11812 8539 11815
rect 8662 11812 8668 11824
rect 8527 11784 8668 11812
rect 8527 11781 8539 11784
rect 8481 11775 8539 11781
rect 8662 11772 8668 11784
rect 8720 11772 8726 11824
rect 8757 11815 8815 11821
rect 8757 11781 8769 11815
rect 8803 11781 8815 11815
rect 8757 11775 8815 11781
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5408 11716 5457 11744
rect 5408 11704 5414 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5445 11707 5503 11713
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 5997 11747 6055 11753
rect 5997 11744 6009 11747
rect 5592 11716 6009 11744
rect 5592 11704 5598 11716
rect 5997 11713 6009 11716
rect 6043 11744 6055 11747
rect 6086 11744 6092 11756
rect 6043 11716 6092 11744
rect 6043 11713 6055 11716
rect 5997 11707 6055 11713
rect 6086 11704 6092 11716
rect 6144 11704 6150 11756
rect 6178 11704 6184 11756
rect 6236 11704 6242 11756
rect 7374 11704 7380 11756
rect 7432 11753 7438 11756
rect 7432 11747 7460 11753
rect 7448 11713 7460 11747
rect 8772 11744 8800 11775
rect 8846 11772 8852 11824
rect 8904 11772 8910 11824
rect 9398 11772 9404 11824
rect 9456 11812 9462 11824
rect 12158 11812 12164 11824
rect 9456 11784 12164 11812
rect 9456 11772 9462 11784
rect 12158 11772 12164 11784
rect 12216 11812 12222 11824
rect 12216 11784 12480 11812
rect 12216 11772 12222 11784
rect 12452 11778 12480 11784
rect 9030 11744 9036 11756
rect 8772 11716 9036 11744
rect 7432 11707 7460 11713
rect 7432 11704 7438 11707
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9214 11704 9220 11756
rect 9272 11704 9278 11756
rect 10227 11747 10285 11753
rect 10227 11713 10239 11747
rect 10273 11744 10285 11747
rect 11606 11744 11612 11756
rect 10273 11716 11612 11744
rect 10273 11713 10285 11716
rect 10227 11707 10285 11713
rect 11606 11704 11612 11716
rect 11664 11704 11670 11756
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12250 11744 12256 11756
rect 11940 11716 12256 11744
rect 11940 11704 11946 11716
rect 12250 11704 12256 11716
rect 12308 11704 12314 11756
rect 12452 11750 12572 11778
rect 12894 11772 12900 11824
rect 12952 11812 12958 11824
rect 15396 11812 15424 11840
rect 16298 11812 16304 11824
rect 12952 11784 13860 11812
rect 15396 11784 16304 11812
rect 12952 11772 12958 11784
rect 12544 11744 12572 11750
rect 12603 11747 12661 11753
rect 12603 11744 12615 11747
rect 12544 11716 12615 11744
rect 12603 11713 12615 11716
rect 12649 11713 12661 11747
rect 12603 11707 12661 11713
rect 13262 11704 13268 11756
rect 13320 11744 13326 11756
rect 13722 11744 13728 11756
rect 13320 11716 13728 11744
rect 13320 11704 13326 11716
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 13832 11744 13860 11784
rect 16298 11772 16304 11784
rect 16356 11772 16362 11824
rect 13999 11747 14057 11753
rect 13999 11744 14011 11747
rect 13832 11716 14011 11744
rect 13999 11713 14011 11716
rect 14045 11744 14057 11747
rect 14090 11744 14096 11756
rect 14045 11716 14096 11744
rect 14045 11713 14057 11716
rect 13999 11707 14057 11713
rect 14090 11704 14096 11716
rect 14148 11704 14154 11756
rect 14826 11744 14832 11756
rect 14384 11716 14832 11744
rect 5718 11636 5724 11688
rect 5776 11676 5782 11688
rect 6196 11676 6224 11704
rect 5776 11648 6224 11676
rect 5776 11636 5782 11648
rect 6362 11636 6368 11688
rect 6420 11636 6426 11688
rect 6549 11679 6607 11685
rect 6549 11645 6561 11679
rect 6595 11645 6607 11679
rect 7285 11679 7343 11685
rect 7285 11676 7297 11679
rect 6549 11639 6607 11645
rect 6932 11648 7297 11676
rect 4998 11580 5210 11608
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 5810 11608 5816 11620
rect 5500 11580 5816 11608
rect 5500 11568 5506 11580
rect 5810 11568 5816 11580
rect 5868 11568 5874 11620
rect 5902 11568 5908 11620
rect 5960 11608 5966 11620
rect 6270 11608 6276 11620
rect 5960 11580 6276 11608
rect 5960 11568 5966 11580
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 6564 11608 6592 11639
rect 6932 11620 6960 11648
rect 7285 11645 7297 11648
rect 7331 11645 7343 11679
rect 7285 11639 7343 11645
rect 7558 11636 7564 11688
rect 7616 11636 7622 11688
rect 7742 11636 7748 11688
rect 7800 11676 7806 11688
rect 9953 11679 10011 11685
rect 7800 11648 8326 11676
rect 7800 11636 7806 11648
rect 9953 11645 9965 11679
rect 9999 11645 10011 11679
rect 9953 11639 10011 11645
rect 6822 11608 6828 11620
rect 6564 11580 6828 11608
rect 6822 11568 6828 11580
rect 6880 11568 6886 11620
rect 6914 11568 6920 11620
rect 6972 11568 6978 11620
rect 7009 11611 7067 11617
rect 7009 11577 7021 11611
rect 7055 11608 7067 11611
rect 7098 11608 7104 11620
rect 7055 11580 7104 11608
rect 7055 11577 7067 11580
rect 7009 11571 7067 11577
rect 7098 11568 7104 11580
rect 7156 11568 7162 11620
rect 2130 11500 2136 11552
rect 2188 11540 2194 11552
rect 3142 11540 3148 11552
rect 2188 11512 3148 11540
rect 2188 11500 2194 11512
rect 3142 11500 3148 11512
rect 3200 11500 3206 11552
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 5261 11543 5319 11549
rect 5261 11540 5273 11543
rect 3292 11512 5273 11540
rect 3292 11500 3298 11512
rect 5261 11509 5273 11512
rect 5307 11509 5319 11543
rect 5261 11503 5319 11509
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 8205 11543 8263 11549
rect 8205 11540 8217 11543
rect 5684 11512 8217 11540
rect 5684 11500 5690 11512
rect 8205 11509 8217 11512
rect 8251 11509 8263 11543
rect 9968 11540 9996 11639
rect 11422 11636 11428 11688
rect 11480 11636 11486 11688
rect 12268 11676 12296 11704
rect 12345 11679 12403 11685
rect 12345 11676 12357 11679
rect 12268 11648 12357 11676
rect 12345 11645 12357 11648
rect 12391 11645 12403 11679
rect 12345 11639 12403 11645
rect 11440 11608 11468 11636
rect 10610 11580 11468 11608
rect 10226 11540 10232 11552
rect 9968 11512 10232 11540
rect 8205 11503 8263 11509
rect 10226 11500 10232 11512
rect 10284 11540 10290 11552
rect 10610 11540 10638 11580
rect 10284 11512 10638 11540
rect 10284 11500 10290 11512
rect 12710 11500 12716 11552
rect 12768 11540 12774 11552
rect 13357 11543 13415 11549
rect 13357 11540 13369 11543
rect 12768 11512 13369 11540
rect 12768 11500 12774 11512
rect 13357 11509 13369 11512
rect 13403 11509 13415 11543
rect 13357 11503 13415 11509
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 14384 11540 14412 11716
rect 14826 11704 14832 11716
rect 14884 11744 14890 11756
rect 15347 11747 15405 11753
rect 15347 11744 15359 11747
rect 14884 11716 15359 11744
rect 14884 11704 14890 11716
rect 15347 11713 15359 11716
rect 15393 11713 15405 11747
rect 15347 11707 15405 11713
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 16546 11744 16574 11852
rect 18064 11812 18092 11852
rect 18509 11849 18521 11883
rect 18555 11880 18567 11883
rect 18782 11880 18788 11892
rect 18555 11852 18788 11880
rect 18555 11849 18567 11852
rect 18509 11843 18567 11849
rect 18782 11840 18788 11852
rect 18840 11840 18846 11892
rect 19981 11883 20039 11889
rect 19981 11849 19993 11883
rect 20027 11880 20039 11883
rect 20530 11880 20536 11892
rect 20027 11852 20536 11880
rect 20027 11849 20039 11852
rect 19981 11843 20039 11849
rect 20530 11840 20536 11852
rect 20588 11840 20594 11892
rect 18868 11815 18926 11821
rect 18868 11812 18880 11815
rect 16776 11784 17540 11812
rect 18064 11784 18880 11812
rect 15528 11716 16574 11744
rect 15528 11704 15534 11716
rect 16666 11704 16672 11756
rect 16724 11744 16730 11756
rect 16776 11753 16804 11784
rect 17512 11756 17540 11784
rect 18868 11781 18880 11784
rect 18914 11781 18926 11815
rect 18868 11775 18926 11781
rect 19794 11772 19800 11824
rect 19852 11812 19858 11824
rect 20165 11815 20223 11821
rect 20165 11812 20177 11815
rect 19852 11784 20177 11812
rect 19852 11772 19858 11784
rect 20165 11781 20177 11784
rect 20211 11781 20223 11815
rect 20165 11775 20223 11781
rect 16761 11747 16819 11753
rect 16761 11744 16773 11747
rect 16724 11716 16773 11744
rect 16724 11704 16730 11716
rect 16761 11713 16773 11716
rect 16807 11713 16819 11747
rect 16761 11707 16819 11713
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17017 11747 17075 11753
rect 17017 11744 17029 11747
rect 16908 11716 17029 11744
rect 16908 11704 16914 11716
rect 17017 11713 17029 11716
rect 17063 11713 17075 11747
rect 17017 11707 17075 11713
rect 17494 11704 17500 11756
rect 17552 11744 17558 11756
rect 17552 11716 17816 11744
rect 17552 11704 17558 11716
rect 15102 11636 15108 11688
rect 15160 11636 15166 11688
rect 17788 11676 17816 11716
rect 18230 11704 18236 11756
rect 18288 11704 18294 11756
rect 18322 11704 18328 11756
rect 18380 11704 18386 11756
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 18432 11716 18613 11744
rect 18432 11676 18460 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 17788 11648 18460 11676
rect 18506 11636 18512 11688
rect 18564 11636 18570 11688
rect 13872 11512 14412 11540
rect 13872 11500 13878 11512
rect 14458 11500 14464 11552
rect 14516 11540 14522 11552
rect 17494 11540 17500 11552
rect 14516 11512 17500 11540
rect 14516 11500 14522 11512
rect 17494 11500 17500 11512
rect 17552 11500 17558 11552
rect 18138 11500 18144 11552
rect 18196 11500 18202 11552
rect 20441 11543 20499 11549
rect 20441 11509 20453 11543
rect 20487 11540 20499 11543
rect 21266 11540 21272 11552
rect 20487 11512 21272 11540
rect 20487 11509 20499 11512
rect 20441 11503 20499 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 1104 11450 20884 11472
rect 14 11364 20 11416
rect 72 11404 78 11416
rect 566 11404 572 11416
rect 72 11376 572 11404
rect 72 11364 78 11376
rect 566 11364 572 11376
rect 624 11364 630 11416
rect 1104 11398 3422 11450
rect 3474 11398 3486 11450
rect 3538 11398 3550 11450
rect 3602 11398 3614 11450
rect 3666 11398 3678 11450
rect 3730 11398 8367 11450
rect 8419 11398 8431 11450
rect 8483 11398 8495 11450
rect 8547 11398 8559 11450
rect 8611 11398 8623 11450
rect 8675 11398 13312 11450
rect 13364 11398 13376 11450
rect 13428 11398 13440 11450
rect 13492 11398 13504 11450
rect 13556 11398 13568 11450
rect 13620 11398 18257 11450
rect 18309 11398 18321 11450
rect 18373 11398 18385 11450
rect 18437 11398 18449 11450
rect 18501 11398 18513 11450
rect 18565 11398 20884 11450
rect 1104 11376 20884 11398
rect 1670 11296 1676 11348
rect 1728 11296 1734 11348
rect 3234 11336 3240 11348
rect 1780 11308 3240 11336
rect 474 11228 480 11280
rect 532 11268 538 11280
rect 1780 11268 1808 11308
rect 3234 11296 3240 11308
rect 3292 11296 3298 11348
rect 3329 11339 3387 11345
rect 3329 11305 3341 11339
rect 3375 11336 3387 11339
rect 4062 11336 4068 11348
rect 3375 11308 4068 11336
rect 3375 11305 3387 11308
rect 3329 11299 3387 11305
rect 4062 11296 4068 11308
rect 4120 11296 4126 11348
rect 4522 11296 4528 11348
rect 4580 11296 4586 11348
rect 4706 11296 4712 11348
rect 4764 11336 4770 11348
rect 5629 11339 5687 11345
rect 5629 11336 5641 11339
rect 4764 11308 5641 11336
rect 4764 11296 4770 11308
rect 5629 11305 5641 11308
rect 5675 11305 5687 11339
rect 5629 11299 5687 11305
rect 5736 11308 6592 11336
rect 2130 11268 2136 11280
rect 532 11240 1808 11268
rect 1964 11240 2136 11268
rect 532 11228 538 11240
rect 1964 11132 1992 11240
rect 2130 11228 2136 11240
rect 2188 11228 2194 11280
rect 3510 11228 3516 11280
rect 3568 11268 3574 11280
rect 4540 11268 4568 11296
rect 5736 11268 5764 11308
rect 6564 11280 6592 11308
rect 6638 11296 6644 11348
rect 6696 11336 6702 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6696 11308 6745 11336
rect 6696 11296 6702 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 9858 11296 9864 11348
rect 9916 11296 9922 11348
rect 10781 11339 10839 11345
rect 10781 11305 10793 11339
rect 10827 11336 10839 11339
rect 11330 11336 11336 11348
rect 10827 11308 11336 11336
rect 10827 11305 10839 11308
rect 10781 11299 10839 11305
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 12250 11296 12256 11348
rect 12308 11296 12314 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 12492 11308 13185 11336
rect 12492 11296 12498 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 13173 11299 13231 11305
rect 13722 11296 13728 11348
rect 13780 11336 13786 11348
rect 15105 11339 15163 11345
rect 15105 11336 15117 11339
rect 13780 11308 15117 11336
rect 13780 11296 13786 11308
rect 15105 11305 15117 11308
rect 15151 11305 15163 11339
rect 15105 11299 15163 11305
rect 15286 11296 15292 11348
rect 15344 11336 15350 11348
rect 15344 11308 17080 11336
rect 15344 11296 15350 11308
rect 3568 11240 4568 11268
rect 5570 11240 5764 11268
rect 3568 11228 3574 11240
rect 2038 11160 2044 11212
rect 2096 11200 2102 11212
rect 2314 11200 2320 11212
rect 2096 11172 2320 11200
rect 2096 11160 2102 11172
rect 2314 11160 2320 11172
rect 2372 11160 2378 11212
rect 3970 11160 3976 11212
rect 4028 11160 4034 11212
rect 4430 11160 4436 11212
rect 4488 11160 4494 11212
rect 4706 11160 4712 11212
rect 4764 11160 4770 11212
rect 4847 11203 4905 11209
rect 4847 11169 4859 11203
rect 4893 11200 4905 11203
rect 5166 11200 5172 11212
rect 4893 11172 5172 11200
rect 4893 11169 4905 11172
rect 4847 11163 4905 11169
rect 5166 11160 5172 11172
rect 5224 11160 5230 11212
rect 2225 11135 2283 11141
rect 2225 11132 2237 11135
rect 1964 11104 2237 11132
rect 2225 11101 2237 11104
rect 2271 11101 2283 11135
rect 2225 11095 2283 11101
rect 2498 11092 2504 11144
rect 2556 11132 2562 11144
rect 2591 11135 2649 11141
rect 2591 11132 2603 11135
rect 2556 11104 2603 11132
rect 2556 11092 2562 11104
rect 2591 11101 2603 11104
rect 2637 11132 2649 11135
rect 2958 11132 2964 11144
rect 2637 11104 2964 11132
rect 2637 11101 2649 11104
rect 2591 11095 2649 11101
rect 2958 11092 2964 11104
rect 3016 11092 3022 11144
rect 3326 11092 3332 11144
rect 3384 11132 3390 11144
rect 3789 11135 3847 11141
rect 3789 11132 3801 11135
rect 3384 11104 3801 11132
rect 3384 11092 3390 11104
rect 3789 11101 3801 11104
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 1581 11067 1639 11073
rect 1581 11033 1593 11067
rect 1627 11064 1639 11067
rect 3602 11064 3608 11076
rect 1627 11036 3608 11064
rect 1627 11033 1639 11036
rect 1581 11027 1639 11033
rect 3602 11024 3608 11036
rect 3660 11024 3666 11076
rect 2038 10956 2044 11008
rect 2096 10956 2102 11008
rect 2130 10956 2136 11008
rect 2188 10996 2194 11008
rect 2406 10996 2412 11008
rect 2188 10968 2412 10996
rect 2188 10956 2194 10968
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 3988 10996 4016 11160
rect 5570 11144 5598 11240
rect 6546 11228 6552 11280
rect 6604 11228 6610 11280
rect 6914 11228 6920 11280
rect 6972 11268 6978 11280
rect 7374 11268 7380 11280
rect 6972 11240 7380 11268
rect 6972 11228 6978 11240
rect 7374 11228 7380 11240
rect 7432 11228 7438 11280
rect 7466 11228 7472 11280
rect 7524 11228 7530 11280
rect 9876 11268 9904 11296
rect 8772 11240 9904 11268
rect 7484 11200 7512 11228
rect 6346 11172 7512 11200
rect 4982 11092 4988 11144
rect 5040 11092 5046 11144
rect 5552 11092 5558 11144
rect 5610 11092 5616 11144
rect 5721 11135 5779 11141
rect 5721 11101 5733 11135
rect 5767 11101 5779 11135
rect 5995 11135 6053 11141
rect 5995 11132 6007 11135
rect 5721 11095 5779 11101
rect 5828 11104 6007 11132
rect 3292 10968 4016 10996
rect 3292 10956 3298 10968
rect 4614 10956 4620 11008
rect 4672 10996 4678 11008
rect 5736 10996 5764 11095
rect 5828 11008 5856 11104
rect 5995 11101 6007 11104
rect 6041 11101 6053 11135
rect 6346 11132 6374 11172
rect 5995 11095 6053 11101
rect 6196 11104 6374 11132
rect 6196 11064 6224 11104
rect 6638 11092 6644 11144
rect 6696 11132 6702 11144
rect 7466 11132 7472 11144
rect 6696 11104 7472 11132
rect 6696 11092 6702 11104
rect 7466 11092 7472 11104
rect 7524 11092 7530 11144
rect 7743 11135 7801 11141
rect 7743 11101 7755 11135
rect 7789 11132 7801 11135
rect 8110 11132 8116 11144
rect 7789 11104 8116 11132
rect 7789 11101 7801 11104
rect 7743 11095 7801 11101
rect 8110 11092 8116 11104
rect 8168 11132 8174 11144
rect 8772 11132 8800 11240
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 12066 11268 12072 11280
rect 10744 11240 12072 11268
rect 10744 11228 10750 11240
rect 12066 11228 12072 11240
rect 12124 11228 12130 11280
rect 12268 11268 12296 11296
rect 12176 11240 12296 11268
rect 9582 11160 9588 11212
rect 9640 11160 9646 11212
rect 11514 11160 11520 11212
rect 11572 11200 11578 11212
rect 12176 11209 12204 11240
rect 13078 11228 13084 11280
rect 13136 11268 13142 11280
rect 14090 11268 14096 11280
rect 13136 11240 14096 11268
rect 13136 11228 13142 11240
rect 14090 11228 14096 11240
rect 14148 11228 14154 11280
rect 14826 11228 14832 11280
rect 14884 11268 14890 11280
rect 15010 11268 15016 11280
rect 14884 11240 15016 11268
rect 14884 11228 14890 11240
rect 15010 11228 15016 11240
rect 15068 11228 15074 11280
rect 17052 11268 17080 11308
rect 17126 11296 17132 11348
rect 17184 11296 17190 11348
rect 17420 11308 18000 11336
rect 17420 11268 17448 11308
rect 17052 11240 17448 11268
rect 17972 11268 18000 11308
rect 18046 11296 18052 11348
rect 18104 11336 18110 11348
rect 18325 11339 18383 11345
rect 18325 11336 18337 11339
rect 18104 11308 18337 11336
rect 18104 11296 18110 11308
rect 18325 11305 18337 11308
rect 18371 11305 18383 11339
rect 18325 11299 18383 11305
rect 18690 11296 18696 11348
rect 18748 11296 18754 11348
rect 20070 11296 20076 11348
rect 20128 11336 20134 11348
rect 20257 11339 20315 11345
rect 20257 11336 20269 11339
rect 20128 11308 20269 11336
rect 20128 11296 20134 11308
rect 20257 11305 20269 11308
rect 20303 11305 20315 11339
rect 20257 11299 20315 11305
rect 18782 11268 18788 11280
rect 17972 11240 18788 11268
rect 18782 11228 18788 11240
rect 18840 11228 18846 11280
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 11572 11172 12173 11200
rect 11572 11160 11578 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 19150 11200 19156 11212
rect 12161 11163 12219 11169
rect 17926 11172 19156 11200
rect 8168 11104 8800 11132
rect 8168 11092 8174 11104
rect 9214 11092 9220 11144
rect 9272 11132 9278 11144
rect 9398 11132 9404 11144
rect 9272 11104 9404 11132
rect 9272 11092 9278 11104
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 9600 11132 9628 11160
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9600 11104 9689 11132
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9677 11095 9735 11101
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 10043 11135 10101 11141
rect 10043 11101 10055 11135
rect 10089 11132 10101 11135
rect 11054 11132 11060 11144
rect 10089 11104 11060 11132
rect 10089 11101 10101 11104
rect 10043 11095 10101 11101
rect 5920 11036 6224 11064
rect 5920 11008 5948 11036
rect 8386 11024 8392 11076
rect 8444 11064 8450 11076
rect 9784 11064 9812 11095
rect 11054 11092 11060 11104
rect 11112 11092 11118 11144
rect 11330 11092 11336 11144
rect 11388 11132 11394 11144
rect 11606 11132 11612 11144
rect 11388 11104 11612 11132
rect 11388 11092 11394 11104
rect 11606 11092 11612 11104
rect 11664 11132 11670 11144
rect 12435 11135 12493 11141
rect 12435 11132 12447 11135
rect 11664 11104 12447 11132
rect 11664 11092 11670 11104
rect 12435 11101 12447 11104
rect 12481 11132 12493 11135
rect 13906 11132 13912 11144
rect 12481 11104 13912 11132
rect 12481 11101 12493 11104
rect 12435 11095 12493 11101
rect 13906 11092 13912 11104
rect 13964 11092 13970 11144
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11101 14151 11135
rect 14366 11132 14372 11144
rect 14327 11104 14372 11132
rect 14093 11095 14151 11101
rect 10226 11064 10232 11076
rect 8444 11036 9628 11064
rect 9784 11036 10232 11064
rect 8444 11024 8450 11036
rect 4672 10968 5764 10996
rect 4672 10956 4678 10968
rect 5810 10956 5816 11008
rect 5868 10956 5874 11008
rect 5902 10956 5908 11008
rect 5960 10956 5966 11008
rect 5994 10956 6000 11008
rect 6052 10996 6058 11008
rect 6362 10996 6368 11008
rect 6052 10968 6368 10996
rect 6052 10956 6058 10968
rect 6362 10956 6368 10968
rect 6420 10956 6426 11008
rect 8018 10956 8024 11008
rect 8076 10996 8082 11008
rect 8294 10996 8300 11008
rect 8076 10968 8300 10996
rect 8076 10956 8082 10968
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 8481 10999 8539 11005
rect 8481 10965 8493 10999
rect 8527 10996 8539 10999
rect 9398 10996 9404 11008
rect 8527 10968 9404 10996
rect 8527 10965 8539 10968
rect 8481 10959 8539 10965
rect 9398 10956 9404 10968
rect 9456 10956 9462 11008
rect 9490 10956 9496 11008
rect 9548 10956 9554 11008
rect 9600 10996 9628 11036
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 14108 11064 14136 11095
rect 14366 11092 14372 11104
rect 14424 11092 14430 11144
rect 15473 11135 15531 11141
rect 15473 11101 15485 11135
rect 15519 11132 15531 11135
rect 15519 11104 15608 11132
rect 15519 11101 15531 11104
rect 15473 11095 15531 11101
rect 15580 11076 15608 11104
rect 15654 11092 15660 11144
rect 15712 11132 15718 11144
rect 15747 11135 15805 11141
rect 15747 11132 15759 11135
rect 15712 11104 15759 11132
rect 15712 11092 15718 11104
rect 15747 11101 15759 11104
rect 15793 11132 15805 11135
rect 16758 11132 16764 11144
rect 15793 11104 16764 11132
rect 15793 11101 15805 11104
rect 15747 11095 15805 11101
rect 16758 11092 16764 11104
rect 16816 11092 16822 11144
rect 17313 11135 17371 11141
rect 17313 11101 17325 11135
rect 17359 11132 17371 11135
rect 17359 11104 17448 11132
rect 17359 11101 17371 11104
rect 17313 11095 17371 11101
rect 17420 11076 17448 11104
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 17587 11135 17645 11141
rect 17587 11132 17599 11135
rect 17552 11104 17599 11132
rect 17552 11092 17558 11104
rect 17587 11101 17599 11104
rect 17633 11101 17645 11135
rect 17926 11132 17954 11172
rect 19150 11160 19156 11172
rect 19208 11200 19214 11212
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 19208 11172 19257 11200
rect 19208 11160 19214 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 19245 11163 19303 11169
rect 17587 11095 17645 11101
rect 17696 11104 17954 11132
rect 10560 11036 13814 11064
rect 14108 11036 15148 11064
rect 10560 11024 10566 11036
rect 11790 10996 11796 11008
rect 9600 10968 11796 10996
rect 11790 10956 11796 10968
rect 11848 10956 11854 11008
rect 12250 10956 12256 11008
rect 12308 10996 12314 11008
rect 12986 10996 12992 11008
rect 12308 10968 12992 10996
rect 12308 10956 12314 10968
rect 12986 10956 12992 10968
rect 13044 10956 13050 11008
rect 13786 10996 13814 11036
rect 15120 11008 15148 11036
rect 15562 11024 15568 11076
rect 15620 11024 15626 11076
rect 16114 11024 16120 11076
rect 16172 11064 16178 11076
rect 17037 11067 17095 11073
rect 16172 11036 16528 11064
rect 16172 11024 16178 11036
rect 13906 10996 13912 11008
rect 13786 10968 13912 10996
rect 13906 10956 13912 10968
rect 13964 10996 13970 11008
rect 14918 10996 14924 11008
rect 13964 10968 14924 10996
rect 13964 10956 13970 10968
rect 14918 10956 14924 10968
rect 14976 10956 14982 11008
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 16206 10996 16212 11008
rect 15160 10968 16212 10996
rect 15160 10956 15166 10968
rect 16206 10956 16212 10968
rect 16264 10956 16270 11008
rect 16500 11005 16528 11036
rect 17037 11033 17049 11067
rect 17083 11064 17095 11067
rect 17218 11064 17224 11076
rect 17083 11036 17224 11064
rect 17083 11033 17095 11036
rect 17037 11027 17095 11033
rect 17218 11024 17224 11036
rect 17276 11024 17282 11076
rect 17402 11024 17408 11076
rect 17460 11064 17466 11076
rect 17696 11064 17724 11104
rect 18874 11092 18880 11144
rect 18932 11092 18938 11144
rect 19487 11135 19545 11141
rect 19487 11101 19499 11135
rect 19533 11101 19545 11135
rect 19487 11095 19545 11101
rect 17460 11036 17724 11064
rect 17460 11024 17466 11036
rect 17770 11024 17776 11076
rect 17828 11064 17834 11076
rect 18598 11064 18604 11076
rect 17828 11036 18604 11064
rect 17828 11024 17834 11036
rect 18598 11024 18604 11036
rect 18656 11024 18662 11076
rect 18782 11024 18788 11076
rect 18840 11064 18846 11076
rect 19502 11064 19530 11095
rect 18840 11036 19530 11064
rect 18840 11024 18846 11036
rect 19610 11024 19616 11076
rect 19668 11064 19674 11076
rect 20070 11064 20076 11076
rect 19668 11036 20076 11064
rect 19668 11024 19674 11036
rect 20070 11024 20076 11036
rect 20128 11024 20134 11076
rect 16485 10999 16543 11005
rect 16485 10965 16497 10999
rect 16531 10965 16543 10999
rect 16485 10959 16543 10965
rect 17678 10956 17684 11008
rect 17736 10996 17742 11008
rect 19628 10996 19656 11024
rect 17736 10968 19656 10996
rect 17736 10956 17742 10968
rect 1104 10906 21043 10928
rect 1104 10854 5894 10906
rect 5946 10854 5958 10906
rect 6010 10854 6022 10906
rect 6074 10854 6086 10906
rect 6138 10854 6150 10906
rect 6202 10854 10839 10906
rect 10891 10854 10903 10906
rect 10955 10854 10967 10906
rect 11019 10854 11031 10906
rect 11083 10854 11095 10906
rect 11147 10854 15784 10906
rect 15836 10854 15848 10906
rect 15900 10854 15912 10906
rect 15964 10854 15976 10906
rect 16028 10854 16040 10906
rect 16092 10854 20729 10906
rect 20781 10854 20793 10906
rect 20845 10854 20857 10906
rect 20909 10854 20921 10906
rect 20973 10854 20985 10906
rect 21037 10854 21043 10906
rect 1104 10832 21043 10854
rect 1026 10752 1032 10804
rect 1084 10792 1090 10804
rect 1394 10792 1400 10804
rect 1084 10764 1400 10792
rect 1084 10752 1090 10764
rect 1394 10752 1400 10764
rect 1452 10752 1458 10804
rect 1578 10752 1584 10804
rect 1636 10752 1642 10804
rect 2498 10792 2504 10804
rect 1688 10764 2504 10792
rect 14 10684 20 10736
rect 72 10724 78 10736
rect 1688 10724 1716 10764
rect 2498 10752 2504 10764
rect 2556 10752 2562 10804
rect 3145 10795 3203 10801
rect 3145 10761 3157 10795
rect 3191 10792 3203 10795
rect 4430 10792 4436 10804
rect 3191 10764 4436 10792
rect 3191 10761 3203 10764
rect 3145 10755 3203 10761
rect 4430 10752 4436 10764
rect 4488 10752 4494 10804
rect 4525 10795 4583 10801
rect 4525 10761 4537 10795
rect 4571 10792 4583 10795
rect 4982 10792 4988 10804
rect 4571 10764 4988 10792
rect 4571 10761 4583 10764
rect 4525 10755 4583 10761
rect 4982 10752 4988 10764
rect 5040 10752 5046 10804
rect 5166 10752 5172 10804
rect 5224 10752 5230 10804
rect 5258 10752 5264 10804
rect 5316 10752 5322 10804
rect 5905 10795 5963 10801
rect 5905 10761 5917 10795
rect 5951 10792 5963 10795
rect 6914 10792 6920 10804
rect 5951 10764 6920 10792
rect 5951 10761 5963 10764
rect 5905 10755 5963 10761
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 7006 10752 7012 10804
rect 7064 10752 7070 10804
rect 7745 10795 7803 10801
rect 7745 10761 7757 10795
rect 7791 10792 7803 10795
rect 8846 10792 8852 10804
rect 7791 10764 8852 10792
rect 7791 10761 7803 10764
rect 7745 10755 7803 10761
rect 8846 10752 8852 10764
rect 8904 10752 8910 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 10042 10792 10048 10804
rect 9171 10764 10048 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 10134 10752 10140 10804
rect 10192 10792 10198 10804
rect 10410 10792 10416 10804
rect 10192 10764 10416 10792
rect 10192 10752 10198 10764
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 10505 10795 10563 10801
rect 10505 10761 10517 10795
rect 10551 10792 10563 10795
rect 10594 10792 10600 10804
rect 10551 10764 10600 10792
rect 10551 10761 10563 10764
rect 10505 10755 10563 10761
rect 10594 10752 10600 10764
rect 10652 10752 10658 10804
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 12342 10792 12348 10804
rect 11204 10764 12348 10792
rect 11204 10752 11210 10764
rect 12342 10752 12348 10764
rect 12400 10752 12406 10804
rect 12526 10752 12532 10804
rect 12584 10752 12590 10804
rect 14829 10795 14887 10801
rect 14829 10792 14841 10795
rect 12636 10764 14841 10792
rect 2222 10724 2228 10736
rect 72 10696 1716 10724
rect 2148 10696 2228 10724
rect 72 10684 78 10696
rect 1486 10616 1492 10668
rect 1544 10616 1550 10668
rect 2148 10665 2176 10696
rect 2222 10684 2228 10696
rect 2280 10684 2286 10736
rect 2866 10724 2872 10736
rect 2700 10696 2872 10724
rect 2391 10689 2449 10695
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10625 2191 10659
rect 2391 10655 2403 10689
rect 2437 10686 2449 10689
rect 2437 10656 2452 10686
rect 2700 10656 2728 10696
rect 2866 10684 2872 10696
rect 2924 10724 2930 10736
rect 4246 10724 4252 10736
rect 2924 10696 4252 10724
rect 2924 10684 2930 10696
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 4338 10684 4344 10736
rect 4396 10684 4402 10736
rect 4890 10684 4896 10736
rect 4948 10724 4954 10736
rect 5184 10724 5212 10752
rect 4948 10696 5212 10724
rect 5276 10724 5304 10752
rect 5276 10696 5948 10724
rect 4948 10684 4954 10696
rect 2437 10655 2728 10656
rect 2391 10649 2728 10655
rect 2424 10628 2728 10649
rect 2133 10619 2191 10625
rect 2148 10452 2176 10619
rect 2774 10616 2780 10668
rect 2832 10656 2838 10668
rect 3142 10656 3148 10668
rect 2832 10628 3148 10656
rect 2832 10616 2838 10628
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3755 10659 3813 10665
rect 3755 10656 3767 10659
rect 3200 10628 3767 10656
rect 3200 10616 3206 10628
rect 3755 10625 3767 10628
rect 3801 10625 3813 10659
rect 4356 10656 4384 10684
rect 5920 10668 5948 10696
rect 5994 10684 6000 10736
rect 6052 10724 6058 10736
rect 7024 10724 7052 10752
rect 6052 10696 6684 10724
rect 6052 10684 6058 10696
rect 6656 10668 6684 10696
rect 6748 10696 7052 10724
rect 5135 10659 5193 10665
rect 5135 10656 5147 10659
rect 4356 10628 5147 10656
rect 3755 10619 3813 10625
rect 5135 10625 5147 10628
rect 5181 10656 5193 10659
rect 5181 10628 5764 10656
rect 5181 10625 5193 10628
rect 5135 10619 5193 10625
rect 3510 10548 3516 10600
rect 3568 10548 3574 10600
rect 4798 10548 4804 10600
rect 4856 10548 4862 10600
rect 4893 10591 4951 10597
rect 4893 10557 4905 10591
rect 4939 10557 4951 10591
rect 4893 10551 4951 10557
rect 3528 10452 3556 10548
rect 2148 10424 3556 10452
rect 3602 10412 3608 10464
rect 3660 10452 3666 10464
rect 4816 10452 4844 10548
rect 3660 10424 4844 10452
rect 4908 10452 4936 10551
rect 5736 10520 5764 10628
rect 5902 10616 5908 10668
rect 5960 10616 5966 10668
rect 6362 10656 6368 10668
rect 6010 10628 6368 10656
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6010 10588 6038 10628
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 5868 10560 6038 10588
rect 5868 10548 5874 10560
rect 6178 10548 6184 10600
rect 6236 10588 6242 10600
rect 6748 10597 6776 10696
rect 8110 10684 8116 10736
rect 8168 10724 8174 10736
rect 8168 10696 8340 10724
rect 8168 10684 8174 10696
rect 8312 10686 8340 10696
rect 8386 10695 8392 10736
rect 8371 10689 8392 10695
rect 8371 10686 8383 10689
rect 6975 10659 7033 10665
rect 6975 10625 6987 10659
rect 7021 10656 7033 10659
rect 7021 10628 7420 10656
rect 7021 10625 7033 10628
rect 6975 10619 7033 10625
rect 6733 10591 6791 10597
rect 6733 10588 6745 10591
rect 6236 10560 6745 10588
rect 6236 10548 6242 10560
rect 6733 10557 6745 10560
rect 6779 10557 6791 10591
rect 7392 10588 7420 10628
rect 7466 10616 7472 10668
rect 7524 10656 7530 10668
rect 8312 10658 8383 10686
rect 8444 10684 8450 10736
rect 9306 10684 9312 10736
rect 9364 10724 9370 10736
rect 12636 10724 12664 10764
rect 14829 10761 14841 10764
rect 14875 10761 14887 10795
rect 14829 10755 14887 10761
rect 14918 10752 14924 10804
rect 14976 10792 14982 10804
rect 16298 10792 16304 10804
rect 14976 10764 16304 10792
rect 14976 10752 14982 10764
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 16390 10752 16396 10804
rect 16448 10752 16454 10804
rect 18874 10792 18880 10804
rect 16500 10764 18880 10792
rect 9364 10696 12664 10724
rect 9364 10684 9370 10696
rect 13170 10684 13176 10736
rect 13228 10684 13234 10736
rect 15378 10684 15384 10736
rect 15436 10684 15442 10736
rect 15930 10684 15936 10736
rect 15988 10724 15994 10736
rect 16408 10724 16436 10752
rect 15988 10696 16436 10724
rect 15988 10684 15994 10696
rect 7524 10628 8156 10656
rect 8371 10655 8383 10658
rect 8417 10658 8432 10684
rect 9735 10659 9793 10665
rect 8417 10655 8429 10658
rect 9735 10656 9747 10659
rect 8371 10649 8429 10655
rect 7524 10616 7530 10628
rect 8018 10588 8024 10600
rect 7392 10560 8024 10588
rect 6733 10551 6791 10557
rect 8018 10548 8024 10560
rect 8076 10548 8082 10600
rect 8128 10597 8156 10628
rect 9324 10628 9747 10656
rect 9324 10600 9352 10628
rect 9735 10625 9747 10628
rect 9781 10625 9793 10659
rect 9735 10619 9793 10625
rect 9858 10616 9864 10668
rect 9916 10656 9922 10668
rect 11759 10659 11817 10665
rect 11759 10656 11771 10659
rect 9916 10628 11771 10656
rect 9916 10616 9922 10628
rect 11759 10625 11771 10628
rect 11805 10625 11817 10659
rect 11759 10619 11817 10625
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12492 10628 13001 10656
rect 12492 10616 12498 10628
rect 12989 10625 13001 10628
rect 13035 10656 13047 10659
rect 13188 10656 13216 10684
rect 15195 10669 15253 10675
rect 15195 10668 15207 10669
rect 15241 10668 15253 10669
rect 13035 10628 13400 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10557 8171 10591
rect 8113 10551 8171 10557
rect 5736 10492 6868 10520
rect 5166 10452 5172 10464
rect 4908 10424 5172 10452
rect 3660 10412 3666 10424
rect 5166 10412 5172 10424
rect 5224 10452 5230 10464
rect 5994 10452 6000 10464
rect 5224 10424 6000 10452
rect 5224 10412 5230 10424
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6840 10452 6868 10492
rect 7466 10452 7472 10464
rect 6840 10424 7472 10452
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 8128 10452 8156 10551
rect 9306 10548 9312 10600
rect 9364 10548 9370 10600
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10557 9551 10591
rect 9493 10551 9551 10557
rect 8570 10452 8576 10464
rect 8128 10424 8576 10452
rect 8570 10412 8576 10424
rect 8628 10452 8634 10464
rect 9508 10452 9536 10551
rect 11514 10548 11520 10600
rect 11572 10548 11578 10600
rect 12894 10548 12900 10600
rect 12952 10548 12958 10600
rect 13170 10548 13176 10600
rect 13228 10548 13234 10600
rect 10318 10480 10324 10532
rect 10376 10520 10382 10532
rect 10962 10520 10968 10532
rect 10376 10492 10968 10520
rect 10376 10480 10382 10492
rect 10962 10480 10968 10492
rect 11020 10480 11026 10532
rect 8628 10424 9536 10452
rect 8628 10412 8634 10424
rect 9766 10412 9772 10464
rect 9824 10452 9830 10464
rect 12912 10452 12940 10548
rect 9824 10424 12940 10452
rect 13372 10452 13400 10628
rect 13906 10616 13912 10668
rect 13964 10616 13970 10668
rect 13998 10616 14004 10668
rect 14056 10665 14062 10668
rect 14056 10659 14084 10665
rect 14072 10625 14084 10659
rect 14056 10619 14084 10625
rect 14921 10659 14979 10665
rect 14921 10625 14933 10659
rect 14967 10656 14979 10659
rect 15102 10656 15108 10668
rect 14967 10628 15108 10656
rect 14967 10625 14979 10628
rect 14921 10619 14979 10625
rect 14056 10616 14062 10619
rect 15102 10616 15108 10628
rect 15160 10616 15166 10668
rect 15194 10616 15200 10668
rect 15252 10616 15258 10668
rect 15396 10656 15424 10684
rect 16114 10656 16120 10668
rect 15396 10628 16120 10656
rect 16114 10616 16120 10628
rect 16172 10616 16178 10668
rect 16500 10665 16528 10764
rect 18874 10752 18880 10764
rect 18932 10752 18938 10804
rect 16927 10689 16985 10695
rect 16485 10659 16543 10665
rect 16485 10625 16497 10659
rect 16531 10625 16543 10659
rect 16485 10619 16543 10625
rect 16574 10616 16580 10668
rect 16632 10656 16638 10668
rect 16927 10656 16939 10689
rect 16632 10655 16939 10656
rect 16973 10686 16985 10689
rect 16973 10655 16986 10686
rect 17126 10684 17132 10736
rect 17184 10724 17190 10736
rect 19242 10724 19248 10736
rect 17184 10696 19248 10724
rect 17184 10684 17190 10696
rect 19242 10684 19248 10696
rect 19300 10684 19306 10736
rect 16632 10628 16986 10655
rect 16632 10616 16638 10628
rect 17034 10616 17040 10668
rect 17092 10656 17098 10668
rect 18291 10659 18349 10665
rect 18291 10656 18303 10659
rect 17092 10628 18303 10656
rect 17092 10616 17098 10628
rect 18291 10625 18303 10628
rect 18337 10625 18349 10659
rect 18291 10619 18349 10625
rect 18690 10616 18696 10668
rect 18748 10656 18754 10668
rect 19797 10659 19855 10665
rect 19797 10656 19809 10659
rect 18748 10628 19809 10656
rect 18748 10616 18754 10628
rect 19797 10625 19809 10628
rect 19843 10625 19855 10659
rect 19797 10619 19855 10625
rect 20254 10616 20260 10668
rect 20312 10616 20318 10668
rect 13633 10591 13691 10597
rect 13633 10557 13645 10591
rect 13679 10588 13691 10591
rect 13722 10588 13728 10600
rect 13679 10560 13728 10588
rect 13679 10557 13691 10560
rect 13633 10551 13691 10557
rect 13722 10548 13728 10560
rect 13780 10548 13786 10600
rect 14185 10591 14243 10597
rect 14185 10557 14197 10591
rect 14231 10588 14243 10591
rect 14231 10560 14872 10588
rect 14231 10557 14243 10560
rect 14185 10551 14243 10557
rect 14844 10520 14872 10560
rect 16022 10548 16028 10600
rect 16080 10588 16086 10600
rect 16669 10591 16727 10597
rect 16669 10588 16681 10591
rect 16080 10560 16681 10588
rect 16080 10548 16086 10560
rect 16669 10557 16681 10560
rect 16715 10557 16727 10591
rect 16669 10551 16727 10557
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 14844 10492 14964 10520
rect 14826 10452 14832 10464
rect 13372 10424 14832 10452
rect 9824 10412 9830 10424
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 14936 10452 14964 10492
rect 15838 10480 15844 10532
rect 15896 10520 15902 10532
rect 15896 10492 16436 10520
rect 15896 10480 15902 10492
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 14936 10424 15945 10452
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 15933 10415 15991 10421
rect 16298 10412 16304 10464
rect 16356 10412 16362 10464
rect 16408 10452 16436 10492
rect 17402 10480 17408 10532
rect 17460 10520 17466 10532
rect 18064 10520 18092 10551
rect 19610 10548 19616 10600
rect 19668 10548 19674 10600
rect 17460 10492 18092 10520
rect 17460 10480 17466 10492
rect 19794 10480 19800 10532
rect 19852 10520 19858 10532
rect 20257 10523 20315 10529
rect 20257 10520 20269 10523
rect 19852 10492 20269 10520
rect 19852 10480 19858 10492
rect 20257 10489 20269 10492
rect 20303 10489 20315 10523
rect 20257 10483 20315 10489
rect 17681 10455 17739 10461
rect 17681 10452 17693 10455
rect 16408 10424 17693 10452
rect 17681 10421 17693 10424
rect 17727 10421 17739 10455
rect 17681 10415 17739 10421
rect 17770 10412 17776 10464
rect 17828 10452 17834 10464
rect 19061 10455 19119 10461
rect 19061 10452 19073 10455
rect 17828 10424 19073 10452
rect 17828 10412 17834 10424
rect 19061 10421 19073 10424
rect 19107 10421 19119 10455
rect 19061 10415 19119 10421
rect 1104 10362 20884 10384
rect 1104 10310 3422 10362
rect 3474 10310 3486 10362
rect 3538 10310 3550 10362
rect 3602 10310 3614 10362
rect 3666 10310 3678 10362
rect 3730 10310 8367 10362
rect 8419 10310 8431 10362
rect 8483 10310 8495 10362
rect 8547 10310 8559 10362
rect 8611 10310 8623 10362
rect 8675 10310 13312 10362
rect 13364 10310 13376 10362
rect 13428 10310 13440 10362
rect 13492 10310 13504 10362
rect 13556 10310 13568 10362
rect 13620 10310 18257 10362
rect 18309 10310 18321 10362
rect 18373 10310 18385 10362
rect 18437 10310 18449 10362
rect 18501 10310 18513 10362
rect 18565 10310 20884 10362
rect 1104 10288 20884 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 1581 10251 1639 10257
rect 1581 10248 1593 10251
rect 1544 10220 1593 10248
rect 1544 10208 1550 10220
rect 1581 10217 1593 10220
rect 1627 10217 1639 10251
rect 3326 10248 3332 10260
rect 1581 10211 1639 10217
rect 1964 10220 3332 10248
rect 1964 10180 1992 10220
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3418 10208 3424 10260
rect 3476 10248 3482 10260
rect 3476 10220 4108 10248
rect 3476 10208 3482 10220
rect 1504 10152 1992 10180
rect 1504 10124 1532 10152
rect 3050 10140 3056 10192
rect 3108 10180 3114 10192
rect 4080 10180 4108 10220
rect 4154 10208 4160 10260
rect 4212 10208 4218 10260
rect 4706 10208 4712 10260
rect 4764 10208 4770 10260
rect 4798 10208 4804 10260
rect 4856 10248 4862 10260
rect 6822 10248 6828 10260
rect 4856 10220 5488 10248
rect 4856 10208 4862 10220
rect 4724 10180 4752 10208
rect 5460 10192 5488 10220
rect 5570 10220 6828 10248
rect 3108 10152 4016 10180
rect 4080 10152 4752 10180
rect 3108 10140 3114 10152
rect 1486 10072 1492 10124
rect 1544 10072 1550 10124
rect 2958 10072 2964 10124
rect 3016 10112 3022 10124
rect 3510 10112 3516 10124
rect 3016 10084 3516 10112
rect 3016 10072 3022 10084
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 3878 10112 3884 10124
rect 3620 10084 3884 10112
rect 1302 10004 1308 10056
rect 1360 10044 1366 10056
rect 1765 10047 1823 10053
rect 1765 10044 1777 10047
rect 1360 10016 1777 10044
rect 1360 10004 1366 10016
rect 1765 10013 1777 10016
rect 1811 10013 1823 10047
rect 1765 10007 1823 10013
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10013 1915 10047
rect 1857 10007 1915 10013
rect 2131 10047 2189 10053
rect 2131 10013 2143 10047
rect 2177 10044 2189 10047
rect 2866 10044 2872 10056
rect 2177 10016 2872 10044
rect 2177 10013 2189 10016
rect 2131 10007 2189 10013
rect 1872 9976 1900 10007
rect 2866 10004 2872 10016
rect 2924 10004 2930 10056
rect 3620 10053 3648 10084
rect 3878 10072 3884 10084
rect 3936 10072 3942 10124
rect 3988 10112 4016 10152
rect 5442 10140 5448 10192
rect 5500 10140 5506 10192
rect 4709 10115 4767 10121
rect 4709 10112 4721 10115
rect 3988 10084 4108 10112
rect 3605 10047 3663 10053
rect 3605 10013 3617 10047
rect 3651 10013 3663 10047
rect 3605 10007 3663 10013
rect 1872 9948 2268 9976
rect 2240 9920 2268 9948
rect 2590 9936 2596 9988
rect 2648 9976 2654 9988
rect 3881 9979 3939 9985
rect 3881 9976 3893 9979
rect 2648 9948 3893 9976
rect 2648 9936 2654 9948
rect 3881 9945 3893 9948
rect 3927 9945 3939 9979
rect 3881 9939 3939 9945
rect 4080 9920 4108 10084
rect 4448 10084 4721 10112
rect 4448 10056 4476 10084
rect 4709 10081 4721 10084
rect 4755 10081 4767 10115
rect 4709 10075 4767 10081
rect 4430 10004 4436 10056
rect 4488 10004 4494 10056
rect 4525 10047 4583 10053
rect 4525 10013 4537 10047
rect 4571 10044 4583 10047
rect 4614 10044 4620 10056
rect 4571 10016 4620 10044
rect 4571 10013 4583 10016
rect 4525 10007 4583 10013
rect 4614 10004 4620 10016
rect 4672 10004 4678 10056
rect 4951 10047 5009 10053
rect 4951 10013 4963 10047
rect 4997 10013 5009 10047
rect 4951 10007 5009 10013
rect 4966 9976 4994 10007
rect 5074 10004 5080 10056
rect 5132 10044 5138 10056
rect 5570 10044 5598 10220
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7101 10251 7159 10257
rect 7101 10248 7113 10251
rect 6932 10220 7113 10248
rect 5994 10072 6000 10124
rect 6052 10112 6058 10124
rect 6089 10115 6147 10121
rect 6089 10112 6101 10115
rect 6052 10084 6101 10112
rect 6052 10072 6058 10084
rect 6089 10081 6101 10084
rect 6135 10081 6147 10115
rect 6932 10112 6960 10220
rect 7101 10217 7113 10220
rect 7147 10217 7159 10251
rect 7101 10211 7159 10217
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 7248 10220 8800 10248
rect 7248 10208 7254 10220
rect 7282 10140 7288 10192
rect 7340 10180 7346 10192
rect 7340 10152 7512 10180
rect 7340 10140 7346 10152
rect 6932 10084 7328 10112
rect 6089 10075 6147 10081
rect 5132 10016 5598 10044
rect 5132 10004 5138 10016
rect 5626 10004 5632 10056
rect 5684 10044 5690 10056
rect 6331 10047 6389 10053
rect 6331 10044 6343 10047
rect 5684 10016 6343 10044
rect 5684 10004 5690 10016
rect 6331 10013 6343 10016
rect 6377 10044 6389 10047
rect 7006 10044 7012 10056
rect 6377 10016 7012 10044
rect 6377 10013 6389 10016
rect 6331 10007 6389 10013
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 7190 9976 7196 9988
rect 4264 9948 7196 9976
rect 2222 9868 2228 9920
rect 2280 9868 2286 9920
rect 2866 9868 2872 9920
rect 2924 9868 2930 9920
rect 2958 9868 2964 9920
rect 3016 9908 3022 9920
rect 3421 9911 3479 9917
rect 3421 9908 3433 9911
rect 3016 9880 3433 9908
rect 3016 9868 3022 9880
rect 3421 9877 3433 9880
rect 3467 9877 3479 9911
rect 3421 9871 3479 9877
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4264 9908 4292 9948
rect 7190 9936 7196 9948
rect 7248 9936 7254 9988
rect 4120 9880 4292 9908
rect 4120 9868 4126 9880
rect 4338 9868 4344 9920
rect 4396 9868 4402 9920
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 5074 9908 5080 9920
rect 4672 9880 5080 9908
rect 4672 9868 4678 9880
rect 5074 9868 5080 9880
rect 5132 9868 5138 9920
rect 5442 9868 5448 9920
rect 5500 9908 5506 9920
rect 5721 9911 5779 9917
rect 5721 9908 5733 9911
rect 5500 9880 5733 9908
rect 5500 9868 5506 9880
rect 5721 9877 5733 9880
rect 5767 9877 5779 9911
rect 5721 9871 5779 9877
rect 6178 9868 6184 9920
rect 6236 9908 6242 9920
rect 6730 9908 6736 9920
rect 6236 9880 6736 9908
rect 6236 9868 6242 9880
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 7300 9908 7328 10084
rect 7484 10053 7512 10152
rect 8772 10124 8800 10220
rect 9306 10208 9312 10260
rect 9364 10248 9370 10260
rect 9766 10248 9772 10260
rect 9364 10220 9772 10248
rect 9364 10208 9370 10220
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 12529 10251 12587 10257
rect 10336 10220 12480 10248
rect 9398 10140 9404 10192
rect 9456 10180 9462 10192
rect 10229 10183 10287 10189
rect 10229 10180 10241 10183
rect 9456 10152 10241 10180
rect 9456 10140 9462 10152
rect 10229 10149 10241 10152
rect 10275 10149 10287 10183
rect 10229 10143 10287 10149
rect 8202 10072 8208 10124
rect 8260 10072 8266 10124
rect 8754 10072 8760 10124
rect 8812 10072 8818 10124
rect 9582 10072 9588 10124
rect 9640 10072 9646 10124
rect 9950 10112 9956 10124
rect 9692 10084 9956 10112
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10044 7527 10047
rect 7743 10047 7801 10053
rect 7515 10016 7696 10044
rect 7515 10013 7527 10016
rect 7469 10007 7527 10013
rect 7558 9908 7564 9920
rect 7300 9880 7564 9908
rect 7558 9868 7564 9880
rect 7616 9868 7622 9920
rect 7668 9908 7696 10016
rect 7743 10013 7755 10047
rect 7789 10044 7801 10047
rect 8110 10044 8116 10056
rect 7789 10016 8116 10044
rect 7789 10013 7801 10016
rect 7743 10007 7801 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 8220 9976 8248 10072
rect 9692 10056 9720 10084
rect 9950 10072 9956 10084
rect 10008 10072 10014 10124
rect 10336 10112 10364 10220
rect 12452 10180 12480 10220
rect 12529 10217 12541 10251
rect 12575 10248 12587 10251
rect 12618 10248 12624 10260
rect 12575 10220 12624 10248
rect 12575 10217 12587 10220
rect 12529 10211 12587 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 13906 10208 13912 10260
rect 13964 10248 13970 10260
rect 14458 10248 14464 10260
rect 13964 10220 14464 10248
rect 13964 10208 13970 10220
rect 14458 10208 14464 10220
rect 14516 10208 14522 10260
rect 15838 10248 15844 10260
rect 14752 10220 15844 10248
rect 14550 10180 14556 10192
rect 12452 10152 14556 10180
rect 14550 10140 14556 10152
rect 14608 10180 14614 10192
rect 14752 10189 14780 10220
rect 15838 10208 15844 10220
rect 15896 10208 15902 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 16040 10220 17049 10248
rect 14737 10183 14795 10189
rect 14608 10152 14688 10180
rect 14608 10140 14614 10152
rect 10502 10112 10508 10124
rect 10336 10084 10508 10112
rect 10502 10072 10508 10084
rect 10560 10072 10566 10124
rect 10594 10072 10600 10124
rect 10652 10121 10658 10124
rect 10652 10115 10680 10121
rect 10668 10081 10680 10115
rect 10652 10075 10680 10081
rect 10652 10072 10658 10075
rect 10962 10072 10968 10124
rect 11020 10112 11026 10124
rect 11425 10115 11483 10121
rect 11425 10112 11437 10115
rect 11020 10084 11437 10112
rect 11020 10072 11026 10084
rect 11425 10081 11437 10084
rect 11471 10081 11483 10115
rect 11425 10075 11483 10081
rect 11514 10072 11520 10124
rect 11572 10072 11578 10124
rect 12894 10072 12900 10124
rect 12952 10112 12958 10124
rect 13170 10112 13176 10124
rect 12952 10084 13176 10112
rect 12952 10072 12958 10084
rect 13170 10072 13176 10084
rect 13228 10112 13234 10124
rect 14274 10112 14280 10124
rect 13228 10084 14280 10112
rect 13228 10072 13234 10084
rect 14274 10072 14280 10084
rect 14332 10072 14338 10124
rect 14660 10112 14688 10152
rect 14737 10149 14749 10183
rect 14783 10149 14795 10183
rect 14737 10143 14795 10149
rect 15013 10115 15071 10121
rect 15013 10112 15025 10115
rect 14660 10084 15025 10112
rect 15013 10081 15025 10084
rect 15059 10081 15071 10115
rect 15013 10075 15071 10081
rect 15102 10072 15108 10124
rect 15160 10121 15166 10124
rect 15160 10115 15188 10121
rect 15176 10081 15188 10115
rect 15160 10075 15188 10081
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10112 15347 10115
rect 16040 10112 16068 10220
rect 17037 10217 17049 10220
rect 17083 10217 17095 10251
rect 18690 10248 18696 10260
rect 17037 10211 17095 10217
rect 17126 10220 18696 10248
rect 16758 10140 16764 10192
rect 16816 10180 16822 10192
rect 17126 10180 17154 10220
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 18782 10208 18788 10260
rect 18840 10208 18846 10260
rect 18874 10208 18880 10260
rect 18932 10248 18938 10260
rect 20257 10251 20315 10257
rect 20257 10248 20269 10251
rect 18932 10220 20269 10248
rect 18932 10208 18938 10220
rect 20257 10217 20269 10220
rect 20303 10217 20315 10251
rect 20257 10211 20315 10217
rect 16816 10152 17154 10180
rect 16816 10140 16822 10152
rect 15335 10084 16068 10112
rect 15335 10081 15347 10084
rect 15289 10075 15347 10081
rect 15160 10072 15166 10075
rect 17218 10072 17224 10124
rect 17276 10112 17282 10124
rect 17402 10112 17408 10124
rect 17276 10084 17408 10112
rect 17276 10072 17282 10084
rect 17402 10072 17408 10084
rect 17460 10072 17466 10124
rect 18782 10072 18788 10124
rect 18840 10112 18846 10124
rect 19150 10112 19156 10124
rect 18840 10084 19156 10112
rect 18840 10072 18846 10084
rect 19150 10072 19156 10084
rect 19208 10112 19214 10124
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 19208 10084 19257 10112
rect 19208 10072 19214 10084
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 19245 10075 19303 10081
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8570 10044 8576 10056
rect 8352 10016 8576 10044
rect 8352 10004 8358 10016
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 9674 10004 9680 10056
rect 9732 10004 9738 10056
rect 9766 10004 9772 10056
rect 9824 10004 9830 10056
rect 10778 10004 10784 10056
rect 10836 10004 10842 10056
rect 11790 10044 11796 10056
rect 11751 10016 11796 10044
rect 11790 10004 11796 10016
rect 11848 10004 11854 10056
rect 12342 10004 12348 10056
rect 12400 10044 12406 10056
rect 13998 10044 14004 10056
rect 12400 10016 14004 10044
rect 12400 10004 12406 10016
rect 13998 10004 14004 10016
rect 14056 10004 14062 10056
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14182 10044 14188 10056
rect 14139 10016 14188 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 14182 10004 14188 10016
rect 14240 10004 14246 10056
rect 14458 10044 14464 10056
rect 14300 10016 14464 10044
rect 8220 9948 9720 9976
rect 8386 9908 8392 9920
rect 7668 9880 8392 9908
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8481 9911 8539 9917
rect 8481 9877 8493 9911
rect 8527 9908 8539 9911
rect 9398 9908 9404 9920
rect 8527 9880 9404 9908
rect 8527 9877 8539 9880
rect 8481 9871 8539 9877
rect 9398 9868 9404 9880
rect 9456 9868 9462 9920
rect 9692 9908 9720 9948
rect 12526 9936 12532 9988
rect 12584 9976 12590 9988
rect 14300 9976 14328 10016
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 15930 10004 15936 10056
rect 15988 10004 15994 10056
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 17678 10053 17684 10056
rect 16267 10047 16325 10053
rect 16267 10044 16279 10047
rect 16132 10016 16279 10044
rect 12584 9948 14328 9976
rect 15948 9976 15976 10004
rect 16132 9976 16160 10016
rect 16267 10013 16279 10016
rect 16313 10013 16325 10047
rect 16267 10007 16325 10013
rect 17647 10047 17684 10053
rect 17647 10013 17659 10047
rect 17647 10007 17684 10013
rect 17678 10004 17684 10007
rect 17736 10004 17742 10056
rect 17770 10004 17776 10056
rect 17828 10004 17834 10056
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 18969 10047 19027 10053
rect 18969 10044 18981 10047
rect 18196 10016 18981 10044
rect 18196 10004 18202 10016
rect 18969 10013 18981 10016
rect 19015 10013 19027 10047
rect 18969 10007 19027 10013
rect 19487 10047 19545 10053
rect 19487 10013 19499 10047
rect 19533 10013 19545 10047
rect 19487 10007 19545 10013
rect 17788 9976 17816 10004
rect 19502 9976 19530 10007
rect 15948 9948 16160 9976
rect 16224 9948 19530 9976
rect 12584 9936 12590 9948
rect 9766 9908 9772 9920
rect 9692 9880 9772 9908
rect 9766 9868 9772 9880
rect 9824 9868 9830 9920
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 15933 9911 15991 9917
rect 15933 9908 15945 9911
rect 10100 9880 15945 9908
rect 10100 9868 10106 9880
rect 15933 9877 15945 9880
rect 15979 9877 15991 9911
rect 15933 9871 15991 9877
rect 16114 9868 16120 9920
rect 16172 9908 16178 9920
rect 16224 9908 16252 9948
rect 19702 9936 19708 9988
rect 19760 9936 19766 9988
rect 16172 9880 16252 9908
rect 16172 9868 16178 9880
rect 16390 9868 16396 9920
rect 16448 9908 16454 9920
rect 18417 9911 18475 9917
rect 18417 9908 18429 9911
rect 16448 9880 18429 9908
rect 16448 9868 16454 9880
rect 18417 9877 18429 9880
rect 18463 9908 18475 9911
rect 19720 9908 19748 9936
rect 18463 9880 19748 9908
rect 18463 9877 18475 9880
rect 18417 9871 18475 9877
rect 1104 9818 21043 9840
rect 1104 9766 5894 9818
rect 5946 9766 5958 9818
rect 6010 9766 6022 9818
rect 6074 9766 6086 9818
rect 6138 9766 6150 9818
rect 6202 9766 10839 9818
rect 10891 9766 10903 9818
rect 10955 9766 10967 9818
rect 11019 9766 11031 9818
rect 11083 9766 11095 9818
rect 11147 9766 15784 9818
rect 15836 9766 15848 9818
rect 15900 9766 15912 9818
rect 15964 9766 15976 9818
rect 16028 9766 16040 9818
rect 16092 9766 20729 9818
rect 20781 9766 20793 9818
rect 20845 9766 20857 9818
rect 20909 9766 20921 9818
rect 20973 9766 20985 9818
rect 21037 9766 21043 9818
rect 1104 9744 21043 9766
rect 1762 9664 1768 9716
rect 1820 9664 1826 9716
rect 2774 9704 2780 9716
rect 2608 9676 2780 9704
rect 1489 9639 1547 9645
rect 1489 9605 1501 9639
rect 1535 9636 1547 9639
rect 2406 9636 2412 9648
rect 1535 9608 2412 9636
rect 1535 9605 1547 9608
rect 1489 9599 1547 9605
rect 2406 9596 2412 9608
rect 2464 9596 2470 9648
rect 106 9528 112 9580
rect 164 9568 170 9580
rect 2608 9577 2636 9676
rect 2774 9664 2780 9676
rect 2832 9704 2838 9716
rect 3234 9704 3240 9716
rect 2832 9676 3240 9704
rect 2832 9664 2838 9676
rect 3234 9664 3240 9676
rect 3292 9664 3298 9716
rect 3326 9664 3332 9716
rect 3384 9704 3390 9716
rect 5350 9704 5356 9716
rect 3384 9676 5356 9704
rect 3384 9664 3390 9676
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 6546 9664 6552 9716
rect 6604 9704 6610 9716
rect 6822 9704 6828 9716
rect 6604 9676 6828 9704
rect 6604 9664 6610 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 7742 9664 7748 9716
rect 7800 9664 7806 9716
rect 8386 9704 8392 9716
rect 8300 9676 8392 9704
rect 4154 9596 4160 9648
rect 4212 9596 4218 9648
rect 6380 9608 7018 9636
rect 3510 9577 3516 9580
rect 2317 9571 2375 9577
rect 164 9540 2268 9568
rect 164 9528 170 9540
rect 2240 9500 2268 9540
rect 2317 9537 2329 9571
rect 2363 9568 2375 9571
rect 2593 9571 2651 9577
rect 2363 9540 2544 9568
rect 2363 9537 2375 9540
rect 2317 9531 2375 9537
rect 2409 9503 2467 9509
rect 2409 9500 2421 9503
rect 2240 9472 2421 9500
rect 2409 9469 2421 9472
rect 2455 9469 2467 9503
rect 2409 9463 2467 9469
rect 2130 9324 2136 9376
rect 2188 9324 2194 9376
rect 2516 9364 2544 9540
rect 2593 9537 2605 9571
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 3467 9571 3516 9577
rect 3467 9537 3479 9571
rect 3513 9537 3516 9571
rect 3467 9531 3516 9537
rect 3510 9528 3516 9531
rect 3568 9528 3574 9580
rect 4172 9568 4200 9596
rect 6380 9580 6408 9608
rect 4341 9571 4399 9577
rect 4341 9568 4353 9571
rect 4172 9540 4353 9568
rect 4341 9537 4353 9540
rect 4387 9537 4399 9571
rect 5279 9571 5337 9577
rect 5279 9546 5291 9571
rect 4341 9531 4399 9537
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 2832 9472 3341 9500
rect 2832 9460 2838 9472
rect 3329 9469 3341 9472
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 4154 9500 4160 9512
rect 3651 9472 4160 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 4154 9460 4160 9472
rect 4212 9460 4218 9512
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 4706 9500 4712 9512
rect 4571 9472 4712 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 4706 9460 4712 9472
rect 4764 9460 4770 9512
rect 4890 9460 4896 9512
rect 4948 9460 4954 9512
rect 5258 9494 5264 9546
rect 5325 9537 5337 9571
rect 5316 9531 5337 9537
rect 5442 9534 5448 9570
rect 5316 9506 5329 9531
rect 5414 9518 5448 9534
rect 5500 9518 5506 9570
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 6546 9528 6552 9580
rect 6604 9528 6610 9580
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 6990 9577 7018 9608
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 7340 9608 7418 9636
rect 7340 9596 7346 9608
rect 6975 9571 7033 9577
rect 6975 9537 6987 9571
rect 7021 9537 7033 9571
rect 6975 9531 7033 9537
rect 5414 9509 5488 9518
rect 5399 9506 5488 9509
rect 5316 9494 5322 9506
rect 5399 9503 5457 9506
rect 5399 9469 5411 9503
rect 5445 9469 5457 9503
rect 5399 9463 5457 9469
rect 5534 9460 5540 9512
rect 5592 9460 5598 9512
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 6748 9500 6776 9528
rect 5960 9472 6776 9500
rect 7390 9500 7418 9608
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 8113 9571 8171 9577
rect 8113 9568 8125 9571
rect 7800 9540 8125 9568
rect 7800 9528 7806 9540
rect 8113 9537 8125 9540
rect 8159 9568 8171 9571
rect 8300 9568 8328 9676
rect 8386 9664 8392 9676
rect 8444 9704 8450 9716
rect 8444 9676 11560 9704
rect 8444 9664 8450 9676
rect 9306 9636 9312 9648
rect 8402 9608 9312 9636
rect 8402 9577 8430 9608
rect 9306 9596 9312 9608
rect 9364 9596 9370 9648
rect 9582 9636 9588 9648
rect 9508 9608 9588 9636
rect 8159 9540 8328 9568
rect 8387 9571 8445 9577
rect 8159 9537 8171 9540
rect 8113 9531 8171 9537
rect 8387 9537 8399 9571
rect 8433 9537 8445 9571
rect 8387 9531 8445 9537
rect 8478 9528 8484 9580
rect 8536 9568 8542 9580
rect 9508 9577 9536 9608
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 9493 9571 9551 9577
rect 8536 9540 8733 9568
rect 8536 9528 8542 9540
rect 8705 9500 8733 9540
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 10410 9528 10416 9580
rect 10468 9528 10474 9580
rect 10594 9577 10600 9580
rect 10551 9571 10600 9577
rect 10551 9537 10563 9571
rect 10597 9537 10600 9571
rect 10551 9531 10600 9537
rect 10594 9528 10600 9531
rect 10652 9528 10658 9580
rect 11532 9512 11560 9676
rect 11698 9664 11704 9716
rect 11756 9664 11762 9716
rect 12342 9664 12348 9716
rect 12400 9704 12406 9716
rect 15749 9707 15807 9713
rect 12400 9676 15700 9704
rect 12400 9664 12406 9676
rect 11716 9636 11744 9664
rect 11716 9608 11986 9636
rect 11958 9577 11986 9608
rect 15672 9580 15700 9676
rect 15749 9673 15761 9707
rect 15795 9704 15807 9707
rect 15795 9676 16252 9704
rect 15795 9673 15807 9676
rect 15749 9667 15807 9673
rect 14918 9577 14924 9580
rect 11943 9571 12001 9577
rect 11943 9537 11955 9571
rect 11989 9537 12001 9571
rect 11943 9531 12001 9537
rect 13817 9571 13875 9577
rect 13817 9537 13829 9571
rect 13863 9568 13875 9571
rect 14875 9571 14924 9577
rect 13863 9540 14228 9568
rect 13863 9537 13875 9540
rect 13817 9531 13875 9537
rect 14200 9512 14228 9540
rect 14875 9537 14887 9571
rect 14921 9537 14924 9571
rect 14875 9531 14924 9537
rect 14918 9528 14924 9531
rect 14976 9528 14982 9580
rect 15654 9528 15660 9580
rect 15712 9528 15718 9580
rect 15933 9571 15991 9577
rect 15933 9537 15945 9571
rect 15979 9568 15991 9571
rect 16022 9568 16028 9580
rect 15979 9540 16028 9568
rect 15979 9537 15991 9540
rect 15933 9531 15991 9537
rect 16022 9528 16028 9540
rect 16080 9528 16086 9580
rect 16224 9577 16252 9676
rect 16298 9664 16304 9716
rect 16356 9704 16362 9716
rect 16393 9707 16451 9713
rect 16393 9704 16405 9707
rect 16356 9676 16405 9704
rect 16356 9664 16362 9676
rect 16393 9673 16405 9676
rect 16439 9673 16451 9707
rect 17218 9704 17224 9716
rect 16393 9667 16451 9673
rect 16500 9676 17224 9704
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 7390 9472 7972 9500
rect 8705 9472 9352 9500
rect 5960 9460 5966 9472
rect 3050 9392 3056 9444
rect 3108 9392 3114 9444
rect 4908 9432 4936 9460
rect 4126 9404 4936 9432
rect 4126 9364 4154 9404
rect 4982 9392 4988 9444
rect 5040 9392 5046 9444
rect 5920 9404 6408 9432
rect 2516 9336 4154 9364
rect 4249 9367 4307 9373
rect 4249 9333 4261 9367
rect 4295 9364 4307 9367
rect 4614 9364 4620 9376
rect 4295 9336 4620 9364
rect 4295 9333 4307 9336
rect 4249 9327 4307 9333
rect 4614 9324 4620 9336
rect 4672 9324 4678 9376
rect 4890 9324 4896 9376
rect 4948 9364 4954 9376
rect 5920 9364 5948 9404
rect 4948 9336 5948 9364
rect 6181 9367 6239 9373
rect 4948 9324 4954 9336
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 6270 9364 6276 9376
rect 6227 9336 6276 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 6270 9324 6276 9336
rect 6328 9324 6334 9376
rect 6380 9373 6408 9404
rect 6365 9367 6423 9373
rect 6365 9333 6377 9367
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 7834 9364 7840 9376
rect 6788 9336 7840 9364
rect 6788 9324 6794 9336
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 7944 9364 7972 9472
rect 9324 9444 9352 9472
rect 9398 9460 9404 9512
rect 9456 9460 9462 9512
rect 9677 9503 9735 9509
rect 9677 9469 9689 9503
rect 9723 9500 9735 9503
rect 9766 9500 9772 9512
rect 9723 9472 9772 9500
rect 9723 9469 9735 9472
rect 9677 9463 9735 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9500 10747 9503
rect 10735 9472 11100 9500
rect 10735 9469 10747 9472
rect 10689 9463 10747 9469
rect 9306 9392 9312 9444
rect 9364 9392 9370 9444
rect 9416 9432 9444 9460
rect 10137 9435 10195 9441
rect 10137 9432 10149 9435
rect 9416 9404 10149 9432
rect 10137 9401 10149 9404
rect 10183 9401 10195 9435
rect 10137 9395 10195 9401
rect 8386 9364 8392 9376
rect 7944 9336 8392 9364
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 9125 9367 9183 9373
rect 9125 9333 9137 9367
rect 9171 9364 9183 9367
rect 11072 9364 11100 9472
rect 11514 9460 11520 9512
rect 11572 9500 11578 9512
rect 11701 9503 11759 9509
rect 11701 9500 11713 9503
rect 11572 9472 11713 9500
rect 11572 9460 11578 9472
rect 11701 9469 11713 9472
rect 11747 9469 11759 9503
rect 11701 9463 11759 9469
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 13170 9500 13176 9512
rect 12676 9472 13176 9500
rect 12676 9460 12682 9472
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 13906 9432 13912 9444
rect 12636 9404 13912 9432
rect 9171 9336 11100 9364
rect 9171 9333 9183 9336
rect 9125 9327 9183 9333
rect 11330 9324 11336 9376
rect 11388 9324 11394 9376
rect 11790 9324 11796 9376
rect 11848 9364 11854 9376
rect 12636 9364 12664 9404
rect 13906 9392 13912 9404
rect 13964 9392 13970 9444
rect 14016 9432 14044 9463
rect 14182 9460 14188 9512
rect 14240 9460 14246 9512
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 14737 9503 14795 9509
rect 14737 9500 14749 9503
rect 14608 9472 14749 9500
rect 14608 9460 14614 9472
rect 14737 9469 14749 9472
rect 14783 9469 14795 9503
rect 14737 9463 14795 9469
rect 15011 9503 15069 9509
rect 15011 9469 15023 9503
rect 15057 9500 15069 9503
rect 16114 9500 16120 9512
rect 15057 9472 16120 9500
rect 15057 9469 15069 9472
rect 15011 9463 15069 9469
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 16224 9500 16252 9531
rect 16298 9528 16304 9580
rect 16356 9528 16362 9580
rect 16500 9577 16528 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 18598 9664 18604 9716
rect 18656 9704 18662 9716
rect 18874 9704 18880 9716
rect 18656 9676 18880 9704
rect 18656 9664 18662 9676
rect 18874 9664 18880 9676
rect 18932 9664 18938 9716
rect 19058 9664 19064 9716
rect 19116 9704 19122 9716
rect 19797 9707 19855 9713
rect 19797 9704 19809 9707
rect 19116 9676 19809 9704
rect 19116 9664 19122 9676
rect 19797 9673 19809 9676
rect 19843 9673 19855 9707
rect 19797 9667 19855 9673
rect 16666 9596 16672 9648
rect 16724 9636 16730 9648
rect 17862 9636 17868 9648
rect 16724 9608 17868 9636
rect 16724 9596 16730 9608
rect 17862 9596 17868 9608
rect 17920 9596 17926 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 20257 9639 20315 9645
rect 20257 9636 20269 9639
rect 19576 9608 20269 9636
rect 19576 9596 19582 9608
rect 20257 9605 20269 9608
rect 20303 9605 20315 9639
rect 20257 9599 20315 9605
rect 16485 9571 16543 9577
rect 16485 9537 16497 9571
rect 16531 9537 16543 9571
rect 16925 9571 16983 9577
rect 16925 9568 16937 9571
rect 16485 9531 16543 9537
rect 16592 9540 16937 9568
rect 16592 9500 16620 9540
rect 16925 9537 16937 9540
rect 16971 9537 16983 9571
rect 16925 9531 16983 9537
rect 18325 9571 18383 9577
rect 18325 9537 18337 9571
rect 18371 9537 18383 9571
rect 18325 9531 18383 9537
rect 16224 9472 16620 9500
rect 16666 9460 16672 9512
rect 16724 9460 16730 9512
rect 14274 9432 14280 9444
rect 14016 9404 14280 9432
rect 14274 9392 14280 9404
rect 14332 9392 14338 9444
rect 14458 9392 14464 9444
rect 14516 9392 14522 9444
rect 18340 9432 18368 9531
rect 18506 9528 18512 9580
rect 18564 9568 18570 9580
rect 19056 9577 19062 9580
rect 19027 9571 19062 9577
rect 19027 9568 19039 9571
rect 18564 9540 19039 9568
rect 18564 9528 18570 9540
rect 19027 9537 19039 9540
rect 19027 9531 19062 9537
rect 19056 9528 19062 9531
rect 19114 9528 19120 9580
rect 20165 9571 20223 9577
rect 20165 9537 20177 9571
rect 20211 9568 20223 9571
rect 21910 9568 21916 9580
rect 20211 9540 21916 9568
rect 20211 9537 20223 9540
rect 20165 9531 20223 9537
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 18601 9503 18659 9509
rect 18601 9469 18613 9503
rect 18647 9500 18659 9503
rect 18690 9500 18696 9512
rect 18647 9472 18696 9500
rect 18647 9469 18659 9472
rect 18601 9463 18659 9469
rect 18690 9460 18696 9472
rect 18748 9460 18754 9512
rect 18782 9460 18788 9512
rect 18840 9460 18846 9512
rect 15396 9404 16710 9432
rect 11848 9336 12664 9364
rect 11848 9324 11854 9336
rect 12710 9324 12716 9376
rect 12768 9324 12774 9376
rect 12802 9324 12808 9376
rect 12860 9364 12866 9376
rect 15396 9364 15424 9404
rect 12860 9336 15424 9364
rect 12860 9324 12866 9336
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 15657 9367 15715 9373
rect 15657 9364 15669 9367
rect 15528 9336 15669 9364
rect 15528 9324 15534 9336
rect 15657 9333 15669 9336
rect 15703 9333 15715 9367
rect 15657 9327 15715 9333
rect 16025 9367 16083 9373
rect 16025 9333 16037 9367
rect 16071 9364 16083 9367
rect 16574 9364 16580 9376
rect 16071 9336 16580 9364
rect 16071 9333 16083 9336
rect 16025 9327 16083 9333
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 16682 9364 16710 9404
rect 17602 9404 18368 9432
rect 17602 9364 17630 9404
rect 19518 9392 19524 9444
rect 19576 9432 19582 9444
rect 19576 9404 19932 9432
rect 19576 9392 19582 9404
rect 16682 9336 17630 9364
rect 18049 9367 18107 9373
rect 18049 9333 18061 9367
rect 18095 9364 18107 9367
rect 18138 9364 18144 9376
rect 18095 9336 18144 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 19904 9364 19932 9404
rect 20070 9364 20076 9376
rect 19904 9336 20076 9364
rect 20070 9324 20076 9336
rect 20128 9324 20134 9376
rect 1104 9274 20884 9296
rect 1104 9222 3422 9274
rect 3474 9222 3486 9274
rect 3538 9222 3550 9274
rect 3602 9222 3614 9274
rect 3666 9222 3678 9274
rect 3730 9222 8367 9274
rect 8419 9222 8431 9274
rect 8483 9222 8495 9274
rect 8547 9222 8559 9274
rect 8611 9222 8623 9274
rect 8675 9222 13312 9274
rect 13364 9222 13376 9274
rect 13428 9222 13440 9274
rect 13492 9222 13504 9274
rect 13556 9222 13568 9274
rect 13620 9222 18257 9274
rect 18309 9222 18321 9274
rect 18373 9222 18385 9274
rect 18437 9222 18449 9274
rect 18501 9222 18513 9274
rect 18565 9222 20884 9274
rect 1104 9200 20884 9222
rect 1762 9120 1768 9172
rect 1820 9120 1826 9172
rect 2314 9120 2320 9172
rect 2372 9160 2378 9172
rect 4157 9163 4215 9169
rect 4157 9160 4169 9163
rect 2372 9132 4169 9160
rect 2372 9120 2378 9132
rect 4157 9129 4169 9132
rect 4203 9129 4215 9163
rect 4157 9123 4215 9129
rect 4246 9120 4252 9172
rect 4304 9160 4310 9172
rect 4525 9163 4583 9169
rect 4525 9160 4537 9163
rect 4304 9132 4537 9160
rect 4304 9120 4310 9132
rect 4525 9129 4537 9132
rect 4571 9129 4583 9163
rect 5166 9160 5172 9172
rect 4525 9123 4583 9129
rect 4908 9132 5172 9160
rect 4908 9092 4936 9132
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 5552 9120 5558 9172
rect 5610 9160 5616 9172
rect 6362 9160 6368 9172
rect 5610 9132 6368 9160
rect 5610 9120 5616 9132
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 11885 9163 11943 9169
rect 11885 9160 11897 9163
rect 6604 9132 11897 9160
rect 6604 9120 6610 9132
rect 11885 9129 11897 9132
rect 11931 9129 11943 9163
rect 11885 9123 11943 9129
rect 12526 9120 12532 9172
rect 12584 9160 12590 9172
rect 13722 9160 13728 9172
rect 12584 9132 13728 9160
rect 12584 9120 12590 9132
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 14458 9120 14464 9172
rect 14516 9160 14522 9172
rect 15105 9163 15163 9169
rect 15105 9160 15117 9163
rect 14516 9132 15117 9160
rect 14516 9120 14522 9132
rect 15105 9129 15117 9132
rect 15151 9129 15163 9163
rect 15562 9160 15568 9172
rect 15105 9123 15163 9129
rect 15488 9132 15568 9160
rect 3252 9064 4936 9092
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8956 1731 8959
rect 2038 8956 2044 8968
rect 1719 8928 2044 8956
rect 1719 8925 1731 8928
rect 1673 8919 1731 8925
rect 2038 8916 2044 8928
rect 2096 8916 2102 8968
rect 2222 8916 2228 8968
rect 2280 8956 2286 8968
rect 2317 8959 2375 8965
rect 2317 8956 2329 8959
rect 2280 8928 2329 8956
rect 2280 8916 2286 8928
rect 2317 8925 2329 8928
rect 2363 8925 2375 8959
rect 2317 8919 2375 8925
rect 2591 8959 2649 8965
rect 2591 8925 2603 8959
rect 2637 8956 2649 8959
rect 3142 8956 3148 8968
rect 2637 8928 3148 8956
rect 2637 8925 2649 8928
rect 2591 8919 2649 8925
rect 2332 8888 2360 8919
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3252 8888 3280 9064
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 4908 9033 4936 9064
rect 5905 9095 5963 9101
rect 5905 9061 5917 9095
rect 5951 9092 5963 9095
rect 5951 9064 6592 9092
rect 5951 9061 5963 9064
rect 5905 9055 5963 9061
rect 6564 9036 6592 9064
rect 6914 9052 6920 9104
rect 6972 9052 6978 9104
rect 9950 9052 9956 9104
rect 10008 9052 10014 9104
rect 10134 9052 10140 9104
rect 10192 9092 10198 9104
rect 12621 9095 12679 9101
rect 10192 9064 10824 9092
rect 10192 9052 10198 9064
rect 4893 9027 4951 9033
rect 3568 8996 4476 9024
rect 3568 8984 3574 8996
rect 3881 8959 3939 8965
rect 3881 8925 3893 8959
rect 3927 8956 3939 8959
rect 4338 8956 4344 8968
rect 3927 8928 4344 8956
rect 3927 8925 3939 8928
rect 3881 8919 3939 8925
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4448 8965 4476 8996
rect 4893 8993 4905 9027
rect 4939 8993 4951 9027
rect 6086 9024 6092 9036
rect 4893 8987 4951 8993
rect 5506 8996 6092 9024
rect 4433 8959 4491 8965
rect 4433 8925 4445 8959
rect 4479 8925 4491 8959
rect 4433 8919 4491 8925
rect 2332 8860 3280 8888
rect 4246 8848 4252 8900
rect 4304 8888 4310 8900
rect 4908 8888 4936 8987
rect 5074 8916 5080 8968
rect 5132 8956 5138 8968
rect 5167 8959 5225 8965
rect 5167 8956 5179 8959
rect 5132 8928 5179 8956
rect 5132 8916 5138 8928
rect 5167 8925 5179 8928
rect 5213 8925 5225 8959
rect 5167 8919 5225 8925
rect 5506 8888 5534 8996
rect 6086 8984 6092 8996
rect 6144 9024 6150 9036
rect 6457 9027 6515 9033
rect 6457 9024 6469 9027
rect 6144 8996 6469 9024
rect 6144 8984 6150 8996
rect 6457 8993 6469 8996
rect 6503 8993 6515 9027
rect 6457 8987 6515 8993
rect 6546 8984 6552 9036
rect 6604 8984 6610 9036
rect 7310 9027 7368 9033
rect 7310 9024 7322 9027
rect 6656 8996 7322 9024
rect 5810 8916 5816 8968
rect 5868 8956 5874 8968
rect 6273 8959 6331 8965
rect 6273 8956 6285 8959
rect 5868 8928 6285 8956
rect 5868 8916 5874 8928
rect 6273 8925 6285 8928
rect 6319 8956 6331 8959
rect 6362 8956 6368 8968
rect 6319 8928 6368 8956
rect 6319 8925 6331 8928
rect 6273 8919 6331 8925
rect 6362 8916 6368 8928
rect 6420 8916 6426 8968
rect 6656 8956 6684 8996
rect 7310 8993 7322 8996
rect 7356 8993 7368 9027
rect 7310 8987 7368 8993
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 7515 8996 8064 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 7208 8965 7214 8968
rect 6472 8928 6684 8956
rect 7193 8959 7214 8965
rect 4304 8860 4936 8888
rect 5276 8860 5534 8888
rect 4304 8848 4310 8860
rect 5276 8832 5304 8860
rect 5994 8848 6000 8900
rect 6052 8888 6058 8900
rect 6472 8888 6500 8928
rect 7193 8925 7205 8959
rect 7193 8919 7214 8925
rect 7208 8916 7214 8919
rect 7266 8916 7272 8968
rect 8036 8956 8064 8996
rect 8202 8984 8208 9036
rect 8260 9024 8266 9036
rect 9674 9024 9680 9036
rect 8260 8996 9680 9024
rect 8260 8984 8266 8996
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9766 8984 9772 9036
rect 9824 9024 9830 9036
rect 9968 9024 9996 9052
rect 10796 9036 10824 9064
rect 12621 9061 12633 9095
rect 12667 9092 12679 9095
rect 12710 9092 12716 9104
rect 12667 9064 12716 9092
rect 12667 9061 12679 9064
rect 12621 9055 12679 9061
rect 12710 9052 12716 9064
rect 12768 9052 12774 9104
rect 14826 9052 14832 9104
rect 14884 9092 14890 9104
rect 15378 9092 15384 9104
rect 14884 9064 15384 9092
rect 14884 9052 14890 9064
rect 15378 9052 15384 9064
rect 15436 9052 15442 9104
rect 10229 9027 10287 9033
rect 10229 9024 10241 9027
rect 9824 8996 10241 9024
rect 9824 8984 9830 8996
rect 10229 8993 10241 8996
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 10594 8984 10600 9036
rect 10652 9024 10658 9036
rect 10689 9027 10747 9033
rect 10689 9024 10701 9027
rect 10652 8996 10701 9024
rect 10652 8984 10658 8996
rect 10689 8993 10701 8996
rect 10735 8993 10747 9027
rect 10689 8987 10747 8993
rect 10778 8984 10784 9036
rect 10836 8984 10842 9036
rect 11103 9027 11161 9033
rect 11103 8993 11115 9027
rect 11149 9024 11161 9027
rect 11422 9024 11428 9036
rect 11149 8996 11428 9024
rect 11149 8993 11161 8996
rect 11103 8987 11161 8993
rect 11422 8984 11428 8996
rect 11480 8984 11486 9036
rect 11974 8984 11980 9036
rect 12032 8984 12038 9036
rect 12250 9024 12256 9036
rect 12176 8996 12256 9024
rect 8478 8956 8484 8968
rect 8036 8928 8484 8956
rect 8478 8916 8484 8928
rect 8536 8916 8542 8968
rect 9692 8956 9720 8984
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 9692 8928 9965 8956
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 10045 8959 10103 8965
rect 10045 8925 10057 8959
rect 10091 8956 10103 8959
rect 10410 8956 10416 8968
rect 10091 8928 10416 8956
rect 10091 8925 10103 8928
rect 10045 8919 10103 8925
rect 9398 8888 9404 8900
rect 6052 8860 6500 8888
rect 8036 8860 9404 8888
rect 6052 8848 6058 8860
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 3142 8820 3148 8832
rect 2556 8792 3148 8820
rect 2556 8780 2562 8792
rect 3142 8780 3148 8792
rect 3200 8780 3206 8832
rect 3329 8823 3387 8829
rect 3329 8789 3341 8823
rect 3375 8820 3387 8823
rect 3694 8820 3700 8832
rect 3375 8792 3700 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 3694 8780 3700 8792
rect 3752 8780 3758 8832
rect 5258 8780 5264 8832
rect 5316 8780 5322 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7374 8820 7380 8832
rect 6972 8792 7380 8820
rect 6972 8780 6978 8792
rect 7374 8780 7380 8792
rect 7432 8820 7438 8832
rect 8036 8820 8064 8860
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 9858 8848 9864 8900
rect 9916 8888 9922 8900
rect 10060 8888 10088 8919
rect 10410 8916 10416 8928
rect 10468 8916 10474 8968
rect 10962 8916 10968 8968
rect 11020 8916 11026 8968
rect 11238 8916 11244 8968
rect 11296 8916 11302 8968
rect 11882 8916 11888 8968
rect 11940 8956 11946 8968
rect 12176 8965 12204 8996
rect 12250 8984 12256 8996
rect 12308 8984 12314 9036
rect 12894 8984 12900 9036
rect 12952 8984 12958 9036
rect 15488 9033 15516 9132
rect 15562 9120 15568 9132
rect 15620 9160 15626 9172
rect 15620 9132 16160 9160
rect 15620 9120 15626 9132
rect 16132 9092 16160 9132
rect 16206 9120 16212 9172
rect 16264 9160 16270 9172
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 16264 9132 16497 9160
rect 16264 9120 16270 9132
rect 16485 9129 16497 9132
rect 16531 9129 16543 9163
rect 16485 9123 16543 9129
rect 16945 9163 17003 9169
rect 16945 9129 16957 9163
rect 16991 9160 17003 9163
rect 17126 9160 17132 9172
rect 16991 9132 17132 9160
rect 16991 9129 17003 9132
rect 16945 9123 17003 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 18969 9163 19027 9169
rect 17236 9132 18911 9160
rect 16132 9064 16436 9092
rect 15473 9027 15531 9033
rect 15473 9024 15485 9027
rect 14732 8996 15485 9024
rect 12161 8959 12219 8965
rect 12161 8956 12173 8959
rect 11940 8928 12173 8956
rect 11940 8916 11946 8928
rect 12161 8925 12173 8928
rect 12207 8925 12219 8959
rect 12161 8919 12219 8925
rect 12986 8916 12992 8968
rect 13044 8965 13050 8968
rect 13044 8959 13072 8965
rect 13060 8925 13072 8959
rect 13044 8919 13072 8925
rect 13044 8916 13050 8919
rect 13170 8916 13176 8968
rect 13228 8916 13234 8968
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8925 14151 8959
rect 14366 8956 14372 8968
rect 14327 8928 14372 8956
rect 14093 8919 14151 8925
rect 9916 8860 10088 8888
rect 9916 8848 9922 8860
rect 13722 8848 13728 8900
rect 13780 8888 13786 8900
rect 14108 8888 14136 8919
rect 14366 8916 14372 8928
rect 14424 8916 14430 8968
rect 14732 8888 14760 8996
rect 15473 8993 15485 8996
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 16408 8968 16436 9064
rect 17236 9024 17264 9132
rect 16940 8996 17264 9024
rect 15194 8916 15200 8968
rect 15252 8956 15258 8968
rect 15715 8959 15773 8965
rect 15715 8956 15727 8959
rect 15252 8928 15727 8956
rect 15252 8916 15258 8928
rect 15715 8925 15727 8928
rect 15761 8925 15773 8959
rect 16114 8956 16120 8968
rect 15715 8919 15773 8925
rect 15856 8928 16120 8956
rect 13780 8860 14760 8888
rect 13780 8848 13786 8860
rect 7432 8792 8064 8820
rect 8113 8823 8171 8829
rect 7432 8780 7438 8792
rect 8113 8789 8125 8823
rect 8159 8820 8171 8823
rect 8386 8820 8392 8832
rect 8159 8792 8392 8820
rect 8159 8789 8171 8792
rect 8113 8783 8171 8789
rect 8386 8780 8392 8792
rect 8444 8780 8450 8832
rect 9582 8780 9588 8832
rect 9640 8820 9646 8832
rect 9769 8823 9827 8829
rect 9769 8820 9781 8823
rect 9640 8792 9781 8820
rect 9640 8780 9646 8792
rect 9769 8789 9781 8792
rect 9815 8789 9827 8823
rect 9769 8783 9827 8789
rect 10410 8780 10416 8832
rect 10468 8820 10474 8832
rect 10870 8820 10876 8832
rect 10468 8792 10876 8820
rect 10468 8780 10474 8792
rect 10870 8780 10876 8792
rect 10928 8780 10934 8832
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 12618 8820 12624 8832
rect 11020 8792 12624 8820
rect 11020 8780 11026 8792
rect 12618 8780 12624 8792
rect 12676 8780 12682 8832
rect 13262 8780 13268 8832
rect 13320 8820 13326 8832
rect 13817 8823 13875 8829
rect 13817 8820 13829 8823
rect 13320 8792 13829 8820
rect 13320 8780 13326 8792
rect 13817 8789 13829 8792
rect 13863 8789 13875 8823
rect 13817 8783 13875 8789
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 15856 8820 15884 8928
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16390 8916 16396 8968
rect 16448 8916 16454 8968
rect 16574 8916 16580 8968
rect 16632 8956 16638 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16632 8928 16865 8956
rect 16632 8916 16638 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 16853 8919 16911 8925
rect 15930 8848 15936 8900
rect 15988 8888 15994 8900
rect 16940 8888 16968 8996
rect 17221 8959 17279 8965
rect 17221 8925 17233 8959
rect 17267 8956 17279 8959
rect 17495 8959 17553 8965
rect 17267 8928 17356 8956
rect 17267 8925 17279 8928
rect 17221 8919 17279 8925
rect 17328 8900 17356 8928
rect 17495 8925 17507 8959
rect 17541 8956 17553 8959
rect 17954 8956 17960 8968
rect 17541 8928 17960 8956
rect 17541 8925 17553 8928
rect 17495 8919 17553 8925
rect 17954 8916 17960 8928
rect 18012 8916 18018 8968
rect 18046 8916 18052 8968
rect 18104 8956 18110 8968
rect 18782 8956 18788 8968
rect 18104 8928 18788 8956
rect 18104 8916 18110 8928
rect 18782 8916 18788 8928
rect 18840 8916 18846 8968
rect 15988 8860 16968 8888
rect 15988 8848 15994 8860
rect 17310 8848 17316 8900
rect 17368 8888 17374 8900
rect 17770 8888 17776 8900
rect 17368 8860 17776 8888
rect 17368 8848 17374 8860
rect 17770 8848 17776 8860
rect 17828 8848 17834 8900
rect 18322 8888 18328 8900
rect 18156 8860 18328 8888
rect 13964 8792 15884 8820
rect 13964 8780 13970 8792
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 18156 8820 18184 8860
rect 18322 8848 18328 8860
rect 18380 8848 18386 8900
rect 18690 8848 18696 8900
rect 18748 8848 18754 8900
rect 16080 8792 18184 8820
rect 18233 8823 18291 8829
rect 16080 8780 16086 8792
rect 18233 8789 18245 8823
rect 18279 8820 18291 8823
rect 18506 8820 18512 8832
rect 18279 8792 18512 8820
rect 18279 8789 18291 8792
rect 18233 8783 18291 8789
rect 18506 8780 18512 8792
rect 18564 8780 18570 8832
rect 18883 8820 18911 9132
rect 18969 9129 18981 9163
rect 19015 9160 19027 9163
rect 20346 9160 20352 9172
rect 19015 9132 20352 9160
rect 19015 9129 19027 9132
rect 18969 9123 19027 9129
rect 20346 9120 20352 9132
rect 20404 9120 20410 9172
rect 20070 9052 20076 9104
rect 20128 9092 20134 9104
rect 20257 9095 20315 9101
rect 20257 9092 20269 9095
rect 20128 9064 20269 9092
rect 20128 9052 20134 9064
rect 20257 9061 20269 9064
rect 20303 9061 20315 9095
rect 20257 9055 20315 9061
rect 19242 8984 19248 9036
rect 19300 8984 19306 9036
rect 19518 8956 19524 8968
rect 19479 8928 19524 8956
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 19610 8820 19616 8832
rect 18883 8792 19616 8820
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 1104 8730 21043 8752
rect 1104 8678 5894 8730
rect 5946 8678 5958 8730
rect 6010 8678 6022 8730
rect 6074 8678 6086 8730
rect 6138 8678 6150 8730
rect 6202 8678 10839 8730
rect 10891 8678 10903 8730
rect 10955 8678 10967 8730
rect 11019 8678 11031 8730
rect 11083 8678 11095 8730
rect 11147 8678 15784 8730
rect 15836 8678 15848 8730
rect 15900 8678 15912 8730
rect 15964 8678 15976 8730
rect 16028 8678 16040 8730
rect 16092 8678 20729 8730
rect 20781 8678 20793 8730
rect 20845 8678 20857 8730
rect 20909 8678 20921 8730
rect 20973 8678 20985 8730
rect 21037 8678 21043 8730
rect 1104 8656 21043 8678
rect 1486 8576 1492 8628
rect 1544 8576 1550 8628
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 1854 8616 1860 8628
rect 1811 8588 1860 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 1854 8576 1860 8588
rect 1912 8576 1918 8628
rect 2958 8616 2964 8628
rect 2056 8588 2964 8616
rect 1504 8548 1532 8576
rect 2056 8557 2084 8588
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 4706 8616 4712 8628
rect 3200 8588 4712 8616
rect 3200 8576 3206 8588
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 4982 8576 4988 8628
rect 5040 8616 5046 8628
rect 5445 8619 5503 8625
rect 5445 8616 5457 8619
rect 5040 8588 5457 8616
rect 5040 8576 5046 8588
rect 5445 8585 5457 8588
rect 5491 8585 5503 8619
rect 8754 8616 8760 8628
rect 5445 8579 5503 8585
rect 6012 8588 8760 8616
rect 2041 8551 2099 8557
rect 1504 8520 1900 8548
rect 1486 8440 1492 8492
rect 1544 8440 1550 8492
rect 1872 8424 1900 8520
rect 2041 8517 2053 8551
rect 2087 8517 2099 8551
rect 2041 8511 2099 8517
rect 2498 8508 2504 8560
rect 2556 8508 2562 8560
rect 4356 8520 4568 8548
rect 2516 8480 2544 8508
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2516 8452 2697 8480
rect 2685 8449 2697 8452
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 3418 8440 3424 8492
rect 3476 8440 3482 8492
rect 3694 8440 3700 8492
rect 3752 8440 3758 8492
rect 1854 8372 1860 8424
rect 1912 8412 1918 8424
rect 2501 8415 2559 8421
rect 2501 8412 2513 8415
rect 1912 8384 2513 8412
rect 1912 8372 1918 8384
rect 2501 8381 2513 8384
rect 2547 8381 2559 8415
rect 2501 8375 2559 8381
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 2924 8384 3157 8412
rect 2924 8372 2930 8384
rect 3145 8381 3157 8384
rect 3191 8381 3203 8415
rect 3145 8375 3203 8381
rect 3559 8415 3617 8421
rect 3559 8381 3571 8415
rect 3605 8412 3617 8415
rect 4062 8412 4068 8424
rect 3605 8384 4068 8412
rect 3605 8381 3617 8384
rect 3559 8375 3617 8381
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4356 8412 4384 8520
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 4540 8480 4568 8520
rect 4707 8483 4765 8489
rect 4707 8480 4719 8483
rect 4540 8452 4719 8480
rect 4707 8449 4719 8452
rect 4753 8480 4765 8483
rect 4753 8452 5212 8480
rect 4753 8449 4765 8452
rect 4707 8443 4765 8449
rect 4264 8384 4384 8412
rect 5184 8412 5212 8452
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 5902 8480 5908 8492
rect 5776 8452 5908 8480
rect 5776 8440 5782 8452
rect 5902 8440 5908 8452
rect 5960 8440 5966 8492
rect 6012 8489 6040 8588
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 9398 8616 9404 8628
rect 9263 8588 9404 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9398 8576 9404 8588
rect 9456 8576 9462 8628
rect 9490 8576 9496 8628
rect 9548 8576 9554 8628
rect 10410 8616 10416 8628
rect 10152 8588 10416 8616
rect 6086 8508 6092 8560
rect 6144 8548 6150 8560
rect 6144 8520 6742 8548
rect 6144 8508 6150 8520
rect 5997 8483 6055 8489
rect 5997 8449 6009 8483
rect 6043 8449 6055 8483
rect 6607 8483 6665 8489
rect 6607 8480 6619 8483
rect 5997 8443 6055 8449
rect 6104 8452 6619 8480
rect 6104 8412 6132 8452
rect 6607 8449 6619 8452
rect 6653 8449 6665 8483
rect 6714 8480 6742 8520
rect 7742 8508 7748 8560
rect 7800 8508 7806 8560
rect 7834 8508 7840 8560
rect 7892 8548 7898 8560
rect 8294 8557 8300 8560
rect 7929 8551 7987 8557
rect 7929 8548 7941 8551
rect 7892 8520 7941 8548
rect 7892 8508 7898 8520
rect 7929 8517 7941 8520
rect 7975 8517 7987 8551
rect 7929 8511 7987 8517
rect 8285 8551 8300 8557
rect 8285 8517 8297 8551
rect 8285 8511 8300 8517
rect 8294 8508 8300 8511
rect 8352 8508 8358 8560
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 9033 8551 9091 8557
rect 9033 8548 9045 8551
rect 8536 8520 9045 8548
rect 8536 8508 8542 8520
rect 9033 8517 9045 8520
rect 9079 8517 9091 8551
rect 9033 8511 9091 8517
rect 7760 8480 7788 8508
rect 6714 8452 7788 8480
rect 8205 8483 8263 8489
rect 6607 8443 6665 8449
rect 8205 8449 8217 8483
rect 8251 8480 8263 8483
rect 8570 8480 8576 8492
rect 8251 8452 8576 8480
rect 8251 8449 8263 8452
rect 8205 8443 8263 8449
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 9508 8480 9536 8576
rect 10152 8519 10180 8588
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 10873 8619 10931 8625
rect 10873 8616 10885 8619
rect 10744 8588 10885 8616
rect 10744 8576 10750 8588
rect 10873 8585 10885 8588
rect 10919 8585 10931 8619
rect 10873 8579 10931 8585
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 15102 8616 15108 8628
rect 11112 8588 15108 8616
rect 11112 8576 11118 8588
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15197 8619 15255 8625
rect 15197 8585 15209 8619
rect 15243 8585 15255 8619
rect 15197 8579 15255 8585
rect 10119 8513 10180 8519
rect 9769 8483 9827 8489
rect 9769 8480 9781 8483
rect 9508 8452 9781 8480
rect 9769 8449 9781 8452
rect 9815 8449 9827 8483
rect 10119 8479 10131 8513
rect 10165 8482 10180 8513
rect 10318 8508 10324 8560
rect 10376 8548 10382 8560
rect 10376 8520 11100 8548
rect 10376 8508 10382 8520
rect 10165 8479 10177 8482
rect 10119 8473 10177 8479
rect 11072 8480 11100 8520
rect 11422 8508 11428 8560
rect 11480 8548 11486 8560
rect 15212 8548 15240 8579
rect 15470 8576 15476 8628
rect 15528 8616 15534 8628
rect 16206 8616 16212 8628
rect 15528 8588 16212 8616
rect 15528 8576 15534 8588
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16393 8619 16451 8625
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 16666 8616 16672 8628
rect 16439 8588 16672 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16666 8576 16672 8588
rect 16724 8576 16730 8628
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8616 16911 8619
rect 16899 8588 17172 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 11480 8520 15240 8548
rect 15304 8520 15792 8548
rect 11480 8508 11486 8520
rect 12066 8480 12072 8492
rect 11072 8452 12072 8480
rect 9769 8443 9827 8449
rect 12066 8440 12072 8452
rect 12124 8440 12130 8492
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12495 8483 12553 8489
rect 12495 8480 12507 8483
rect 12216 8452 12507 8480
rect 12216 8440 12222 8452
rect 12495 8449 12507 8452
rect 12541 8449 12553 8483
rect 12495 8443 12553 8449
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 13538 8480 13544 8492
rect 12676 8452 13544 8480
rect 12676 8440 12682 8452
rect 13004 8424 13032 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8449 13691 8483
rect 13633 8443 13691 8449
rect 5184 8384 6132 8412
rect 566 8304 572 8356
rect 624 8344 630 8356
rect 624 8316 2544 8344
rect 624 8304 630 8316
rect 2516 8288 2544 8316
rect 1026 8236 1032 8288
rect 1084 8276 1090 8288
rect 2133 8279 2191 8285
rect 2133 8276 2145 8279
rect 1084 8248 2145 8276
rect 1084 8236 1090 8248
rect 2133 8245 2145 8248
rect 2179 8245 2191 8279
rect 2133 8239 2191 8245
rect 2498 8236 2504 8288
rect 2556 8236 2562 8288
rect 2866 8236 2872 8288
rect 2924 8276 2930 8288
rect 4264 8276 4292 8384
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6236 8384 6377 8412
rect 6236 8372 6242 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5092 8316 5825 8344
rect 2924 8248 4292 8276
rect 2924 8236 2930 8248
rect 4338 8236 4344 8288
rect 4396 8236 4402 8288
rect 4522 8236 4528 8288
rect 4580 8276 4586 8288
rect 5092 8276 5120 8316
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 5813 8307 5871 8313
rect 7377 8347 7435 8353
rect 7377 8313 7389 8347
rect 7423 8344 7435 8347
rect 7760 8344 7788 8398
rect 9306 8372 9312 8424
rect 9364 8412 9370 8424
rect 9861 8415 9919 8421
rect 9861 8412 9873 8415
rect 9364 8384 9873 8412
rect 9364 8372 9370 8384
rect 9861 8381 9873 8384
rect 9907 8381 9919 8415
rect 9861 8375 9919 8381
rect 7423 8316 7788 8344
rect 7423 8313 7435 8316
rect 7377 8307 7435 8313
rect 4580 8248 5120 8276
rect 4580 8236 4586 8248
rect 5166 8236 5172 8288
rect 5224 8276 5230 8288
rect 7742 8276 7748 8288
rect 5224 8248 7748 8276
rect 5224 8236 5230 8248
rect 7742 8236 7748 8248
rect 7800 8236 7806 8288
rect 9582 8236 9588 8288
rect 9640 8236 9646 8288
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 9876 8276 9904 8375
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 11606 8412 11612 8424
rect 10744 8384 11612 8412
rect 10744 8372 10750 8384
rect 11606 8372 11612 8384
rect 11664 8372 11670 8424
rect 12253 8415 12311 8421
rect 12253 8381 12265 8415
rect 12299 8381 12311 8415
rect 12253 8375 12311 8381
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 11882 8344 11888 8356
rect 11204 8316 11888 8344
rect 11204 8304 11210 8316
rect 11882 8304 11888 8316
rect 11940 8304 11946 8356
rect 12066 8304 12072 8356
rect 12124 8344 12130 8356
rect 12268 8344 12296 8375
rect 12986 8372 12992 8424
rect 13044 8372 13050 8424
rect 13170 8372 13176 8424
rect 13228 8372 13234 8424
rect 12124 8316 12296 8344
rect 13188 8344 13216 8372
rect 13648 8356 13676 8443
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 13907 8483 13965 8489
rect 13907 8480 13919 8483
rect 13872 8452 13919 8480
rect 13872 8440 13878 8452
rect 13907 8449 13919 8452
rect 13953 8449 13965 8483
rect 13907 8443 13965 8449
rect 14366 8440 14372 8492
rect 14424 8480 14430 8492
rect 15194 8480 15200 8492
rect 14424 8452 15200 8480
rect 14424 8440 14430 8452
rect 15194 8440 15200 8452
rect 15252 8440 15258 8492
rect 13265 8347 13323 8353
rect 13265 8344 13277 8347
rect 13188 8316 13277 8344
rect 12124 8304 12130 8316
rect 13265 8313 13277 8316
rect 13311 8313 13323 8347
rect 13630 8344 13636 8356
rect 13265 8307 13323 8313
rect 13370 8316 13636 8344
rect 13370 8276 13398 8316
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 9824 8248 13398 8276
rect 9824 8236 9830 8248
rect 13446 8236 13452 8288
rect 13504 8276 13510 8288
rect 14645 8279 14703 8285
rect 14645 8276 14657 8279
rect 13504 8248 14657 8276
rect 13504 8236 13510 8248
rect 14645 8245 14657 8248
rect 14691 8245 14703 8279
rect 15304 8276 15332 8520
rect 15381 8483 15439 8489
rect 15381 8449 15393 8483
rect 15427 8449 15439 8483
rect 15381 8443 15439 8449
rect 15396 8344 15424 8443
rect 15470 8440 15476 8492
rect 15528 8480 15534 8492
rect 15764 8489 15792 8520
rect 15838 8508 15844 8560
rect 15896 8508 15902 8560
rect 16114 8508 16120 8560
rect 16172 8548 16178 8560
rect 17144 8548 17172 8588
rect 17218 8576 17224 8628
rect 17276 8616 17282 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 17276 8588 17325 8616
rect 17276 8576 17282 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 20533 8619 20591 8625
rect 20533 8616 20545 8619
rect 17460 8588 20545 8616
rect 17460 8576 17466 8588
rect 20533 8585 20545 8588
rect 20579 8585 20591 8619
rect 20533 8579 20591 8585
rect 17586 8548 17592 8560
rect 16172 8520 16988 8548
rect 17144 8520 17592 8548
rect 16172 8508 16178 8520
rect 15657 8483 15715 8489
rect 15657 8480 15669 8483
rect 15528 8452 15669 8480
rect 15528 8440 15534 8452
rect 15657 8449 15669 8452
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15856 8480 15884 8508
rect 16209 8483 16267 8489
rect 16209 8480 16221 8483
rect 15856 8452 16221 8480
rect 15749 8443 15807 8449
rect 16209 8449 16221 8452
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 16298 8440 16304 8492
rect 16356 8440 16362 8492
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8480 16727 8483
rect 16758 8480 16764 8492
rect 16715 8452 16764 8480
rect 16715 8449 16727 8452
rect 16669 8443 16727 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 16960 8489 16988 8520
rect 17586 8508 17592 8520
rect 17644 8508 17650 8560
rect 17862 8508 17868 8560
rect 17920 8548 17926 8560
rect 19426 8557 19432 8560
rect 19420 8548 19432 8557
rect 17920 8520 19196 8548
rect 19387 8520 19432 8548
rect 17920 8508 17926 8520
rect 16853 8483 16911 8489
rect 16853 8449 16865 8483
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 16945 8483 17003 8489
rect 16945 8449 16957 8483
rect 16991 8449 17003 8483
rect 16945 8443 17003 8449
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 15838 8372 15844 8424
rect 15896 8412 15902 8424
rect 16868 8412 16896 8443
rect 15896 8384 16896 8412
rect 17037 8415 17095 8421
rect 15896 8372 15902 8384
rect 17037 8381 17049 8415
rect 17083 8412 17095 8415
rect 17126 8412 17132 8424
rect 17083 8384 17132 8412
rect 17083 8381 17095 8384
rect 17037 8375 17095 8381
rect 17126 8372 17132 8384
rect 17184 8372 17190 8424
rect 17402 8372 17408 8424
rect 17460 8372 17466 8424
rect 17420 8344 17448 8372
rect 15396 8316 17448 8344
rect 17512 8344 17540 8443
rect 17770 8440 17776 8492
rect 17828 8440 17834 8492
rect 18015 8483 18073 8489
rect 18015 8449 18027 8483
rect 18061 8480 18073 8483
rect 18598 8480 18604 8492
rect 18061 8452 18604 8480
rect 18061 8449 18073 8452
rect 18015 8443 18073 8449
rect 18598 8440 18604 8452
rect 18656 8440 18662 8492
rect 19168 8489 19196 8520
rect 19420 8511 19432 8520
rect 19426 8508 19432 8511
rect 19484 8508 19490 8560
rect 19702 8508 19708 8560
rect 19760 8508 19766 8560
rect 19153 8483 19211 8489
rect 18708 8452 18900 8480
rect 18506 8372 18512 8424
rect 18564 8412 18570 8424
rect 18708 8412 18736 8452
rect 18564 8384 18736 8412
rect 18872 8412 18900 8452
rect 19153 8449 19165 8483
rect 19199 8449 19211 8483
rect 19720 8480 19748 8508
rect 19153 8443 19211 8449
rect 19260 8452 19748 8480
rect 19260 8412 19288 8452
rect 18872 8384 19288 8412
rect 18564 8372 18570 8384
rect 17512 8316 17816 8344
rect 15473 8279 15531 8285
rect 15473 8276 15485 8279
rect 15304 8248 15485 8276
rect 14645 8239 14703 8245
rect 15473 8245 15485 8248
rect 15519 8245 15531 8279
rect 15473 8239 15531 8245
rect 15654 8236 15660 8288
rect 15712 8276 15718 8288
rect 15841 8279 15899 8285
rect 15841 8276 15853 8279
rect 15712 8248 15853 8276
rect 15712 8236 15718 8248
rect 15841 8245 15853 8248
rect 15887 8245 15899 8279
rect 15841 8239 15899 8245
rect 16025 8279 16083 8285
rect 16025 8245 16037 8279
rect 16071 8276 16083 8279
rect 17126 8276 17132 8288
rect 16071 8248 17132 8276
rect 16071 8245 16083 8248
rect 16025 8239 16083 8245
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 17402 8236 17408 8288
rect 17460 8276 17466 8288
rect 17678 8276 17684 8288
rect 17460 8248 17684 8276
rect 17460 8236 17466 8248
rect 17678 8236 17684 8248
rect 17736 8236 17742 8288
rect 17788 8276 17816 8316
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 18840 8316 19196 8344
rect 18840 8304 18846 8316
rect 18138 8276 18144 8288
rect 17788 8248 18144 8276
rect 18138 8236 18144 8248
rect 18196 8236 18202 8288
rect 19168 8276 19196 8316
rect 19518 8276 19524 8288
rect 19168 8248 19524 8276
rect 19518 8236 19524 8248
rect 19576 8236 19582 8288
rect 1104 8186 20884 8208
rect 1104 8134 3422 8186
rect 3474 8134 3486 8186
rect 3538 8134 3550 8186
rect 3602 8134 3614 8186
rect 3666 8134 3678 8186
rect 3730 8134 8367 8186
rect 8419 8134 8431 8186
rect 8483 8134 8495 8186
rect 8547 8134 8559 8186
rect 8611 8134 8623 8186
rect 8675 8134 13312 8186
rect 13364 8134 13376 8186
rect 13428 8134 13440 8186
rect 13492 8134 13504 8186
rect 13556 8134 13568 8186
rect 13620 8134 18257 8186
rect 18309 8134 18321 8186
rect 18373 8134 18385 8186
rect 18437 8134 18449 8186
rect 18501 8134 18513 8186
rect 18565 8134 20884 8186
rect 1104 8112 20884 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 1946 8072 1952 8084
rect 1811 8044 1952 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 3329 8075 3387 8081
rect 2332 8044 3004 8072
rect 1394 7896 1400 7948
rect 1452 7936 1458 7948
rect 2332 7945 2360 8044
rect 2317 7939 2375 7945
rect 1452 7908 2176 7936
rect 1452 7896 1458 7908
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7868 1547 7871
rect 2038 7868 2044 7880
rect 1535 7840 2044 7868
rect 1535 7837 1547 7840
rect 1489 7831 1547 7837
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2148 7877 2176 7908
rect 2317 7905 2329 7939
rect 2363 7905 2375 7939
rect 2976 7936 3004 8044
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 4154 8072 4160 8084
rect 3375 8044 4160 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 5166 8032 5172 8084
rect 5224 8072 5230 8084
rect 5224 8044 5534 8072
rect 5224 8032 5230 8044
rect 3510 7964 3516 8016
rect 3568 8004 3574 8016
rect 3878 8004 3884 8016
rect 3568 7976 3884 8004
rect 3568 7964 3574 7976
rect 3878 7964 3884 7976
rect 3936 7964 3942 8016
rect 4126 7976 4292 8004
rect 4126 7936 4154 7976
rect 4264 7948 4292 7976
rect 2976 7908 4154 7936
rect 2317 7899 2375 7905
rect 3252 7880 3280 7908
rect 4246 7896 4252 7948
rect 4304 7936 4310 7948
rect 4709 7939 4767 7945
rect 4709 7936 4721 7939
rect 4304 7908 4721 7936
rect 4304 7896 4310 7908
rect 4709 7905 4721 7908
rect 4755 7905 4767 7939
rect 5506 7936 5534 8044
rect 5718 8032 5724 8084
rect 5776 8032 5782 8084
rect 6178 8032 6184 8084
rect 6236 8072 6242 8084
rect 6546 8072 6552 8084
rect 6236 8044 6552 8072
rect 6236 8032 6242 8044
rect 6546 8032 6552 8044
rect 6604 8072 6610 8084
rect 6604 8044 7328 8072
rect 6604 8032 6610 8044
rect 5506 7908 5672 7936
rect 4709 7899 4767 7905
rect 5644 7880 5672 7908
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6086 7936 6092 7948
rect 5868 7908 6092 7936
rect 5868 7896 5874 7908
rect 6086 7896 6092 7908
rect 6144 7896 6150 7948
rect 7300 7936 7328 8044
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 8481 8075 8539 8081
rect 8481 8072 8493 8075
rect 8352 8044 8493 8072
rect 8352 8032 8358 8044
rect 8481 8041 8493 8044
rect 8527 8041 8539 8075
rect 9214 8072 9220 8084
rect 8481 8035 8539 8041
rect 8956 8044 9220 8072
rect 8956 7945 8984 8044
rect 9214 8032 9220 8044
rect 9272 8032 9278 8084
rect 9674 8032 9680 8084
rect 9732 8072 9738 8084
rect 9950 8072 9956 8084
rect 9732 8044 9956 8072
rect 9732 8032 9738 8044
rect 9950 8032 9956 8044
rect 10008 8032 10014 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10836 8044 11192 8072
rect 10836 8032 10842 8044
rect 11164 8004 11192 8044
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 11517 8075 11575 8081
rect 11517 8072 11529 8075
rect 11296 8044 11529 8072
rect 11296 8032 11302 8044
rect 11517 8041 11529 8044
rect 11563 8041 11575 8075
rect 13906 8072 13912 8084
rect 11517 8035 11575 8041
rect 11624 8044 13912 8072
rect 11624 8004 11652 8044
rect 13906 8032 13912 8044
rect 13964 8032 13970 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 13998 8044 15117 8072
rect 11164 7976 11652 8004
rect 11826 7976 12570 8004
rect 7469 7939 7527 7945
rect 7469 7936 7481 7939
rect 7300 7908 7481 7936
rect 7469 7905 7481 7908
rect 7515 7905 7527 7939
rect 8941 7939 8999 7945
rect 7469 7899 7527 7905
rect 2133 7871 2191 7877
rect 2133 7837 2145 7871
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2591 7871 2649 7877
rect 2591 7837 2603 7871
rect 2637 7868 2649 7871
rect 2637 7840 3188 7868
rect 2637 7837 2649 7840
rect 2591 7831 2649 7837
rect 1394 7760 1400 7812
rect 1452 7760 1458 7812
rect 1854 7760 1860 7812
rect 1912 7800 1918 7812
rect 3160 7800 3188 7840
rect 3234 7828 3240 7880
rect 3292 7828 3298 7880
rect 4890 7868 4896 7880
rect 4172 7840 4896 7868
rect 3510 7800 3516 7812
rect 1912 7772 2820 7800
rect 3160 7772 3516 7800
rect 1912 7760 1918 7772
rect 1412 7732 1440 7760
rect 1949 7735 2007 7741
rect 1949 7732 1961 7735
rect 1412 7704 1961 7732
rect 1949 7701 1961 7704
rect 1995 7701 2007 7735
rect 2792 7732 2820 7772
rect 3510 7760 3516 7772
rect 3568 7760 3574 7812
rect 3881 7803 3939 7809
rect 3881 7769 3893 7803
rect 3927 7800 3939 7803
rect 4172 7800 4200 7840
rect 4890 7828 4896 7840
rect 4948 7828 4954 7880
rect 4983 7871 5041 7877
rect 4983 7837 4995 7871
rect 5029 7868 5041 7871
rect 5534 7868 5540 7880
rect 5029 7840 5540 7868
rect 5029 7837 5041 7840
rect 4983 7831 5041 7837
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 6363 7871 6421 7877
rect 5736 7840 6316 7868
rect 3927 7772 4200 7800
rect 4249 7803 4307 7809
rect 3927 7769 3939 7772
rect 3881 7763 3939 7769
rect 4249 7769 4261 7803
rect 4295 7800 4307 7803
rect 5736 7800 5764 7840
rect 5994 7800 6000 7812
rect 4295 7772 5764 7800
rect 5828 7772 6000 7800
rect 4295 7769 4307 7772
rect 4249 7763 4307 7769
rect 2866 7732 2872 7744
rect 2792 7704 2872 7732
rect 1949 7695 2007 7701
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 3973 7735 4031 7741
rect 3973 7732 3985 7735
rect 3384 7704 3985 7732
rect 3384 7692 3390 7704
rect 3973 7701 3985 7704
rect 4019 7701 4031 7735
rect 3973 7695 4031 7701
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 4341 7735 4399 7741
rect 4341 7732 4353 7735
rect 4120 7704 4353 7732
rect 4120 7692 4126 7704
rect 4341 7701 4353 7704
rect 4387 7701 4399 7735
rect 4341 7695 4399 7701
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 5828 7732 5856 7772
rect 5994 7760 6000 7772
rect 6052 7760 6058 7812
rect 6288 7800 6316 7840
rect 6363 7837 6375 7871
rect 6409 7868 6421 7871
rect 7006 7868 7012 7880
rect 6409 7840 7012 7868
rect 6409 7837 6421 7840
rect 6363 7831 6421 7837
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7742 7877 7748 7880
rect 7711 7871 7748 7877
rect 7711 7837 7723 7871
rect 7711 7831 7748 7837
rect 7742 7828 7748 7831
rect 7800 7828 7806 7880
rect 8110 7862 8116 7914
rect 8168 7868 8174 7914
rect 8941 7905 8953 7939
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 9766 7896 9772 7948
rect 9824 7936 9830 7948
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 9824 7908 10517 7936
rect 9824 7896 9830 7908
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 10505 7899 10563 7905
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 11826 7936 11854 7976
rect 11572 7908 11854 7936
rect 11572 7896 11578 7908
rect 11882 7896 11888 7948
rect 11940 7936 11946 7948
rect 12069 7939 12127 7945
rect 12069 7936 12081 7939
rect 11940 7908 12081 7936
rect 11940 7896 11946 7908
rect 12069 7905 12081 7908
rect 12115 7936 12127 7939
rect 12434 7936 12440 7948
rect 12115 7908 12440 7936
rect 12115 7905 12127 7908
rect 12069 7899 12127 7905
rect 12434 7896 12440 7908
rect 12492 7896 12498 7948
rect 12542 7936 12570 7976
rect 12710 7964 12716 8016
rect 12768 7964 12774 8016
rect 13998 8004 14026 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 15838 8032 15844 8084
rect 15896 8072 15902 8084
rect 15933 8075 15991 8081
rect 15933 8072 15945 8075
rect 15896 8044 15945 8072
rect 15896 8032 15902 8044
rect 15933 8041 15945 8044
rect 15979 8041 15991 8075
rect 15933 8035 15991 8041
rect 16114 8032 16120 8084
rect 16172 8072 16178 8084
rect 16209 8075 16267 8081
rect 16209 8072 16221 8075
rect 16172 8044 16221 8072
rect 16172 8032 16178 8044
rect 16209 8041 16221 8044
rect 16255 8041 16267 8075
rect 16666 8072 16672 8084
rect 16209 8035 16267 8041
rect 16500 8044 16672 8072
rect 16500 8004 16528 8044
rect 16666 8032 16672 8044
rect 16724 8032 16730 8084
rect 16758 8032 16764 8084
rect 16816 8072 16822 8084
rect 16816 8044 17540 8072
rect 16816 8032 16822 8044
rect 13740 7976 14026 8004
rect 14936 7976 16528 8004
rect 12802 7936 12808 7948
rect 12542 7908 12808 7936
rect 12802 7896 12808 7908
rect 12860 7936 12866 7948
rect 13106 7939 13164 7945
rect 13106 7936 13118 7939
rect 12860 7908 13118 7936
rect 12860 7896 12866 7908
rect 13106 7905 13118 7908
rect 13152 7905 13164 7939
rect 13106 7899 13164 7905
rect 13265 7939 13323 7945
rect 13265 7905 13277 7939
rect 13311 7936 13323 7939
rect 13740 7936 13768 7976
rect 13311 7908 13768 7936
rect 13311 7905 13323 7908
rect 13265 7899 13323 7905
rect 13814 7896 13820 7948
rect 13872 7936 13878 7948
rect 14093 7939 14151 7945
rect 14093 7936 14105 7939
rect 13872 7908 14105 7936
rect 13872 7896 13878 7908
rect 14093 7905 14105 7908
rect 14139 7905 14151 7939
rect 14093 7899 14151 7905
rect 8294 7868 8300 7880
rect 8168 7862 8300 7868
rect 8128 7840 8300 7862
rect 8294 7828 8300 7840
rect 8352 7828 8358 7880
rect 9215 7871 9273 7877
rect 9215 7837 9227 7871
rect 9261 7868 9273 7871
rect 9306 7868 9312 7880
rect 9261 7840 9312 7868
rect 9261 7837 9273 7840
rect 9215 7831 9273 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 10686 7868 10692 7880
rect 9416 7840 10692 7868
rect 7834 7800 7840 7812
rect 6288 7772 7840 7800
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 7926 7760 7932 7812
rect 7984 7800 7990 7812
rect 8110 7800 8116 7812
rect 7984 7772 8116 7800
rect 7984 7760 7990 7772
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 9416 7800 9444 7840
rect 10686 7828 10692 7840
rect 10744 7828 10750 7880
rect 12158 7868 12164 7880
rect 10779 7861 10837 7867
rect 10779 7827 10791 7861
rect 10825 7858 10837 7861
rect 10888 7858 12164 7868
rect 10825 7840 12164 7858
rect 10825 7830 10916 7840
rect 10825 7827 10837 7830
rect 12158 7828 12164 7840
rect 12216 7828 12222 7880
rect 12253 7871 12311 7877
rect 12253 7837 12265 7871
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 10779 7821 10837 7827
rect 8220 7772 9444 7800
rect 4948 7704 5856 7732
rect 4948 7692 4954 7704
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 7006 7732 7012 7744
rect 5960 7704 7012 7732
rect 5960 7692 5966 7704
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 7101 7735 7159 7741
rect 7101 7701 7113 7735
rect 7147 7732 7159 7735
rect 7466 7732 7472 7744
rect 7147 7704 7472 7732
rect 7147 7701 7159 7704
rect 7101 7695 7159 7701
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 7650 7692 7656 7744
rect 7708 7732 7714 7744
rect 8220 7732 8248 7772
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 9732 7772 10070 7800
rect 9732 7760 9738 7772
rect 7708 7704 8248 7732
rect 7708 7692 7714 7704
rect 9214 7692 9220 7744
rect 9272 7732 9278 7744
rect 9953 7735 10011 7741
rect 9953 7732 9965 7735
rect 9272 7704 9965 7732
rect 9272 7692 9278 7704
rect 9953 7701 9965 7704
rect 9999 7701 10011 7735
rect 10042 7732 10070 7772
rect 11790 7760 11796 7812
rect 11848 7800 11854 7812
rect 12268 7800 12296 7831
rect 12986 7828 12992 7880
rect 13044 7828 13050 7880
rect 14367 7871 14425 7877
rect 14367 7837 14379 7871
rect 14413 7868 14425 7871
rect 14734 7868 14740 7880
rect 14413 7840 14740 7868
rect 14413 7837 14425 7840
rect 14367 7831 14425 7837
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 14936 7800 14964 7976
rect 15010 7896 15016 7948
rect 15068 7936 15074 7948
rect 15068 7908 16436 7936
rect 15068 7896 15074 7908
rect 15470 7828 15476 7880
rect 15528 7828 15534 7880
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7868 15715 7871
rect 15930 7868 15936 7880
rect 15703 7840 15936 7868
rect 15703 7837 15715 7840
rect 15657 7831 15715 7837
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 16408 7877 16436 7908
rect 16482 7896 16488 7948
rect 16540 7896 16546 7948
rect 16117 7871 16175 7877
rect 16117 7837 16129 7871
rect 16163 7837 16175 7871
rect 16117 7831 16175 7837
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7868 16451 7871
rect 16741 7871 16799 7877
rect 16741 7868 16753 7871
rect 16439 7840 16753 7868
rect 16439 7837 16451 7840
rect 16393 7831 16451 7837
rect 16741 7837 16753 7840
rect 16787 7837 16799 7871
rect 17512 7868 17540 8044
rect 18874 7964 18880 8016
rect 18932 7964 18938 8016
rect 19886 7964 19892 8016
rect 19944 8004 19950 8016
rect 20073 8007 20131 8013
rect 20073 8004 20085 8007
rect 19944 7976 20085 8004
rect 19944 7964 19950 7976
rect 20073 7973 20085 7976
rect 20119 7973 20131 8007
rect 20073 7967 20131 7973
rect 17586 7896 17592 7948
rect 17644 7936 17650 7948
rect 19429 7939 19487 7945
rect 17644 7908 18828 7936
rect 17644 7896 17650 7908
rect 17678 7868 17684 7880
rect 17512 7840 17684 7868
rect 16741 7831 16799 7837
rect 11848 7772 12296 7800
rect 13832 7772 14964 7800
rect 16132 7800 16160 7831
rect 17678 7828 17684 7840
rect 17736 7868 17742 7880
rect 17957 7871 18015 7877
rect 17957 7868 17969 7871
rect 17736 7840 17969 7868
rect 17736 7828 17742 7840
rect 17957 7837 17969 7840
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 18230 7828 18236 7880
rect 18288 7868 18294 7880
rect 18800 7877 18828 7908
rect 19429 7905 19441 7939
rect 19475 7936 19487 7939
rect 19518 7936 19524 7948
rect 19475 7908 19524 7936
rect 19475 7905 19487 7908
rect 19429 7899 19487 7905
rect 19518 7896 19524 7908
rect 19576 7896 19582 7948
rect 18325 7871 18383 7877
rect 18325 7868 18337 7871
rect 18288 7840 18337 7868
rect 18288 7828 18294 7840
rect 18325 7837 18337 7840
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18785 7871 18843 7877
rect 18785 7837 18797 7871
rect 18831 7837 18843 7871
rect 18785 7831 18843 7837
rect 19610 7828 19616 7880
rect 19668 7828 19674 7880
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19944 7840 20085 7868
rect 19944 7828 19950 7840
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 16132 7772 18000 7800
rect 11848 7760 11854 7772
rect 11054 7732 11060 7744
rect 10042 7704 11060 7732
rect 9953 7695 10011 7701
rect 11054 7692 11060 7704
rect 11112 7692 11118 7744
rect 11974 7692 11980 7744
rect 12032 7732 12038 7744
rect 13832 7732 13860 7772
rect 12032 7704 13860 7732
rect 13909 7735 13967 7741
rect 12032 7692 12038 7704
rect 13909 7701 13921 7735
rect 13955 7732 13967 7735
rect 13998 7732 14004 7744
rect 13955 7704 14004 7732
rect 13955 7701 13967 7704
rect 13909 7695 13967 7701
rect 13998 7692 14004 7704
rect 14056 7692 14062 7744
rect 15654 7692 15660 7744
rect 15712 7692 15718 7744
rect 15746 7692 15752 7744
rect 15804 7732 15810 7744
rect 16298 7732 16304 7744
rect 15804 7704 16304 7732
rect 15804 7692 15810 7704
rect 16298 7692 16304 7704
rect 16356 7692 16362 7744
rect 16666 7692 16672 7744
rect 16724 7732 16730 7744
rect 17770 7732 17776 7744
rect 16724 7704 17776 7732
rect 16724 7692 16730 7704
rect 17770 7692 17776 7704
rect 17828 7692 17834 7744
rect 17865 7735 17923 7741
rect 17865 7701 17877 7735
rect 17911 7732 17923 7735
rect 17972 7732 18000 7772
rect 17911 7704 18000 7732
rect 17911 7701 17923 7704
rect 17865 7695 17923 7701
rect 18046 7692 18052 7744
rect 18104 7732 18110 7744
rect 18782 7732 18788 7744
rect 18104 7704 18788 7732
rect 18104 7692 18110 7704
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19610 7732 19616 7744
rect 19392 7704 19616 7732
rect 19392 7692 19398 7704
rect 19610 7692 19616 7704
rect 19668 7692 19674 7744
rect 1104 7642 21043 7664
rect 290 7556 296 7608
rect 348 7596 354 7608
rect 658 7596 664 7608
rect 348 7568 664 7596
rect 348 7556 354 7568
rect 658 7556 664 7568
rect 716 7556 722 7608
rect 1104 7590 5894 7642
rect 5946 7590 5958 7642
rect 6010 7590 6022 7642
rect 6074 7590 6086 7642
rect 6138 7590 6150 7642
rect 6202 7590 10839 7642
rect 10891 7590 10903 7642
rect 10955 7590 10967 7642
rect 11019 7590 11031 7642
rect 11083 7590 11095 7642
rect 11147 7590 15784 7642
rect 15836 7590 15848 7642
rect 15900 7590 15912 7642
rect 15964 7590 15976 7642
rect 16028 7590 16040 7642
rect 16092 7590 20729 7642
rect 20781 7590 20793 7642
rect 20845 7590 20857 7642
rect 20909 7590 20921 7642
rect 20973 7590 20985 7642
rect 21037 7590 21043 7642
rect 21358 7624 21364 7676
rect 21416 7664 21422 7676
rect 21416 7636 21496 7664
rect 21416 7624 21422 7636
rect 1104 7568 21043 7590
rect 750 7488 756 7540
rect 808 7528 814 7540
rect 1118 7528 1124 7540
rect 808 7500 1124 7528
rect 808 7488 814 7500
rect 1118 7488 1124 7500
rect 1176 7488 1182 7540
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 2590 7528 2596 7540
rect 1443 7500 2596 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 2590 7488 2596 7500
rect 2648 7488 2654 7540
rect 2685 7531 2743 7537
rect 2685 7497 2697 7531
rect 2731 7528 2743 7531
rect 3050 7528 3056 7540
rect 2731 7500 3056 7528
rect 2731 7497 2743 7500
rect 2685 7491 2743 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 3142 7488 3148 7540
rect 3200 7528 3206 7540
rect 3973 7531 4031 7537
rect 3973 7528 3985 7531
rect 3200 7500 3985 7528
rect 3200 7488 3206 7500
rect 3973 7497 3985 7500
rect 4019 7497 4031 7531
rect 3973 7491 4031 7497
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 4396 7500 6592 7528
rect 4396 7488 4402 7500
rect 2222 7460 2228 7472
rect 1596 7432 2228 7460
rect 1596 7401 1624 7432
rect 2222 7420 2228 7432
rect 2280 7420 2286 7472
rect 3329 7463 3387 7469
rect 3329 7429 3341 7463
rect 3375 7460 3387 7463
rect 4522 7460 4528 7472
rect 3375 7432 4528 7460
rect 3375 7429 3387 7432
rect 3329 7423 3387 7429
rect 4522 7420 4528 7432
rect 4580 7420 4586 7472
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7361 1639 7395
rect 1581 7355 1639 7361
rect 1854 7352 1860 7404
rect 1912 7392 1918 7404
rect 1947 7395 2005 7401
rect 1947 7392 1959 7395
rect 1912 7364 1959 7392
rect 1912 7352 1918 7364
rect 1947 7361 1959 7364
rect 1993 7361 2005 7395
rect 1947 7355 2005 7361
rect 3878 7352 3884 7404
rect 3936 7352 3942 7404
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4341 7395 4399 7401
rect 4341 7392 4353 7395
rect 4212 7364 4353 7392
rect 4212 7352 4218 7364
rect 4341 7361 4353 7364
rect 4387 7361 4399 7395
rect 4341 7355 4399 7361
rect 5258 7352 5264 7404
rect 5316 7352 5322 7404
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 6178 7352 6184 7404
rect 6236 7392 6242 7404
rect 6454 7392 6460 7404
rect 6236 7364 6460 7392
rect 6236 7352 6242 7364
rect 6454 7352 6460 7364
rect 6512 7352 6518 7404
rect 6564 7401 6592 7500
rect 7006 7488 7012 7540
rect 7064 7528 7070 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7064 7500 7665 7528
rect 7064 7488 7070 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 7098 7352 7104 7404
rect 7156 7352 7162 7404
rect 7668 7392 7696 7491
rect 7834 7488 7840 7540
rect 7892 7528 7898 7540
rect 7892 7500 9720 7528
rect 7892 7488 7898 7500
rect 8202 7420 8208 7472
rect 8260 7420 8266 7472
rect 9692 7460 9720 7500
rect 10594 7488 10600 7540
rect 10652 7528 10658 7540
rect 10965 7531 11023 7537
rect 10965 7528 10977 7531
rect 10652 7500 10977 7528
rect 10652 7488 10658 7500
rect 10965 7497 10977 7500
rect 11011 7497 11023 7531
rect 10965 7491 11023 7497
rect 11517 7531 11575 7537
rect 11517 7497 11529 7531
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 11532 7460 11560 7491
rect 12618 7488 12624 7540
rect 12676 7528 12682 7540
rect 12676 7500 16068 7528
rect 12676 7488 12682 7500
rect 9692 7432 11560 7460
rect 13998 7420 14004 7472
rect 14056 7420 14062 7472
rect 14182 7420 14188 7472
rect 14240 7460 14246 7472
rect 14240 7432 14378 7460
rect 14240 7420 14246 7432
rect 14350 7431 14378 7432
rect 14350 7425 14409 7431
rect 7834 7392 7840 7404
rect 7668 7364 7840 7392
rect 7834 7352 7840 7364
rect 7892 7392 7898 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7892 7364 8033 7392
rect 7892 7352 7898 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8220 7392 8248 7420
rect 8220 7364 8328 7392
rect 8021 7355 8079 7361
rect 1118 7284 1124 7336
rect 1176 7324 1182 7336
rect 1673 7327 1731 7333
rect 1673 7324 1685 7327
rect 1176 7296 1685 7324
rect 1176 7284 1182 7296
rect 1673 7293 1685 7296
rect 1719 7293 1731 7327
rect 1673 7287 1731 7293
rect 2866 7284 2872 7336
rect 2924 7324 2930 7336
rect 3970 7324 3976 7336
rect 2924 7296 3976 7324
rect 2924 7284 2930 7296
rect 3970 7284 3976 7296
rect 4028 7284 4034 7336
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 4525 7327 4583 7333
rect 4525 7324 4537 7327
rect 4304 7296 4537 7324
rect 4304 7284 4310 7296
rect 4525 7293 4537 7296
rect 4571 7324 4583 7327
rect 4890 7324 4896 7336
rect 4571 7296 4896 7324
rect 4571 7293 4583 7296
rect 4525 7287 4583 7293
rect 4890 7284 4896 7296
rect 4948 7284 4954 7336
rect 5399 7327 5457 7333
rect 5399 7293 5411 7327
rect 5445 7324 5457 7327
rect 6086 7324 6092 7336
rect 5445 7296 6092 7324
rect 5445 7293 5457 7296
rect 5399 7287 5457 7293
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 7116 7324 7144 7352
rect 7926 7324 7932 7336
rect 7116 7296 7932 7324
rect 7926 7284 7932 7296
rect 7984 7324 7990 7336
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 7984 7296 8217 7324
rect 7984 7284 7990 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8300 7324 8328 7364
rect 9030 7352 9036 7404
rect 9088 7401 9094 7404
rect 9088 7395 9116 7401
rect 9104 7361 9116 7395
rect 9088 7355 9116 7361
rect 9088 7352 9094 7355
rect 9214 7352 9220 7404
rect 9272 7352 9278 7404
rect 10227 7395 10285 7401
rect 10227 7361 10239 7395
rect 10273 7392 10285 7395
rect 11514 7392 11520 7404
rect 10273 7364 11520 7392
rect 10273 7361 10285 7364
rect 10227 7355 10285 7361
rect 11514 7352 11520 7364
rect 11572 7352 11578 7404
rect 11698 7352 11704 7404
rect 11756 7352 11762 7404
rect 11793 7395 11851 7401
rect 11793 7361 11805 7395
rect 11839 7392 11851 7395
rect 11882 7392 11888 7404
rect 11839 7364 11888 7392
rect 11839 7361 11851 7364
rect 11793 7355 11851 7361
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12710 7352 12716 7404
rect 12768 7352 12774 7404
rect 12802 7352 12808 7404
rect 12860 7401 12866 7404
rect 12860 7395 12888 7401
rect 12876 7361 12888 7395
rect 12860 7355 12888 7361
rect 12860 7352 12866 7355
rect 12986 7352 12992 7404
rect 13044 7352 13050 7404
rect 13725 7395 13783 7401
rect 13725 7361 13737 7395
rect 13771 7392 13783 7395
rect 14016 7392 14044 7420
rect 14350 7394 14363 7425
rect 13771 7364 14044 7392
rect 14351 7391 14363 7394
rect 14397 7391 14409 7425
rect 14550 7420 14556 7472
rect 14608 7460 14614 7472
rect 14608 7432 15700 7460
rect 14608 7420 14614 7432
rect 14351 7385 14409 7391
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 15672 7401 15700 7432
rect 15746 7420 15752 7472
rect 15804 7420 15810 7472
rect 16040 7460 16068 7500
rect 16114 7488 16120 7540
rect 16172 7488 16178 7540
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 16264 7500 17632 7528
rect 16264 7488 16270 7500
rect 16758 7460 16764 7472
rect 16040 7432 16764 7460
rect 16758 7420 16764 7432
rect 16816 7420 16822 7472
rect 17126 7420 17132 7472
rect 17184 7420 17190 7472
rect 17218 7420 17224 7472
rect 17276 7460 17282 7472
rect 17604 7460 17632 7500
rect 17678 7488 17684 7540
rect 17736 7488 17742 7540
rect 19518 7528 19524 7540
rect 17926 7500 19524 7528
rect 17926 7460 17954 7500
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 19797 7531 19855 7537
rect 19797 7497 19809 7531
rect 19843 7528 19855 7531
rect 20254 7528 20260 7540
rect 19843 7500 20260 7528
rect 19843 7497 19855 7500
rect 19797 7491 19855 7497
rect 20254 7488 20260 7500
rect 20312 7488 20318 7540
rect 20441 7531 20499 7537
rect 20441 7497 20453 7531
rect 20487 7528 20499 7531
rect 20530 7528 20536 7540
rect 20487 7500 20536 7528
rect 20487 7497 20499 7500
rect 20441 7491 20499 7497
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 21468 7472 21496 7636
rect 17276 7432 17506 7460
rect 17604 7432 17954 7460
rect 17276 7420 17282 7432
rect 15657 7395 15715 7401
rect 14516 7364 15608 7392
rect 14516 7352 14522 7364
rect 8941 7327 8999 7333
rect 8941 7324 8953 7327
rect 8300 7296 8953 7324
rect 2774 7216 2780 7268
rect 2832 7256 2838 7268
rect 4706 7256 4712 7268
rect 2832 7228 4712 7256
rect 2832 7216 2838 7228
rect 4706 7216 4712 7228
rect 4764 7216 4770 7268
rect 4982 7216 4988 7268
rect 5040 7216 5046 7268
rect 7098 7216 7104 7268
rect 7156 7256 7162 7268
rect 8300 7256 8328 7296
rect 8941 7293 8953 7296
rect 8987 7293 8999 7327
rect 8941 7287 8999 7293
rect 9766 7284 9772 7336
rect 9824 7324 9830 7336
rect 9953 7327 10011 7333
rect 9953 7324 9965 7327
rect 9824 7296 9965 7324
rect 9824 7284 9830 7296
rect 9953 7293 9965 7296
rect 9999 7293 10011 7327
rect 9953 7287 10011 7293
rect 10962 7284 10968 7336
rect 11020 7324 11026 7336
rect 11606 7324 11612 7336
rect 11020 7296 11612 7324
rect 11020 7284 11026 7296
rect 11606 7284 11612 7296
rect 11664 7324 11670 7336
rect 11977 7327 12035 7333
rect 11977 7324 11989 7327
rect 11664 7296 11989 7324
rect 11664 7284 11670 7296
rect 11977 7293 11989 7296
rect 12023 7293 12035 7327
rect 12820 7324 12848 7352
rect 11977 7287 12035 7293
rect 12082 7296 12848 7324
rect 14093 7327 14151 7333
rect 7156 7228 8328 7256
rect 8665 7259 8723 7265
rect 7156 7216 7162 7228
rect 8665 7225 8677 7259
rect 8711 7225 8723 7259
rect 8665 7219 8723 7225
rect 1762 7148 1768 7200
rect 1820 7188 1826 7200
rect 3421 7191 3479 7197
rect 3421 7188 3433 7191
rect 1820 7160 3433 7188
rect 1820 7148 1826 7160
rect 3421 7157 3433 7160
rect 3467 7157 3479 7191
rect 3421 7151 3479 7157
rect 3694 7148 3700 7200
rect 3752 7188 3758 7200
rect 3878 7188 3884 7200
rect 3752 7160 3884 7188
rect 3752 7148 3758 7160
rect 3878 7148 3884 7160
rect 3936 7188 3942 7200
rect 5258 7188 5264 7200
rect 3936 7160 5264 7188
rect 3936 7148 3942 7160
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 6181 7191 6239 7197
rect 6181 7188 6193 7191
rect 5776 7160 6193 7188
rect 5776 7148 5782 7160
rect 6181 7157 6193 7160
rect 6227 7157 6239 7191
rect 6181 7151 6239 7157
rect 6362 7148 6368 7200
rect 6420 7148 6426 7200
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8680 7188 8708 7219
rect 8260 7160 8708 7188
rect 8260 7148 8266 7160
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9784 7188 9812 7284
rect 11146 7216 11152 7268
rect 11204 7256 11210 7268
rect 12082 7256 12110 7296
rect 14093 7293 14105 7327
rect 14139 7293 14151 7327
rect 15470 7324 15476 7336
rect 14093 7287 14151 7293
rect 15120 7296 15476 7324
rect 11204 7228 12110 7256
rect 11204 7216 11210 7228
rect 12434 7216 12440 7268
rect 12492 7216 12498 7268
rect 13556 7228 13768 7256
rect 9088 7160 9812 7188
rect 9088 7148 9094 7160
rect 9858 7148 9864 7200
rect 9916 7148 9922 7200
rect 10778 7148 10784 7200
rect 10836 7188 10842 7200
rect 11514 7188 11520 7200
rect 10836 7160 11520 7188
rect 10836 7148 10842 7160
rect 11514 7148 11520 7160
rect 11572 7148 11578 7200
rect 11606 7148 11612 7200
rect 11664 7188 11670 7200
rect 13556 7188 13584 7228
rect 11664 7160 13584 7188
rect 11664 7148 11670 7160
rect 13630 7148 13636 7200
rect 13688 7148 13694 7200
rect 13740 7188 13768 7228
rect 13906 7216 13912 7268
rect 13964 7216 13970 7268
rect 13998 7216 14004 7268
rect 14056 7256 14062 7268
rect 14108 7256 14136 7287
rect 15120 7265 15148 7296
rect 15470 7284 15476 7296
rect 15528 7284 15534 7336
rect 15580 7324 15608 7364
rect 15657 7361 15669 7395
rect 15703 7361 15715 7395
rect 15764 7392 15792 7420
rect 16025 7395 16083 7401
rect 16025 7392 16037 7395
rect 15764 7364 16037 7392
rect 15657 7355 15715 7361
rect 16025 7361 16037 7364
rect 16071 7361 16083 7395
rect 16025 7355 16083 7361
rect 16298 7352 16304 7404
rect 16356 7352 16362 7404
rect 16850 7392 16856 7404
rect 16390 7364 16856 7392
rect 16390 7324 16418 7364
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17144 7392 17172 7420
rect 17000 7364 17043 7392
rect 17144 7364 17356 7392
rect 17000 7352 17006 7364
rect 15580 7296 16418 7324
rect 16482 7284 16488 7336
rect 16540 7284 16546 7336
rect 16666 7284 16672 7336
rect 16724 7284 16730 7336
rect 14056 7228 14136 7256
rect 15105 7259 15163 7265
rect 14056 7216 14062 7228
rect 15105 7225 15117 7259
rect 15151 7225 15163 7259
rect 15105 7219 15163 7225
rect 15378 7216 15384 7268
rect 15436 7256 15442 7268
rect 15657 7259 15715 7265
rect 15657 7256 15669 7259
rect 15436 7228 15669 7256
rect 15436 7216 15442 7228
rect 15657 7225 15669 7228
rect 15703 7225 15715 7259
rect 15657 7219 15715 7225
rect 15746 7216 15752 7268
rect 15804 7256 15810 7268
rect 16500 7256 16528 7284
rect 15804 7228 16528 7256
rect 17328 7256 17356 7364
rect 17478 7324 17506 7432
rect 18046 7420 18052 7472
rect 18104 7460 18110 7472
rect 18104 7432 19840 7460
rect 18104 7420 18110 7432
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 18012 7364 18153 7392
rect 18012 7352 18018 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18230 7352 18236 7404
rect 18288 7352 18294 7404
rect 18397 7395 18455 7401
rect 18397 7361 18409 7395
rect 18443 7392 18455 7395
rect 18966 7392 18972 7404
rect 18443 7364 18972 7392
rect 18443 7361 18455 7364
rect 18397 7355 18455 7361
rect 18966 7352 18972 7364
rect 19024 7352 19030 7404
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 19702 7392 19708 7404
rect 19659 7364 19708 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 19702 7352 19708 7364
rect 19760 7352 19766 7404
rect 19812 7401 19840 7432
rect 19886 7420 19892 7472
rect 19944 7460 19950 7472
rect 20165 7463 20223 7469
rect 20165 7460 20177 7463
rect 19944 7432 20177 7460
rect 19944 7420 19950 7432
rect 20165 7429 20177 7432
rect 20211 7429 20223 7463
rect 20165 7423 20223 7429
rect 21450 7420 21456 7472
rect 21508 7420 21514 7472
rect 19797 7395 19855 7401
rect 19797 7361 19809 7395
rect 19843 7361 19855 7395
rect 19797 7355 19855 7361
rect 18248 7324 18276 7352
rect 17478 7296 18276 7324
rect 18046 7256 18052 7268
rect 17328 7228 18052 7256
rect 15804 7216 15810 7228
rect 18046 7216 18052 7228
rect 18104 7216 18110 7268
rect 16206 7188 16212 7200
rect 13740 7160 16212 7188
rect 16206 7148 16212 7160
rect 16264 7148 16270 7200
rect 16390 7148 16396 7200
rect 16448 7188 16454 7200
rect 19521 7191 19579 7197
rect 19521 7188 19533 7191
rect 16448 7160 19533 7188
rect 16448 7148 16454 7160
rect 19521 7157 19533 7160
rect 19567 7157 19579 7191
rect 19521 7151 19579 7157
rect 1104 7098 20884 7120
rect 1104 7046 3422 7098
rect 3474 7046 3486 7098
rect 3538 7046 3550 7098
rect 3602 7046 3614 7098
rect 3666 7046 3678 7098
rect 3730 7046 8367 7098
rect 8419 7046 8431 7098
rect 8483 7046 8495 7098
rect 8547 7046 8559 7098
rect 8611 7046 8623 7098
rect 8675 7046 13312 7098
rect 13364 7046 13376 7098
rect 13428 7046 13440 7098
rect 13492 7046 13504 7098
rect 13556 7046 13568 7098
rect 13620 7046 18257 7098
rect 18309 7046 18321 7098
rect 18373 7046 18385 7098
rect 18437 7046 18449 7098
rect 18501 7046 18513 7098
rect 18565 7046 20884 7098
rect 1104 7024 20884 7046
rect 1486 6944 1492 6996
rect 1544 6944 1550 6996
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 1949 6987 2007 6993
rect 1949 6984 1961 6987
rect 1636 6956 1961 6984
rect 1636 6944 1642 6956
rect 1949 6953 1961 6956
rect 1995 6953 2007 6987
rect 1949 6947 2007 6953
rect 2038 6944 2044 6996
rect 2096 6984 2102 6996
rect 3973 6987 4031 6993
rect 3973 6984 3985 6987
rect 2096 6956 3985 6984
rect 2096 6944 2102 6956
rect 3973 6953 3985 6956
rect 4019 6953 4031 6987
rect 3973 6947 4031 6953
rect 4126 6956 5304 6984
rect 1118 6808 1124 6860
rect 1176 6848 1182 6860
rect 2222 6848 2228 6860
rect 1176 6820 2228 6848
rect 1176 6808 1182 6820
rect 2222 6808 2228 6820
rect 2280 6848 2286 6860
rect 2317 6851 2375 6857
rect 2317 6848 2329 6851
rect 2280 6820 2329 6848
rect 2280 6808 2286 6820
rect 2317 6817 2329 6820
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 4126 6848 4154 6956
rect 5276 6916 5304 6956
rect 5534 6944 5540 6996
rect 5592 6984 5598 6996
rect 5629 6987 5687 6993
rect 5629 6984 5641 6987
rect 5592 6956 5641 6984
rect 5592 6944 5598 6956
rect 5629 6953 5641 6956
rect 5675 6953 5687 6987
rect 5629 6947 5687 6953
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 6972 6956 7077 6984
rect 6972 6944 6978 6956
rect 6362 6916 6368 6928
rect 5276 6888 6368 6916
rect 6362 6876 6368 6888
rect 6420 6876 6426 6928
rect 3108 6820 4154 6848
rect 3108 6808 3114 6820
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 4617 6851 4675 6857
rect 4617 6848 4629 6851
rect 4396 6820 4629 6848
rect 4396 6808 4402 6820
rect 4617 6817 4629 6820
rect 4663 6817 4675 6851
rect 4617 6811 4675 6817
rect 5626 6808 5632 6860
rect 5684 6848 5690 6860
rect 6457 6851 6515 6857
rect 6457 6848 6469 6851
rect 5684 6820 6469 6848
rect 5684 6808 5690 6820
rect 6457 6817 6469 6820
rect 6503 6817 6515 6851
rect 6822 6848 6828 6860
rect 6457 6811 6515 6817
rect 6656 6820 6828 6848
rect 474 6740 480 6792
rect 532 6780 538 6792
rect 2590 6789 2596 6792
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 532 6752 1685 6780
rect 532 6740 538 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 1673 6743 1731 6749
rect 1857 6783 1915 6789
rect 1857 6749 1869 6783
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 2559 6783 2596 6789
rect 2559 6749 2571 6783
rect 2559 6743 2596 6749
rect 1872 6712 1900 6743
rect 2590 6740 2596 6743
rect 2648 6740 2654 6792
rect 2976 6752 4476 6780
rect 2976 6712 3004 6752
rect 1872 6684 3004 6712
rect 3881 6715 3939 6721
rect 3881 6681 3893 6715
rect 3927 6712 3939 6715
rect 3927 6684 4384 6712
rect 3927 6681 3939 6684
rect 3881 6675 3939 6681
rect 1762 6604 1768 6656
rect 1820 6644 1826 6656
rect 3050 6644 3056 6656
rect 1820 6616 3056 6644
rect 1820 6604 1826 6616
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 3786 6644 3792 6656
rect 3375 6616 3792 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4356 6653 4384 6684
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6613 4399 6647
rect 4448 6644 4476 6752
rect 4522 6740 4528 6792
rect 4580 6740 4586 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5258 6780 5264 6792
rect 4948 6752 5264 6780
rect 4948 6740 4954 6752
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 5994 6780 6000 6792
rect 5868 6752 6000 6780
rect 5868 6740 5874 6752
rect 5994 6740 6000 6752
rect 6052 6740 6058 6792
rect 6178 6740 6184 6792
rect 6236 6740 6242 6792
rect 6273 6783 6331 6789
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 6273 6743 6331 6749
rect 6288 6712 6316 6743
rect 6362 6740 6368 6792
rect 6420 6780 6426 6792
rect 6656 6780 6684 6820
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 6914 6808 6920 6860
rect 6972 6808 6978 6860
rect 7049 6848 7077 6956
rect 7834 6944 7840 6996
rect 7892 6984 7898 6996
rect 9306 6984 9312 6996
rect 7892 6956 9312 6984
rect 7892 6944 7898 6956
rect 9306 6944 9312 6956
rect 9364 6944 9370 6996
rect 9398 6944 9404 6996
rect 9456 6984 9462 6996
rect 11977 6987 12035 6993
rect 11977 6984 11989 6987
rect 9456 6956 10898 6984
rect 9456 6944 9462 6956
rect 7926 6876 7932 6928
rect 7984 6916 7990 6928
rect 9766 6916 9772 6928
rect 7984 6888 9772 6916
rect 7984 6876 7990 6888
rect 9766 6876 9772 6888
rect 9824 6876 9830 6928
rect 7193 6851 7251 6857
rect 7193 6848 7205 6851
rect 7049 6820 7205 6848
rect 7193 6817 7205 6820
rect 7239 6848 7251 6851
rect 8478 6848 8484 6860
rect 7239 6820 8484 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10321 6851 10379 6857
rect 10321 6848 10333 6851
rect 10008 6820 10333 6848
rect 10008 6808 10014 6820
rect 10321 6817 10333 6820
rect 10367 6817 10379 6851
rect 10321 6811 10379 6817
rect 10502 6808 10508 6860
rect 10560 6808 10566 6860
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10781 6851 10839 6857
rect 10781 6848 10793 6851
rect 10744 6820 10793 6848
rect 10744 6808 10750 6820
rect 10781 6817 10793 6820
rect 10827 6817 10839 6851
rect 10870 6848 10898 6956
rect 11958 6953 11989 6984
rect 12023 6953 12035 6987
rect 11958 6947 12035 6953
rect 11808 6876 11814 6928
rect 11866 6916 11872 6928
rect 11958 6916 11986 6947
rect 12158 6944 12164 6996
rect 12216 6944 12222 6996
rect 12342 6944 12348 6996
rect 12400 6984 12406 6996
rect 12400 6956 12940 6984
rect 12400 6944 12406 6956
rect 12176 6916 12204 6944
rect 11866 6888 11986 6916
rect 12082 6888 12204 6916
rect 12912 6916 12940 6956
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 13044 6956 13093 6984
rect 13044 6944 13050 6956
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 13081 6947 13139 6953
rect 13817 6987 13875 6993
rect 13817 6953 13829 6987
rect 13863 6984 13875 6987
rect 14550 6984 14556 6996
rect 13863 6956 14556 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 14700 6956 17816 6984
rect 14700 6944 14706 6956
rect 13906 6916 13912 6928
rect 12912 6888 13912 6916
rect 11866 6876 11872 6888
rect 12082 6848 12110 6888
rect 13906 6876 13912 6888
rect 13964 6876 13970 6928
rect 14090 6876 14096 6928
rect 14148 6876 14154 6928
rect 10870 6820 12110 6848
rect 10781 6811 10839 6817
rect 6420 6752 6684 6780
rect 6420 6740 6426 6752
rect 7282 6740 7288 6792
rect 7340 6789 7346 6792
rect 7340 6783 7368 6789
rect 7356 6749 7368 6783
rect 7340 6743 7368 6749
rect 7340 6740 7346 6743
rect 7466 6740 7472 6792
rect 7524 6740 7530 6792
rect 9214 6740 9220 6792
rect 9272 6740 9278 6792
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6780 10195 6783
rect 10520 6780 10548 6808
rect 10183 6752 10548 6780
rect 10183 6749 10195 6752
rect 10137 6743 10195 6749
rect 11054 6740 11060 6792
rect 11112 6740 11118 6792
rect 11146 6740 11152 6792
rect 11204 6789 11210 6792
rect 11204 6783 11232 6789
rect 11220 6749 11232 6783
rect 11204 6743 11232 6749
rect 11204 6740 11210 6743
rect 11330 6740 11336 6792
rect 11388 6740 11394 6792
rect 6454 6712 6460 6724
rect 5092 6684 6040 6712
rect 6288 6684 6460 6712
rect 5092 6644 5120 6684
rect 4448 6616 5120 6644
rect 4341 6607 4399 6613
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5902 6644 5908 6656
rect 5316 6616 5908 6644
rect 5316 6604 5322 6616
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6012 6653 6040 6684
rect 6454 6672 6460 6684
rect 6512 6672 6518 6724
rect 9490 6672 9496 6724
rect 9548 6712 9554 6724
rect 11992 6712 12020 6820
rect 13354 6808 13360 6860
rect 13412 6848 13418 6860
rect 14108 6848 14136 6876
rect 13412 6820 14136 6848
rect 13412 6808 13418 6820
rect 15378 6808 15384 6860
rect 15436 6848 15442 6860
rect 15654 6848 15660 6860
rect 15436 6820 15660 6848
rect 15436 6808 15442 6820
rect 15654 6808 15660 6820
rect 15712 6808 15718 6860
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 17129 6851 17187 6857
rect 17129 6848 17141 6851
rect 16724 6820 17141 6848
rect 16724 6808 16730 6820
rect 17129 6817 17141 6820
rect 17175 6817 17187 6851
rect 17788 6848 17816 6956
rect 18598 6944 18604 6996
rect 18656 6984 18662 6996
rect 19242 6984 19248 6996
rect 18656 6956 19248 6984
rect 18656 6944 18662 6956
rect 19242 6944 19248 6956
rect 19300 6944 19306 6996
rect 20070 6876 20076 6928
rect 20128 6876 20134 6928
rect 17788 6820 20116 6848
rect 17129 6811 17187 6817
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 12327 6783 12385 6789
rect 12327 6749 12339 6783
rect 12373 6749 12385 6783
rect 12327 6743 12385 6749
rect 12342 6712 12370 6743
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 13262 6780 13268 6792
rect 12768 6752 13268 6780
rect 12768 6740 12774 6752
rect 13262 6740 13268 6752
rect 13320 6740 13326 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 13630 6780 13636 6792
rect 13495 6752 13636 6780
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 13630 6740 13636 6752
rect 13688 6740 13694 6792
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 13998 6740 14004 6792
rect 14056 6780 14062 6792
rect 14277 6783 14335 6789
rect 14277 6780 14289 6783
rect 14056 6752 14289 6780
rect 14056 6740 14062 6752
rect 14277 6749 14289 6752
rect 14323 6749 14335 6783
rect 14277 6743 14335 6749
rect 14551 6783 14609 6789
rect 14551 6749 14563 6783
rect 14597 6780 14609 6783
rect 14918 6780 14924 6792
rect 14597 6752 14924 6780
rect 14597 6749 14609 6752
rect 14551 6743 14609 6749
rect 14918 6740 14924 6752
rect 14976 6740 14982 6792
rect 15470 6740 15476 6792
rect 15528 6780 15534 6792
rect 15913 6783 15971 6789
rect 15913 6780 15925 6783
rect 15528 6752 15925 6780
rect 15528 6740 15534 6752
rect 15913 6749 15925 6752
rect 15959 6749 15971 6783
rect 17034 6780 17040 6792
rect 15913 6743 15971 6749
rect 16036 6752 17040 6780
rect 9548 6684 10088 6712
rect 11992 6684 12370 6712
rect 9548 6672 9554 6684
rect 10060 6656 10088 6684
rect 12618 6672 12624 6724
rect 12676 6712 12682 6724
rect 16036 6712 16064 6752
rect 17034 6740 17040 6752
rect 17092 6780 17098 6792
rect 17371 6783 17429 6789
rect 17371 6780 17383 6783
rect 17092 6752 17383 6780
rect 17092 6740 17098 6752
rect 17371 6749 17383 6752
rect 17417 6749 17429 6783
rect 17371 6743 17429 6749
rect 18046 6740 18052 6792
rect 18104 6780 18110 6792
rect 18414 6780 18420 6792
rect 18104 6752 18420 6780
rect 18104 6740 18110 6752
rect 18414 6740 18420 6752
rect 18472 6740 18478 6792
rect 18509 6783 18567 6789
rect 18509 6749 18521 6783
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 18524 6712 18552 6743
rect 18598 6740 18604 6792
rect 18656 6780 18662 6792
rect 18693 6783 18751 6789
rect 18693 6780 18705 6783
rect 18656 6752 18705 6780
rect 18656 6740 18662 6752
rect 18693 6749 18705 6752
rect 18739 6749 18751 6783
rect 18693 6743 18751 6749
rect 18785 6783 18843 6789
rect 18785 6749 18797 6783
rect 18831 6749 18843 6783
rect 18785 6743 18843 6749
rect 18800 6712 18828 6743
rect 18874 6740 18880 6792
rect 18932 6780 18938 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18932 6752 18981 6780
rect 18932 6740 18938 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 19337 6783 19395 6789
rect 19337 6749 19349 6783
rect 19383 6749 19395 6783
rect 19337 6743 19395 6749
rect 12676 6684 16064 6712
rect 16408 6684 18552 6712
rect 18708 6684 18828 6712
rect 12676 6672 12682 6684
rect 5997 6647 6055 6653
rect 5997 6613 6009 6647
rect 6043 6613 6055 6647
rect 5997 6607 6055 6613
rect 6822 6604 6828 6656
rect 6880 6644 6886 6656
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 6880 6616 8125 6644
rect 6880 6604 6886 6616
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8113 6607 8171 6613
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 9858 6644 9864 6656
rect 9732 6616 9864 6644
rect 9732 6604 9738 6616
rect 9858 6604 9864 6616
rect 9916 6604 9922 6656
rect 10042 6604 10048 6656
rect 10100 6604 10106 6656
rect 10502 6604 10508 6656
rect 10560 6644 10566 6656
rect 13633 6647 13691 6653
rect 13633 6644 13645 6647
rect 10560 6616 13645 6644
rect 10560 6604 10566 6616
rect 13633 6613 13645 6616
rect 13679 6613 13691 6647
rect 13633 6607 13691 6613
rect 13998 6604 14004 6656
rect 14056 6644 14062 6656
rect 15194 6644 15200 6656
rect 14056 6616 15200 6644
rect 14056 6604 14062 6616
rect 15194 6604 15200 6616
rect 15252 6604 15258 6656
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6644 15347 6647
rect 15654 6644 15660 6656
rect 15335 6616 15660 6644
rect 15335 6613 15347 6616
rect 15289 6607 15347 6613
rect 15654 6604 15660 6616
rect 15712 6644 15718 6656
rect 16408 6644 16436 6684
rect 18708 6656 18736 6684
rect 15712 6616 16436 6644
rect 17037 6647 17095 6653
rect 15712 6604 15718 6616
rect 17037 6613 17049 6647
rect 17083 6644 17095 6647
rect 17770 6644 17776 6656
rect 17083 6616 17776 6644
rect 17083 6613 17095 6616
rect 17037 6607 17095 6613
rect 17770 6604 17776 6616
rect 17828 6604 17834 6656
rect 18138 6604 18144 6656
rect 18196 6604 18202 6656
rect 18598 6604 18604 6656
rect 18656 6604 18662 6656
rect 18690 6604 18696 6656
rect 18748 6604 18754 6656
rect 18874 6604 18880 6656
rect 18932 6604 18938 6656
rect 19352 6644 19380 6743
rect 19610 6740 19616 6792
rect 19668 6740 19674 6792
rect 20088 6789 20116 6820
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6749 20131 6783
rect 20073 6743 20131 6749
rect 19886 6644 19892 6656
rect 19352 6616 19892 6644
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 20530 6604 20536 6656
rect 20588 6644 20594 6656
rect 20990 6644 20996 6656
rect 20588 6616 20996 6644
rect 20588 6604 20594 6616
rect 20990 6604 20996 6616
rect 21048 6604 21054 6656
rect 1104 6554 21043 6576
rect 1104 6502 5894 6554
rect 5946 6502 5958 6554
rect 6010 6502 6022 6554
rect 6074 6502 6086 6554
rect 6138 6502 6150 6554
rect 6202 6502 10839 6554
rect 10891 6502 10903 6554
rect 10955 6502 10967 6554
rect 11019 6502 11031 6554
rect 11083 6502 11095 6554
rect 11147 6502 15784 6554
rect 15836 6502 15848 6554
rect 15900 6502 15912 6554
rect 15964 6502 15976 6554
rect 16028 6502 16040 6554
rect 16092 6502 20729 6554
rect 20781 6502 20793 6554
rect 20845 6502 20857 6554
rect 20909 6502 20921 6554
rect 20973 6502 20985 6554
rect 21037 6502 21043 6554
rect 1104 6480 21043 6502
rect 1578 6400 1584 6452
rect 1636 6400 1642 6452
rect 2314 6400 2320 6452
rect 2372 6400 2378 6452
rect 3878 6440 3884 6452
rect 2792 6412 3884 6440
rect 1489 6375 1547 6381
rect 1489 6341 1501 6375
rect 1535 6372 1547 6375
rect 2130 6372 2136 6384
rect 1535 6344 2136 6372
rect 1535 6341 1547 6344
rect 1489 6335 1547 6341
rect 2130 6332 2136 6344
rect 2188 6332 2194 6384
rect 106 6264 112 6316
rect 164 6264 170 6316
rect 2038 6264 2044 6316
rect 2096 6264 2102 6316
rect 2792 6313 2820 6412
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 4433 6443 4491 6449
rect 4433 6409 4445 6443
rect 4479 6440 4491 6443
rect 4522 6440 4528 6452
rect 4479 6412 4528 6440
rect 4479 6409 4491 6412
rect 4433 6403 4491 6409
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4982 6400 4988 6452
rect 5040 6440 5046 6452
rect 5537 6443 5595 6449
rect 5537 6440 5549 6443
rect 5040 6412 5549 6440
rect 5040 6400 5046 6412
rect 5537 6409 5549 6412
rect 5583 6409 5595 6443
rect 5537 6403 5595 6409
rect 5626 6400 5632 6452
rect 5684 6440 5690 6452
rect 5684 6412 6224 6440
rect 5684 6400 5690 6412
rect 4338 6332 4344 6384
rect 4396 6372 4402 6384
rect 4396 6344 5856 6372
rect 4396 6332 4402 6344
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6273 2835 6307
rect 2777 6267 2835 6273
rect 3786 6264 3792 6316
rect 3844 6264 3850 6316
rect 4540 6313 4568 6344
rect 5828 6316 5856 6344
rect 4525 6307 4583 6313
rect 4525 6273 4537 6307
rect 4571 6273 4583 6307
rect 4525 6267 4583 6273
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 4799 6307 4857 6313
rect 4799 6304 4811 6307
rect 4764 6276 4811 6304
rect 4764 6264 4770 6276
rect 4799 6273 4811 6276
rect 4845 6273 4857 6307
rect 4799 6267 4857 6273
rect 5166 6264 5172 6316
rect 5224 6304 5230 6316
rect 5626 6304 5632 6316
rect 5224 6276 5632 6304
rect 5224 6264 5230 6276
rect 5626 6264 5632 6276
rect 5684 6264 5690 6316
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 6086 6264 6092 6316
rect 6144 6264 6150 6316
rect 124 6236 152 6264
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 124 6208 2605 6236
rect 2593 6205 2605 6208
rect 2639 6205 2651 6239
rect 2593 6199 2651 6205
rect 2608 6168 2636 6199
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 3513 6239 3571 6245
rect 3513 6236 3525 6239
rect 2924 6208 3525 6236
rect 2924 6196 2930 6208
rect 3513 6205 3525 6208
rect 3559 6205 3571 6239
rect 3513 6199 3571 6205
rect 3651 6239 3709 6245
rect 3651 6205 3663 6239
rect 3697 6236 3709 6239
rect 6196 6236 6224 6412
rect 6270 6400 6276 6452
rect 6328 6440 6334 6452
rect 6328 6412 6592 6440
rect 6328 6400 6334 6412
rect 6564 6313 6592 6412
rect 8202 6400 8208 6452
rect 8260 6400 8266 6452
rect 8478 6400 8484 6452
rect 8536 6440 8542 6452
rect 8536 6412 8800 6440
rect 8536 6400 8542 6412
rect 7282 6372 7288 6384
rect 7208 6344 7288 6372
rect 7208 6313 7236 6344
rect 7282 6332 7288 6344
rect 7340 6332 7346 6384
rect 8772 6381 8800 6412
rect 8956 6412 9812 6440
rect 8757 6375 8815 6381
rect 8757 6341 8769 6375
rect 8803 6341 8815 6375
rect 8757 6335 8815 6341
rect 7467 6317 7525 6323
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 7193 6307 7251 6313
rect 7193 6273 7205 6307
rect 7239 6273 7251 6307
rect 7467 6283 7479 6317
rect 7513 6314 7525 6317
rect 7513 6304 7604 6314
rect 8956 6304 8984 6412
rect 9033 6375 9091 6381
rect 9033 6341 9045 6375
rect 9079 6372 9091 6375
rect 9214 6372 9220 6384
rect 9079 6344 9220 6372
rect 9079 6341 9091 6344
rect 9033 6335 9091 6341
rect 9214 6332 9220 6344
rect 9272 6332 9278 6384
rect 9306 6332 9312 6384
rect 9364 6372 9370 6384
rect 9493 6375 9551 6381
rect 9493 6372 9505 6375
rect 9364 6344 9505 6372
rect 9364 6332 9370 6344
rect 9493 6341 9505 6344
rect 9539 6341 9551 6375
rect 9784 6372 9812 6412
rect 9858 6400 9864 6452
rect 9916 6400 9922 6452
rect 10045 6443 10103 6449
rect 10045 6409 10057 6443
rect 10091 6440 10103 6443
rect 10134 6440 10140 6452
rect 10091 6412 10140 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10134 6400 10140 6412
rect 10192 6400 10198 6452
rect 11790 6440 11796 6452
rect 11026 6412 11796 6440
rect 11026 6372 11054 6412
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 12066 6440 12072 6452
rect 11900 6412 12072 6440
rect 11900 6372 11928 6412
rect 12066 6400 12072 6412
rect 12124 6440 12130 6452
rect 12124 6412 12296 6440
rect 12124 6400 12130 6412
rect 9784 6344 11054 6372
rect 11532 6344 11928 6372
rect 12268 6372 12296 6412
rect 12342 6400 12348 6452
rect 12400 6440 12406 6452
rect 12529 6443 12587 6449
rect 12529 6440 12541 6443
rect 12400 6412 12541 6440
rect 12400 6400 12406 6412
rect 12529 6409 12541 6412
rect 12575 6409 12587 6443
rect 12529 6403 12587 6409
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 14458 6440 14464 6452
rect 12768 6412 14464 6440
rect 12768 6400 12774 6412
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 15746 6440 15752 6452
rect 14792 6412 15752 6440
rect 14792 6400 14798 6412
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15838 6400 15844 6452
rect 15896 6400 15902 6452
rect 15933 6443 15991 6449
rect 15933 6409 15945 6443
rect 15979 6409 15991 6443
rect 15933 6403 15991 6409
rect 12268 6344 13492 6372
rect 9493 6335 9551 6341
rect 7513 6286 8984 6304
rect 7513 6283 7525 6286
rect 7467 6277 7525 6283
rect 7576 6276 8984 6286
rect 9125 6307 9183 6313
rect 7193 6267 7251 6273
rect 9125 6273 9137 6307
rect 9171 6304 9183 6307
rect 9171 6276 9904 6304
rect 9171 6273 9183 6276
rect 9125 6267 9183 6273
rect 3697 6208 4568 6236
rect 6196 6208 7254 6236
rect 3697 6205 3709 6208
rect 3651 6199 3709 6205
rect 3050 6168 3056 6180
rect 2608 6140 3056 6168
rect 3050 6128 3056 6140
rect 3108 6128 3114 6180
rect 3234 6128 3240 6180
rect 3292 6128 3298 6180
rect 2590 6060 2596 6112
rect 2648 6100 2654 6112
rect 3326 6100 3332 6112
rect 2648 6072 3332 6100
rect 2648 6060 2654 6072
rect 3326 6060 3332 6072
rect 3384 6060 3390 6112
rect 4540 6100 4568 6208
rect 7098 6168 7104 6180
rect 5828 6140 7104 6168
rect 5828 6100 5856 6140
rect 7098 6128 7104 6140
rect 7156 6128 7162 6180
rect 4540 6072 5856 6100
rect 5902 6060 5908 6112
rect 5960 6060 5966 6112
rect 6362 6060 6368 6112
rect 6420 6060 6426 6112
rect 7226 6100 7254 6208
rect 9398 6196 9404 6248
rect 9456 6196 9462 6248
rect 9876 6236 9904 6276
rect 10226 6264 10232 6316
rect 10284 6264 10290 6316
rect 11054 6264 11060 6316
rect 11112 6264 11118 6316
rect 11146 6264 11152 6316
rect 11204 6264 11210 6316
rect 11532 6313 11560 6344
rect 11333 6307 11391 6313
rect 11333 6273 11345 6307
rect 11379 6273 11391 6307
rect 11333 6267 11391 6273
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 11790 6304 11796 6316
rect 11751 6276 11796 6304
rect 11517 6267 11575 6273
rect 9950 6236 9956 6248
rect 9876 6208 9956 6236
rect 9950 6196 9956 6208
rect 10008 6196 10014 6248
rect 11348 6236 11376 6267
rect 11790 6264 11796 6276
rect 11848 6304 11854 6316
rect 11848 6276 12204 6304
rect 11848 6264 11854 6276
rect 11422 6236 11428 6248
rect 11348 6208 11428 6236
rect 11422 6196 11428 6208
rect 11480 6196 11486 6248
rect 12176 6168 12204 6276
rect 12342 6264 12348 6316
rect 12400 6304 12406 6316
rect 13354 6313 13360 6316
rect 13323 6307 13360 6313
rect 13323 6304 13335 6307
rect 12400 6276 13335 6304
rect 12400 6264 12406 6276
rect 13323 6273 13335 6276
rect 13323 6267 13360 6273
rect 13354 6264 13360 6267
rect 13412 6264 13418 6316
rect 13464 6304 13492 6344
rect 13722 6332 13728 6384
rect 13780 6372 13786 6384
rect 15102 6372 15108 6384
rect 13780 6344 15108 6372
rect 13780 6332 13786 6344
rect 15102 6332 15108 6344
rect 15160 6332 15166 6384
rect 14182 6304 14188 6316
rect 13464 6276 14188 6304
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 14734 6313 14740 6316
rect 14728 6304 14740 6313
rect 14695 6276 14740 6304
rect 14728 6267 14740 6276
rect 14734 6264 14740 6267
rect 14792 6264 14798 6316
rect 15194 6264 15200 6316
rect 15252 6304 15258 6316
rect 15252 6276 15516 6304
rect 15252 6264 15258 6276
rect 13081 6239 13139 6245
rect 13081 6205 13093 6239
rect 13127 6205 13139 6239
rect 13081 6199 13139 6205
rect 14461 6239 14519 6245
rect 14461 6205 14473 6239
rect 14507 6205 14519 6239
rect 14461 6199 14519 6205
rect 12526 6168 12532 6180
rect 12176 6140 12532 6168
rect 12526 6128 12532 6140
rect 12584 6128 12590 6180
rect 7558 6100 7564 6112
rect 7226 6072 7564 6100
rect 7558 6060 7564 6072
rect 7616 6060 7622 6112
rect 10134 6060 10140 6112
rect 10192 6100 10198 6112
rect 10413 6103 10471 6109
rect 10413 6100 10425 6103
rect 10192 6072 10425 6100
rect 10192 6060 10198 6072
rect 10413 6069 10425 6072
rect 10459 6069 10471 6103
rect 10413 6063 10471 6069
rect 10594 6060 10600 6112
rect 10652 6100 10658 6112
rect 10873 6103 10931 6109
rect 10873 6100 10885 6103
rect 10652 6072 10885 6100
rect 10652 6060 10658 6072
rect 10873 6069 10885 6072
rect 10919 6069 10931 6103
rect 10873 6063 10931 6069
rect 11241 6103 11299 6109
rect 11241 6069 11253 6103
rect 11287 6100 11299 6103
rect 12434 6100 12440 6112
rect 11287 6072 12440 6100
rect 11287 6069 11299 6072
rect 11241 6063 11299 6069
rect 12434 6060 12440 6072
rect 12492 6060 12498 6112
rect 12618 6060 12624 6112
rect 12676 6100 12682 6112
rect 12986 6100 12992 6112
rect 12676 6072 12992 6100
rect 12676 6060 12682 6072
rect 12986 6060 12992 6072
rect 13044 6060 13050 6112
rect 13096 6100 13124 6199
rect 13745 6128 13751 6180
rect 13803 6168 13809 6180
rect 14093 6171 14151 6177
rect 14093 6168 14105 6171
rect 13803 6140 14105 6168
rect 13803 6128 13809 6140
rect 14093 6137 14105 6140
rect 14139 6137 14151 6171
rect 14093 6131 14151 6137
rect 14476 6112 14504 6199
rect 15488 6168 15516 6276
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 15948 6304 15976 6403
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 16298 6440 16304 6452
rect 16080 6412 16304 6440
rect 16080 6400 16086 6412
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 16408 6412 18184 6440
rect 15896 6276 15976 6304
rect 15896 6264 15902 6276
rect 16022 6264 16028 6316
rect 16080 6304 16086 6316
rect 16117 6307 16175 6313
rect 16117 6304 16129 6307
rect 16080 6276 16129 6304
rect 16080 6264 16086 6276
rect 16117 6273 16129 6276
rect 16163 6273 16175 6307
rect 16117 6267 16175 6273
rect 16206 6264 16212 6316
rect 16264 6304 16270 6316
rect 16301 6307 16359 6313
rect 16301 6304 16313 6307
rect 16264 6276 16313 6304
rect 16264 6264 16270 6276
rect 16301 6273 16313 6276
rect 16347 6304 16359 6307
rect 16408 6304 16436 6412
rect 18156 6384 18184 6412
rect 18248 6412 19334 6440
rect 18248 6384 18276 6412
rect 18046 6372 18052 6384
rect 16500 6344 18052 6372
rect 16500 6313 16528 6344
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 18138 6332 18144 6384
rect 18196 6332 18202 6384
rect 18230 6332 18236 6384
rect 18288 6332 18294 6384
rect 18506 6332 18512 6384
rect 18564 6372 18570 6384
rect 18785 6375 18843 6381
rect 18785 6372 18797 6375
rect 18564 6344 18797 6372
rect 18564 6332 18570 6344
rect 18785 6341 18797 6344
rect 18831 6341 18843 6375
rect 18785 6335 18843 6341
rect 16347 6276 16436 6304
rect 16485 6307 16543 6313
rect 16347 6273 16359 6276
rect 16301 6267 16359 6273
rect 16485 6273 16497 6307
rect 16531 6273 16543 6307
rect 16485 6267 16543 6273
rect 16574 6264 16580 6316
rect 16632 6264 16638 6316
rect 16666 6264 16672 6316
rect 16724 6304 16730 6316
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16724 6276 16865 6304
rect 16724 6264 16730 6276
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17126 6264 17132 6316
rect 17184 6264 17190 6316
rect 17678 6264 17684 6316
rect 17736 6304 17742 6316
rect 18417 6307 18475 6313
rect 18417 6304 18429 6307
rect 17736 6276 18429 6304
rect 17736 6264 17742 6276
rect 18417 6273 18429 6276
rect 18463 6273 18475 6307
rect 18417 6267 18475 6273
rect 18601 6307 18659 6313
rect 18601 6273 18613 6307
rect 18647 6304 18659 6307
rect 18690 6304 18696 6316
rect 18647 6276 18696 6304
rect 18647 6273 18659 6276
rect 18601 6267 18659 6273
rect 18690 6264 18696 6276
rect 18748 6264 18754 6316
rect 19133 6307 19191 6313
rect 19133 6304 19145 6307
rect 18800 6276 19145 6304
rect 16390 6196 16396 6248
rect 16448 6196 16454 6248
rect 16592 6236 16620 6264
rect 16592 6208 16896 6236
rect 16758 6168 16764 6180
rect 15488 6140 16764 6168
rect 16758 6128 16764 6140
rect 16816 6128 16822 6180
rect 13998 6100 14004 6112
rect 13096 6072 14004 6100
rect 13998 6060 14004 6072
rect 14056 6060 14062 6112
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 15378 6100 15384 6112
rect 14516 6072 15384 6100
rect 14516 6060 14522 6072
rect 15378 6060 15384 6072
rect 15436 6060 15442 6112
rect 15562 6060 15568 6112
rect 15620 6100 15626 6112
rect 16574 6100 16580 6112
rect 15620 6072 16580 6100
rect 15620 6060 15626 6072
rect 16574 6060 16580 6072
rect 16632 6060 16638 6112
rect 16868 6100 16896 6208
rect 17862 6196 17868 6248
rect 17920 6236 17926 6248
rect 18138 6236 18144 6248
rect 17920 6208 18144 6236
rect 17920 6196 17926 6208
rect 18138 6196 18144 6208
rect 18196 6196 18202 6248
rect 18800 6236 18828 6276
rect 19133 6273 19145 6276
rect 19179 6273 19191 6307
rect 19306 6304 19334 6412
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 20257 6443 20315 6449
rect 20257 6440 20269 6443
rect 19668 6412 20269 6440
rect 19668 6400 19674 6412
rect 20257 6409 20269 6412
rect 20303 6409 20315 6443
rect 20257 6403 20315 6409
rect 19702 6304 19708 6316
rect 19306 6276 19708 6304
rect 19133 6267 19191 6273
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 20346 6264 20352 6316
rect 20404 6264 20410 6316
rect 18248 6208 18828 6236
rect 17678 6128 17684 6180
rect 17736 6168 17742 6180
rect 18248 6168 18276 6208
rect 18874 6196 18880 6248
rect 18932 6196 18938 6248
rect 17736 6140 18276 6168
rect 17736 6128 17742 6140
rect 18414 6128 18420 6180
rect 18472 6128 18478 6180
rect 17865 6103 17923 6109
rect 17865 6100 17877 6103
rect 16868 6072 17877 6100
rect 17865 6069 17877 6072
rect 17911 6100 17923 6103
rect 19886 6100 19892 6112
rect 17911 6072 19892 6100
rect 17911 6069 17923 6072
rect 17865 6063 17923 6069
rect 19886 6060 19892 6072
rect 19944 6060 19950 6112
rect 20438 6060 20444 6112
rect 20496 6060 20502 6112
rect 1104 6010 20884 6032
rect 1104 5958 3422 6010
rect 3474 5958 3486 6010
rect 3538 5958 3550 6010
rect 3602 5958 3614 6010
rect 3666 5958 3678 6010
rect 3730 5958 8367 6010
rect 8419 5958 8431 6010
rect 8483 5958 8495 6010
rect 8547 5958 8559 6010
rect 8611 5958 8623 6010
rect 8675 5958 13312 6010
rect 13364 5958 13376 6010
rect 13428 5958 13440 6010
rect 13492 5958 13504 6010
rect 13556 5958 13568 6010
rect 13620 5958 18257 6010
rect 18309 5958 18321 6010
rect 18373 5958 18385 6010
rect 18437 5958 18449 6010
rect 18501 5958 18513 6010
rect 18565 5958 20884 6010
rect 1104 5936 20884 5958
rect 2774 5896 2780 5908
rect 1504 5868 2780 5896
rect 1118 5720 1124 5772
rect 1176 5720 1182 5772
rect 1136 5624 1164 5720
rect 1504 5701 1532 5868
rect 2774 5856 2780 5868
rect 2832 5856 2838 5908
rect 3053 5899 3111 5905
rect 3053 5865 3065 5899
rect 3099 5896 3111 5899
rect 3234 5896 3240 5908
rect 3099 5868 3240 5896
rect 3099 5865 3111 5868
rect 3053 5859 3111 5865
rect 3234 5856 3240 5868
rect 3292 5856 3298 5908
rect 3970 5856 3976 5908
rect 4028 5856 4034 5908
rect 6822 5896 6828 5908
rect 4540 5868 6828 5896
rect 2041 5763 2099 5769
rect 2041 5760 2053 5763
rect 1780 5732 2053 5760
rect 1489 5695 1547 5701
rect 1489 5661 1501 5695
rect 1535 5661 1547 5695
rect 1489 5655 1547 5661
rect 1670 5624 1676 5636
rect 1136 5596 1676 5624
rect 1670 5584 1676 5596
rect 1728 5624 1734 5636
rect 1780 5624 1808 5732
rect 2041 5729 2053 5732
rect 2087 5729 2099 5763
rect 4154 5760 4160 5772
rect 2041 5723 2099 5729
rect 3620 5732 4160 5760
rect 1857 5695 1915 5701
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2315 5695 2373 5701
rect 2315 5661 2327 5695
rect 2361 5692 2373 5695
rect 2406 5692 2412 5704
rect 2361 5664 2412 5692
rect 2361 5661 2373 5664
rect 2315 5655 2373 5661
rect 1728 5596 1808 5624
rect 1872 5624 1900 5655
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 3620 5701 3648 5732
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5661 3663 5695
rect 4430 5692 4436 5704
rect 3605 5655 3663 5661
rect 3712 5664 4436 5692
rect 3712 5624 3740 5664
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4540 5701 4568 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7009 5899 7067 5905
rect 7009 5896 7021 5899
rect 6972 5868 7021 5896
rect 6972 5856 6978 5868
rect 7009 5865 7021 5868
rect 7055 5865 7067 5899
rect 9214 5896 9220 5908
rect 7009 5859 7067 5865
rect 8956 5868 9220 5896
rect 7190 5828 7196 5840
rect 6840 5800 7196 5828
rect 5810 5720 5816 5772
rect 5868 5760 5874 5772
rect 5997 5763 6055 5769
rect 5997 5760 6009 5763
rect 5868 5732 6009 5760
rect 5868 5720 5874 5732
rect 5997 5729 6009 5732
rect 6043 5729 6055 5763
rect 5997 5723 6055 5729
rect 4525 5695 4583 5701
rect 4525 5661 4537 5695
rect 4571 5661 4583 5695
rect 4525 5655 4583 5661
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5661 4675 5695
rect 4617 5655 4675 5661
rect 4891 5695 4949 5701
rect 4891 5661 4903 5695
rect 4937 5692 4949 5695
rect 5534 5692 5540 5704
rect 4937 5664 5540 5692
rect 4937 5661 4949 5664
rect 4891 5655 4949 5661
rect 1872 5596 3740 5624
rect 1728 5584 1734 5596
rect 1780 5556 1808 5596
rect 3878 5584 3884 5636
rect 3936 5584 3942 5636
rect 4632 5624 4660 5655
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 5074 5624 5080 5636
rect 4632 5596 5080 5624
rect 5074 5584 5080 5596
rect 5132 5624 5138 5636
rect 5828 5624 5856 5720
rect 6271 5695 6329 5701
rect 6271 5661 6283 5695
rect 6317 5692 6329 5695
rect 6840 5692 6868 5800
rect 7190 5788 7196 5800
rect 7248 5788 7254 5840
rect 8386 5720 8392 5772
rect 8444 5760 8450 5772
rect 8956 5769 8984 5868
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9950 5856 9956 5908
rect 10008 5856 10014 5908
rect 11330 5856 11336 5908
rect 11388 5856 11394 5908
rect 12250 5856 12256 5908
rect 12308 5896 12314 5908
rect 12621 5899 12679 5905
rect 12308 5868 12570 5896
rect 12308 5856 12314 5868
rect 9766 5828 9772 5840
rect 9600 5800 9772 5828
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 8444 5732 8953 5760
rect 8444 5720 8450 5732
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 6317 5664 6868 5692
rect 9214 5671 9220 5704
rect 9199 5665 9220 5671
rect 6317 5661 6329 5664
rect 6271 5655 6329 5661
rect 5132 5596 5856 5624
rect 5132 5584 5138 5596
rect 6362 5584 6368 5636
rect 6420 5624 6426 5636
rect 8754 5624 8760 5636
rect 6420 5596 8760 5624
rect 6420 5584 6426 5596
rect 8754 5584 8760 5596
rect 8812 5584 8818 5636
rect 9199 5631 9211 5665
rect 9272 5652 9278 5704
rect 9600 5692 9628 5800
rect 9766 5788 9772 5800
rect 9824 5788 9830 5840
rect 12437 5831 12495 5837
rect 12437 5828 12449 5831
rect 12176 5800 12449 5828
rect 12176 5772 12204 5800
rect 12437 5797 12449 5800
rect 12483 5797 12495 5831
rect 12542 5828 12570 5868
rect 12621 5865 12633 5899
rect 12667 5896 12679 5899
rect 12710 5896 12716 5908
rect 12667 5868 12716 5896
rect 12667 5865 12679 5868
rect 12621 5859 12679 5865
rect 12710 5856 12716 5868
rect 12768 5856 12774 5908
rect 12897 5899 12955 5905
rect 12897 5865 12909 5899
rect 12943 5896 12955 5899
rect 12943 5868 15332 5896
rect 12943 5865 12955 5868
rect 12897 5859 12955 5865
rect 12542 5800 12572 5828
rect 12437 5791 12495 5797
rect 12158 5720 12164 5772
rect 12216 5720 12222 5772
rect 9324 5664 9628 5692
rect 9245 5634 9260 5652
rect 9245 5631 9257 5634
rect 9199 5625 9257 5631
rect 2498 5556 2504 5568
rect 1780 5528 2504 5556
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 3418 5516 3424 5568
rect 3476 5516 3482 5568
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4341 5559 4399 5565
rect 4341 5556 4353 5559
rect 4120 5528 4353 5556
rect 4120 5516 4126 5528
rect 4341 5525 4353 5528
rect 4387 5525 4399 5559
rect 4341 5519 4399 5525
rect 5534 5516 5540 5568
rect 5592 5556 5598 5568
rect 5629 5559 5687 5565
rect 5629 5556 5641 5559
rect 5592 5528 5641 5556
rect 5592 5516 5598 5528
rect 5629 5525 5641 5528
rect 5675 5525 5687 5559
rect 5629 5519 5687 5525
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 9324 5556 9352 5664
rect 9766 5652 9772 5704
rect 9824 5692 9830 5704
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 9824 5664 10333 5692
rect 9824 5652 9830 5664
rect 10321 5661 10333 5664
rect 10367 5661 10379 5695
rect 10321 5655 10379 5661
rect 10595 5695 10653 5701
rect 10595 5661 10607 5695
rect 10641 5692 10653 5695
rect 11790 5692 11796 5704
rect 10641 5664 11796 5692
rect 10641 5661 10653 5664
rect 10595 5655 10653 5661
rect 11790 5652 11796 5664
rect 11848 5652 11854 5704
rect 11977 5695 12035 5701
rect 11977 5661 11989 5695
rect 12023 5692 12035 5695
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 12023 5664 12265 5692
rect 12023 5661 12035 5664
rect 11977 5655 12035 5661
rect 12253 5661 12265 5664
rect 12299 5692 12311 5695
rect 12434 5692 12440 5704
rect 12299 5664 12440 5692
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 12544 5701 12572 5800
rect 12618 5800 13032 5828
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5661 12587 5695
rect 12529 5655 12587 5661
rect 10226 5584 10232 5636
rect 10284 5624 10290 5636
rect 12618 5624 12646 5800
rect 13004 5760 13032 5800
rect 13078 5788 13084 5840
rect 13136 5828 13142 5840
rect 13541 5831 13599 5837
rect 13541 5828 13553 5831
rect 13136 5800 13553 5828
rect 13136 5788 13142 5800
rect 13541 5797 13553 5800
rect 13587 5797 13599 5831
rect 13541 5791 13599 5797
rect 13648 5800 13952 5828
rect 13648 5760 13676 5800
rect 13924 5772 13952 5800
rect 13998 5788 14004 5840
rect 14056 5828 14062 5840
rect 15304 5828 15332 5868
rect 15378 5856 15384 5908
rect 15436 5896 15442 5908
rect 18509 5899 18567 5905
rect 18509 5896 18521 5899
rect 15436 5868 18521 5896
rect 15436 5856 15442 5868
rect 18509 5865 18521 5868
rect 18555 5865 18567 5899
rect 18509 5859 18567 5865
rect 18782 5856 18788 5908
rect 18840 5896 18846 5908
rect 20070 5896 20076 5908
rect 18840 5868 20076 5896
rect 18840 5856 18846 5868
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 15562 5828 15568 5840
rect 14056 5800 14136 5828
rect 15304 5800 15568 5828
rect 14056 5788 14062 5800
rect 13004 5732 13676 5760
rect 13722 5720 13728 5772
rect 13780 5760 13786 5772
rect 13780 5732 13860 5760
rect 13780 5720 13786 5732
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 12894 5692 12900 5704
rect 12851 5664 12900 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 12894 5652 12900 5664
rect 12952 5652 12958 5704
rect 13541 5695 13599 5701
rect 13081 5689 13139 5695
rect 13081 5682 13093 5689
rect 13004 5655 13093 5682
rect 13127 5655 13139 5689
rect 13541 5661 13553 5695
rect 13587 5661 13599 5695
rect 13832 5692 13860 5732
rect 13906 5720 13912 5772
rect 13964 5720 13970 5772
rect 14108 5769 14136 5800
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 15746 5788 15752 5840
rect 15804 5828 15810 5840
rect 16301 5831 16359 5837
rect 16301 5828 16313 5831
rect 15804 5800 16313 5828
rect 15804 5788 15810 5800
rect 16301 5797 16313 5800
rect 16347 5797 16359 5831
rect 16301 5791 16359 5797
rect 16669 5831 16727 5837
rect 16669 5797 16681 5831
rect 16715 5828 16727 5831
rect 17126 5828 17132 5840
rect 16715 5800 17132 5828
rect 16715 5797 16727 5800
rect 16669 5791 16727 5797
rect 17126 5788 17132 5800
rect 17184 5788 17190 5840
rect 14093 5763 14151 5769
rect 14093 5729 14105 5763
rect 14139 5729 14151 5763
rect 14093 5723 14151 5729
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 15528 5732 16896 5760
rect 15528 5720 15534 5732
rect 14366 5692 14372 5704
rect 13832 5664 14136 5692
rect 14327 5664 14372 5692
rect 13541 5655 13599 5661
rect 13004 5654 13139 5655
rect 10284 5596 12646 5624
rect 10284 5584 10290 5596
rect 13004 5568 13032 5654
rect 13081 5649 13139 5654
rect 13556 5624 13584 5655
rect 14108 5636 14136 5664
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 15378 5692 15384 5704
rect 14458 5664 15384 5692
rect 13188 5596 13584 5624
rect 7156 5528 9352 5556
rect 7156 5516 7162 5528
rect 10042 5516 10048 5568
rect 10100 5556 10106 5568
rect 10778 5556 10784 5568
rect 10100 5528 10784 5556
rect 10100 5516 10106 5528
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 12986 5516 12992 5568
rect 13044 5516 13050 5568
rect 13188 5565 13216 5596
rect 13630 5584 13636 5636
rect 13688 5624 13694 5636
rect 13688 5596 13860 5624
rect 13688 5584 13694 5596
rect 13173 5559 13231 5565
rect 13173 5525 13185 5559
rect 13219 5525 13231 5559
rect 13173 5519 13231 5525
rect 13446 5516 13452 5568
rect 13504 5556 13510 5568
rect 13722 5556 13728 5568
rect 13504 5528 13728 5556
rect 13504 5516 13510 5528
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 13832 5556 13860 5596
rect 13906 5584 13912 5636
rect 13964 5584 13970 5636
rect 14090 5584 14096 5636
rect 14148 5584 14154 5636
rect 14458 5556 14486 5664
rect 15378 5652 15384 5664
rect 15436 5652 15442 5704
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5661 15715 5695
rect 15657 5655 15715 5661
rect 16025 5695 16083 5701
rect 16025 5661 16037 5695
rect 16071 5694 16083 5695
rect 16071 5692 16160 5694
rect 16206 5692 16212 5704
rect 16071 5666 16212 5692
rect 16071 5661 16083 5666
rect 16132 5664 16212 5666
rect 16025 5655 16083 5661
rect 14826 5584 14832 5636
rect 14884 5624 14890 5636
rect 15672 5624 15700 5655
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 16482 5692 16488 5704
rect 16439 5664 16488 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 16868 5701 16896 5732
rect 18138 5720 18144 5772
rect 18196 5760 18202 5772
rect 19061 5763 19119 5769
rect 19061 5760 19073 5763
rect 18196 5732 19073 5760
rect 18196 5720 18202 5732
rect 19061 5729 19073 5732
rect 19107 5760 19119 5763
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 19107 5732 19257 5760
rect 19107 5729 19119 5732
rect 19061 5723 19119 5729
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 16853 5695 16911 5701
rect 16853 5661 16865 5695
rect 16899 5661 16911 5695
rect 16853 5655 16911 5661
rect 17129 5695 17187 5701
rect 17129 5661 17141 5695
rect 17175 5692 17187 5695
rect 17954 5692 17960 5704
rect 17175 5664 17960 5692
rect 17175 5661 17187 5664
rect 17129 5655 17187 5661
rect 17954 5652 17960 5664
rect 18012 5692 18018 5704
rect 18782 5692 18788 5704
rect 18012 5664 18788 5692
rect 18012 5652 18018 5664
rect 18782 5652 18788 5664
rect 18840 5652 18846 5704
rect 19519 5695 19577 5701
rect 19519 5661 19531 5695
rect 19565 5692 19577 5695
rect 20162 5692 20168 5704
rect 19565 5664 20168 5692
rect 19565 5661 19577 5664
rect 19519 5655 19577 5661
rect 20162 5652 20168 5664
rect 20220 5652 20226 5704
rect 16114 5624 16120 5636
rect 14884 5596 15611 5624
rect 15672 5596 16120 5624
rect 14884 5584 14890 5596
rect 13832 5528 14486 5556
rect 14642 5516 14648 5568
rect 14700 5556 14706 5568
rect 15105 5559 15163 5565
rect 15105 5556 15117 5559
rect 14700 5528 15117 5556
rect 14700 5516 14706 5528
rect 15105 5525 15117 5528
rect 15151 5525 15163 5559
rect 15105 5519 15163 5525
rect 15194 5516 15200 5568
rect 15252 5556 15258 5568
rect 15378 5556 15384 5568
rect 15252 5528 15384 5556
rect 15252 5516 15258 5528
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 15583 5556 15611 5596
rect 16114 5584 16120 5596
rect 16172 5584 16178 5636
rect 16666 5584 16672 5636
rect 16724 5624 16730 5636
rect 17374 5627 17432 5633
rect 17374 5624 17386 5627
rect 16724 5596 17386 5624
rect 16724 5584 16730 5596
rect 17374 5593 17386 5596
rect 17420 5593 17432 5627
rect 17374 5587 17432 5593
rect 17862 5584 17868 5636
rect 17920 5624 17926 5636
rect 18877 5627 18935 5633
rect 18877 5624 18889 5627
rect 17920 5596 18889 5624
rect 17920 5584 17926 5596
rect 18877 5593 18889 5596
rect 18923 5593 18935 5627
rect 18877 5587 18935 5593
rect 19610 5584 19616 5636
rect 19668 5624 19674 5636
rect 19794 5624 19800 5636
rect 19668 5596 19800 5624
rect 19668 5584 19674 5596
rect 19794 5584 19800 5596
rect 19852 5584 19858 5636
rect 16850 5556 16856 5568
rect 15583 5528 16856 5556
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 16942 5516 16948 5568
rect 17000 5556 17006 5568
rect 20257 5559 20315 5565
rect 20257 5556 20269 5559
rect 17000 5528 20269 5556
rect 17000 5516 17006 5528
rect 20257 5525 20269 5528
rect 20303 5525 20315 5559
rect 20257 5519 20315 5525
rect 1104 5466 21043 5488
rect 1104 5414 5894 5466
rect 5946 5414 5958 5466
rect 6010 5414 6022 5466
rect 6074 5414 6086 5466
rect 6138 5414 6150 5466
rect 6202 5414 10839 5466
rect 10891 5414 10903 5466
rect 10955 5414 10967 5466
rect 11019 5414 11031 5466
rect 11083 5414 11095 5466
rect 11147 5414 15784 5466
rect 15836 5414 15848 5466
rect 15900 5414 15912 5466
rect 15964 5414 15976 5466
rect 16028 5414 16040 5466
rect 16092 5414 20729 5466
rect 20781 5414 20793 5466
rect 20845 5414 20857 5466
rect 20909 5414 20921 5466
rect 20973 5414 20985 5466
rect 21037 5414 21043 5466
rect 1104 5392 21043 5414
rect 1302 5312 1308 5364
rect 1360 5352 1366 5364
rect 1581 5355 1639 5361
rect 1581 5352 1593 5355
rect 1360 5324 1593 5352
rect 1360 5312 1366 5324
rect 1581 5321 1593 5324
rect 1627 5321 1639 5355
rect 1581 5315 1639 5321
rect 1949 5355 2007 5361
rect 1949 5321 1961 5355
rect 1995 5352 2007 5355
rect 3878 5352 3884 5364
rect 1995 5324 3884 5352
rect 1995 5321 2007 5324
rect 1949 5315 2007 5321
rect 3878 5312 3884 5324
rect 3936 5312 3942 5364
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 5442 5352 5448 5364
rect 4028 5324 5448 5352
rect 4028 5312 4034 5324
rect 5442 5312 5448 5324
rect 5500 5312 5506 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6270 5352 6276 5364
rect 6227 5324 6276 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 6270 5312 6276 5324
rect 6328 5312 6334 5364
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 7006 5352 7012 5364
rect 6788 5324 7012 5352
rect 6788 5312 6794 5324
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7834 5312 7840 5364
rect 7892 5312 7898 5364
rect 7926 5312 7932 5364
rect 7984 5352 7990 5364
rect 9214 5352 9220 5364
rect 7984 5324 9220 5352
rect 7984 5312 7990 5324
rect 9214 5312 9220 5324
rect 9272 5312 9278 5364
rect 9398 5312 9404 5364
rect 9456 5312 9462 5364
rect 10042 5312 10048 5364
rect 10100 5312 10106 5364
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 10781 5355 10839 5361
rect 10781 5352 10793 5355
rect 10744 5324 10793 5352
rect 10744 5312 10750 5324
rect 10781 5321 10793 5324
rect 10827 5321 10839 5355
rect 10781 5315 10839 5321
rect 11149 5355 11207 5361
rect 11149 5321 11161 5355
rect 11195 5352 11207 5355
rect 11238 5352 11244 5364
rect 11195 5324 11244 5352
rect 11195 5321 11207 5324
rect 11149 5315 11207 5321
rect 11238 5312 11244 5324
rect 11296 5312 11302 5364
rect 11698 5312 11704 5364
rect 11756 5312 11762 5364
rect 11790 5312 11796 5364
rect 11848 5312 11854 5364
rect 12069 5355 12127 5361
rect 12069 5321 12081 5355
rect 12115 5352 12127 5355
rect 12250 5352 12256 5364
rect 12115 5324 12256 5352
rect 12115 5321 12127 5324
rect 12069 5315 12127 5321
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 12529 5355 12587 5361
rect 12529 5321 12541 5355
rect 12575 5352 12587 5355
rect 13354 5352 13360 5364
rect 12575 5324 13360 5352
rect 12575 5321 12587 5324
rect 12529 5315 12587 5321
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 13630 5352 13636 5364
rect 13554 5324 13636 5352
rect 6549 5287 6607 5293
rect 6549 5253 6561 5287
rect 6595 5284 6607 5287
rect 6595 5256 7604 5284
rect 6595 5253 6607 5256
rect 6549 5247 6607 5253
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5216 1547 5219
rect 1946 5216 1952 5228
rect 1535 5188 1952 5216
rect 1535 5185 1547 5188
rect 1489 5179 1547 5185
rect 1946 5176 1952 5188
rect 2004 5176 2010 5228
rect 2130 5176 2136 5228
rect 2188 5176 2194 5228
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5216 2283 5219
rect 2314 5216 2320 5228
rect 2271 5188 2320 5216
rect 2271 5185 2283 5188
rect 2225 5179 2283 5185
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 2406 5176 2412 5228
rect 2464 5176 2470 5228
rect 2590 5176 2596 5228
rect 2648 5176 2654 5228
rect 3372 5176 3378 5228
rect 3430 5225 3436 5228
rect 3430 5219 3479 5225
rect 3430 5185 3433 5219
rect 3467 5185 3479 5219
rect 3430 5179 3479 5185
rect 3430 5176 3436 5179
rect 4430 5176 4436 5228
rect 4488 5176 4494 5228
rect 4522 5176 4528 5228
rect 4580 5176 4586 5228
rect 5350 5222 5356 5228
rect 5294 5188 5356 5222
rect 5408 5225 5414 5228
rect 5408 5219 5436 5225
rect 5350 5176 5356 5188
rect 5424 5185 5436 5219
rect 5408 5179 5436 5185
rect 5408 5176 5414 5179
rect 5534 5176 5540 5228
rect 5592 5176 5598 5228
rect 6822 5176 6828 5228
rect 6880 5176 6886 5228
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 7190 5216 7196 5228
rect 6963 5188 7196 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 7285 5219 7343 5225
rect 7285 5185 7297 5219
rect 7331 5216 7343 5219
rect 7374 5216 7380 5228
rect 7331 5188 7380 5216
rect 7331 5185 7343 5188
rect 7285 5179 7343 5185
rect 7374 5176 7380 5188
rect 7432 5176 7438 5228
rect 7576 5216 7604 5256
rect 7650 5244 7656 5296
rect 7708 5244 7714 5296
rect 10060 5284 10088 5312
rect 7760 5256 10088 5284
rect 7760 5216 7788 5256
rect 10318 5244 10324 5296
rect 10376 5284 10382 5296
rect 10376 5256 10456 5284
rect 10376 5244 10382 5256
rect 7576 5188 7788 5216
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 8662 5216 8668 5228
rect 8623 5188 8668 5216
rect 8662 5176 8668 5188
rect 8720 5176 8726 5228
rect 9030 5176 9036 5228
rect 9088 5176 9094 5228
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 10011 5219 10069 5225
rect 10011 5216 10023 5219
rect 9272 5188 10023 5216
rect 9272 5176 9278 5188
rect 10011 5185 10023 5188
rect 10057 5185 10069 5219
rect 10428 5216 10456 5256
rect 11716 5225 11744 5312
rect 11790 5256 12110 5284
rect 11333 5219 11391 5225
rect 11333 5216 11345 5219
rect 10428 5188 11345 5216
rect 10011 5179 10069 5185
rect 11333 5185 11345 5188
rect 11379 5185 11391 5219
rect 11333 5179 11391 5185
rect 11701 5219 11759 5225
rect 11701 5185 11713 5219
rect 11747 5185 11759 5219
rect 11701 5179 11759 5185
rect 2608 5148 2636 5176
rect 2240 5120 2636 5148
rect 2240 5092 2268 5120
rect 2774 5108 2780 5160
rect 2832 5148 2838 5160
rect 3145 5151 3203 5157
rect 3145 5148 3157 5151
rect 2832 5120 3157 5148
rect 2832 5108 2838 5120
rect 3145 5117 3157 5120
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 3283 5151 3341 5157
rect 3283 5117 3295 5151
rect 3329 5148 3341 5151
rect 3329 5120 3832 5148
rect 3329 5117 3341 5120
rect 3283 5111 3341 5117
rect 2222 5040 2228 5092
rect 2280 5040 2286 5092
rect 2590 5040 2596 5092
rect 2648 5080 2654 5092
rect 2869 5083 2927 5089
rect 2869 5080 2881 5083
rect 2648 5052 2881 5080
rect 2648 5040 2654 5052
rect 2869 5049 2881 5052
rect 2915 5049 2927 5083
rect 3804 5080 3832 5120
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 4341 5151 4399 5157
rect 4341 5148 4353 5151
rect 4212 5120 4353 5148
rect 4212 5108 4218 5120
rect 4341 5117 4353 5120
rect 4387 5117 4399 5151
rect 4448 5148 4476 5176
rect 6368 5160 6420 5166
rect 5261 5151 5319 5157
rect 5261 5148 5273 5151
rect 4448 5120 5273 5148
rect 4341 5111 4399 5117
rect 5261 5117 5273 5120
rect 5307 5117 5319 5151
rect 5261 5111 5319 5117
rect 9048 5148 9076 5176
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9048 5120 9781 5148
rect 9769 5117 9781 5120
rect 9815 5117 9827 5151
rect 9769 5111 9827 5117
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 11514 5148 11520 5160
rect 11020 5120 11520 5148
rect 11020 5108 11026 5120
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 6368 5102 6420 5108
rect 3970 5080 3976 5092
rect 3804 5052 3976 5080
rect 2869 5043 2927 5049
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 4985 5083 5043 5089
rect 4985 5049 4997 5083
rect 5031 5049 5043 5083
rect 4985 5043 5043 5049
rect 2774 4972 2780 5024
rect 2832 5012 2838 5024
rect 4065 5015 4123 5021
rect 4065 5012 4077 5015
rect 2832 4984 4077 5012
rect 2832 4972 2838 4984
rect 4065 4981 4077 4984
rect 4111 4981 4123 5015
rect 5000 5012 5028 5043
rect 10686 5040 10692 5092
rect 10744 5080 10750 5092
rect 11790 5080 11818 5256
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 11900 5148 11928 5179
rect 12082 5148 12110 5256
rect 12158 5244 12164 5296
rect 12216 5244 12222 5296
rect 13554 5284 13582 5324
rect 13630 5312 13636 5324
rect 13688 5312 13694 5364
rect 13722 5312 13728 5364
rect 13780 5352 13786 5364
rect 14182 5352 14188 5364
rect 13780 5324 14188 5352
rect 13780 5312 13786 5324
rect 14182 5312 14188 5324
rect 14240 5312 14246 5364
rect 14734 5352 14740 5364
rect 14292 5324 14740 5352
rect 14292 5296 14320 5324
rect 14734 5312 14740 5324
rect 14792 5352 14798 5364
rect 14918 5352 14924 5364
rect 14792 5324 14924 5352
rect 14792 5312 14798 5324
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15102 5312 15108 5364
rect 15160 5352 15166 5364
rect 15197 5355 15255 5361
rect 15197 5352 15209 5355
rect 15160 5324 15209 5352
rect 15160 5312 15166 5324
rect 15197 5321 15209 5324
rect 15243 5321 15255 5355
rect 15197 5315 15255 5321
rect 15378 5312 15384 5364
rect 15436 5352 15442 5364
rect 15746 5352 15752 5364
rect 15436 5324 15752 5352
rect 15436 5312 15442 5324
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 16206 5312 16212 5364
rect 16264 5352 16270 5364
rect 17497 5355 17555 5361
rect 16264 5324 17448 5352
rect 16264 5312 16270 5324
rect 13970 5287 14028 5293
rect 13970 5284 13982 5287
rect 12820 5256 13582 5284
rect 13648 5256 13982 5284
rect 12176 5216 12204 5244
rect 12253 5219 12311 5225
rect 12253 5216 12265 5219
rect 12176 5188 12265 5216
rect 12253 5185 12265 5188
rect 12299 5185 12311 5219
rect 12253 5179 12311 5185
rect 12345 5219 12403 5225
rect 12345 5185 12357 5219
rect 12391 5216 12403 5219
rect 12710 5216 12716 5228
rect 12391 5188 12716 5216
rect 12391 5185 12403 5188
rect 12345 5179 12403 5185
rect 12710 5176 12716 5188
rect 12768 5176 12774 5228
rect 12820 5225 12848 5256
rect 13648 5228 13676 5256
rect 13970 5253 13982 5256
rect 14016 5253 14028 5287
rect 13970 5247 14028 5253
rect 14274 5244 14280 5296
rect 14332 5244 14338 5296
rect 15010 5244 15016 5296
rect 15068 5284 15074 5296
rect 16021 5287 16079 5293
rect 15068 5256 15884 5284
rect 15068 5244 15074 5256
rect 12805 5219 12863 5225
rect 12805 5185 12817 5219
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 13078 5176 13084 5228
rect 13136 5176 13142 5228
rect 13262 5176 13268 5228
rect 13320 5176 13326 5228
rect 13354 5176 13360 5228
rect 13412 5176 13418 5228
rect 13541 5219 13599 5225
rect 13541 5185 13553 5219
rect 13587 5185 13599 5219
rect 13541 5179 13599 5185
rect 12526 5148 12532 5160
rect 11900 5120 12002 5148
rect 12082 5120 12532 5148
rect 10744 5052 11818 5080
rect 11974 5080 12002 5120
rect 12526 5108 12532 5120
rect 12584 5108 12590 5160
rect 12621 5083 12679 5089
rect 12621 5080 12633 5083
rect 11974 5052 12633 5080
rect 10744 5040 10750 5052
rect 12621 5049 12633 5052
rect 12667 5049 12679 5083
rect 12621 5043 12679 5049
rect 12710 5040 12716 5092
rect 12768 5080 12774 5092
rect 13078 5080 13084 5092
rect 12768 5052 13084 5080
rect 12768 5040 12774 5052
rect 13078 5040 13084 5052
rect 13136 5040 13142 5092
rect 13280 5089 13308 5176
rect 13370 5148 13398 5176
rect 13556 5148 13584 5179
rect 13630 5176 13636 5228
rect 13688 5176 13694 5228
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 13832 5188 14872 5216
rect 13832 5148 13860 5188
rect 13370 5120 13860 5148
rect 14844 5148 14872 5188
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 14976 5188 15393 5216
rect 14976 5176 14982 5188
rect 15381 5185 15393 5188
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 15470 5176 15476 5228
rect 15528 5176 15534 5228
rect 15657 5219 15715 5225
rect 15657 5185 15669 5219
rect 15703 5216 15715 5219
rect 15703 5188 15792 5216
rect 15703 5185 15715 5188
rect 15657 5179 15715 5185
rect 15194 5148 15200 5160
rect 14844 5120 15200 5148
rect 15194 5108 15200 5120
rect 15252 5108 15258 5160
rect 13265 5083 13323 5089
rect 13265 5049 13277 5083
rect 13311 5049 13323 5083
rect 13265 5043 13323 5049
rect 13357 5083 13415 5089
rect 13357 5049 13369 5083
rect 13403 5080 13415 5083
rect 13538 5080 13544 5092
rect 13403 5052 13544 5080
rect 13403 5049 13415 5052
rect 13357 5043 13415 5049
rect 13538 5040 13544 5052
rect 13596 5040 13602 5092
rect 15102 5040 15108 5092
rect 15160 5040 15166 5092
rect 15378 5040 15384 5092
rect 15436 5080 15442 5092
rect 15657 5083 15715 5089
rect 15657 5080 15669 5083
rect 15436 5052 15669 5080
rect 15436 5040 15442 5052
rect 15657 5049 15669 5052
rect 15703 5049 15715 5083
rect 15764 5080 15792 5188
rect 15856 5148 15884 5256
rect 16021 5253 16033 5287
rect 16067 5284 16079 5287
rect 16758 5284 16764 5296
rect 16067 5256 16764 5284
rect 16067 5253 16079 5256
rect 16021 5247 16079 5253
rect 16758 5244 16764 5256
rect 16816 5244 16822 5296
rect 17420 5284 17448 5324
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 17586 5352 17592 5364
rect 17543 5324 17592 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 17678 5312 17684 5364
rect 17736 5352 17742 5364
rect 19978 5352 19984 5364
rect 17736 5324 19984 5352
rect 17736 5312 17742 5324
rect 19978 5312 19984 5324
rect 20036 5312 20042 5364
rect 17420 5256 20484 5284
rect 20456 5228 20484 5256
rect 16117 5219 16175 5225
rect 16117 5185 16129 5219
rect 16163 5216 16175 5219
rect 16298 5216 16304 5228
rect 16163 5188 16304 5216
rect 16163 5185 16175 5188
rect 16117 5179 16175 5185
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 16482 5176 16488 5228
rect 16540 5216 16546 5228
rect 16853 5219 16911 5225
rect 16853 5216 16865 5219
rect 16540 5188 16865 5216
rect 16540 5176 16546 5188
rect 16853 5185 16865 5188
rect 16899 5185 16911 5219
rect 16853 5179 16911 5185
rect 17034 5176 17040 5228
rect 17092 5176 17098 5228
rect 17405 5219 17463 5225
rect 17405 5185 17417 5219
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 17420 5148 17448 5179
rect 17494 5176 17500 5228
rect 17552 5176 17558 5228
rect 17678 5176 17684 5228
rect 17736 5176 17742 5228
rect 17955 5219 18013 5225
rect 17955 5185 17967 5219
rect 18001 5216 18013 5219
rect 18782 5216 18788 5228
rect 18001 5188 18788 5216
rect 18001 5185 18013 5188
rect 17955 5179 18013 5185
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 18874 5176 18880 5228
rect 18932 5216 18938 5228
rect 19426 5225 19432 5228
rect 19153 5219 19211 5225
rect 19153 5216 19165 5219
rect 18932 5188 19165 5216
rect 18932 5176 18938 5188
rect 19153 5185 19165 5188
rect 19199 5185 19211 5219
rect 19153 5179 19211 5185
rect 19420 5179 19432 5225
rect 19426 5176 19432 5179
rect 19484 5176 19490 5228
rect 20438 5176 20444 5228
rect 20496 5176 20502 5228
rect 15856 5120 16252 5148
rect 16114 5080 16120 5092
rect 15764 5052 16120 5080
rect 15657 5043 15715 5049
rect 16114 5040 16120 5052
rect 16172 5040 16178 5092
rect 16224 5080 16252 5120
rect 16390 5120 17448 5148
rect 16390 5080 16418 5120
rect 16224 5052 16418 5080
rect 17221 5083 17279 5089
rect 17221 5049 17233 5083
rect 17267 5080 17279 5083
rect 17512 5080 17540 5176
rect 18598 5108 18604 5160
rect 18656 5108 18662 5160
rect 17267 5052 17540 5080
rect 17267 5049 17279 5052
rect 17221 5043 17279 5049
rect 5350 5012 5356 5024
rect 5000 4984 5356 5012
rect 4065 4975 4123 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 13446 5012 13452 5024
rect 9916 4984 13452 5012
rect 9916 4972 9922 4984
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 13722 4972 13728 5024
rect 13780 5012 13786 5024
rect 14366 5012 14372 5024
rect 13780 4984 14372 5012
rect 13780 4972 13786 4984
rect 14366 4972 14372 4984
rect 14424 4972 14430 5024
rect 14458 4972 14464 5024
rect 14516 5012 14522 5024
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 14516 4984 16221 5012
rect 14516 4972 14522 4984
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16209 4975 16267 4981
rect 16482 4972 16488 5024
rect 16540 5012 16546 5024
rect 16669 5015 16727 5021
rect 16669 5012 16681 5015
rect 16540 4984 16681 5012
rect 16540 4972 16546 4984
rect 16669 4981 16681 4984
rect 16715 4981 16727 5015
rect 16669 4975 16727 4981
rect 16758 4972 16764 5024
rect 16816 5012 16822 5024
rect 18616 5012 18644 5108
rect 18690 5040 18696 5092
rect 18748 5040 18754 5092
rect 16816 4984 18644 5012
rect 16816 4972 16822 4984
rect 18782 4972 18788 5024
rect 18840 5012 18846 5024
rect 20533 5015 20591 5021
rect 20533 5012 20545 5015
rect 18840 4984 20545 5012
rect 18840 4972 18846 4984
rect 20533 4981 20545 4984
rect 20579 4981 20591 5015
rect 20533 4975 20591 4981
rect 1104 4922 20884 4944
rect 1104 4870 3422 4922
rect 3474 4870 3486 4922
rect 3538 4870 3550 4922
rect 3602 4870 3614 4922
rect 3666 4870 3678 4922
rect 3730 4870 8367 4922
rect 8419 4870 8431 4922
rect 8483 4870 8495 4922
rect 8547 4870 8559 4922
rect 8611 4870 8623 4922
rect 8675 4870 13312 4922
rect 13364 4870 13376 4922
rect 13428 4870 13440 4922
rect 13492 4870 13504 4922
rect 13556 4870 13568 4922
rect 13620 4870 18257 4922
rect 18309 4870 18321 4922
rect 18373 4870 18385 4922
rect 18437 4870 18449 4922
rect 18501 4870 18513 4922
rect 18565 4870 20884 4922
rect 1104 4848 20884 4870
rect 1210 4768 1216 4820
rect 1268 4808 1274 4820
rect 1581 4811 1639 4817
rect 1581 4808 1593 4811
rect 1268 4780 1593 4808
rect 1268 4768 1274 4780
rect 1581 4777 1593 4780
rect 1627 4777 1639 4811
rect 1581 4771 1639 4777
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2038 4808 2044 4820
rect 1995 4780 2044 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 2682 4808 2688 4820
rect 2148 4780 2688 4808
rect 566 4564 572 4616
rect 624 4564 630 4616
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4604 1547 4607
rect 1762 4604 1768 4616
rect 1535 4576 1768 4604
rect 1535 4573 1547 4576
rect 1489 4567 1547 4573
rect 1762 4564 1768 4576
rect 1820 4564 1826 4616
rect 2148 4613 2176 4780
rect 2682 4768 2688 4780
rect 2740 4768 2746 4820
rect 3326 4768 3332 4820
rect 3384 4768 3390 4820
rect 3510 4768 3516 4820
rect 3568 4808 3574 4820
rect 3970 4808 3976 4820
rect 3568 4780 3976 4808
rect 3568 4768 3574 4780
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 4126 4780 4537 4808
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 4126 4740 4154 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4525 4771 4583 4777
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 5040 4780 5181 4808
rect 5040 4768 5046 4780
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 5169 4771 5227 4777
rect 5276 4780 6316 4808
rect 3108 4712 4154 4740
rect 3108 4700 3114 4712
rect 3326 4632 3332 4684
rect 3384 4672 3390 4684
rect 5276 4672 5304 4780
rect 6288 4740 6316 4780
rect 6362 4768 6368 4820
rect 6420 4768 6426 4820
rect 7098 4808 7104 4820
rect 6472 4780 7104 4808
rect 6472 4740 6500 4780
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 7248 4780 7757 4808
rect 7248 4768 7254 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 7745 4771 7803 4777
rect 9858 4768 9864 4820
rect 9916 4768 9922 4820
rect 10502 4768 10508 4820
rect 10560 4808 10566 4820
rect 10781 4811 10839 4817
rect 10781 4808 10793 4811
rect 10560 4780 10793 4808
rect 10560 4768 10566 4780
rect 10781 4777 10793 4780
rect 10827 4777 10839 4811
rect 10781 4771 10839 4777
rect 10870 4768 10876 4820
rect 10928 4808 10934 4820
rect 11149 4811 11207 4817
rect 10928 4780 11098 4808
rect 10928 4768 10934 4780
rect 6288 4712 6500 4740
rect 7558 4700 7564 4752
rect 7616 4740 7622 4752
rect 9401 4743 9459 4749
rect 9401 4740 9413 4743
rect 7616 4712 9413 4740
rect 7616 4700 7622 4712
rect 9401 4709 9413 4712
rect 9447 4709 9459 4743
rect 9401 4703 9459 4709
rect 9490 4700 9496 4752
rect 9548 4740 9554 4752
rect 10321 4743 10379 4749
rect 10321 4740 10333 4743
rect 9548 4712 10333 4740
rect 9548 4700 9554 4712
rect 10321 4709 10333 4712
rect 10367 4709 10379 4743
rect 10321 4703 10379 4709
rect 10410 4700 10416 4752
rect 10468 4700 10474 4752
rect 10965 4743 11023 4749
rect 10965 4740 10977 4743
rect 10796 4712 10977 4740
rect 3384 4644 5304 4672
rect 3384 4632 3390 4644
rect 6730 4632 6736 4684
rect 6788 4632 6794 4684
rect 10042 4632 10048 4684
rect 10100 4632 10106 4684
rect 10428 4672 10456 4700
rect 10796 4684 10824 4712
rect 10965 4709 10977 4712
rect 11011 4709 11023 4743
rect 11070 4740 11098 4780
rect 11149 4777 11161 4811
rect 11195 4808 11207 4811
rect 11422 4808 11428 4820
rect 11195 4780 11428 4808
rect 11195 4777 11207 4780
rect 11149 4771 11207 4777
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 11606 4768 11612 4820
rect 11664 4808 11670 4820
rect 12437 4811 12495 4817
rect 12437 4808 12449 4811
rect 11664 4780 12449 4808
rect 11664 4768 11670 4780
rect 12437 4777 12449 4780
rect 12483 4777 12495 4811
rect 12437 4771 12495 4777
rect 12621 4811 12679 4817
rect 12621 4777 12633 4811
rect 12667 4808 12679 4811
rect 13078 4808 13084 4820
rect 12667 4780 13084 4808
rect 12667 4777 12679 4780
rect 12621 4771 12679 4777
rect 13078 4768 13084 4780
rect 13136 4768 13142 4820
rect 13173 4811 13231 4817
rect 13173 4777 13185 4811
rect 13219 4777 13231 4811
rect 13173 4771 13231 4777
rect 11793 4743 11851 4749
rect 11793 4740 11805 4743
rect 11070 4712 11805 4740
rect 10965 4703 11023 4709
rect 11793 4709 11805 4712
rect 11839 4709 11851 4743
rect 12897 4743 12955 4749
rect 12897 4740 12909 4743
rect 11793 4703 11851 4709
rect 12728 4712 12909 4740
rect 10428 4644 10640 4672
rect 2133 4607 2191 4613
rect 2133 4573 2145 4607
rect 2179 4573 2191 4607
rect 2133 4567 2191 4573
rect 2317 4607 2375 4613
rect 2317 4573 2329 4607
rect 2363 4604 2375 4607
rect 2498 4604 2504 4616
rect 2363 4576 2504 4604
rect 2363 4573 2375 4576
rect 2317 4567 2375 4573
rect 2498 4564 2504 4576
rect 2556 4564 2562 4616
rect 2591 4607 2649 4613
rect 2591 4573 2603 4607
rect 2637 4604 2649 4607
rect 3602 4604 3608 4616
rect 2637 4576 3608 4604
rect 2637 4573 2649 4576
rect 2591 4567 2649 4573
rect 3602 4564 3608 4576
rect 3660 4564 3666 4616
rect 3881 4607 3939 4613
rect 3881 4573 3893 4607
rect 3927 4604 3939 4607
rect 4062 4604 4068 4616
rect 3927 4576 4068 4604
rect 3927 4573 3939 4576
rect 3881 4567 3939 4573
rect 4062 4564 4068 4576
rect 4120 4564 4126 4616
rect 4522 4564 4528 4616
rect 4580 4564 4586 4616
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4573 5411 4607
rect 5595 4607 5653 4613
rect 5595 4604 5607 4607
rect 5353 4567 5411 4573
rect 5460 4576 5607 4604
rect 584 4468 612 4564
rect 1946 4496 1952 4548
rect 2004 4536 2010 4548
rect 4338 4536 4344 4548
rect 2004 4508 4344 4536
rect 2004 4496 2010 4508
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 4430 4496 4436 4548
rect 4488 4496 4494 4548
rect 4540 4536 4568 4564
rect 5077 4539 5135 4545
rect 5077 4536 5089 4539
rect 4540 4508 5089 4536
rect 5077 4505 5089 4508
rect 5123 4505 5135 4539
rect 5077 4499 5135 4505
rect 3973 4471 4031 4477
rect 3973 4468 3985 4471
rect 584 4440 3985 4468
rect 3973 4437 3985 4440
rect 4019 4437 4031 4471
rect 5368 4468 5396 4567
rect 5460 4548 5488 4576
rect 5595 4573 5607 4576
rect 5641 4573 5653 4607
rect 6748 4604 6776 4632
rect 5595 4567 5653 4573
rect 6564 4576 6776 4604
rect 10060 4604 10088 4632
rect 10612 4613 10640 4644
rect 10778 4632 10784 4684
rect 10836 4632 10842 4684
rect 11146 4632 11152 4684
rect 11204 4672 11210 4684
rect 11422 4672 11428 4684
rect 11204 4644 11428 4672
rect 11204 4632 11210 4644
rect 11422 4632 11428 4644
rect 11480 4632 11486 4684
rect 11882 4632 11888 4684
rect 11940 4632 11946 4684
rect 12161 4675 12219 4681
rect 12161 4641 12173 4675
rect 12207 4672 12219 4675
rect 12250 4672 12256 4684
rect 12207 4644 12256 4672
rect 12207 4641 12219 4644
rect 12161 4635 12219 4641
rect 12250 4632 12256 4644
rect 12308 4632 12314 4684
rect 12618 4672 12624 4684
rect 12360 4644 12624 4672
rect 10505 4607 10563 4613
rect 10505 4604 10517 4607
rect 6991 4577 7049 4583
rect 5442 4496 5448 4548
rect 5500 4496 5506 4548
rect 6564 4468 6592 4576
rect 6991 4574 7003 4577
rect 6730 4496 6736 4548
rect 6788 4536 6794 4548
rect 6886 4546 7003 4574
rect 6886 4536 6914 4546
rect 6991 4543 7003 4546
rect 7037 4543 7049 4577
rect 10060 4576 10517 4604
rect 10505 4573 10517 4576
rect 10551 4573 10563 4607
rect 10505 4567 10563 4573
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4573 10655 4607
rect 10597 4567 10655 4573
rect 10686 4564 10692 4616
rect 10744 4564 10750 4616
rect 10873 4607 10931 4613
rect 10873 4573 10885 4607
rect 10919 4573 10931 4607
rect 10873 4567 10931 4573
rect 6991 4537 7049 4543
rect 10704 4536 10732 4564
rect 6788 4508 6914 4536
rect 7114 4508 10732 4536
rect 10888 4536 10916 4567
rect 10962 4564 10968 4616
rect 11020 4604 11026 4616
rect 11333 4607 11391 4613
rect 11333 4604 11345 4607
rect 11020 4576 11345 4604
rect 11020 4564 11026 4576
rect 11333 4573 11345 4576
rect 11379 4573 11391 4607
rect 11333 4567 11391 4573
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4604 11759 4607
rect 11900 4604 11928 4632
rect 11747 4576 11928 4604
rect 11747 4573 11759 4576
rect 11701 4567 11759 4573
rect 11974 4564 11980 4616
rect 12032 4564 12038 4616
rect 12360 4613 12388 4644
rect 12618 4632 12624 4644
rect 12676 4632 12682 4684
rect 12069 4607 12127 4613
rect 12069 4573 12081 4607
rect 12115 4573 12127 4607
rect 12069 4567 12127 4573
rect 12345 4607 12403 4613
rect 12345 4573 12357 4607
rect 12391 4573 12403 4607
rect 12345 4567 12403 4573
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 12728 4604 12756 4712
rect 12897 4709 12909 4712
rect 12943 4709 12955 4743
rect 12897 4703 12955 4709
rect 12986 4700 12992 4752
rect 13044 4740 13050 4752
rect 13188 4740 13216 4771
rect 13814 4768 13820 4820
rect 13872 4768 13878 4820
rect 14090 4768 14096 4820
rect 14148 4808 14154 4820
rect 14921 4811 14979 4817
rect 14148 4780 14688 4808
rect 14148 4768 14154 4780
rect 13044 4712 13216 4740
rect 13044 4700 13050 4712
rect 13262 4700 13268 4752
rect 13320 4740 13326 4752
rect 14277 4743 14335 4749
rect 14277 4740 14289 4743
rect 13320 4712 14289 4740
rect 13320 4700 13326 4712
rect 14277 4709 14289 4712
rect 14323 4709 14335 4743
rect 14550 4740 14556 4752
rect 14277 4703 14335 4709
rect 14364 4712 14556 4740
rect 13170 4672 13176 4684
rect 13096 4644 13176 4672
rect 13096 4613 13124 4644
rect 13170 4632 13176 4644
rect 13228 4632 13234 4684
rect 13446 4632 13452 4684
rect 13504 4672 13510 4684
rect 14364 4672 14392 4712
rect 14550 4700 14556 4712
rect 14608 4700 14614 4752
rect 14660 4740 14688 4780
rect 14921 4777 14933 4811
rect 14967 4808 14979 4811
rect 15286 4808 15292 4820
rect 14967 4780 15292 4808
rect 14967 4777 14979 4780
rect 14921 4771 14979 4777
rect 15286 4768 15292 4780
rect 15344 4768 15350 4820
rect 15562 4808 15568 4820
rect 15396 4780 15568 4808
rect 15194 4740 15200 4752
rect 14660 4712 15200 4740
rect 15194 4700 15200 4712
rect 15252 4700 15258 4752
rect 13504 4644 14392 4672
rect 14461 4675 14519 4681
rect 13504 4632 13510 4644
rect 14461 4641 14473 4675
rect 14507 4672 14519 4675
rect 14642 4672 14648 4684
rect 14507 4644 14648 4672
rect 14507 4641 14519 4644
rect 14461 4635 14519 4641
rect 14642 4632 14648 4644
rect 14700 4672 14706 4684
rect 15105 4675 15163 4681
rect 14700 4644 15056 4672
rect 15105 4650 15117 4675
rect 15151 4650 15163 4675
rect 15396 4672 15424 4780
rect 15562 4768 15568 4780
rect 15620 4768 15626 4820
rect 15654 4768 15660 4820
rect 15712 4808 15718 4820
rect 18782 4808 18788 4820
rect 15712 4780 18788 4808
rect 15712 4768 15718 4780
rect 18782 4768 18788 4780
rect 18840 4768 18846 4820
rect 17310 4700 17316 4752
rect 17368 4740 17374 4752
rect 17589 4743 17647 4749
rect 17589 4740 17601 4743
rect 17368 4712 17601 4740
rect 17368 4700 17374 4712
rect 17589 4709 17601 4712
rect 17635 4709 17647 4743
rect 17589 4703 17647 4709
rect 17770 4700 17776 4752
rect 17828 4740 17834 4752
rect 19794 4740 19800 4752
rect 17828 4712 19800 4740
rect 17828 4700 17834 4712
rect 19794 4700 19800 4712
rect 19852 4700 19858 4752
rect 20070 4700 20076 4752
rect 20128 4700 20134 4752
rect 16666 4672 16672 4684
rect 14700 4632 14706 4644
rect 12575 4576 12756 4604
rect 12805 4607 12863 4613
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 12805 4573 12817 4607
rect 12851 4573 12863 4607
rect 12805 4567 12863 4573
rect 13081 4607 13139 4613
rect 13081 4573 13093 4607
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 10888 4508 11560 4536
rect 6788 4496 6794 4508
rect 5368 4440 6592 4468
rect 3973 4431 4031 4437
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 7114 4468 7142 4508
rect 6880 4440 7142 4468
rect 6880 4428 6886 4440
rect 10042 4428 10048 4480
rect 10100 4468 10106 4480
rect 11532 4477 11560 4508
rect 10137 4471 10195 4477
rect 10137 4468 10149 4471
rect 10100 4440 10149 4468
rect 10100 4428 10106 4440
rect 10137 4437 10149 4440
rect 10183 4437 10195 4471
rect 10137 4431 10195 4437
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4437 11575 4471
rect 11517 4431 11575 4437
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 12084 4468 12112 4567
rect 12434 4496 12440 4548
rect 12492 4536 12498 4548
rect 12820 4536 12848 4567
rect 13354 4564 13360 4616
rect 13412 4564 13418 4616
rect 13538 4564 13544 4616
rect 13596 4604 13602 4616
rect 13633 4607 13691 4613
rect 13633 4604 13645 4607
rect 13596 4576 13645 4604
rect 13596 4564 13602 4576
rect 13633 4573 13645 4576
rect 13679 4573 13691 4607
rect 13633 4567 13691 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4573 13783 4607
rect 13725 4567 13783 4573
rect 13909 4607 13967 4613
rect 13909 4573 13921 4607
rect 13955 4604 13967 4607
rect 13955 4576 14231 4604
rect 13955 4573 13967 4576
rect 13909 4567 13967 4573
rect 13372 4536 13400 4564
rect 12492 4508 12848 4536
rect 12912 4508 13400 4536
rect 13740 4536 13768 4567
rect 13998 4536 14004 4548
rect 13740 4508 14004 4536
rect 12492 4496 12498 4508
rect 11940 4440 12112 4468
rect 11940 4428 11946 4440
rect 12158 4428 12164 4480
rect 12216 4468 12222 4480
rect 12912 4468 12940 4508
rect 13998 4496 14004 4508
rect 14056 4496 14062 4548
rect 14203 4536 14231 4576
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 14734 4564 14740 4616
rect 14792 4564 14798 4616
rect 14826 4564 14832 4616
rect 14884 4564 14890 4616
rect 15028 4613 15056 4644
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4573 15071 4607
rect 15102 4598 15108 4650
rect 15160 4598 15166 4650
rect 15304 4644 15424 4672
rect 16390 4644 16672 4672
rect 15205 4607 15263 4613
rect 15013 4567 15071 4573
rect 15205 4573 15217 4607
rect 15251 4604 15263 4607
rect 15304 4604 15332 4644
rect 15251 4576 15332 4604
rect 15381 4607 15439 4613
rect 15251 4573 15263 4576
rect 15205 4567 15263 4573
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 16390 4604 16418 4644
rect 16666 4632 16672 4644
rect 16724 4632 16730 4684
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17405 4675 17463 4681
rect 17405 4672 17417 4675
rect 17000 4644 17417 4672
rect 17000 4632 17006 4644
rect 17405 4641 17417 4644
rect 17451 4641 17463 4675
rect 17405 4635 17463 4641
rect 18138 4632 18144 4684
rect 18196 4672 18202 4684
rect 20438 4672 20444 4684
rect 18196 4644 20444 4672
rect 18196 4632 18202 4644
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 15427 4576 16418 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 16574 4564 16580 4616
rect 16632 4604 16638 4616
rect 17589 4607 17647 4613
rect 17589 4604 17601 4607
rect 16632 4576 17601 4604
rect 16632 4564 16638 4576
rect 17589 4573 17601 4576
rect 17635 4573 17647 4607
rect 18049 4607 18107 4613
rect 18049 4604 18061 4607
rect 17589 4567 17647 4573
rect 17696 4576 18061 4604
rect 14645 4539 14703 4545
rect 14203 4508 14594 4536
rect 12216 4440 12940 4468
rect 12216 4428 12222 4440
rect 12986 4428 12992 4480
rect 13044 4468 13050 4480
rect 13449 4471 13507 4477
rect 13449 4468 13461 4471
rect 13044 4440 13461 4468
rect 13044 4428 13050 4440
rect 13449 4437 13461 4440
rect 13495 4437 13507 4471
rect 13449 4431 13507 4437
rect 14182 4428 14188 4480
rect 14240 4468 14246 4480
rect 14458 4468 14464 4480
rect 14240 4440 14464 4468
rect 14240 4428 14246 4440
rect 14458 4428 14464 4440
rect 14516 4428 14522 4480
rect 14566 4468 14594 4508
rect 14645 4505 14657 4539
rect 14691 4536 14703 4539
rect 14844 4536 14872 4564
rect 14691 4508 14872 4536
rect 14691 4505 14703 4508
rect 14645 4499 14703 4505
rect 14918 4496 14924 4548
rect 14976 4536 14982 4548
rect 15626 4539 15684 4545
rect 15626 4536 15638 4539
rect 14976 4508 15638 4536
rect 14976 4496 14982 4508
rect 15626 4505 15638 4508
rect 15672 4505 15684 4539
rect 15626 4499 15684 4505
rect 15746 4496 15752 4548
rect 15804 4536 15810 4548
rect 16945 4539 17003 4545
rect 16945 4536 16957 4539
rect 15804 4508 16957 4536
rect 15804 4496 15810 4508
rect 16945 4505 16957 4508
rect 16991 4505 17003 4539
rect 16945 4499 17003 4505
rect 17126 4496 17132 4548
rect 17184 4536 17190 4548
rect 17696 4536 17724 4576
rect 18049 4573 18061 4576
rect 18095 4573 18107 4607
rect 18049 4567 18107 4573
rect 18230 4564 18236 4616
rect 18288 4604 18294 4616
rect 18877 4607 18935 4613
rect 18877 4604 18889 4607
rect 18288 4576 18889 4604
rect 18288 4564 18294 4576
rect 18877 4573 18889 4576
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 19242 4564 19248 4616
rect 19300 4564 19306 4616
rect 19610 4564 19616 4616
rect 19668 4564 19674 4616
rect 20073 4607 20131 4613
rect 20073 4573 20085 4607
rect 20119 4573 20131 4607
rect 20073 4567 20131 4573
rect 17184 4508 17724 4536
rect 17184 4496 17190 4508
rect 17770 4496 17776 4548
rect 17828 4536 17834 4548
rect 17957 4539 18015 4545
rect 17957 4536 17969 4539
rect 17828 4508 17969 4536
rect 17828 4496 17834 4508
rect 17957 4505 17969 4508
rect 18003 4505 18015 4539
rect 19058 4536 19064 4548
rect 17957 4499 18015 4505
rect 18708 4508 19064 4536
rect 16482 4468 16488 4480
rect 14566 4440 16488 4468
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 16758 4428 16764 4480
rect 16816 4428 16822 4480
rect 17034 4428 17040 4480
rect 17092 4428 17098 4480
rect 17218 4428 17224 4480
rect 17276 4468 17282 4480
rect 18708 4468 18736 4508
rect 19058 4496 19064 4508
rect 19116 4496 19122 4548
rect 19426 4496 19432 4548
rect 19484 4536 19490 4548
rect 20088 4536 20116 4567
rect 19484 4508 20116 4536
rect 19484 4496 19490 4508
rect 17276 4440 18736 4468
rect 17276 4428 17282 4440
rect 18782 4428 18788 4480
rect 18840 4468 18846 4480
rect 21450 4468 21456 4480
rect 18840 4440 21456 4468
rect 18840 4428 18846 4440
rect 21450 4428 21456 4440
rect 21508 4428 21514 4480
rect 1104 4378 21043 4400
rect 1104 4326 5894 4378
rect 5946 4326 5958 4378
rect 6010 4326 6022 4378
rect 6074 4326 6086 4378
rect 6138 4326 6150 4378
rect 6202 4326 10839 4378
rect 10891 4326 10903 4378
rect 10955 4326 10967 4378
rect 11019 4326 11031 4378
rect 11083 4326 11095 4378
rect 11147 4326 15784 4378
rect 15836 4326 15848 4378
rect 15900 4326 15912 4378
rect 15964 4326 15976 4378
rect 16028 4326 16040 4378
rect 16092 4326 20729 4378
rect 20781 4326 20793 4378
rect 20845 4326 20857 4378
rect 20909 4326 20921 4378
rect 20973 4326 20985 4378
rect 21037 4326 21043 4378
rect 1104 4304 21043 4326
rect 1780 4236 4384 4264
rect 1780 4205 1808 4236
rect 1765 4199 1823 4205
rect 1765 4165 1777 4199
rect 1811 4165 1823 4199
rect 4356 4196 4384 4236
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 5629 4267 5687 4273
rect 5629 4264 5641 4267
rect 5408 4236 5641 4264
rect 5408 4224 5414 4236
rect 5629 4233 5641 4236
rect 5675 4233 5687 4267
rect 5629 4227 5687 4233
rect 9585 4267 9643 4273
rect 9585 4233 9597 4267
rect 9631 4264 9643 4267
rect 10226 4264 10232 4276
rect 9631 4236 10232 4264
rect 9631 4233 9643 4236
rect 9585 4227 9643 4233
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 10410 4224 10416 4276
rect 10468 4264 10474 4276
rect 10505 4267 10563 4273
rect 10505 4264 10517 4267
rect 10468 4236 10517 4264
rect 10468 4224 10474 4236
rect 10505 4233 10517 4236
rect 10551 4233 10563 4267
rect 10505 4227 10563 4233
rect 10594 4224 10600 4276
rect 10652 4224 10658 4276
rect 10873 4267 10931 4273
rect 10873 4233 10885 4267
rect 10919 4264 10931 4267
rect 11146 4264 11152 4276
rect 10919 4236 11152 4264
rect 10919 4233 10931 4236
rect 10873 4227 10931 4233
rect 11146 4224 11152 4236
rect 11204 4224 11210 4276
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 11756 4236 12173 4264
rect 11756 4224 11762 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 12437 4267 12495 4273
rect 12437 4233 12449 4267
rect 12483 4264 12495 4267
rect 13354 4264 13360 4276
rect 12483 4236 13360 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 13354 4224 13360 4236
rect 13412 4224 13418 4276
rect 13449 4267 13507 4273
rect 13449 4233 13461 4267
rect 13495 4264 13507 4267
rect 13722 4264 13728 4276
rect 13495 4236 13728 4264
rect 13495 4233 13507 4236
rect 13449 4227 13507 4233
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 13909 4267 13967 4273
rect 13909 4233 13921 4267
rect 13955 4264 13967 4267
rect 14090 4264 14096 4276
rect 13955 4236 14096 4264
rect 13955 4233 13967 4236
rect 13909 4227 13967 4233
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 14300 4236 15792 4264
rect 5810 4196 5816 4208
rect 4356 4168 5816 4196
rect 1765 4159 1823 4165
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 7282 4156 7288 4208
rect 7340 4196 7346 4208
rect 10134 4196 10140 4208
rect 7340 4168 10140 4196
rect 7340 4156 7346 4168
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 10244 4196 10272 4224
rect 10612 4196 10640 4224
rect 13538 4196 13544 4208
rect 10244 4168 10364 4196
rect 10612 4168 10824 4196
rect 1581 4131 1639 4137
rect 1581 4097 1593 4131
rect 1627 4128 1639 4131
rect 1627 4100 2452 4128
rect 1627 4097 1639 4100
rect 1581 4091 1639 4097
rect 2314 4020 2320 4072
rect 2372 4020 2378 4072
rect 2424 4060 2452 4100
rect 2498 4088 2504 4140
rect 2556 4088 2562 4140
rect 3418 4137 3424 4140
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3375 4131 3424 4137
rect 3375 4097 3387 4131
rect 3421 4097 3424 4131
rect 3375 4091 3424 4097
rect 2682 4060 2688 4072
rect 2424 4032 2688 4060
rect 2682 4020 2688 4032
rect 2740 4020 2746 4072
rect 2866 4020 2872 4072
rect 2924 4060 2930 4072
rect 3252 4060 3280 4091
rect 3418 4088 3424 4091
rect 3476 4088 3482 4140
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4128 4215 4131
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4203 4100 4445 4128
rect 4203 4097 4215 4100
rect 4157 4091 4215 4097
rect 4433 4097 4445 4100
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 4891 4131 4949 4137
rect 4891 4097 4903 4131
rect 4937 4128 4949 4131
rect 8754 4128 8760 4140
rect 4937 4100 8760 4128
rect 4937 4097 4949 4100
rect 4891 4091 4949 4097
rect 2924 4032 3280 4060
rect 3513 4063 3571 4069
rect 2924 4020 2930 4032
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 3878 4060 3884 4072
rect 3559 4032 3884 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 1397 3995 1455 4001
rect 1397 3961 1409 3995
rect 1443 3992 1455 3995
rect 2222 3992 2228 4004
rect 1443 3964 2228 3992
rect 1443 3961 1455 3964
rect 1397 3955 1455 3961
rect 2222 3952 2228 3964
rect 2280 3952 2286 4004
rect 2774 3952 2780 4004
rect 2832 3952 2838 4004
rect 2958 3952 2964 4004
rect 3016 3952 3022 4004
rect 4126 3964 4292 3992
rect 1854 3884 1860 3936
rect 1912 3884 1918 3936
rect 2792 3924 2820 3952
rect 4126 3924 4154 3964
rect 4264 3933 4292 3964
rect 2792 3896 4154 3924
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3893 4307 3927
rect 4632 3924 4660 4091
rect 8754 4088 8760 4100
rect 8812 4088 8818 4140
rect 10226 4088 10232 4140
rect 10284 4088 10290 4140
rect 10336 4137 10364 4168
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 10594 4088 10600 4140
rect 10652 4088 10658 4140
rect 10796 4137 10824 4168
rect 10980 4168 13544 4196
rect 10781 4131 10839 4137
rect 10781 4097 10793 4131
rect 10827 4097 10839 4131
rect 10781 4091 10839 4097
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 7466 4060 7472 4072
rect 5868 4032 7472 4060
rect 5868 4020 5874 4032
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 9953 4063 10011 4069
rect 9953 4029 9965 4063
rect 9999 4060 10011 4063
rect 10980 4060 11008 4168
rect 11057 4131 11115 4137
rect 11057 4097 11069 4131
rect 11103 4097 11115 4131
rect 11057 4091 11115 4097
rect 9999 4032 11008 4060
rect 11072 4060 11100 4091
rect 11330 4088 11336 4140
rect 11388 4088 11394 4140
rect 11514 4088 11520 4140
rect 11572 4128 11578 4140
rect 11609 4131 11667 4137
rect 11609 4128 11621 4131
rect 11572 4100 11621 4128
rect 11572 4088 11578 4100
rect 11609 4097 11621 4100
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 11698 4088 11704 4140
rect 11756 4128 11762 4140
rect 11756 4100 11986 4128
rect 11756 4088 11762 4100
rect 11958 4060 11986 4100
rect 12066 4088 12072 4140
rect 12124 4088 12130 4140
rect 12342 4088 12348 4140
rect 12400 4088 12406 4140
rect 12636 4137 12664 4168
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 13814 4196 13820 4208
rect 13648 4168 13820 4196
rect 12621 4131 12679 4137
rect 12621 4097 12633 4131
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 12713 4131 12771 4137
rect 12713 4097 12725 4131
rect 12759 4097 12771 4131
rect 12713 4091 12771 4097
rect 12897 4131 12955 4137
rect 12897 4097 12909 4131
rect 12943 4097 12955 4131
rect 12897 4091 12955 4097
rect 12526 4060 12532 4072
rect 11072 4032 11928 4060
rect 11958 4032 12532 4060
rect 9999 4029 10011 4032
rect 9953 4023 10011 4029
rect 10594 3952 10600 4004
rect 10652 3992 10658 4004
rect 11790 3992 11796 4004
rect 10652 3964 11796 3992
rect 10652 3952 10658 3964
rect 11790 3952 11796 3964
rect 11848 3952 11854 4004
rect 11900 3992 11928 4032
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 11900 3964 12002 3992
rect 5074 3924 5080 3936
rect 4632 3896 5080 3924
rect 4249 3887 4307 3893
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 6730 3924 6736 3936
rect 5684 3896 6736 3924
rect 5684 3884 5690 3896
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 8849 3927 8907 3933
rect 8849 3893 8861 3927
rect 8895 3924 8907 3927
rect 9030 3924 9036 3936
rect 8895 3896 9036 3924
rect 8895 3893 8907 3896
rect 8849 3887 8907 3893
rect 9030 3884 9036 3896
rect 9088 3884 9094 3936
rect 9214 3884 9220 3936
rect 9272 3884 9278 3936
rect 10042 3884 10048 3936
rect 10100 3884 10106 3936
rect 10686 3884 10692 3936
rect 10744 3884 10750 3936
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11330 3924 11336 3936
rect 11195 3896 11336 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11330 3884 11336 3896
rect 11388 3884 11394 3936
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 11701 3927 11759 3933
rect 11701 3924 11713 3927
rect 11664 3896 11713 3924
rect 11664 3884 11670 3896
rect 11701 3893 11713 3896
rect 11747 3893 11759 3927
rect 11701 3887 11759 3893
rect 11882 3884 11888 3936
rect 11940 3884 11946 3936
rect 11974 3924 12002 3964
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 12728 3992 12756 4091
rect 12912 4060 12940 4091
rect 13078 4088 13084 4140
rect 13136 4088 13142 4140
rect 13648 4137 13676 4168
rect 13814 4156 13820 4168
rect 13872 4156 13878 4208
rect 14300 4196 14328 4236
rect 13932 4168 14328 4196
rect 14360 4199 14418 4205
rect 13173 4131 13231 4137
rect 13173 4097 13185 4131
rect 13219 4128 13231 4131
rect 13633 4131 13691 4137
rect 13219 4100 13584 4128
rect 13219 4097 13231 4100
rect 13173 4091 13231 4097
rect 12986 4060 12992 4072
rect 12912 4032 12992 4060
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13096 4060 13124 4088
rect 13354 4060 13360 4072
rect 13096 4032 13360 4060
rect 13354 4020 13360 4032
rect 13412 4020 13418 4072
rect 12400 3964 12756 3992
rect 12805 3995 12863 4001
rect 12400 3952 12406 3964
rect 12805 3961 12817 3995
rect 12851 3992 12863 3995
rect 13170 3992 13176 4004
rect 12851 3964 13176 3992
rect 12851 3961 12863 3964
rect 12805 3955 12863 3961
rect 13170 3952 13176 3964
rect 13228 3952 13234 4004
rect 13556 3992 13584 4100
rect 13633 4097 13645 4131
rect 13679 4097 13691 4131
rect 13633 4091 13691 4097
rect 13725 4131 13783 4137
rect 13725 4097 13737 4131
rect 13771 4128 13783 4131
rect 13932 4128 13960 4168
rect 14360 4165 14372 4199
rect 14406 4196 14418 4199
rect 14826 4196 14832 4208
rect 14406 4168 14832 4196
rect 14406 4165 14418 4168
rect 14360 4159 14418 4165
rect 14826 4156 14832 4168
rect 14884 4156 14890 4208
rect 14918 4156 14924 4208
rect 14976 4196 14982 4208
rect 15654 4196 15660 4208
rect 14976 4168 15660 4196
rect 14976 4156 14982 4168
rect 15654 4156 15660 4168
rect 15712 4156 15718 4208
rect 15764 4196 15792 4236
rect 15838 4224 15844 4276
rect 15896 4264 15902 4276
rect 15896 4236 16344 4264
rect 15896 4224 15902 4236
rect 16316 4205 16344 4236
rect 16390 4224 16396 4276
rect 16448 4264 16454 4276
rect 17218 4264 17224 4276
rect 16448 4236 17224 4264
rect 16448 4224 16454 4236
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 19150 4264 19156 4276
rect 17328 4236 19156 4264
rect 16301 4199 16359 4205
rect 15764 4168 16252 4196
rect 15749 4131 15807 4137
rect 15749 4128 15761 4131
rect 13771 4100 13960 4128
rect 14016 4100 15761 4128
rect 13771 4097 13783 4100
rect 13725 4091 13783 4097
rect 13814 4020 13820 4072
rect 13872 4060 13878 4072
rect 14016 4060 14044 4100
rect 15749 4097 15761 4100
rect 15795 4097 15807 4131
rect 15749 4091 15807 4097
rect 16114 4088 16120 4140
rect 16172 4088 16178 4140
rect 16224 4128 16252 4168
rect 16301 4165 16313 4199
rect 16347 4165 16359 4199
rect 16301 4159 16359 4165
rect 16850 4156 16856 4208
rect 16908 4156 16914 4208
rect 17328 4196 17356 4236
rect 19150 4224 19156 4236
rect 19208 4224 19214 4276
rect 19886 4224 19892 4276
rect 19944 4224 19950 4276
rect 20438 4224 20444 4276
rect 20496 4224 20502 4276
rect 17052 4168 17356 4196
rect 16390 4128 16396 4140
rect 16224 4100 16396 4128
rect 16390 4088 16396 4100
rect 16448 4088 16454 4140
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 17052 4128 17080 4168
rect 17494 4156 17500 4208
rect 17552 4196 17558 4208
rect 18874 4196 18880 4208
rect 17552 4168 18184 4196
rect 17552 4156 17558 4168
rect 16531 4100 17080 4128
rect 17129 4131 17187 4137
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 17129 4097 17141 4131
rect 17175 4128 17187 4131
rect 17310 4128 17316 4140
rect 17175 4100 17316 4128
rect 17175 4097 17187 4100
rect 17129 4091 17187 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 17402 4088 17408 4140
rect 17460 4088 17466 4140
rect 13872 4032 14044 4060
rect 14093 4063 14151 4069
rect 13872 4020 13878 4032
rect 14093 4029 14105 4063
rect 14139 4029 14151 4063
rect 14093 4023 14151 4029
rect 13906 3992 13912 4004
rect 13556 3964 13912 3992
rect 13906 3952 13912 3964
rect 13964 3952 13970 4004
rect 13998 3952 14004 4004
rect 14056 3952 14062 4004
rect 13357 3927 13415 3933
rect 13357 3924 13369 3927
rect 11974 3896 13369 3924
rect 13357 3893 13369 3896
rect 13403 3924 13415 3927
rect 14016 3924 14044 3952
rect 13403 3896 14044 3924
rect 14108 3924 14136 4023
rect 15654 4020 15660 4072
rect 15712 4060 15718 4072
rect 16022 4060 16028 4072
rect 15712 4032 16028 4060
rect 15712 4020 15718 4032
rect 16022 4020 16028 4032
rect 16080 4020 16086 4072
rect 15473 3995 15531 4001
rect 15473 3961 15485 3995
rect 15519 3992 15531 3995
rect 16132 3992 16160 4088
rect 18156 4072 18184 4168
rect 18524 4168 18880 4196
rect 18524 4137 18552 4168
rect 18874 4156 18880 4168
rect 18932 4156 18938 4208
rect 19058 4156 19064 4208
rect 19116 4156 19122 4208
rect 19306 4168 20392 4196
rect 18509 4131 18567 4137
rect 18509 4097 18521 4131
rect 18555 4097 18567 4131
rect 18509 4091 18567 4097
rect 18598 4088 18604 4140
rect 18656 4128 18662 4140
rect 18765 4131 18823 4137
rect 18765 4128 18777 4131
rect 18656 4100 18777 4128
rect 18656 4088 18662 4100
rect 18765 4097 18777 4100
rect 18811 4097 18823 4131
rect 19076 4128 19104 4156
rect 19306 4128 19334 4168
rect 19076 4100 19334 4128
rect 18765 4091 18823 4097
rect 19702 4088 19708 4140
rect 19760 4128 19766 4140
rect 20364 4137 20392 4168
rect 20073 4131 20131 4137
rect 20073 4128 20085 4131
rect 19760 4100 20085 4128
rect 19760 4088 19766 4100
rect 20073 4097 20085 4100
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 20349 4131 20407 4137
rect 20349 4097 20361 4131
rect 20395 4097 20407 4131
rect 20349 4091 20407 4097
rect 17954 4020 17960 4072
rect 18012 4020 18018 4072
rect 18138 4020 18144 4072
rect 18196 4020 18202 4072
rect 20257 4063 20315 4069
rect 20257 4029 20269 4063
rect 20303 4060 20315 4063
rect 21174 4060 21180 4072
rect 20303 4032 21180 4060
rect 20303 4029 20315 4032
rect 20257 4023 20315 4029
rect 21174 4020 21180 4032
rect 21232 4020 21238 4072
rect 15519 3964 16160 3992
rect 17972 3992 18000 4020
rect 17972 3964 18552 3992
rect 15519 3961 15531 3964
rect 15473 3955 15531 3961
rect 14458 3924 14464 3936
rect 14108 3896 14464 3924
rect 13403 3893 13415 3896
rect 13357 3887 13415 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 15194 3884 15200 3936
rect 15252 3924 15258 3936
rect 15841 3927 15899 3933
rect 15841 3924 15853 3927
rect 15252 3896 15853 3924
rect 15252 3884 15258 3896
rect 15841 3893 15853 3896
rect 15887 3893 15899 3927
rect 15841 3887 15899 3893
rect 16942 3884 16948 3936
rect 17000 3884 17006 3936
rect 17954 3884 17960 3936
rect 18012 3924 18018 3936
rect 18141 3927 18199 3933
rect 18141 3924 18153 3927
rect 18012 3896 18153 3924
rect 18012 3884 18018 3896
rect 18141 3893 18153 3896
rect 18187 3893 18199 3927
rect 18524 3924 18552 3964
rect 19150 3924 19156 3936
rect 18524 3896 19156 3924
rect 18141 3887 18199 3893
rect 19150 3884 19156 3896
rect 19208 3884 19214 3936
rect 1104 3834 20884 3856
rect 1104 3782 3422 3834
rect 3474 3782 3486 3834
rect 3538 3782 3550 3834
rect 3602 3782 3614 3834
rect 3666 3782 3678 3834
rect 3730 3782 8367 3834
rect 8419 3782 8431 3834
rect 8483 3782 8495 3834
rect 8547 3782 8559 3834
rect 8611 3782 8623 3834
rect 8675 3782 13312 3834
rect 13364 3782 13376 3834
rect 13428 3782 13440 3834
rect 13492 3782 13504 3834
rect 13556 3782 13568 3834
rect 13620 3782 18257 3834
rect 18309 3782 18321 3834
rect 18373 3782 18385 3834
rect 18437 3782 18449 3834
rect 18501 3782 18513 3834
rect 18565 3782 20884 3834
rect 1104 3760 20884 3782
rect 2590 3680 2596 3732
rect 2648 3680 2654 3732
rect 3142 3680 3148 3732
rect 3200 3680 3206 3732
rect 3970 3680 3976 3732
rect 4028 3680 4034 3732
rect 4338 3680 4344 3732
rect 4396 3680 4402 3732
rect 4430 3680 4436 3732
rect 4488 3720 4494 3732
rect 4617 3723 4675 3729
rect 4617 3720 4629 3723
rect 4488 3692 4629 3720
rect 4488 3680 4494 3692
rect 4617 3689 4629 3692
rect 4663 3689 4675 3723
rect 4617 3683 4675 3689
rect 6362 3680 6368 3732
rect 6420 3720 6426 3732
rect 7469 3723 7527 3729
rect 7469 3720 7481 3723
rect 6420 3692 7481 3720
rect 6420 3680 6426 3692
rect 7469 3689 7481 3692
rect 7515 3689 7527 3723
rect 7469 3683 7527 3689
rect 7742 3680 7748 3732
rect 7800 3680 7806 3732
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 8297 3723 8355 3729
rect 8297 3720 8309 3723
rect 7892 3692 8309 3720
rect 7892 3680 7898 3692
rect 8297 3689 8309 3692
rect 8343 3689 8355 3723
rect 8297 3683 8355 3689
rect 8941 3723 8999 3729
rect 8941 3689 8953 3723
rect 8987 3720 8999 3723
rect 9766 3720 9772 3732
rect 8987 3692 9772 3720
rect 8987 3689 8999 3692
rect 8941 3683 8999 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 9858 3680 9864 3732
rect 9916 3680 9922 3732
rect 10778 3680 10784 3732
rect 10836 3680 10842 3732
rect 11241 3723 11299 3729
rect 11241 3689 11253 3723
rect 11287 3720 11299 3723
rect 11422 3720 11428 3732
rect 11287 3692 11428 3720
rect 11287 3689 11299 3692
rect 11241 3683 11299 3689
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 11514 3680 11520 3732
rect 11572 3680 11578 3732
rect 12069 3723 12127 3729
rect 12069 3689 12081 3723
rect 12115 3720 12127 3723
rect 12250 3720 12256 3732
rect 12115 3692 12256 3720
rect 12115 3689 12127 3692
rect 12069 3683 12127 3689
rect 12250 3680 12256 3692
rect 12308 3680 12314 3732
rect 18690 3720 18696 3732
rect 12452 3692 13860 3720
rect 5442 3652 5448 3664
rect 4126 3624 5448 3652
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 1762 3516 1768 3528
rect 1627 3488 1768 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 1762 3476 1768 3488
rect 1820 3476 1826 3528
rect 1855 3519 1913 3525
rect 1855 3485 1867 3519
rect 1901 3516 1913 3519
rect 4126 3516 4154 3624
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 6549 3655 6607 3661
rect 6549 3621 6561 3655
rect 6595 3652 6607 3655
rect 7190 3652 7196 3664
rect 6595 3624 7196 3652
rect 6595 3621 6607 3624
rect 6549 3615 6607 3621
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 7760 3584 7788 3680
rect 4724 3556 7788 3584
rect 9876 3584 9904 3680
rect 10321 3655 10379 3661
rect 10321 3621 10333 3655
rect 10367 3652 10379 3655
rect 11146 3652 11152 3664
rect 10367 3624 11152 3652
rect 10367 3621 10379 3624
rect 10321 3615 10379 3621
rect 11146 3612 11152 3624
rect 11204 3612 11210 3664
rect 9876 3556 10180 3584
rect 1901 3488 4154 3516
rect 1901 3485 1913 3488
rect 1855 3479 1913 3485
rect 4522 3476 4528 3528
rect 4580 3476 4586 3528
rect 3053 3451 3111 3457
rect 3053 3417 3065 3451
rect 3099 3448 3111 3451
rect 3326 3448 3332 3460
rect 3099 3420 3332 3448
rect 3099 3417 3111 3420
rect 3053 3411 3111 3417
rect 3326 3408 3332 3420
rect 3384 3408 3390 3460
rect 3881 3451 3939 3457
rect 3881 3417 3893 3451
rect 3927 3448 3939 3451
rect 3970 3448 3976 3460
rect 3927 3420 3976 3448
rect 3927 3417 3939 3420
rect 3881 3411 3939 3417
rect 3970 3408 3976 3420
rect 4028 3408 4034 3460
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 4724 3380 4752 3556
rect 4801 3519 4859 3525
rect 4801 3485 4813 3519
rect 4847 3516 4859 3519
rect 5718 3516 5724 3528
rect 4847 3488 5724 3516
rect 4847 3485 4859 3488
rect 4801 3479 4859 3485
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 6730 3476 6736 3528
rect 6788 3476 6794 3528
rect 7006 3476 7012 3528
rect 7064 3476 7070 3528
rect 7098 3476 7104 3528
rect 7156 3516 7162 3528
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7156 3488 7297 3516
rect 7156 3476 7162 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 9122 3476 9128 3528
rect 9180 3476 9186 3528
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9493 3519 9551 3525
rect 9493 3516 9505 3519
rect 9456 3488 9505 3516
rect 9456 3476 9462 3488
rect 9493 3485 9505 3488
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 9858 3476 9864 3528
rect 9916 3476 9922 3528
rect 10152 3525 10180 3556
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 11532 3584 11560 3680
rect 12452 3664 12480 3692
rect 13832 3664 13860 3692
rect 13932 3692 18696 3720
rect 11701 3655 11759 3661
rect 11701 3621 11713 3655
rect 11747 3621 11759 3655
rect 11701 3615 11759 3621
rect 11793 3655 11851 3661
rect 11793 3621 11805 3655
rect 11839 3652 11851 3655
rect 12158 3652 12164 3664
rect 11839 3624 12164 3652
rect 11839 3621 11851 3624
rect 11793 3615 11851 3621
rect 11112 3556 11192 3584
rect 11112 3544 11118 3556
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3485 10103 3519
rect 10045 3479 10103 3485
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3485 10195 3519
rect 10137 3479 10195 3485
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 8757 3451 8815 3457
rect 5500 3420 7144 3448
rect 5500 3408 5506 3420
rect 1728 3352 4752 3380
rect 1728 3340 1734 3352
rect 5350 3340 5356 3392
rect 5408 3380 5414 3392
rect 6270 3380 6276 3392
rect 5408 3352 6276 3380
rect 5408 3340 5414 3352
rect 6270 3340 6276 3352
rect 6328 3340 6334 3392
rect 6822 3340 6828 3392
rect 6880 3340 6886 3392
rect 7116 3389 7144 3420
rect 8757 3417 8769 3451
rect 8803 3448 8815 3451
rect 10060 3448 10088 3479
rect 10594 3476 10600 3528
rect 10652 3476 10658 3528
rect 11164 3525 11192 3556
rect 11256 3556 11560 3584
rect 11716 3584 11744 3615
rect 12158 3612 12164 3624
rect 12216 3612 12222 3664
rect 12434 3612 12440 3664
rect 12492 3612 12498 3664
rect 12621 3655 12679 3661
rect 12621 3621 12633 3655
rect 12667 3652 12679 3655
rect 12894 3652 12900 3664
rect 12667 3624 12900 3652
rect 12667 3621 12679 3624
rect 12621 3615 12679 3621
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 13814 3612 13820 3664
rect 13872 3612 13878 3664
rect 11716 3556 12646 3584
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3485 11207 3519
rect 11149 3479 11207 3485
rect 8803 3420 9444 3448
rect 10060 3420 10640 3448
rect 8803 3417 8815 3420
rect 8757 3411 8815 3417
rect 9416 3392 9444 3420
rect 10612 3392 10640 3420
rect 7101 3383 7159 3389
rect 7101 3349 7113 3383
rect 7147 3349 7159 3383
rect 7101 3343 7159 3349
rect 7742 3340 7748 3392
rect 7800 3340 7806 3392
rect 9306 3340 9312 3392
rect 9364 3340 9370 3392
rect 9398 3340 9404 3392
rect 9456 3340 9462 3392
rect 10045 3383 10103 3389
rect 10045 3349 10057 3383
rect 10091 3380 10103 3383
rect 10318 3380 10324 3392
rect 10091 3352 10324 3380
rect 10091 3349 10103 3352
rect 10045 3343 10103 3349
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 10594 3340 10600 3392
rect 10652 3340 10658 3392
rect 10965 3383 11023 3389
rect 10965 3349 10977 3383
rect 11011 3380 11023 3383
rect 11256 3380 11284 3556
rect 11425 3519 11483 3525
rect 11425 3485 11437 3519
rect 11471 3485 11483 3519
rect 11425 3479 11483 3485
rect 11517 3519 11575 3525
rect 11517 3485 11529 3519
rect 11563 3516 11575 3519
rect 11790 3516 11796 3528
rect 11563 3488 11796 3516
rect 11563 3485 11575 3488
rect 11517 3479 11575 3485
rect 11440 3448 11468 3479
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 11974 3476 11980 3528
rect 12032 3476 12038 3528
rect 12250 3476 12256 3528
rect 12308 3476 12314 3528
rect 12526 3476 12532 3528
rect 12584 3476 12590 3528
rect 12618 3448 12646 3556
rect 12710 3544 12716 3596
rect 12768 3584 12774 3596
rect 13932 3584 13960 3692
rect 18690 3680 18696 3692
rect 18748 3680 18754 3732
rect 19334 3680 19340 3732
rect 19392 3680 19398 3732
rect 14090 3612 14096 3664
rect 14148 3612 14154 3664
rect 14918 3612 14924 3664
rect 14976 3652 14982 3664
rect 15378 3652 15384 3664
rect 14976 3624 15384 3652
rect 14976 3612 14982 3624
rect 15378 3612 15384 3624
rect 15436 3612 15442 3664
rect 15473 3655 15531 3661
rect 15473 3621 15485 3655
rect 15519 3652 15531 3655
rect 16206 3652 16212 3664
rect 15519 3624 16212 3652
rect 15519 3621 15531 3624
rect 15473 3615 15531 3621
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 17218 3612 17224 3664
rect 17276 3652 17282 3664
rect 17405 3655 17463 3661
rect 17405 3652 17417 3655
rect 17276 3624 17417 3652
rect 17276 3612 17282 3624
rect 17405 3621 17417 3624
rect 17451 3621 17463 3655
rect 17405 3615 17463 3621
rect 12768 3556 12848 3584
rect 12768 3544 12774 3556
rect 12820 3525 12848 3556
rect 13464 3556 13960 3584
rect 13464 3525 13492 3556
rect 12805 3519 12863 3525
rect 12805 3485 12817 3519
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 13081 3519 13139 3525
rect 13081 3485 13093 3519
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13449 3519 13507 3525
rect 13449 3485 13461 3519
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 13725 3519 13783 3525
rect 13725 3485 13737 3519
rect 13771 3516 13783 3519
rect 13814 3516 13820 3528
rect 13771 3488 13820 3516
rect 13771 3485 13783 3488
rect 13725 3479 13783 3485
rect 13096 3448 13124 3479
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 14108 3525 14136 3612
rect 14826 3544 14832 3596
rect 14884 3584 14890 3596
rect 15194 3584 15200 3596
rect 14884 3556 15200 3584
rect 14884 3544 14890 3556
rect 15194 3544 15200 3556
rect 15252 3544 15258 3596
rect 17420 3584 17448 3615
rect 18138 3612 18144 3664
rect 18196 3652 18202 3664
rect 19352 3652 19380 3680
rect 18196 3624 19380 3652
rect 18196 3612 18202 3624
rect 17865 3587 17923 3593
rect 17865 3584 17877 3587
rect 15746 3556 16344 3584
rect 17420 3556 17877 3584
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 14367 3519 14425 3525
rect 14367 3485 14379 3519
rect 14413 3516 14425 3519
rect 15513 3516 15611 3518
rect 14413 3490 15611 3516
rect 14413 3488 15541 3490
rect 14413 3485 14425 3488
rect 14367 3479 14425 3485
rect 14826 3448 14832 3460
rect 11440 3420 12572 3448
rect 12618 3420 14832 3448
rect 11011 3352 11284 3380
rect 11011 3349 11023 3352
rect 10965 3343 11023 3349
rect 12250 3340 12256 3392
rect 12308 3380 12314 3392
rect 12345 3383 12403 3389
rect 12345 3380 12357 3383
rect 12308 3352 12357 3380
rect 12308 3340 12314 3352
rect 12345 3349 12357 3352
rect 12391 3349 12403 3383
rect 12544 3380 12572 3420
rect 14826 3408 14832 3420
rect 14884 3408 14890 3460
rect 15583 3448 15611 3490
rect 15654 3476 15660 3528
rect 15712 3476 15718 3528
rect 15746 3448 15774 3556
rect 16316 3528 16344 3556
rect 17865 3553 17877 3556
rect 17911 3553 17923 3587
rect 19337 3587 19395 3593
rect 19337 3584 19349 3587
rect 17865 3547 17923 3553
rect 17972 3556 19349 3584
rect 17972 3528 18000 3556
rect 19337 3553 19349 3556
rect 19383 3553 19395 3587
rect 19337 3547 19395 3553
rect 20162 3544 20168 3596
rect 20220 3544 20226 3596
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 15933 3519 15991 3525
rect 15933 3516 15945 3519
rect 15896 3488 15945 3516
rect 15896 3476 15902 3488
rect 15933 3485 15945 3488
rect 15979 3485 15991 3519
rect 15933 3479 15991 3485
rect 16298 3476 16304 3528
rect 16356 3476 16362 3528
rect 16393 3519 16451 3525
rect 16393 3485 16405 3519
rect 16439 3485 16451 3519
rect 16393 3479 16451 3485
rect 16667 3519 16725 3525
rect 16667 3485 16679 3519
rect 16713 3516 16725 3519
rect 16713 3488 17908 3516
rect 16713 3485 16725 3488
rect 16667 3479 16725 3485
rect 16408 3448 16436 3479
rect 16850 3448 16856 3460
rect 15038 3420 15541 3448
rect 15583 3420 15774 3448
rect 15948 3420 16344 3448
rect 16408 3420 16856 3448
rect 12618 3380 12624 3392
rect 12544 3352 12624 3380
rect 12345 3343 12403 3349
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 12897 3383 12955 3389
rect 12897 3380 12909 3383
rect 12860 3352 12909 3380
rect 12860 3340 12866 3352
rect 12897 3349 12909 3352
rect 12943 3349 12955 3383
rect 12897 3343 12955 3349
rect 12986 3340 12992 3392
rect 13044 3380 13050 3392
rect 13265 3383 13323 3389
rect 13265 3380 13277 3383
rect 13044 3352 13277 3380
rect 13044 3340 13050 3352
rect 13265 3349 13277 3352
rect 13311 3349 13323 3383
rect 13265 3343 13323 3349
rect 13352 3340 13358 3392
rect 13410 3380 13416 3392
rect 13541 3383 13599 3389
rect 13541 3380 13553 3383
rect 13410 3352 13553 3380
rect 13410 3340 13416 3352
rect 13541 3349 13553 3352
rect 13587 3349 13599 3383
rect 13541 3343 13599 3349
rect 13630 3340 13636 3392
rect 13688 3380 13694 3392
rect 15038 3380 15066 3420
rect 13688 3352 15066 3380
rect 15105 3383 15163 3389
rect 13688 3340 13694 3352
rect 15105 3349 15117 3383
rect 15151 3380 15163 3383
rect 15378 3380 15384 3392
rect 15151 3352 15384 3380
rect 15151 3349 15163 3352
rect 15105 3343 15163 3349
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 15513 3380 15541 3420
rect 15948 3380 15976 3420
rect 15513 3352 15976 3380
rect 16025 3383 16083 3389
rect 16025 3349 16037 3383
rect 16071 3380 16083 3383
rect 16114 3380 16120 3392
rect 16071 3352 16120 3380
rect 16071 3349 16083 3352
rect 16025 3343 16083 3349
rect 16114 3340 16120 3352
rect 16172 3340 16178 3392
rect 16316 3380 16344 3420
rect 16850 3408 16856 3420
rect 16908 3448 16914 3460
rect 17310 3448 17316 3460
rect 16908 3420 17316 3448
rect 16908 3408 16914 3420
rect 17310 3408 17316 3420
rect 17368 3408 17374 3460
rect 17880 3448 17908 3488
rect 17954 3476 17960 3528
rect 18012 3476 18018 3528
rect 18138 3476 18144 3528
rect 18196 3476 18202 3528
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18380 3488 18613 3516
rect 18380 3476 18386 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3516 18935 3519
rect 19058 3516 19064 3528
rect 18923 3488 19064 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 19058 3476 19064 3488
rect 19116 3476 19122 3528
rect 19610 3476 19616 3528
rect 19668 3476 19674 3528
rect 20070 3476 20076 3528
rect 20128 3476 20134 3528
rect 18966 3448 18972 3460
rect 17880 3420 18972 3448
rect 18966 3408 18972 3420
rect 19024 3408 19030 3460
rect 21266 3380 21272 3392
rect 16316 3352 21272 3380
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 1104 3290 21043 3312
rect 1104 3238 5894 3290
rect 5946 3238 5958 3290
rect 6010 3238 6022 3290
rect 6074 3238 6086 3290
rect 6138 3238 6150 3290
rect 6202 3238 10839 3290
rect 10891 3238 10903 3290
rect 10955 3238 10967 3290
rect 11019 3238 11031 3290
rect 11083 3238 11095 3290
rect 11147 3238 15784 3290
rect 15836 3238 15848 3290
rect 15900 3238 15912 3290
rect 15964 3238 15976 3290
rect 16028 3238 16040 3290
rect 16092 3238 20729 3290
rect 20781 3238 20793 3290
rect 20845 3238 20857 3290
rect 20909 3238 20921 3290
rect 20973 3238 20985 3290
rect 21037 3238 21043 3290
rect 1104 3216 21043 3238
rect 1578 3136 1584 3188
rect 1636 3136 1642 3188
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3176 2375 3179
rect 3050 3176 3056 3188
rect 2363 3148 3056 3176
rect 2363 3145 2375 3148
rect 2317 3139 2375 3145
rect 3050 3136 3056 3148
rect 3108 3136 3114 3188
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 3878 3176 3884 3188
rect 3743 3148 3884 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4154 3136 4160 3188
rect 4212 3176 4218 3188
rect 4249 3179 4307 3185
rect 4249 3176 4261 3179
rect 4212 3148 4261 3176
rect 4212 3136 4218 3148
rect 4249 3145 4261 3148
rect 4295 3145 4307 3179
rect 4249 3139 4307 3145
rect 5813 3179 5871 3185
rect 5813 3145 5825 3179
rect 5859 3176 5871 3179
rect 7374 3176 7380 3188
rect 5859 3148 7380 3176
rect 5859 3145 5871 3148
rect 5813 3139 5871 3145
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 8294 3136 8300 3188
rect 8352 3176 8358 3188
rect 8352 3148 9536 3176
rect 8352 3136 8358 3148
rect 1489 3111 1547 3117
rect 1489 3077 1501 3111
rect 1535 3108 1547 3111
rect 2774 3108 2780 3120
rect 1535 3080 2780 3108
rect 1535 3077 1547 3080
rect 1489 3071 1547 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 3234 3108 3240 3120
rect 2884 3080 3240 3108
rect 1762 3000 1768 3052
rect 1820 3000 1826 3052
rect 2041 3043 2099 3049
rect 2041 3009 2053 3043
rect 2087 3040 2099 3043
rect 2884 3040 2912 3080
rect 3234 3068 3240 3080
rect 3292 3068 3298 3120
rect 5534 3068 5540 3120
rect 5592 3108 5598 3120
rect 5592 3080 7236 3108
rect 5592 3068 5598 3080
rect 2087 3012 2912 3040
rect 2943 3043 3001 3049
rect 2087 3009 2099 3012
rect 2041 3003 2099 3009
rect 2943 3009 2955 3043
rect 2989 3040 3001 3043
rect 3050 3040 3056 3052
rect 2989 3012 3056 3040
rect 2989 3009 3001 3012
rect 2943 3003 3001 3009
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 5718 3000 5724 3052
rect 5776 3040 5782 3052
rect 5997 3043 6055 3049
rect 5997 3040 6009 3043
rect 5776 3012 6009 3040
rect 5776 3000 5782 3012
rect 5997 3009 6009 3012
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6638 3000 6644 3052
rect 6696 3000 6702 3052
rect 7208 3049 7236 3080
rect 8386 3068 8392 3120
rect 8444 3108 8450 3120
rect 8444 3080 9444 3108
rect 8444 3068 8450 3080
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 7193 3043 7251 3049
rect 7193 3009 7205 3043
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 1780 2972 1808 3000
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 1780 2944 2697 2972
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 2685 2935 2743 2941
rect 4614 2932 4620 2984
rect 4672 2972 4678 2984
rect 5810 2972 5816 2984
rect 4672 2944 5816 2972
rect 4672 2932 4678 2944
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 6932 2972 6960 3003
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 7926 3040 7932 3052
rect 7791 3012 7932 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 8018 3000 8024 3052
rect 8076 3000 8082 3052
rect 8294 3000 8300 3052
rect 8352 3000 8358 3052
rect 8570 3000 8576 3052
rect 8628 3000 8634 3052
rect 8846 3000 8852 3052
rect 8904 3000 8910 3052
rect 9122 3000 9128 3052
rect 9180 3000 9186 3052
rect 9416 3049 9444 3080
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9214 2972 9220 2984
rect 6932 2944 7420 2972
rect 7392 2916 7420 2944
rect 7484 2944 9220 2972
rect 6546 2864 6552 2916
rect 6604 2904 6610 2916
rect 7285 2907 7343 2913
rect 7285 2904 7297 2907
rect 6604 2876 7297 2904
rect 6604 2864 6610 2876
rect 7285 2873 7297 2876
rect 7331 2873 7343 2907
rect 7285 2867 7343 2873
rect 7374 2864 7380 2916
rect 7432 2864 7438 2916
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 3050 2836 3056 2848
rect 716 2808 3056 2836
rect 716 2796 722 2808
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 4890 2796 4896 2848
rect 4948 2836 4954 2848
rect 5626 2836 5632 2848
rect 4948 2808 5632 2836
rect 4948 2796 4954 2808
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 6457 2839 6515 2845
rect 6457 2805 6469 2839
rect 6503 2836 6515 2839
rect 6638 2836 6644 2848
rect 6503 2808 6644 2836
rect 6503 2805 6515 2808
rect 6457 2799 6515 2805
rect 6638 2796 6644 2808
rect 6696 2796 6702 2848
rect 6730 2796 6736 2848
rect 6788 2796 6794 2848
rect 7009 2839 7067 2845
rect 7009 2805 7021 2839
rect 7055 2836 7067 2839
rect 7484 2836 7512 2944
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9508 2972 9536 3148
rect 10962 3136 10968 3188
rect 11020 3176 11026 3188
rect 12437 3179 12495 3185
rect 12437 3176 12449 3179
rect 11020 3148 12449 3176
rect 11020 3136 11026 3148
rect 12437 3145 12449 3148
rect 12483 3145 12495 3179
rect 12437 3139 12495 3145
rect 12710 3136 12716 3188
rect 12768 3136 12774 3188
rect 12802 3136 12808 3188
rect 12860 3136 12866 3188
rect 13354 3136 13360 3188
rect 13412 3136 13418 3188
rect 13449 3179 13507 3185
rect 13449 3145 13461 3179
rect 13495 3176 13507 3179
rect 13495 3148 13860 3176
rect 13495 3145 13507 3148
rect 13449 3139 13507 3145
rect 12728 3108 12756 3136
rect 10336 3080 12570 3108
rect 9674 3000 9680 3052
rect 9732 3000 9738 3052
rect 9950 3000 9956 3052
rect 10008 3000 10014 3052
rect 10045 3043 10103 3049
rect 10045 3009 10057 3043
rect 10091 3040 10103 3043
rect 10226 3040 10232 3052
rect 10091 3012 10232 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 10336 3049 10364 3080
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3009 10379 3043
rect 10321 3003 10379 3009
rect 10778 3000 10784 3052
rect 10836 3000 10842 3052
rect 11054 3000 11060 3052
rect 11112 3000 11118 3052
rect 11146 3000 11152 3052
rect 11204 3000 11210 3052
rect 11698 3000 11704 3052
rect 11756 3000 11762 3052
rect 11793 3027 11851 3033
rect 10410 2972 10416 2984
rect 9508 2944 10416 2972
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 11606 2972 11612 2984
rect 11072 2944 11612 2972
rect 10042 2904 10048 2916
rect 8680 2876 10048 2904
rect 7055 2808 7512 2836
rect 7055 2805 7067 2808
rect 7009 2799 7067 2805
rect 7558 2796 7564 2848
rect 7616 2796 7622 2848
rect 7834 2796 7840 2848
rect 7892 2796 7898 2848
rect 8110 2796 8116 2848
rect 8168 2796 8174 2848
rect 8386 2796 8392 2848
rect 8444 2796 8450 2848
rect 8680 2845 8708 2876
rect 10042 2864 10048 2876
rect 10100 2864 10106 2916
rect 10229 2907 10287 2913
rect 10229 2873 10241 2907
rect 10275 2904 10287 2907
rect 11072 2904 11100 2944
rect 11606 2932 11612 2944
rect 11664 2932 11670 2984
rect 10275 2876 11100 2904
rect 11333 2907 11391 2913
rect 10275 2873 10287 2876
rect 10229 2867 10287 2873
rect 11333 2873 11345 2907
rect 11379 2904 11391 2907
rect 11716 2904 11744 3000
rect 11793 2993 11805 3027
rect 11839 2993 11851 3027
rect 11882 3000 11888 3052
rect 11940 3049 11946 3052
rect 11940 3043 11969 3049
rect 11957 3009 11969 3043
rect 11940 3003 11969 3009
rect 11940 3000 11946 3003
rect 12066 3000 12072 3052
rect 12124 3000 12130 3052
rect 12161 3043 12219 3049
rect 12161 3009 12173 3043
rect 12207 3040 12219 3043
rect 12434 3040 12440 3052
rect 12207 3012 12440 3040
rect 12207 3009 12219 3012
rect 12161 3003 12219 3009
rect 12434 3000 12440 3012
rect 12492 3000 12498 3052
rect 11793 2987 11851 2993
rect 11379 2876 11744 2904
rect 11808 2904 11836 2987
rect 12084 2972 12112 3000
rect 12542 2972 12570 3080
rect 12628 3080 12756 3108
rect 12820 3108 12848 3136
rect 12820 3080 13318 3108
rect 12628 3049 12656 3080
rect 12613 3043 12671 3049
rect 12613 3009 12625 3043
rect 12659 3009 12671 3043
rect 12613 3003 12671 3009
rect 12713 3043 12771 3049
rect 12713 3009 12725 3043
rect 12759 3040 12771 3043
rect 12802 3040 12808 3052
rect 12759 3012 12808 3040
rect 12759 3009 12771 3012
rect 12713 3003 12771 3009
rect 12802 3000 12808 3012
rect 12860 3000 12866 3052
rect 13078 3000 13084 3052
rect 13136 3040 13142 3052
rect 13173 3043 13231 3049
rect 13173 3040 13185 3043
rect 13136 3012 13185 3040
rect 13136 3000 13142 3012
rect 13173 3009 13185 3012
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 13290 2972 13318 3080
rect 13372 3049 13400 3136
rect 13832 3108 13860 3148
rect 13906 3136 13912 3188
rect 13964 3176 13970 3188
rect 14274 3176 14280 3188
rect 13964 3148 14280 3176
rect 13964 3136 13970 3148
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 14366 3136 14372 3188
rect 14424 3136 14430 3188
rect 14642 3136 14648 3188
rect 14700 3176 14706 3188
rect 14700 3148 15056 3176
rect 14700 3136 14706 3148
rect 14382 3108 14410 3136
rect 13464 3080 13768 3108
rect 13832 3080 14410 3108
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3009 13415 3043
rect 13357 3003 13415 3009
rect 13464 2972 13492 3080
rect 13633 3043 13691 3049
rect 13633 3009 13645 3043
rect 13679 3009 13691 3043
rect 13740 3040 13768 3080
rect 14826 3068 14832 3120
rect 14884 3068 14890 3120
rect 15028 3117 15056 3148
rect 15194 3136 15200 3188
rect 15252 3176 15258 3188
rect 16758 3176 16764 3188
rect 15252 3148 16764 3176
rect 15252 3136 15258 3148
rect 16758 3136 16764 3148
rect 16816 3136 16822 3188
rect 16942 3136 16948 3188
rect 17000 3136 17006 3188
rect 17310 3136 17316 3188
rect 17368 3176 17374 3188
rect 17770 3176 17776 3188
rect 17368 3148 17776 3176
rect 17368 3136 17374 3148
rect 17770 3136 17776 3148
rect 17828 3136 17834 3188
rect 18230 3136 18236 3188
rect 18288 3136 18294 3188
rect 18509 3179 18567 3185
rect 18509 3145 18521 3179
rect 18555 3176 18567 3179
rect 18782 3176 18788 3188
rect 18555 3148 18788 3176
rect 18555 3145 18567 3148
rect 18509 3139 18567 3145
rect 18782 3136 18788 3148
rect 18840 3136 18846 3188
rect 20349 3179 20407 3185
rect 20349 3145 20361 3179
rect 20395 3176 20407 3179
rect 21818 3176 21824 3188
rect 20395 3148 21824 3176
rect 20395 3145 20407 3148
rect 20349 3139 20407 3145
rect 21818 3136 21824 3148
rect 21876 3136 21882 3188
rect 15013 3111 15071 3117
rect 15013 3077 15025 3111
rect 15059 3077 15071 3111
rect 15013 3071 15071 3077
rect 15102 3068 15108 3120
rect 15160 3108 15166 3120
rect 15160 3080 15332 3108
rect 15160 3068 15166 3080
rect 13817 3043 13875 3049
rect 13817 3040 13829 3043
rect 13740 3012 13829 3040
rect 13633 3003 13691 3009
rect 13817 3009 13829 3012
rect 13863 3009 13875 3043
rect 14093 3043 14151 3049
rect 14093 3040 14105 3043
rect 13817 3003 13875 3009
rect 13922 3012 14105 3040
rect 12084 2944 12388 2972
rect 12542 2944 12940 2972
rect 13290 2944 13492 2972
rect 13648 2972 13676 3003
rect 13722 2972 13728 2984
rect 13648 2944 13728 2972
rect 11882 2904 11888 2916
rect 11808 2876 11888 2904
rect 11379 2873 11391 2876
rect 11333 2867 11391 2873
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 12069 2907 12127 2913
rect 12069 2873 12081 2907
rect 12115 2904 12127 2907
rect 12158 2904 12164 2916
rect 12115 2876 12164 2904
rect 12115 2873 12127 2876
rect 12069 2867 12127 2873
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 12360 2913 12388 2944
rect 12912 2913 12940 2944
rect 13722 2932 13728 2944
rect 13780 2932 13786 2984
rect 12345 2907 12403 2913
rect 12345 2873 12357 2907
rect 12391 2873 12403 2907
rect 12345 2867 12403 2873
rect 12897 2907 12955 2913
rect 12897 2873 12909 2907
rect 12943 2873 12955 2907
rect 12897 2867 12955 2873
rect 12986 2864 12992 2916
rect 13044 2904 13050 2916
rect 13265 2907 13323 2913
rect 13265 2904 13277 2907
rect 13044 2876 13277 2904
rect 13044 2864 13050 2876
rect 13265 2873 13277 2876
rect 13311 2873 13323 2907
rect 13265 2867 13323 2873
rect 13354 2864 13360 2916
rect 13412 2904 13418 2916
rect 13922 2904 13950 3012
rect 14093 3009 14105 3012
rect 14139 3009 14151 3043
rect 14093 3003 14151 3009
rect 14357 3000 14363 3052
rect 14415 3038 14421 3052
rect 14458 3038 14504 3040
rect 14415 3010 14504 3038
rect 14415 3000 14421 3010
rect 13998 2932 14004 2984
rect 14056 2932 14062 2984
rect 14476 2981 14504 3010
rect 14642 3000 14648 3052
rect 14700 3000 14706 3052
rect 14844 3040 14872 3068
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14844 3012 15209 3040
rect 15197 3009 15209 3012
rect 15243 3009 15255 3043
rect 15304 3040 15332 3080
rect 15470 3068 15476 3120
rect 15528 3108 15534 3120
rect 15749 3111 15807 3117
rect 15749 3108 15761 3111
rect 15528 3080 15761 3108
rect 15528 3068 15534 3080
rect 15749 3077 15761 3080
rect 15795 3077 15807 3111
rect 15749 3071 15807 3077
rect 16298 3068 16304 3120
rect 16356 3068 16362 3120
rect 16960 3108 16988 3136
rect 18322 3108 18328 3120
rect 16960 3080 18328 3108
rect 18322 3068 18328 3080
rect 18380 3068 18386 3120
rect 18598 3068 18604 3120
rect 18656 3108 18662 3120
rect 18938 3111 18996 3117
rect 18938 3108 18950 3111
rect 18656 3080 18950 3108
rect 18656 3068 18662 3080
rect 18938 3077 18950 3080
rect 18984 3077 18996 3111
rect 18938 3071 18996 3077
rect 19518 3068 19524 3120
rect 19576 3108 19582 3120
rect 20257 3111 20315 3117
rect 20257 3108 20269 3111
rect 19576 3080 20269 3108
rect 19576 3068 19582 3080
rect 20257 3077 20269 3080
rect 20303 3077 20315 3111
rect 20257 3071 20315 3077
rect 15304 3012 15884 3040
rect 15197 3003 15255 3009
rect 15856 2984 15884 3012
rect 16482 3000 16488 3052
rect 16540 3000 16546 3052
rect 16574 3000 16580 3052
rect 16632 3040 16638 3052
rect 17109 3043 17167 3049
rect 17109 3040 17121 3043
rect 16632 3012 17121 3040
rect 16632 3000 16638 3012
rect 17109 3009 17121 3012
rect 17155 3009 17167 3043
rect 17109 3003 17167 3009
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 18417 3043 18475 3049
rect 18417 3040 18429 3043
rect 17460 3012 18429 3040
rect 17460 3000 17466 3012
rect 18417 3009 18429 3012
rect 18463 3009 18475 3043
rect 18417 3003 18475 3009
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3040 18751 3043
rect 18782 3040 18788 3052
rect 18739 3012 18788 3040
rect 18739 3009 18751 3012
rect 18693 3003 18751 3009
rect 18782 3000 18788 3012
rect 18840 3000 18846 3052
rect 14461 2975 14519 2981
rect 14461 2941 14473 2975
rect 14507 2941 14519 2975
rect 14461 2935 14519 2941
rect 13412 2876 13950 2904
rect 14016 2904 14044 2932
rect 14476 2904 14504 2935
rect 14918 2932 14924 2984
rect 14976 2932 14982 2984
rect 15286 2972 15292 2984
rect 15145 2944 15292 2972
rect 15145 2904 15173 2944
rect 15286 2932 15292 2944
rect 15344 2932 15350 2984
rect 15838 2932 15844 2984
rect 15896 2972 15902 2984
rect 16666 2972 16672 2984
rect 15896 2944 16672 2972
rect 15896 2932 15902 2944
rect 16666 2932 16672 2944
rect 16724 2972 16730 2984
rect 16853 2975 16911 2981
rect 16853 2972 16865 2975
rect 16724 2944 16865 2972
rect 16724 2932 16730 2944
rect 16853 2941 16865 2944
rect 16899 2941 16911 2975
rect 16853 2935 16911 2941
rect 15930 2904 15936 2916
rect 14016 2876 14394 2904
rect 14476 2876 15173 2904
rect 15220 2876 15936 2904
rect 13412 2864 13418 2876
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2805 8723 2839
rect 8665 2799 8723 2805
rect 8938 2796 8944 2848
rect 8996 2796 9002 2848
rect 9214 2796 9220 2848
rect 9272 2796 9278 2848
rect 9493 2839 9551 2845
rect 9493 2805 9505 2839
rect 9539 2836 9551 2839
rect 9674 2836 9680 2848
rect 9539 2808 9680 2836
rect 9539 2805 9551 2808
rect 9493 2799 9551 2805
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 9766 2796 9772 2848
rect 9824 2796 9830 2848
rect 10410 2796 10416 2848
rect 10468 2796 10474 2848
rect 10597 2839 10655 2845
rect 10597 2805 10609 2839
rect 10643 2836 10655 2839
rect 10686 2836 10692 2848
rect 10643 2808 10692 2836
rect 10643 2805 10655 2808
rect 10597 2799 10655 2805
rect 10686 2796 10692 2808
rect 10744 2796 10750 2848
rect 10870 2796 10876 2848
rect 10928 2796 10934 2848
rect 11422 2796 11428 2848
rect 11480 2836 11486 2848
rect 11609 2839 11667 2845
rect 11609 2836 11621 2839
rect 11480 2808 11621 2836
rect 11480 2796 11486 2808
rect 11609 2805 11621 2808
rect 11655 2805 11667 2839
rect 11609 2799 11667 2805
rect 13170 2796 13176 2848
rect 13228 2836 13234 2848
rect 13814 2836 13820 2848
rect 13228 2808 13820 2836
rect 13228 2796 13234 2808
rect 13814 2796 13820 2808
rect 13872 2796 13878 2848
rect 13906 2796 13912 2848
rect 13964 2796 13970 2848
rect 14274 2796 14280 2848
rect 14332 2796 14338 2848
rect 14366 2836 14394 2876
rect 15220 2836 15248 2876
rect 15930 2864 15936 2876
rect 15988 2864 15994 2916
rect 20073 2907 20131 2913
rect 20073 2873 20085 2907
rect 20119 2873 20131 2907
rect 20073 2867 20131 2873
rect 14366 2808 15248 2836
rect 15286 2796 15292 2848
rect 15344 2796 15350 2848
rect 15470 2796 15476 2848
rect 15528 2836 15534 2848
rect 15841 2839 15899 2845
rect 15841 2836 15853 2839
rect 15528 2808 15853 2836
rect 15528 2796 15534 2808
rect 15841 2805 15853 2808
rect 15887 2805 15899 2839
rect 15841 2799 15899 2805
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 16850 2836 16856 2848
rect 16172 2808 16856 2836
rect 16172 2796 16178 2808
rect 16850 2796 16856 2808
rect 16908 2796 16914 2848
rect 17218 2796 17224 2848
rect 17276 2836 17282 2848
rect 20088 2836 20116 2867
rect 17276 2808 20116 2836
rect 17276 2796 17282 2808
rect 1104 2746 20884 2768
rect 1104 2694 3422 2746
rect 3474 2694 3486 2746
rect 3538 2694 3550 2746
rect 3602 2694 3614 2746
rect 3666 2694 3678 2746
rect 3730 2694 8367 2746
rect 8419 2694 8431 2746
rect 8483 2694 8495 2746
rect 8547 2694 8559 2746
rect 8611 2694 8623 2746
rect 8675 2694 13312 2746
rect 13364 2694 13376 2746
rect 13428 2694 13440 2746
rect 13492 2694 13504 2746
rect 13556 2694 13568 2746
rect 13620 2694 18257 2746
rect 18309 2694 18321 2746
rect 18373 2694 18385 2746
rect 18437 2694 18449 2746
rect 18501 2694 18513 2746
rect 18565 2694 20884 2746
rect 1104 2672 20884 2694
rect 1670 2592 1676 2644
rect 1728 2592 1734 2644
rect 2869 2635 2927 2641
rect 2869 2601 2881 2635
rect 2915 2632 2927 2635
rect 2958 2632 2964 2644
rect 2915 2604 2964 2632
rect 2915 2601 2927 2604
rect 2869 2595 2927 2601
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 3786 2632 3792 2644
rect 3651 2604 3792 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4341 2635 4399 2641
rect 4341 2601 4353 2635
rect 4387 2632 4399 2635
rect 4430 2632 4436 2644
rect 4387 2604 4436 2632
rect 4387 2601 4399 2604
rect 4341 2595 4399 2601
rect 4430 2592 4436 2604
rect 4488 2592 4494 2644
rect 4801 2635 4859 2641
rect 4801 2601 4813 2635
rect 4847 2632 4859 2635
rect 5166 2632 5172 2644
rect 4847 2604 5172 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5350 2592 5356 2644
rect 5408 2592 5414 2644
rect 6181 2635 6239 2641
rect 6181 2601 6193 2635
rect 6227 2632 6239 2635
rect 6454 2632 6460 2644
rect 6227 2604 6460 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 7006 2592 7012 2644
rect 7064 2592 7070 2644
rect 7466 2592 7472 2644
rect 7524 2632 7530 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7524 2604 7849 2632
rect 7524 2592 7530 2604
rect 7837 2601 7849 2604
rect 7883 2632 7895 2635
rect 8386 2632 8392 2644
rect 7883 2604 8392 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 8386 2592 8392 2604
rect 8444 2592 8450 2644
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 11422 2632 11428 2644
rect 9088 2604 11428 2632
rect 9088 2592 9094 2604
rect 11422 2592 11428 2604
rect 11480 2592 11486 2644
rect 11514 2592 11520 2644
rect 11572 2632 11578 2644
rect 14093 2635 14151 2641
rect 14093 2632 14105 2635
rect 11572 2604 14105 2632
rect 11572 2592 11578 2604
rect 14093 2601 14105 2604
rect 14139 2601 14151 2635
rect 14093 2595 14151 2601
rect 14752 2604 16344 2632
rect 5721 2567 5779 2573
rect 5721 2533 5733 2567
rect 5767 2564 5779 2567
rect 6270 2564 6276 2576
rect 5767 2536 6276 2564
rect 5767 2533 5779 2536
rect 5721 2527 5779 2533
rect 6270 2524 6276 2536
rect 6328 2524 6334 2576
rect 7377 2567 7435 2573
rect 7377 2533 7389 2567
rect 7423 2564 7435 2567
rect 7423 2536 8156 2564
rect 7423 2533 7435 2536
rect 7377 2527 7435 2533
rect 1762 2456 1768 2508
rect 1820 2496 1826 2508
rect 1857 2499 1915 2505
rect 1857 2496 1869 2499
rect 1820 2468 1869 2496
rect 1820 2456 1826 2468
rect 1857 2465 1869 2468
rect 1903 2465 1915 2499
rect 4062 2496 4068 2508
rect 1857 2459 1915 2465
rect 3344 2468 4068 2496
rect 1489 2431 1547 2437
rect 1489 2397 1501 2431
rect 1535 2397 1547 2431
rect 1489 2391 1547 2397
rect 2131 2431 2189 2437
rect 2131 2397 2143 2431
rect 2177 2428 2189 2431
rect 3344 2428 3372 2468
rect 4062 2456 4068 2468
rect 4120 2456 4126 2508
rect 6380 2468 6868 2496
rect 6380 2440 6408 2468
rect 2177 2400 3372 2428
rect 2177 2397 2189 2400
rect 2131 2391 2189 2397
rect 1504 2360 1532 2391
rect 3418 2388 3424 2440
rect 3476 2388 3482 2440
rect 3786 2388 3792 2440
rect 3844 2388 3850 2440
rect 4522 2388 4528 2440
rect 4580 2388 4586 2440
rect 4617 2431 4675 2437
rect 4617 2397 4629 2431
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5169 2431 5227 2437
rect 5169 2397 5181 2431
rect 5215 2428 5227 2431
rect 5626 2428 5632 2440
rect 5215 2400 5632 2428
rect 5215 2397 5227 2400
rect 5169 2391 5227 2397
rect 2958 2360 2964 2372
rect 1504 2332 2964 2360
rect 2958 2320 2964 2332
rect 3016 2320 3022 2372
rect 4062 2320 4068 2372
rect 4120 2360 4126 2372
rect 4632 2360 4660 2391
rect 5626 2388 5632 2400
rect 5684 2388 5690 2440
rect 6362 2388 6368 2440
rect 6420 2388 6426 2440
rect 6638 2388 6644 2440
rect 6696 2388 6702 2440
rect 6840 2437 6868 2468
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 7340 2400 7573 2428
rect 7340 2388 7346 2400
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 8128 2428 8156 2536
rect 9306 2524 9312 2576
rect 9364 2564 9370 2576
rect 10505 2567 10563 2573
rect 9364 2536 9720 2564
rect 9364 2524 9370 2536
rect 9692 2496 9720 2536
rect 10505 2533 10517 2567
rect 10551 2564 10563 2567
rect 11698 2564 11704 2576
rect 10551 2536 11704 2564
rect 10551 2533 10563 2536
rect 10505 2527 10563 2533
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 11793 2567 11851 2573
rect 11793 2533 11805 2567
rect 11839 2564 11851 2567
rect 11839 2536 14143 2564
rect 11839 2533 11851 2536
rect 11793 2527 11851 2533
rect 13817 2499 13875 2505
rect 8312 2468 9628 2496
rect 9692 2468 11008 2496
rect 8312 2428 8340 2468
rect 8128 2400 8340 2428
rect 7561 2391 7619 2397
rect 8386 2388 8392 2440
rect 8444 2388 8450 2440
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2397 8539 2431
rect 8481 2391 8539 2397
rect 4120 2332 4660 2360
rect 4120 2320 4126 2332
rect 5534 2320 5540 2372
rect 5592 2320 5598 2372
rect 6089 2363 6147 2369
rect 6089 2329 6101 2363
rect 6135 2329 6147 2363
rect 6089 2323 6147 2329
rect 3970 2252 3976 2304
rect 4028 2252 4034 2304
rect 5902 2252 5908 2304
rect 5960 2292 5966 2304
rect 6104 2292 6132 2323
rect 6270 2320 6276 2372
rect 6328 2360 6334 2372
rect 6549 2363 6607 2369
rect 6549 2360 6561 2363
rect 6328 2332 6561 2360
rect 6328 2320 6334 2332
rect 6549 2329 6561 2332
rect 6595 2329 6607 2363
rect 6656 2360 6684 2388
rect 8496 2360 8524 2391
rect 9122 2388 9128 2440
rect 9180 2428 9186 2440
rect 9217 2431 9275 2437
rect 9217 2428 9229 2431
rect 9180 2400 9229 2428
rect 9180 2388 9186 2400
rect 9217 2397 9229 2400
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 9490 2388 9496 2440
rect 9548 2388 9554 2440
rect 9600 2437 9628 2468
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 10134 2388 10140 2440
rect 10192 2388 10198 2440
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2397 10471 2431
rect 10413 2391 10471 2397
rect 10428 2360 10456 2391
rect 10686 2388 10692 2440
rect 10744 2388 10750 2440
rect 10980 2437 11008 2468
rect 11164 2468 13584 2496
rect 11164 2440 11192 2468
rect 10965 2431 11023 2437
rect 10965 2397 10977 2431
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11333 2431 11391 2437
rect 11333 2428 11345 2431
rect 11296 2400 11345 2428
rect 11296 2388 11302 2400
rect 11333 2397 11345 2400
rect 11379 2397 11391 2431
rect 11333 2391 11391 2397
rect 11422 2388 11428 2440
rect 11480 2388 11486 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11716 2400 11989 2428
rect 6656 2332 8524 2360
rect 9508 2332 10364 2360
rect 10428 2332 11468 2360
rect 6549 2323 6607 2329
rect 9508 2304 9536 2332
rect 5960 2264 6132 2292
rect 5960 2252 5966 2264
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6236 2264 6653 2292
rect 6236 2252 6242 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 8205 2295 8263 2301
rect 8205 2261 8217 2295
rect 8251 2292 8263 2295
rect 8570 2292 8576 2304
rect 8251 2264 8576 2292
rect 8251 2261 8263 2264
rect 8205 2255 8263 2261
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 8665 2295 8723 2301
rect 8665 2261 8677 2295
rect 8711 2292 8723 2295
rect 8938 2292 8944 2304
rect 8711 2264 8944 2292
rect 8711 2261 8723 2264
rect 8665 2255 8723 2261
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 9030 2252 9036 2304
rect 9088 2252 9094 2304
rect 9306 2252 9312 2304
rect 9364 2252 9370 2304
rect 9490 2252 9496 2304
rect 9548 2252 9554 2304
rect 9769 2295 9827 2301
rect 9769 2261 9781 2295
rect 9815 2292 9827 2295
rect 9858 2292 9864 2304
rect 9815 2264 9864 2292
rect 9815 2261 9827 2264
rect 9769 2255 9827 2261
rect 9858 2252 9864 2264
rect 9916 2252 9922 2304
rect 9950 2252 9956 2304
rect 10008 2252 10014 2304
rect 10226 2252 10232 2304
rect 10284 2252 10290 2304
rect 10336 2292 10364 2332
rect 11440 2304 11468 2332
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10336 2264 10793 2292
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 11149 2295 11207 2301
rect 11149 2261 11161 2295
rect 11195 2292 11207 2295
rect 11238 2292 11244 2304
rect 11195 2264 11244 2292
rect 11195 2261 11207 2264
rect 11149 2255 11207 2261
rect 11238 2252 11244 2264
rect 11296 2252 11302 2304
rect 11422 2252 11428 2304
rect 11480 2252 11486 2304
rect 11606 2252 11612 2304
rect 11664 2252 11670 2304
rect 11716 2292 11744 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12250 2388 12256 2440
rect 12308 2388 12314 2440
rect 12526 2388 12532 2440
rect 12584 2388 12590 2440
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2428 12863 2431
rect 12894 2428 12900 2440
rect 12851 2400 12900 2428
rect 12851 2397 12863 2400
rect 12805 2391 12863 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2428 13231 2431
rect 13354 2428 13360 2440
rect 13219 2400 13360 2428
rect 13219 2397 13231 2400
rect 13173 2391 13231 2397
rect 13354 2388 13360 2400
rect 13412 2388 13418 2440
rect 13556 2437 13584 2468
rect 13817 2465 13829 2499
rect 13863 2496 13875 2499
rect 13906 2496 13912 2508
rect 13863 2468 13912 2496
rect 13863 2465 13875 2468
rect 13817 2459 13875 2465
rect 13906 2456 13912 2468
rect 13964 2456 13970 2508
rect 14115 2496 14143 2536
rect 14366 2524 14372 2576
rect 14424 2564 14430 2576
rect 14642 2564 14648 2576
rect 14424 2536 14648 2564
rect 14424 2524 14430 2536
rect 14642 2524 14648 2536
rect 14700 2524 14706 2576
rect 14752 2496 14780 2604
rect 14115 2468 14780 2496
rect 13541 2431 13599 2437
rect 13541 2397 13553 2431
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 13630 2388 13636 2440
rect 13688 2428 13694 2440
rect 14182 2428 14188 2440
rect 13688 2400 14188 2428
rect 13688 2388 13694 2400
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 14277 2431 14335 2437
rect 14277 2397 14289 2431
rect 14323 2428 14335 2431
rect 14737 2431 14795 2437
rect 14323 2400 14688 2428
rect 14323 2397 14335 2400
rect 14277 2391 14335 2397
rect 11790 2320 11796 2372
rect 11848 2360 11854 2372
rect 12636 2360 12664 2388
rect 14366 2360 14372 2372
rect 11848 2332 12388 2360
rect 12636 2332 14372 2360
rect 11848 2320 11854 2332
rect 11974 2292 11980 2304
rect 11716 2264 11980 2292
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 12066 2252 12072 2304
rect 12124 2252 12130 2304
rect 12360 2301 12388 2332
rect 14366 2320 14372 2332
rect 14424 2320 14430 2372
rect 12345 2295 12403 2301
rect 12345 2261 12357 2295
rect 12391 2261 12403 2295
rect 12345 2255 12403 2261
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 12621 2295 12679 2301
rect 12621 2292 12633 2295
rect 12492 2264 12633 2292
rect 12492 2252 12498 2264
rect 12621 2261 12633 2264
rect 12667 2261 12679 2295
rect 12621 2255 12679 2261
rect 12986 2252 12992 2304
rect 13044 2252 13050 2304
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 14458 2292 14464 2304
rect 13780 2264 14464 2292
rect 13780 2252 13786 2264
rect 14458 2252 14464 2264
rect 14516 2252 14522 2304
rect 14660 2301 14688 2400
rect 14737 2397 14749 2431
rect 14783 2397 14795 2431
rect 14737 2391 14795 2397
rect 14752 2360 14780 2391
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 16316 2437 16344 2604
rect 16390 2592 16396 2644
rect 16448 2592 16454 2644
rect 16574 2592 16580 2644
rect 16632 2632 16638 2644
rect 20070 2632 20076 2644
rect 16632 2604 20076 2632
rect 16632 2592 16638 2604
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 16482 2524 16488 2576
rect 16540 2564 16546 2576
rect 18877 2567 18935 2573
rect 18877 2564 18889 2567
rect 16540 2536 18889 2564
rect 16540 2524 16546 2536
rect 18877 2533 18889 2536
rect 18923 2533 18935 2567
rect 18877 2527 18935 2533
rect 19242 2524 19248 2576
rect 19300 2524 19306 2576
rect 17218 2496 17224 2508
rect 16408 2468 17224 2496
rect 15004 2431 15062 2437
rect 15004 2428 15016 2431
rect 14884 2400 15016 2428
rect 14884 2388 14890 2400
rect 15004 2397 15016 2400
rect 15050 2397 15062 2431
rect 15004 2391 15062 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2397 16359 2431
rect 16301 2391 16359 2397
rect 15654 2360 15660 2372
rect 14752 2332 15660 2360
rect 15654 2320 15660 2332
rect 15712 2360 15718 2372
rect 15838 2360 15844 2372
rect 15712 2332 15844 2360
rect 15712 2320 15718 2332
rect 15838 2320 15844 2332
rect 15896 2320 15902 2372
rect 15930 2320 15936 2372
rect 15988 2360 15994 2372
rect 16408 2360 16436 2468
rect 17218 2456 17224 2468
rect 17276 2456 17282 2508
rect 17494 2456 17500 2508
rect 17552 2456 17558 2508
rect 18509 2499 18567 2505
rect 18509 2465 18521 2499
rect 18555 2496 18567 2499
rect 18690 2496 18696 2508
rect 18555 2468 18696 2496
rect 18555 2465 18567 2468
rect 18509 2459 18567 2465
rect 18690 2456 18696 2468
rect 18748 2496 18754 2508
rect 19260 2496 19288 2524
rect 18748 2468 19288 2496
rect 18748 2456 18754 2468
rect 16482 2388 16488 2440
rect 16540 2388 16546 2440
rect 16666 2388 16672 2440
rect 16724 2388 16730 2440
rect 19076 2437 19104 2468
rect 19061 2431 19119 2437
rect 19061 2397 19073 2431
rect 19107 2428 19119 2431
rect 20254 2428 20260 2440
rect 19107 2400 19141 2428
rect 19996 2400 20260 2428
rect 19107 2397 19119 2400
rect 19061 2391 19119 2397
rect 15988 2332 16436 2360
rect 16500 2360 16528 2388
rect 17865 2363 17923 2369
rect 17865 2360 17877 2363
rect 16500 2332 17877 2360
rect 15988 2320 15994 2332
rect 17865 2329 17877 2332
rect 17911 2329 17923 2363
rect 17865 2323 17923 2329
rect 19150 2320 19156 2372
rect 19208 2360 19214 2372
rect 19337 2363 19395 2369
rect 19337 2360 19349 2363
rect 19208 2332 19349 2360
rect 19208 2320 19214 2332
rect 19337 2329 19349 2332
rect 19383 2329 19395 2363
rect 19337 2323 19395 2329
rect 19996 2304 20024 2400
rect 20254 2388 20260 2400
rect 20312 2428 20318 2440
rect 20533 2431 20591 2437
rect 20533 2428 20545 2431
rect 20312 2400 20545 2428
rect 20312 2388 20318 2400
rect 20533 2397 20545 2400
rect 20579 2397 20591 2431
rect 20533 2391 20591 2397
rect 14645 2295 14703 2301
rect 14645 2261 14657 2295
rect 14691 2292 14703 2295
rect 14734 2292 14740 2304
rect 14691 2264 14740 2292
rect 14691 2261 14703 2264
rect 14645 2255 14703 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 14918 2252 14924 2304
rect 14976 2292 14982 2304
rect 16117 2295 16175 2301
rect 16117 2292 16129 2295
rect 14976 2264 16129 2292
rect 14976 2252 14982 2264
rect 16117 2261 16129 2264
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 16482 2252 16488 2304
rect 16540 2292 16546 2304
rect 17034 2292 17040 2304
rect 16540 2264 17040 2292
rect 16540 2252 16546 2264
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 17957 2295 18015 2301
rect 17957 2292 17969 2295
rect 17276 2264 17969 2292
rect 17276 2252 17282 2264
rect 17957 2261 17969 2264
rect 18003 2261 18015 2295
rect 17957 2255 18015 2261
rect 19242 2252 19248 2304
rect 19300 2292 19306 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 19300 2264 19441 2292
rect 19300 2252 19306 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 19978 2252 19984 2304
rect 20036 2252 20042 2304
rect 20346 2252 20352 2304
rect 20404 2252 20410 2304
rect 1104 2202 21043 2224
rect 1104 2150 5894 2202
rect 5946 2150 5958 2202
rect 6010 2150 6022 2202
rect 6074 2150 6086 2202
rect 6138 2150 6150 2202
rect 6202 2150 10839 2202
rect 10891 2150 10903 2202
rect 10955 2150 10967 2202
rect 11019 2150 11031 2202
rect 11083 2150 11095 2202
rect 11147 2150 15784 2202
rect 15836 2150 15848 2202
rect 15900 2150 15912 2202
rect 15964 2150 15976 2202
rect 16028 2150 16040 2202
rect 16092 2150 20729 2202
rect 20781 2150 20793 2202
rect 20845 2150 20857 2202
rect 20909 2150 20921 2202
rect 20973 2150 20985 2202
rect 21037 2150 21043 2202
rect 1104 2128 21043 2150
rect 1394 2048 1400 2100
rect 1452 2088 1458 2100
rect 1765 2091 1823 2097
rect 1765 2088 1777 2091
rect 1452 2060 1777 2088
rect 1452 2048 1458 2060
rect 1765 2057 1777 2060
rect 1811 2057 1823 2091
rect 2685 2091 2743 2097
rect 2685 2088 2697 2091
rect 1765 2051 1823 2057
rect 1964 2060 2697 2088
rect 1302 1980 1308 2032
rect 1360 2020 1366 2032
rect 1964 2020 1992 2060
rect 2685 2057 2697 2060
rect 2731 2057 2743 2091
rect 2685 2051 2743 2057
rect 3789 2091 3847 2097
rect 3789 2057 3801 2091
rect 3835 2088 3847 2091
rect 4154 2088 4160 2100
rect 3835 2060 4160 2088
rect 3835 2057 3847 2060
rect 3789 2051 3847 2057
rect 4154 2048 4160 2060
rect 4212 2048 4218 2100
rect 4890 2088 4896 2100
rect 4264 2060 4896 2088
rect 1360 1992 1992 2020
rect 1360 1980 1366 1992
rect 2406 1980 2412 2032
rect 2464 1980 2470 2032
rect 2590 1980 2596 2032
rect 2648 1980 2654 2032
rect 1673 1955 1731 1961
rect 1673 1921 1685 1955
rect 1719 1952 1731 1955
rect 2424 1952 2452 1980
rect 1719 1924 2452 1952
rect 1719 1921 1731 1924
rect 1673 1915 1731 1921
rect 3234 1912 3240 1964
rect 3292 1912 3298 1964
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1921 3755 1955
rect 3697 1915 3755 1921
rect 750 1844 756 1896
rect 808 1844 814 1896
rect 2774 1844 2780 1896
rect 2832 1884 2838 1896
rect 3712 1884 3740 1915
rect 3970 1912 3976 1964
rect 4028 1912 4034 1964
rect 4154 1912 4160 1964
rect 4212 1952 4218 1964
rect 4264 1952 4292 2060
rect 4890 2048 4896 2060
rect 4948 2048 4954 2100
rect 6546 2088 6552 2100
rect 6012 2060 6552 2088
rect 6012 2029 6040 2060
rect 6546 2048 6552 2060
rect 6604 2048 6610 2100
rect 6822 2048 6828 2100
rect 6880 2048 6886 2100
rect 7006 2048 7012 2100
rect 7064 2048 7070 2100
rect 7834 2048 7840 2100
rect 7892 2088 7898 2100
rect 7892 2060 8800 2088
rect 7892 2048 7898 2060
rect 5997 2023 6055 2029
rect 4632 1992 5948 2020
rect 4632 1961 4660 1992
rect 4212 1924 4292 1952
rect 4617 1955 4675 1961
rect 4212 1912 4218 1924
rect 4617 1921 4629 1955
rect 4663 1921 4675 1955
rect 4617 1915 4675 1921
rect 4982 1912 4988 1964
rect 5040 1912 5046 1964
rect 5534 1912 5540 1964
rect 5592 1952 5598 1964
rect 5813 1955 5871 1961
rect 5813 1952 5825 1955
rect 5592 1924 5825 1952
rect 5592 1912 5598 1924
rect 5813 1921 5825 1924
rect 5859 1921 5871 1955
rect 5920 1952 5948 1992
rect 5997 1989 6009 2023
rect 6043 1989 6055 2023
rect 6840 2020 6868 2048
rect 5997 1983 6055 1989
rect 6472 1992 6868 2020
rect 7653 2023 7711 2029
rect 6472 1961 6500 1992
rect 7653 1989 7665 2023
rect 7699 2020 7711 2023
rect 8110 2020 8116 2032
rect 7699 1992 8116 2020
rect 7699 1989 7711 1992
rect 7653 1983 7711 1989
rect 8110 1980 8116 1992
rect 8168 1980 8174 2032
rect 8478 1980 8484 2032
rect 8536 1980 8542 2032
rect 8570 1980 8576 2032
rect 8628 1980 8634 2032
rect 8772 2029 8800 2060
rect 9306 2048 9312 2100
rect 9364 2048 9370 2100
rect 9950 2048 9956 2100
rect 10008 2088 10014 2100
rect 10008 2060 13676 2088
rect 10008 2048 10014 2060
rect 8757 2023 8815 2029
rect 8757 1989 8769 2023
rect 8803 1989 8815 2023
rect 9324 2020 9352 2048
rect 10965 2023 11023 2029
rect 10965 2020 10977 2023
rect 9324 1992 10977 2020
rect 8757 1983 8815 1989
rect 10965 1989 10977 1992
rect 11011 1989 11023 2023
rect 10965 1983 11023 1989
rect 11330 1980 11336 2032
rect 11388 2020 11394 2032
rect 12345 2023 12403 2029
rect 12345 2020 12357 2023
rect 11388 1992 12357 2020
rect 11388 1980 11394 1992
rect 12345 1989 12357 1992
rect 12391 1989 12403 2023
rect 12345 1983 12403 1989
rect 12897 2023 12955 2029
rect 12897 1989 12909 2023
rect 12943 2020 12955 2023
rect 13538 2020 13544 2032
rect 12943 1992 13544 2020
rect 12943 1989 12955 1992
rect 12897 1983 12955 1989
rect 13538 1980 13544 1992
rect 13596 1980 13602 2032
rect 13648 2020 13676 2060
rect 14458 2048 14464 2100
rect 14516 2088 14522 2100
rect 15197 2091 15255 2097
rect 15197 2088 15209 2091
rect 14516 2060 15209 2088
rect 14516 2048 14522 2060
rect 15197 2057 15209 2060
rect 15243 2057 15255 2091
rect 15197 2051 15255 2057
rect 15286 2048 15292 2100
rect 15344 2088 15350 2100
rect 16206 2088 16212 2100
rect 15344 2060 16212 2088
rect 15344 2048 15350 2060
rect 16206 2048 16212 2060
rect 16264 2048 16270 2100
rect 16390 2048 16396 2100
rect 16448 2088 16454 2100
rect 16574 2088 16580 2100
rect 16448 2060 16580 2088
rect 16448 2048 16454 2060
rect 16574 2048 16580 2060
rect 16632 2048 16638 2100
rect 19797 2091 19855 2097
rect 19797 2088 19809 2091
rect 19306 2060 19809 2088
rect 13983 2023 14041 2029
rect 13983 2020 13995 2023
rect 13648 1992 13995 2020
rect 13983 1989 13995 1992
rect 14029 1989 14041 2023
rect 14274 2020 14280 2032
rect 13983 1983 14041 1989
rect 14115 1992 14280 2020
rect 6457 1955 6515 1961
rect 5920 1924 6408 1952
rect 5813 1915 5871 1921
rect 2832 1856 3740 1884
rect 2832 1844 2838 1856
rect 4706 1844 4712 1896
rect 4764 1844 4770 1896
rect 5166 1844 5172 1896
rect 5224 1884 5230 1896
rect 6181 1887 6239 1893
rect 6181 1884 6193 1887
rect 5224 1856 6193 1884
rect 5224 1844 5230 1856
rect 6181 1853 6193 1856
rect 6227 1853 6239 1887
rect 6181 1847 6239 1853
rect 768 1816 796 1844
rect 3421 1819 3479 1825
rect 3421 1816 3433 1819
rect 768 1788 3433 1816
rect 3421 1785 3433 1788
rect 3467 1785 3479 1819
rect 3421 1779 3479 1785
rect 4433 1819 4491 1825
rect 4433 1785 4445 1819
rect 4479 1816 4491 1819
rect 6270 1816 6276 1828
rect 4479 1788 6276 1816
rect 4479 1785 4491 1788
rect 4433 1779 4491 1785
rect 6270 1776 6276 1788
rect 6328 1776 6334 1828
rect 4157 1751 4215 1757
rect 4157 1717 4169 1751
rect 4203 1748 4215 1751
rect 4522 1748 4528 1760
rect 4203 1720 4528 1748
rect 4203 1717 4215 1720
rect 4157 1711 4215 1717
rect 4522 1708 4528 1720
rect 4580 1708 4586 1760
rect 5629 1751 5687 1757
rect 5629 1717 5641 1751
rect 5675 1748 5687 1751
rect 5994 1748 6000 1760
rect 5675 1720 6000 1748
rect 5675 1717 5687 1720
rect 5629 1711 5687 1717
rect 5994 1708 6000 1720
rect 6052 1708 6058 1760
rect 6380 1748 6408 1924
rect 6457 1921 6469 1955
rect 6503 1921 6515 1955
rect 6457 1915 6515 1921
rect 6825 1955 6883 1961
rect 6825 1921 6837 1955
rect 6871 1921 6883 1955
rect 6825 1915 6883 1921
rect 6840 1884 6868 1915
rect 6914 1912 6920 1964
rect 6972 1952 6978 1964
rect 7193 1955 7251 1961
rect 7193 1952 7205 1955
rect 6972 1924 7205 1952
rect 6972 1912 6978 1924
rect 7193 1921 7205 1924
rect 7239 1921 7251 1955
rect 7193 1915 7251 1921
rect 7558 1912 7564 1964
rect 7616 1912 7622 1964
rect 7742 1912 7748 1964
rect 7800 1952 7806 1964
rect 7929 1955 7987 1961
rect 7929 1952 7941 1955
rect 7800 1924 7941 1952
rect 7800 1912 7806 1924
rect 7929 1921 7941 1924
rect 7975 1921 7987 1955
rect 7929 1915 7987 1921
rect 8202 1912 8208 1964
rect 8260 1952 8266 1964
rect 8297 1955 8355 1961
rect 8297 1952 8309 1955
rect 8260 1924 8309 1952
rect 8260 1912 8266 1924
rect 8297 1921 8309 1924
rect 8343 1921 8355 1955
rect 8297 1915 8355 1921
rect 7576 1884 7604 1912
rect 8496 1884 8524 1980
rect 6840 1856 7604 1884
rect 7760 1856 8524 1884
rect 8588 1884 8616 1980
rect 9306 1912 9312 1964
rect 9364 1912 9370 1964
rect 9582 1912 9588 1964
rect 9640 1952 9646 1964
rect 9861 1955 9919 1961
rect 9861 1952 9873 1955
rect 9640 1924 9873 1952
rect 9640 1912 9646 1924
rect 9861 1921 9873 1924
rect 9907 1921 9919 1955
rect 9861 1915 9919 1921
rect 10413 1955 10471 1961
rect 10413 1921 10425 1955
rect 10459 1921 10471 1955
rect 11793 1955 11851 1961
rect 11793 1952 11805 1955
rect 10413 1915 10471 1921
rect 10520 1924 11805 1952
rect 10428 1884 10456 1915
rect 8588 1856 10456 1884
rect 6641 1819 6699 1825
rect 6641 1785 6653 1819
rect 6687 1816 6699 1819
rect 7466 1816 7472 1828
rect 6687 1788 7472 1816
rect 6687 1785 6699 1788
rect 6641 1779 6699 1785
rect 7466 1776 7472 1788
rect 7524 1776 7530 1828
rect 7760 1816 7788 1856
rect 7576 1788 7788 1816
rect 6914 1748 6920 1760
rect 6380 1720 6920 1748
rect 6914 1708 6920 1720
rect 6972 1708 6978 1760
rect 7377 1751 7435 1757
rect 7377 1717 7389 1751
rect 7423 1748 7435 1751
rect 7576 1748 7604 1788
rect 7834 1776 7840 1828
rect 7892 1816 7898 1828
rect 8846 1816 8852 1828
rect 7892 1788 8852 1816
rect 7892 1776 7898 1788
rect 8846 1776 8852 1788
rect 8904 1776 8910 1828
rect 9674 1776 9680 1828
rect 9732 1816 9738 1828
rect 10520 1816 10548 1924
rect 11793 1921 11805 1924
rect 11839 1921 11851 1955
rect 11793 1915 11851 1921
rect 11882 1912 11888 1964
rect 11940 1952 11946 1964
rect 12618 1952 12624 1964
rect 11940 1924 12624 1952
rect 11940 1912 11946 1924
rect 12618 1912 12624 1924
rect 12676 1912 12682 1964
rect 13449 1955 13507 1961
rect 13449 1921 13461 1955
rect 13495 1952 13507 1955
rect 14115 1952 14143 1992
rect 14274 1980 14280 1992
rect 14332 1980 14338 2032
rect 14366 1980 14372 2032
rect 14424 2020 14430 2032
rect 14553 2023 14611 2029
rect 14553 2020 14565 2023
rect 14424 1992 14565 2020
rect 14424 1980 14430 1992
rect 14553 1989 14565 1992
rect 14599 1989 14611 2023
rect 14553 1983 14611 1989
rect 14918 1980 14924 2032
rect 14976 2020 14982 2032
rect 19306 2020 19334 2060
rect 19797 2057 19809 2060
rect 19843 2057 19855 2091
rect 19797 2051 19855 2057
rect 14976 1992 19334 2020
rect 14976 1980 14982 1992
rect 15013 1955 15071 1961
rect 15013 1952 15025 1955
rect 13495 1924 14143 1952
rect 14200 1924 15025 1952
rect 13495 1921 13507 1924
rect 13449 1915 13507 1921
rect 11146 1844 11152 1896
rect 11204 1884 11210 1896
rect 12434 1884 12440 1896
rect 11204 1856 12440 1884
rect 11204 1844 11210 1856
rect 12434 1844 12440 1856
rect 12492 1844 12498 1896
rect 12894 1844 12900 1896
rect 12952 1884 12958 1896
rect 12952 1856 13768 1884
rect 12952 1844 12958 1856
rect 9732 1788 10548 1816
rect 9732 1776 9738 1788
rect 10870 1776 10876 1828
rect 10928 1816 10934 1828
rect 10928 1788 12002 1816
rect 10928 1776 10934 1788
rect 7423 1720 7604 1748
rect 7423 1717 7435 1720
rect 7377 1711 7435 1717
rect 7650 1708 7656 1760
rect 7708 1748 7714 1760
rect 7745 1751 7803 1757
rect 7745 1748 7757 1751
rect 7708 1720 7757 1748
rect 7708 1708 7714 1720
rect 7745 1717 7757 1720
rect 7791 1717 7803 1751
rect 7745 1711 7803 1717
rect 8110 1708 8116 1760
rect 8168 1708 8174 1760
rect 8202 1708 8208 1760
rect 8260 1748 8266 1760
rect 8481 1751 8539 1757
rect 8481 1748 8493 1751
rect 8260 1720 8493 1748
rect 8260 1708 8266 1720
rect 8481 1717 8493 1720
rect 8527 1717 8539 1751
rect 8481 1711 8539 1717
rect 9033 1751 9091 1757
rect 9033 1717 9045 1751
rect 9079 1748 9091 1751
rect 9398 1748 9404 1760
rect 9079 1720 9404 1748
rect 9079 1717 9091 1720
rect 9033 1711 9091 1717
rect 9398 1708 9404 1720
rect 9456 1708 9462 1760
rect 9582 1708 9588 1760
rect 9640 1708 9646 1760
rect 10134 1708 10140 1760
rect 10192 1708 10198 1760
rect 10502 1708 10508 1760
rect 10560 1708 10566 1760
rect 10686 1708 10692 1760
rect 10744 1748 10750 1760
rect 11057 1751 11115 1757
rect 11057 1748 11069 1751
rect 10744 1720 11069 1748
rect 10744 1708 10750 1720
rect 11057 1717 11069 1720
rect 11103 1717 11115 1751
rect 11057 1711 11115 1717
rect 11882 1708 11888 1760
rect 11940 1708 11946 1760
rect 11974 1748 12002 1788
rect 12158 1776 12164 1828
rect 12216 1816 12222 1828
rect 12802 1816 12808 1828
rect 12216 1788 12808 1816
rect 12216 1776 12222 1788
rect 12802 1776 12808 1788
rect 12860 1776 12866 1828
rect 13630 1816 13636 1828
rect 12912 1788 13636 1816
rect 12526 1748 12532 1760
rect 11974 1720 12532 1748
rect 12526 1708 12532 1720
rect 12584 1708 12590 1760
rect 12621 1751 12679 1757
rect 12621 1717 12633 1751
rect 12667 1748 12679 1751
rect 12912 1748 12940 1788
rect 13630 1776 13636 1788
rect 13688 1776 13694 1828
rect 13740 1816 13768 1856
rect 14090 1844 14096 1896
rect 14148 1884 14154 1896
rect 14200 1884 14228 1924
rect 15013 1921 15025 1924
rect 15059 1921 15071 1955
rect 15013 1915 15071 1921
rect 15657 1955 15715 1961
rect 15657 1921 15669 1955
rect 15703 1952 15715 1955
rect 15703 1924 16160 1952
rect 15703 1921 15715 1924
rect 15657 1915 15715 1921
rect 14148 1856 14228 1884
rect 14148 1844 14154 1856
rect 14274 1844 14280 1896
rect 14332 1884 14338 1896
rect 14332 1856 14872 1884
rect 14332 1844 14338 1856
rect 14458 1816 14464 1828
rect 13740 1788 14464 1816
rect 14458 1776 14464 1788
rect 14516 1776 14522 1828
rect 14734 1776 14740 1828
rect 14792 1776 14798 1828
rect 14844 1816 14872 1856
rect 14918 1844 14924 1896
rect 14976 1884 14982 1896
rect 15286 1884 15292 1896
rect 14976 1856 15292 1884
rect 14976 1844 14982 1856
rect 15286 1844 15292 1856
rect 15344 1844 15350 1896
rect 16022 1844 16028 1896
rect 16080 1844 16086 1896
rect 16132 1884 16160 1924
rect 16298 1912 16304 1964
rect 16356 1952 16362 1964
rect 16669 1955 16727 1961
rect 16669 1952 16681 1955
rect 16356 1924 16681 1952
rect 16356 1912 16362 1924
rect 16669 1921 16681 1924
rect 16715 1921 16727 1955
rect 16669 1915 16727 1921
rect 17034 1912 17040 1964
rect 17092 1952 17098 1964
rect 18509 1955 18567 1961
rect 18509 1952 18521 1955
rect 17092 1924 18521 1952
rect 17092 1912 17098 1924
rect 18509 1921 18521 1924
rect 18555 1921 18567 1955
rect 18509 1915 18567 1921
rect 20530 1912 20536 1964
rect 20588 1912 20594 1964
rect 17494 1884 17500 1896
rect 16132 1856 17500 1884
rect 17494 1844 17500 1856
rect 17552 1844 17558 1896
rect 20349 1819 20407 1825
rect 20349 1816 20361 1819
rect 14844 1788 20361 1816
rect 20349 1785 20361 1788
rect 20395 1785 20407 1819
rect 20349 1779 20407 1785
rect 12667 1720 12940 1748
rect 12667 1717 12679 1720
rect 12621 1711 12679 1717
rect 12986 1708 12992 1760
rect 13044 1708 13050 1760
rect 13078 1708 13084 1760
rect 13136 1748 13142 1760
rect 13541 1751 13599 1757
rect 13541 1748 13553 1751
rect 13136 1720 13553 1748
rect 13136 1708 13142 1720
rect 13541 1717 13553 1720
rect 13587 1717 13599 1751
rect 13541 1711 13599 1717
rect 13722 1708 13728 1760
rect 13780 1748 13786 1760
rect 14093 1751 14151 1757
rect 14093 1748 14105 1751
rect 13780 1720 14105 1748
rect 13780 1708 13786 1720
rect 14093 1717 14105 1720
rect 14139 1717 14151 1751
rect 14093 1711 14151 1717
rect 14182 1708 14188 1760
rect 14240 1748 14246 1760
rect 16390 1748 16396 1760
rect 14240 1720 16396 1748
rect 14240 1708 14246 1720
rect 16390 1708 16396 1720
rect 16448 1708 16454 1760
rect 16482 1708 16488 1760
rect 16540 1748 16546 1760
rect 17957 1751 18015 1757
rect 17957 1748 17969 1751
rect 16540 1720 17969 1748
rect 16540 1708 16546 1720
rect 17957 1717 17969 1720
rect 18003 1717 18015 1751
rect 17957 1711 18015 1717
rect 1104 1658 20884 1680
rect 1104 1606 3422 1658
rect 3474 1606 3486 1658
rect 3538 1606 3550 1658
rect 3602 1606 3614 1658
rect 3666 1606 3678 1658
rect 3730 1606 8367 1658
rect 8419 1606 8431 1658
rect 8483 1606 8495 1658
rect 8547 1606 8559 1658
rect 8611 1606 8623 1658
rect 8675 1606 13312 1658
rect 13364 1606 13376 1658
rect 13428 1606 13440 1658
rect 13492 1606 13504 1658
rect 13556 1606 13568 1658
rect 13620 1606 18257 1658
rect 18309 1606 18321 1658
rect 18373 1606 18385 1658
rect 18437 1606 18449 1658
rect 18501 1606 18513 1658
rect 18565 1606 20884 1658
rect 1104 1584 20884 1606
rect 1854 1504 1860 1556
rect 1912 1504 1918 1556
rect 2409 1547 2467 1553
rect 2409 1513 2421 1547
rect 2455 1544 2467 1547
rect 2498 1544 2504 1556
rect 2455 1516 2504 1544
rect 2455 1513 2467 1516
rect 2409 1507 2467 1513
rect 2498 1504 2504 1516
rect 2556 1504 2562 1556
rect 2777 1547 2835 1553
rect 2777 1513 2789 1547
rect 2823 1544 2835 1547
rect 4154 1544 4160 1556
rect 2823 1516 4160 1544
rect 2823 1513 2835 1516
rect 2777 1507 2835 1513
rect 4154 1504 4160 1516
rect 4212 1504 4218 1556
rect 4338 1504 4344 1556
rect 4396 1544 4402 1556
rect 4617 1547 4675 1553
rect 4617 1544 4629 1547
rect 4396 1516 4629 1544
rect 4396 1504 4402 1516
rect 4617 1513 4629 1516
rect 4663 1513 4675 1547
rect 4617 1507 4675 1513
rect 4982 1504 4988 1556
rect 5040 1504 5046 1556
rect 5074 1504 5080 1556
rect 5132 1544 5138 1556
rect 5353 1547 5411 1553
rect 5353 1544 5365 1547
rect 5132 1516 5365 1544
rect 5132 1504 5138 1516
rect 5353 1513 5365 1516
rect 5399 1513 5411 1547
rect 5353 1507 5411 1513
rect 5721 1547 5779 1553
rect 5721 1513 5733 1547
rect 5767 1513 5779 1547
rect 5721 1507 5779 1513
rect 474 1436 480 1488
rect 532 1476 538 1488
rect 3237 1479 3295 1485
rect 3237 1476 3249 1479
rect 532 1448 3249 1476
rect 532 1436 538 1448
rect 3237 1445 3249 1448
rect 3283 1445 3295 1479
rect 3237 1439 3295 1445
rect 3605 1479 3663 1485
rect 3605 1445 3617 1479
rect 3651 1445 3663 1479
rect 4890 1476 4896 1488
rect 3605 1439 3663 1445
rect 3804 1448 4896 1476
rect 1026 1368 1032 1420
rect 1084 1408 1090 1420
rect 3620 1408 3648 1439
rect 1084 1380 3648 1408
rect 1084 1368 1090 1380
rect 14 1300 20 1352
rect 72 1340 78 1352
rect 3694 1340 3700 1352
rect 72 1312 2820 1340
rect 72 1300 78 1312
rect 1762 1232 1768 1284
rect 1820 1232 1826 1284
rect 2133 1275 2191 1281
rect 2133 1241 2145 1275
rect 2179 1272 2191 1275
rect 2179 1244 2360 1272
rect 2179 1241 2191 1244
rect 2133 1235 2191 1241
rect 2332 1204 2360 1244
rect 2406 1232 2412 1284
rect 2464 1272 2470 1284
rect 2685 1275 2743 1281
rect 2685 1272 2697 1275
rect 2464 1244 2697 1272
rect 2464 1232 2470 1244
rect 2685 1241 2697 1244
rect 2731 1241 2743 1275
rect 2685 1235 2743 1241
rect 2590 1204 2596 1216
rect 2332 1176 2596 1204
rect 2590 1164 2596 1176
rect 2648 1164 2654 1216
rect 2792 1204 2820 1312
rect 3068 1312 3700 1340
rect 3068 1281 3096 1312
rect 3694 1300 3700 1312
rect 3752 1300 3758 1352
rect 3804 1349 3832 1448
rect 4890 1436 4896 1448
rect 4948 1436 4954 1488
rect 5258 1436 5264 1488
rect 5316 1476 5322 1488
rect 5736 1476 5764 1507
rect 6086 1504 6092 1556
rect 6144 1504 6150 1556
rect 6638 1504 6644 1556
rect 6696 1504 6702 1556
rect 6822 1504 6828 1556
rect 6880 1544 6886 1556
rect 7009 1547 7067 1553
rect 7009 1544 7021 1547
rect 6880 1516 7021 1544
rect 6880 1504 6886 1516
rect 7009 1513 7021 1516
rect 7055 1513 7067 1547
rect 7009 1507 7067 1513
rect 9306 1504 9312 1556
rect 9364 1504 9370 1556
rect 9766 1504 9772 1556
rect 9824 1504 9830 1556
rect 10594 1504 10600 1556
rect 10652 1544 10658 1556
rect 10652 1516 12388 1544
rect 10652 1504 10658 1516
rect 5316 1448 5764 1476
rect 5316 1436 5322 1448
rect 5994 1436 6000 1488
rect 6052 1436 6058 1488
rect 9324 1476 9352 1504
rect 8404 1448 9352 1476
rect 5166 1408 5172 1420
rect 4080 1380 5172 1408
rect 4080 1349 4108 1380
rect 5166 1368 5172 1380
rect 5224 1368 5230 1420
rect 6012 1408 6040 1436
rect 6012 1380 7512 1408
rect 3789 1343 3847 1349
rect 3789 1309 3801 1343
rect 3835 1309 3847 1343
rect 3789 1303 3847 1309
rect 4065 1343 4123 1349
rect 4065 1309 4077 1343
rect 4111 1309 4123 1343
rect 4065 1303 4123 1309
rect 5350 1300 5356 1352
rect 5408 1300 5414 1352
rect 6362 1340 6368 1352
rect 5644 1312 6368 1340
rect 3053 1275 3111 1281
rect 3053 1241 3065 1275
rect 3099 1241 3111 1275
rect 3053 1235 3111 1241
rect 3421 1275 3479 1281
rect 3421 1241 3433 1275
rect 3467 1272 3479 1275
rect 4430 1272 4436 1284
rect 3467 1244 4436 1272
rect 3467 1241 3479 1244
rect 3421 1235 3479 1241
rect 4430 1232 4436 1244
rect 4488 1232 4494 1284
rect 4522 1232 4528 1284
rect 4580 1232 4586 1284
rect 4890 1232 4896 1284
rect 4948 1232 4954 1284
rect 5258 1232 5264 1284
rect 5316 1232 5322 1284
rect 3973 1207 4031 1213
rect 3973 1204 3985 1207
rect 2792 1176 3985 1204
rect 3973 1173 3985 1176
rect 4019 1173 4031 1207
rect 3973 1167 4031 1173
rect 4249 1207 4307 1213
rect 4249 1173 4261 1207
rect 4295 1204 4307 1207
rect 5074 1204 5080 1216
rect 4295 1176 5080 1204
rect 4295 1173 4307 1176
rect 4249 1167 4307 1173
rect 5074 1164 5080 1176
rect 5132 1164 5138 1216
rect 5368 1204 5396 1300
rect 5644 1281 5672 1312
rect 6362 1300 6368 1312
rect 6420 1300 6426 1352
rect 6457 1343 6515 1349
rect 6457 1309 6469 1343
rect 6503 1340 6515 1343
rect 6546 1340 6552 1352
rect 6503 1312 6552 1340
rect 6503 1309 6515 1312
rect 6457 1303 6515 1309
rect 6546 1300 6552 1312
rect 6604 1300 6610 1352
rect 6730 1300 6736 1352
rect 6788 1340 6794 1352
rect 7484 1349 7512 1380
rect 6917 1343 6975 1349
rect 6917 1340 6929 1343
rect 6788 1312 6929 1340
rect 6788 1300 6794 1312
rect 6917 1309 6929 1312
rect 6963 1309 6975 1343
rect 6917 1303 6975 1309
rect 7469 1343 7527 1349
rect 7469 1309 7481 1343
rect 7515 1309 7527 1343
rect 7469 1303 7527 1309
rect 7834 1300 7840 1352
rect 7892 1300 7898 1352
rect 8404 1349 8432 1448
rect 9784 1408 9812 1504
rect 9858 1436 9864 1488
rect 9916 1476 9922 1488
rect 10318 1476 10324 1488
rect 9916 1448 10324 1476
rect 9916 1436 9922 1448
rect 10318 1436 10324 1448
rect 10376 1436 10382 1488
rect 11701 1479 11759 1485
rect 11701 1445 11713 1479
rect 11747 1476 11759 1479
rect 11974 1476 11980 1488
rect 11747 1448 11980 1476
rect 11747 1445 11759 1448
rect 11701 1439 11759 1445
rect 11974 1436 11980 1448
rect 12032 1436 12038 1488
rect 9232 1380 9812 1408
rect 8389 1343 8447 1349
rect 8389 1309 8401 1343
rect 8435 1309 8447 1343
rect 8389 1303 8447 1309
rect 8941 1343 8999 1349
rect 8941 1309 8953 1343
rect 8987 1340 8999 1343
rect 9232 1340 9260 1380
rect 10042 1354 10048 1406
rect 10100 1354 10106 1406
rect 11606 1354 11612 1406
rect 11664 1354 11670 1406
rect 11790 1368 11796 1420
rect 11848 1408 11854 1420
rect 12250 1408 12256 1420
rect 11848 1380 12256 1408
rect 11848 1368 11854 1380
rect 12250 1368 12256 1380
rect 12308 1368 12314 1420
rect 12360 1408 12388 1516
rect 12434 1504 12440 1556
rect 12492 1544 12498 1556
rect 13173 1547 13231 1553
rect 13173 1544 13185 1547
rect 12492 1516 13185 1544
rect 12492 1504 12498 1516
rect 13173 1513 13185 1516
rect 13219 1513 13231 1547
rect 13173 1507 13231 1513
rect 13280 1516 14318 1544
rect 12618 1436 12624 1488
rect 12676 1476 12682 1488
rect 13280 1476 13308 1516
rect 12676 1448 13308 1476
rect 12676 1436 12682 1448
rect 13354 1436 13360 1488
rect 13412 1436 13418 1488
rect 13630 1436 13636 1488
rect 13688 1476 13694 1488
rect 13688 1448 14044 1476
rect 13688 1436 13694 1448
rect 13262 1408 13268 1420
rect 12360 1380 13268 1408
rect 13262 1368 13268 1380
rect 13320 1368 13326 1420
rect 13372 1408 13400 1436
rect 14016 1408 14044 1448
rect 14090 1436 14096 1488
rect 14148 1436 14154 1488
rect 14182 1408 14188 1420
rect 13372 1380 13768 1408
rect 14016 1380 14188 1408
rect 9766 1340 9772 1352
rect 8987 1312 9260 1340
rect 9324 1312 9772 1340
rect 8987 1309 8999 1312
rect 8941 1303 8999 1309
rect 5629 1275 5687 1281
rect 5629 1241 5641 1275
rect 5675 1241 5687 1275
rect 5629 1235 5687 1241
rect 5997 1275 6055 1281
rect 5997 1241 6009 1275
rect 6043 1241 6055 1275
rect 5997 1235 6055 1241
rect 8205 1275 8263 1281
rect 8205 1241 8217 1275
rect 8251 1241 8263 1275
rect 8205 1235 8263 1241
rect 8757 1275 8815 1281
rect 8757 1241 8769 1275
rect 8803 1272 8815 1275
rect 9324 1272 9352 1312
rect 9766 1300 9772 1312
rect 9824 1300 9830 1352
rect 8803 1244 9352 1272
rect 9401 1275 9459 1281
rect 8803 1241 8815 1244
rect 8757 1235 8815 1241
rect 9401 1241 9413 1275
rect 9447 1272 9459 1275
rect 9490 1272 9496 1284
rect 9447 1244 9496 1272
rect 9447 1241 9459 1244
rect 9401 1235 9459 1241
rect 6012 1204 6040 1235
rect 5368 1176 6040 1204
rect 7558 1164 7564 1216
rect 7616 1164 7622 1216
rect 8220 1204 8248 1235
rect 9490 1232 9496 1244
rect 9548 1232 9554 1284
rect 9953 1275 10011 1281
rect 9953 1241 9965 1275
rect 9999 1272 10011 1275
rect 10060 1272 10088 1354
rect 10597 1343 10655 1349
rect 10597 1309 10609 1343
rect 10643 1309 10655 1343
rect 10597 1303 10655 1309
rect 9999 1244 10088 1272
rect 10612 1272 10640 1303
rect 11054 1300 11060 1352
rect 11112 1300 11118 1352
rect 11238 1300 11244 1352
rect 11296 1300 11302 1352
rect 11514 1300 11520 1352
rect 11572 1300 11578 1352
rect 11256 1272 11284 1300
rect 10612 1244 11284 1272
rect 9999 1241 10011 1244
rect 9953 1235 10011 1241
rect 11422 1232 11428 1284
rect 11480 1272 11486 1284
rect 11624 1272 11652 1354
rect 11698 1300 11704 1352
rect 11756 1340 11762 1352
rect 12529 1343 12587 1349
rect 12529 1340 12541 1343
rect 11756 1312 12541 1340
rect 11756 1300 11762 1312
rect 12529 1309 12541 1312
rect 12575 1309 12587 1343
rect 12529 1303 12587 1309
rect 12710 1300 12716 1352
rect 12768 1340 12774 1352
rect 12768 1312 13308 1340
rect 12768 1300 12774 1312
rect 11480 1244 11652 1272
rect 11480 1232 11486 1244
rect 11882 1232 11888 1284
rect 11940 1232 11946 1284
rect 11977 1275 12035 1281
rect 11977 1241 11989 1275
rect 12023 1272 12035 1275
rect 12250 1272 12256 1284
rect 12023 1244 12256 1272
rect 12023 1241 12035 1244
rect 11977 1235 12035 1241
rect 12250 1232 12256 1244
rect 12308 1232 12314 1284
rect 12345 1275 12403 1281
rect 12345 1241 12357 1275
rect 12391 1272 12403 1275
rect 12434 1272 12440 1284
rect 12391 1244 12440 1272
rect 12391 1241 12403 1244
rect 12345 1235 12403 1241
rect 12434 1232 12440 1244
rect 12492 1232 12498 1284
rect 12894 1232 12900 1284
rect 12952 1272 12958 1284
rect 13081 1275 13139 1281
rect 13081 1272 13093 1275
rect 12952 1244 13093 1272
rect 12952 1232 12958 1244
rect 13081 1241 13093 1244
rect 13127 1241 13139 1275
rect 13280 1272 13308 1312
rect 13538 1300 13544 1352
rect 13596 1300 13602 1352
rect 13740 1340 13768 1380
rect 14182 1368 14188 1380
rect 14240 1368 14246 1420
rect 14290 1408 14318 1516
rect 14642 1504 14648 1556
rect 14700 1544 14706 1556
rect 14700 1516 14872 1544
rect 14700 1504 14706 1516
rect 14844 1476 14872 1516
rect 15010 1504 15016 1556
rect 15068 1544 15074 1556
rect 15378 1544 15384 1556
rect 15068 1516 15384 1544
rect 15068 1504 15074 1516
rect 15378 1504 15384 1516
rect 15436 1504 15442 1556
rect 15470 1504 15476 1556
rect 15528 1544 15534 1556
rect 16574 1544 16580 1556
rect 15528 1516 16580 1544
rect 15528 1504 15534 1516
rect 16574 1504 16580 1516
rect 16632 1504 16638 1556
rect 17402 1544 17408 1556
rect 16776 1516 17408 1544
rect 16482 1476 16488 1488
rect 14844 1448 16488 1476
rect 16482 1436 16488 1448
rect 16540 1436 16546 1488
rect 14737 1411 14795 1417
rect 14737 1408 14749 1411
rect 14290 1380 14749 1408
rect 14737 1377 14749 1380
rect 14783 1377 14795 1411
rect 14737 1371 14795 1377
rect 15010 1368 15016 1420
rect 15068 1408 15074 1420
rect 16776 1408 16804 1516
rect 17402 1504 17408 1516
rect 17460 1504 17466 1556
rect 18046 1504 18052 1556
rect 18104 1544 18110 1556
rect 20349 1547 20407 1553
rect 20349 1544 20361 1547
rect 18104 1516 20361 1544
rect 18104 1504 18110 1516
rect 20349 1513 20361 1516
rect 20395 1513 20407 1547
rect 20349 1507 20407 1513
rect 16850 1436 16856 1488
rect 16908 1476 16914 1488
rect 17126 1476 17132 1488
rect 16908 1448 17132 1476
rect 16908 1436 16914 1448
rect 17126 1436 17132 1448
rect 17184 1436 17190 1488
rect 15068 1380 16804 1408
rect 15068 1368 15074 1380
rect 16942 1368 16948 1420
rect 17000 1408 17006 1420
rect 17037 1411 17095 1417
rect 17037 1408 17049 1411
rect 17000 1380 17049 1408
rect 17000 1368 17006 1380
rect 17037 1377 17049 1380
rect 17083 1377 17095 1411
rect 17037 1371 17095 1377
rect 17310 1368 17316 1420
rect 17368 1408 17374 1420
rect 17368 1380 19380 1408
rect 17368 1368 17374 1380
rect 14277 1343 14335 1349
rect 13740 1312 14143 1340
rect 13814 1272 13820 1284
rect 13280 1244 13820 1272
rect 13081 1235 13139 1241
rect 13814 1232 13820 1244
rect 13872 1232 13878 1284
rect 9030 1204 9036 1216
rect 8220 1176 9036 1204
rect 9030 1164 9036 1176
rect 9088 1164 9094 1216
rect 9122 1164 9128 1216
rect 9180 1164 9186 1216
rect 9674 1164 9680 1216
rect 9732 1164 9738 1216
rect 9766 1164 9772 1216
rect 9824 1204 9830 1216
rect 10045 1207 10103 1213
rect 10045 1204 10057 1207
rect 9824 1176 10057 1204
rect 9824 1164 9830 1176
rect 10045 1173 10057 1176
rect 10091 1173 10103 1207
rect 10045 1167 10103 1173
rect 10594 1164 10600 1216
rect 10652 1204 10658 1216
rect 10689 1207 10747 1213
rect 10689 1204 10701 1207
rect 10652 1176 10701 1204
rect 10652 1164 10658 1176
rect 10689 1173 10701 1176
rect 10735 1173 10747 1207
rect 10689 1167 10747 1173
rect 11241 1207 11299 1213
rect 11241 1173 11253 1207
rect 11287 1204 11299 1207
rect 11514 1204 11520 1216
rect 11287 1176 11520 1204
rect 11287 1173 11299 1176
rect 11241 1167 11299 1173
rect 11514 1164 11520 1176
rect 11572 1164 11578 1216
rect 11698 1164 11704 1216
rect 11756 1204 11762 1216
rect 11900 1204 11928 1232
rect 11756 1176 11928 1204
rect 11756 1164 11762 1176
rect 12158 1164 12164 1216
rect 12216 1204 12222 1216
rect 12621 1207 12679 1213
rect 12621 1204 12633 1207
rect 12216 1176 12633 1204
rect 12216 1164 12222 1176
rect 12621 1173 12633 1176
rect 12667 1173 12679 1207
rect 12621 1167 12679 1173
rect 12710 1164 12716 1216
rect 12768 1204 12774 1216
rect 13725 1207 13783 1213
rect 13725 1204 13737 1207
rect 12768 1176 13737 1204
rect 12768 1164 12774 1176
rect 13725 1173 13737 1176
rect 13771 1173 13783 1207
rect 14115 1204 14143 1312
rect 14277 1309 14289 1343
rect 14323 1340 14335 1343
rect 14553 1343 14611 1349
rect 14323 1316 14412 1340
rect 14323 1312 14504 1316
rect 14323 1309 14335 1312
rect 14277 1303 14335 1309
rect 14384 1288 14504 1312
rect 14553 1309 14565 1343
rect 14599 1336 14611 1343
rect 15657 1343 15715 1349
rect 14743 1336 15611 1340
rect 14599 1312 15611 1336
rect 14599 1309 14771 1312
rect 14553 1308 14771 1309
rect 14553 1303 14611 1308
rect 14476 1272 14504 1288
rect 15583 1272 15611 1312
rect 15657 1309 15669 1343
rect 15703 1340 15715 1343
rect 16114 1340 16120 1352
rect 15703 1312 16120 1340
rect 15703 1309 15715 1312
rect 15657 1303 15715 1309
rect 16114 1300 16120 1312
rect 16172 1300 16178 1352
rect 16298 1300 16304 1352
rect 16356 1300 16362 1352
rect 16574 1300 16580 1352
rect 16632 1340 16638 1352
rect 16669 1343 16727 1349
rect 16669 1340 16681 1343
rect 16632 1312 16681 1340
rect 16632 1300 16638 1312
rect 16669 1309 16681 1312
rect 16715 1309 16727 1343
rect 16669 1303 16727 1309
rect 17126 1300 17132 1352
rect 17184 1300 17190 1352
rect 17954 1300 17960 1352
rect 18012 1300 18018 1352
rect 18049 1343 18107 1349
rect 18049 1309 18061 1343
rect 18095 1309 18107 1343
rect 18049 1303 18107 1309
rect 17144 1272 17172 1300
rect 18064 1272 18092 1303
rect 18874 1300 18880 1352
rect 18932 1300 18938 1352
rect 19352 1349 19380 1380
rect 19610 1368 19616 1420
rect 19668 1368 19674 1420
rect 19337 1343 19395 1349
rect 19337 1309 19349 1343
rect 19383 1309 19395 1343
rect 19337 1303 19395 1309
rect 19794 1300 19800 1352
rect 19852 1340 19858 1352
rect 20533 1343 20591 1349
rect 20533 1340 20545 1343
rect 19852 1312 20545 1340
rect 19852 1300 19858 1312
rect 20533 1309 20545 1312
rect 20579 1309 20591 1343
rect 20533 1303 20591 1309
rect 14476 1244 15516 1272
rect 15583 1244 17172 1272
rect 17236 1244 18092 1272
rect 15010 1204 15016 1216
rect 14115 1176 15016 1204
rect 13725 1167 13783 1173
rect 15010 1164 15016 1176
rect 15068 1164 15074 1216
rect 15488 1204 15516 1244
rect 16298 1204 16304 1216
rect 15488 1176 16304 1204
rect 16298 1164 16304 1176
rect 16356 1164 16362 1216
rect 16482 1164 16488 1216
rect 16540 1204 16546 1216
rect 17236 1204 17264 1244
rect 16540 1176 17264 1204
rect 16540 1164 16546 1176
rect 17770 1164 17776 1216
rect 17828 1164 17834 1216
rect 1104 1114 21043 1136
rect 1104 1062 5894 1114
rect 5946 1062 5958 1114
rect 6010 1062 6022 1114
rect 6074 1062 6086 1114
rect 6138 1062 6150 1114
rect 6202 1062 10839 1114
rect 10891 1062 10903 1114
rect 10955 1062 10967 1114
rect 11019 1062 11031 1114
rect 11083 1062 11095 1114
rect 11147 1062 15784 1114
rect 15836 1062 15848 1114
rect 15900 1062 15912 1114
rect 15964 1062 15976 1114
rect 16028 1062 16040 1114
rect 16092 1062 20729 1114
rect 20781 1062 20793 1114
rect 20845 1062 20857 1114
rect 20909 1062 20921 1114
rect 20973 1062 20985 1114
rect 21037 1062 21043 1114
rect 1104 1040 21043 1062
rect 5350 960 5356 1012
rect 5408 1000 5414 1012
rect 7650 1000 7656 1012
rect 5408 972 7656 1000
rect 5408 960 5414 972
rect 7650 960 7656 972
rect 7708 960 7714 1012
rect 9306 960 9312 1012
rect 9364 1000 9370 1012
rect 9364 972 9674 1000
rect 9364 960 9370 972
rect 9646 932 9674 972
rect 10594 960 10600 1012
rect 10652 1000 10658 1012
rect 11238 1000 11244 1012
rect 10652 972 11244 1000
rect 10652 960 10658 972
rect 11238 960 11244 972
rect 11296 960 11302 1012
rect 11514 960 11520 1012
rect 11572 1000 11578 1012
rect 11790 1000 11796 1012
rect 11572 972 11796 1000
rect 11572 960 11578 972
rect 11790 960 11796 972
rect 11848 960 11854 1012
rect 13998 960 14004 1012
rect 14056 1000 14062 1012
rect 14458 1000 14464 1012
rect 14056 972 14464 1000
rect 14056 960 14062 972
rect 14458 960 14464 972
rect 14516 960 14522 1012
rect 14550 960 14556 1012
rect 14608 960 14614 1012
rect 14826 960 14832 1012
rect 14884 960 14890 1012
rect 15010 960 15016 1012
rect 15068 1000 15074 1012
rect 17218 1000 17224 1012
rect 15068 972 17224 1000
rect 15068 960 15074 972
rect 17218 960 17224 972
rect 17276 960 17282 1012
rect 18046 960 18052 1012
rect 18104 960 18110 1012
rect 14568 932 14596 960
rect 9646 904 14596 932
rect 14844 932 14872 960
rect 17770 932 17776 944
rect 14844 904 17776 932
rect 17770 892 17776 904
rect 17828 892 17834 944
rect 10226 824 10232 876
rect 10284 864 10290 876
rect 10962 864 10968 876
rect 10284 836 10968 864
rect 10284 824 10290 836
rect 10962 824 10968 836
rect 11020 824 11026 876
rect 13262 824 13268 876
rect 13320 864 13326 876
rect 13320 836 13860 864
rect 13320 824 13326 836
rect 10042 756 10048 808
rect 10100 796 10106 808
rect 13538 796 13544 808
rect 10100 768 13544 796
rect 10100 756 10106 768
rect 13538 756 13544 768
rect 13596 756 13602 808
rect 13832 796 13860 836
rect 13906 824 13912 876
rect 13964 864 13970 876
rect 15746 864 15752 876
rect 13964 836 14897 864
rect 13964 824 13970 836
rect 14734 796 14740 808
rect 13832 768 14740 796
rect 14734 756 14740 768
rect 14792 756 14798 808
rect 14869 796 14897 836
rect 15053 836 15752 864
rect 15053 796 15081 836
rect 15746 824 15752 836
rect 15804 824 15810 876
rect 15838 824 15844 876
rect 15896 864 15902 876
rect 18064 864 18092 960
rect 15896 836 18092 864
rect 15896 824 15902 836
rect 20346 796 20352 808
rect 14869 768 15081 796
rect 15120 768 20352 796
rect 4522 688 4528 740
rect 4580 728 4586 740
rect 6086 728 6092 740
rect 4580 700 6092 728
rect 4580 688 4586 700
rect 6086 688 6092 700
rect 6144 688 6150 740
rect 10226 688 10232 740
rect 10284 728 10290 740
rect 10284 700 11192 728
rect 10284 688 10290 700
rect 1762 620 1768 672
rect 1820 660 1826 672
rect 3326 660 3332 672
rect 1820 632 3332 660
rect 1820 620 1826 632
rect 3326 620 3332 632
rect 3384 620 3390 672
rect 5258 620 5264 672
rect 5316 660 5322 672
rect 6638 660 6644 672
rect 5316 632 6644 660
rect 5316 620 5322 632
rect 6638 620 6644 632
rect 6696 620 6702 672
rect 9674 620 9680 672
rect 9732 660 9738 672
rect 11054 660 11060 672
rect 9732 632 11060 660
rect 9732 620 9738 632
rect 11054 620 11060 632
rect 11112 620 11118 672
rect 11164 660 11192 700
rect 12526 688 12532 740
rect 12584 728 12590 740
rect 12584 700 13860 728
rect 12584 688 12590 700
rect 13262 660 13268 672
rect 11164 632 13268 660
rect 13262 620 13268 632
rect 13320 620 13326 672
rect 9122 552 9128 604
rect 9180 592 9186 604
rect 10594 592 10600 604
rect 9180 564 10600 592
rect 9180 552 9186 564
rect 10594 552 10600 564
rect 10652 552 10658 604
rect 12250 552 12256 604
rect 12308 592 12314 604
rect 13722 592 13728 604
rect 12308 564 13728 592
rect 12308 552 12314 564
rect 13722 552 13728 564
rect 13780 552 13786 604
rect 13832 592 13860 700
rect 13906 688 13912 740
rect 13964 728 13970 740
rect 15120 728 15148 768
rect 20346 756 20352 768
rect 20404 756 20410 808
rect 13964 700 15148 728
rect 13964 688 13970 700
rect 15378 688 15384 740
rect 15436 728 15442 740
rect 15838 728 15844 740
rect 15436 700 15844 728
rect 15436 688 15442 700
rect 15838 688 15844 700
rect 15896 688 15902 740
rect 16022 688 16028 740
rect 16080 728 16086 740
rect 16574 728 16580 740
rect 16080 700 16580 728
rect 16080 688 16086 700
rect 16574 688 16580 700
rect 16632 688 16638 740
rect 16758 688 16764 740
rect 16816 728 16822 740
rect 19978 728 19984 740
rect 16816 700 19984 728
rect 16816 688 16822 700
rect 19978 688 19984 700
rect 20036 688 20042 740
rect 14274 620 14280 672
rect 14332 660 14338 672
rect 20162 660 20168 672
rect 14332 632 20168 660
rect 14332 620 14338 632
rect 20162 620 20168 632
rect 20220 620 20226 672
rect 17862 592 17868 604
rect 13832 564 17868 592
rect 17862 552 17868 564
rect 17920 552 17926 604
rect 18690 552 18696 604
rect 18748 552 18754 604
rect 11146 484 11152 536
rect 11204 524 11210 536
rect 18708 524 18736 552
rect 11204 496 18736 524
rect 11204 484 11210 496
rect 2314 416 2320 468
rect 2372 456 2378 468
rect 14274 456 14280 468
rect 2372 428 14280 456
rect 2372 416 2378 428
rect 14274 416 14280 428
rect 14332 416 14338 468
rect 14366 416 14372 468
rect 14424 456 14430 468
rect 14826 456 14832 468
rect 14424 428 14832 456
rect 14424 416 14430 428
rect 14826 416 14832 428
rect 14884 416 14890 468
rect 14918 416 14924 468
rect 14976 456 14982 468
rect 15102 456 15108 468
rect 14976 428 15108 456
rect 14976 416 14982 428
rect 15102 416 15108 428
rect 15160 416 15166 468
rect 15286 416 15292 468
rect 15344 456 15350 468
rect 18230 456 18236 468
rect 15344 428 18236 456
rect 15344 416 15350 428
rect 18230 416 18236 428
rect 18288 416 18294 468
rect 11514 348 11520 400
rect 11572 388 11578 400
rect 11572 360 13860 388
rect 11572 348 11578 360
rect 12434 280 12440 332
rect 12492 320 12498 332
rect 13722 320 13728 332
rect 12492 292 13728 320
rect 12492 280 12498 292
rect 13722 280 13728 292
rect 13780 280 13786 332
rect 13832 320 13860 360
rect 14182 348 14188 400
rect 14240 388 14246 400
rect 19242 388 19248 400
rect 14240 360 19248 388
rect 14240 348 14246 360
rect 19242 348 19248 360
rect 19300 348 19306 400
rect 19426 320 19432 332
rect 13832 292 19432 320
rect 19426 280 19432 292
rect 19484 280 19490 332
rect 13354 212 13360 264
rect 13412 252 13418 264
rect 19150 252 19156 264
rect 13412 224 19156 252
rect 13412 212 13418 224
rect 19150 212 19156 224
rect 19208 212 19214 264
rect 10410 144 10416 196
rect 10468 184 10474 196
rect 21174 184 21180 196
rect 10468 156 21180 184
rect 10468 144 10474 156
rect 21174 144 21180 156
rect 21232 144 21238 196
rect 10962 76 10968 128
rect 11020 116 11026 128
rect 20438 116 20444 128
rect 11020 88 20444 116
rect 11020 76 11026 88
rect 20438 76 20444 88
rect 20496 76 20502 128
rect 5074 8 5080 60
rect 5132 48 5138 60
rect 20622 48 20628 60
rect 5132 20 20628 48
rect 5132 8 5138 20
rect 20622 8 20628 20
rect 20680 8 20686 60
<< via1 >>
rect 1308 43800 1360 43852
rect 11520 43936 11572 43988
rect 17776 43936 17828 43988
rect 19432 43936 19484 43988
rect 2320 43732 2372 43784
rect 12072 43868 12124 43920
rect 13544 43868 13596 43920
rect 14924 43868 14976 43920
rect 18512 43868 18564 43920
rect 19248 43868 19300 43920
rect 9864 43800 9916 43852
rect 10140 43800 10192 43852
rect 5632 43664 5684 43716
rect 9680 43664 9732 43716
rect 19708 43800 19760 43852
rect 12440 43732 12492 43784
rect 13820 43664 13872 43716
rect 15200 43664 15252 43716
rect 19064 43664 19116 43716
rect 1492 43596 1544 43648
rect 10140 43596 10192 43648
rect 11704 43596 11756 43648
rect 13636 43596 13688 43648
rect 14188 43596 14240 43648
rect 14832 43596 14884 43648
rect 19800 43596 19852 43648
rect 5894 43494 5946 43546
rect 5958 43494 6010 43546
rect 6022 43494 6074 43546
rect 6086 43494 6138 43546
rect 6150 43494 6202 43546
rect 10839 43494 10891 43546
rect 10903 43494 10955 43546
rect 10967 43494 11019 43546
rect 11031 43494 11083 43546
rect 11095 43494 11147 43546
rect 15784 43494 15836 43546
rect 15848 43494 15900 43546
rect 15912 43494 15964 43546
rect 15976 43494 16028 43546
rect 16040 43494 16092 43546
rect 20729 43494 20781 43546
rect 20793 43494 20845 43546
rect 20857 43494 20909 43546
rect 20921 43494 20973 43546
rect 20985 43494 21037 43546
rect 2412 43392 2464 43444
rect 2780 43392 2832 43444
rect 3516 43392 3568 43444
rect 4160 43435 4212 43444
rect 4160 43401 4169 43435
rect 4169 43401 4203 43435
rect 4203 43401 4212 43435
rect 4160 43392 4212 43401
rect 4528 43435 4580 43444
rect 4528 43401 4537 43435
rect 4537 43401 4571 43435
rect 4571 43401 4580 43435
rect 4528 43392 4580 43401
rect 5540 43392 5592 43444
rect 7380 43392 7432 43444
rect 8668 43392 8720 43444
rect 1492 43299 1544 43308
rect 1492 43265 1501 43299
rect 1501 43265 1535 43299
rect 1535 43265 1544 43299
rect 1492 43256 1544 43265
rect 2136 43256 2188 43308
rect 2504 43299 2556 43308
rect 2504 43265 2513 43299
rect 2513 43265 2547 43299
rect 2547 43265 2556 43299
rect 2504 43256 2556 43265
rect 3056 43299 3108 43308
rect 3056 43265 3065 43299
rect 3065 43265 3099 43299
rect 3099 43265 3108 43299
rect 3056 43256 3108 43265
rect 4160 43256 4212 43308
rect 4344 43256 4396 43308
rect 7196 43324 7248 43376
rect 8392 43324 8444 43376
rect 8576 43324 8628 43376
rect 10600 43392 10652 43444
rect 5264 43299 5316 43308
rect 5264 43265 5273 43299
rect 5273 43265 5307 43299
rect 5307 43265 5316 43299
rect 5264 43256 5316 43265
rect 5448 43256 5500 43308
rect 3148 43188 3200 43240
rect 6736 43299 6788 43308
rect 6736 43265 6745 43299
rect 6745 43265 6779 43299
rect 6779 43265 6788 43299
rect 6736 43256 6788 43265
rect 7380 43188 7432 43240
rect 5816 43120 5868 43172
rect 6920 43120 6972 43172
rect 9036 43256 9088 43308
rect 9404 43256 9456 43308
rect 9496 43299 9548 43308
rect 9496 43265 9505 43299
rect 9505 43265 9539 43299
rect 9539 43265 9548 43299
rect 9496 43256 9548 43265
rect 9864 43256 9916 43308
rect 10416 43324 10468 43376
rect 11520 43392 11572 43444
rect 13268 43392 13320 43444
rect 10784 43299 10836 43308
rect 10784 43265 10793 43299
rect 10793 43265 10827 43299
rect 10827 43265 10836 43299
rect 10784 43256 10836 43265
rect 11704 43324 11756 43376
rect 11796 43367 11848 43376
rect 11796 43333 11805 43367
rect 11805 43333 11839 43367
rect 11839 43333 11848 43367
rect 11796 43324 11848 43333
rect 12900 43324 12952 43376
rect 11980 43256 12032 43308
rect 12256 43299 12308 43308
rect 12256 43265 12265 43299
rect 12265 43265 12299 43299
rect 12299 43265 12308 43299
rect 12256 43256 12308 43265
rect 12348 43256 12400 43308
rect 12716 43256 12768 43308
rect 14464 43392 14516 43444
rect 14188 43324 14240 43376
rect 16120 43392 16172 43444
rect 16212 43392 16264 43444
rect 8760 43188 8812 43240
rect 9680 43188 9732 43240
rect 14832 43256 14884 43308
rect 14924 43299 14976 43308
rect 14924 43265 14933 43299
rect 14933 43265 14967 43299
rect 14967 43265 14976 43299
rect 14924 43256 14976 43265
rect 15108 43256 15160 43308
rect 16304 43324 16356 43376
rect 16396 43324 16448 43376
rect 17500 43392 17552 43444
rect 19432 43435 19484 43444
rect 19432 43401 19441 43435
rect 19441 43401 19475 43435
rect 19475 43401 19484 43435
rect 19432 43392 19484 43401
rect 19800 43435 19852 43444
rect 19800 43401 19809 43435
rect 19809 43401 19843 43435
rect 19843 43401 19852 43435
rect 19800 43392 19852 43401
rect 15476 43299 15528 43308
rect 15476 43265 15485 43299
rect 15485 43265 15519 43299
rect 15519 43265 15528 43299
rect 15476 43256 15528 43265
rect 15660 43299 15712 43308
rect 15660 43265 15669 43299
rect 15669 43265 15703 43299
rect 15703 43265 15712 43299
rect 15660 43256 15712 43265
rect 16120 43299 16172 43308
rect 16120 43265 16129 43299
rect 16129 43265 16163 43299
rect 16163 43265 16172 43299
rect 16120 43256 16172 43265
rect 17224 43256 17276 43308
rect 17500 43256 17552 43308
rect 17960 43256 18012 43308
rect 18144 43256 18196 43308
rect 18604 43256 18656 43308
rect 18696 43299 18748 43308
rect 18696 43265 18705 43299
rect 18705 43265 18739 43299
rect 18739 43265 18748 43299
rect 18696 43256 18748 43265
rect 19064 43256 19116 43308
rect 19984 43299 20036 43308
rect 19984 43265 19993 43299
rect 19993 43265 20027 43299
rect 20027 43265 20036 43299
rect 19984 43256 20036 43265
rect 20168 43299 20220 43308
rect 20168 43265 20177 43299
rect 20177 43265 20211 43299
rect 20211 43265 20220 43299
rect 20168 43256 20220 43265
rect 8944 43120 8996 43172
rect 5908 43052 5960 43104
rect 6000 43052 6052 43104
rect 8576 43052 8628 43104
rect 9036 43052 9088 43104
rect 9680 43095 9732 43104
rect 9680 43061 9689 43095
rect 9689 43061 9723 43095
rect 9723 43061 9732 43095
rect 9680 43052 9732 43061
rect 9864 43052 9916 43104
rect 11612 43120 11664 43172
rect 12716 43120 12768 43172
rect 11152 43052 11204 43104
rect 11980 43052 12032 43104
rect 12992 43052 13044 43104
rect 13636 43120 13688 43172
rect 16948 43120 17000 43172
rect 13544 43095 13596 43104
rect 13544 43061 13553 43095
rect 13553 43061 13587 43095
rect 13587 43061 13596 43095
rect 13544 43052 13596 43061
rect 13728 43095 13780 43104
rect 13728 43061 13737 43095
rect 13737 43061 13771 43095
rect 13771 43061 13780 43095
rect 13728 43052 13780 43061
rect 14280 43095 14332 43104
rect 14280 43061 14289 43095
rect 14289 43061 14323 43095
rect 14323 43061 14332 43095
rect 14280 43052 14332 43061
rect 14464 43095 14516 43104
rect 14464 43061 14473 43095
rect 14473 43061 14507 43095
rect 14507 43061 14516 43095
rect 14464 43052 14516 43061
rect 14924 43052 14976 43104
rect 16396 43052 16448 43104
rect 16580 43052 16632 43104
rect 18052 43052 18104 43104
rect 18604 43052 18656 43104
rect 21272 43052 21324 43104
rect 3422 42950 3474 43002
rect 3486 42950 3538 43002
rect 3550 42950 3602 43002
rect 3614 42950 3666 43002
rect 3678 42950 3730 43002
rect 8367 42950 8419 43002
rect 8431 42950 8483 43002
rect 8495 42950 8547 43002
rect 8559 42950 8611 43002
rect 8623 42950 8675 43002
rect 13312 42950 13364 43002
rect 13376 42950 13428 43002
rect 13440 42950 13492 43002
rect 13504 42950 13556 43002
rect 13568 42950 13620 43002
rect 18257 42950 18309 43002
rect 18321 42950 18373 43002
rect 18385 42950 18437 43002
rect 18449 42950 18501 43002
rect 18513 42950 18565 43002
rect 3700 42848 3752 42900
rect 5264 42848 5316 42900
rect 6368 42848 6420 42900
rect 7288 42891 7340 42900
rect 7288 42857 7297 42891
rect 7297 42857 7331 42891
rect 7331 42857 7340 42891
rect 7288 42848 7340 42857
rect 7472 42848 7524 42900
rect 3608 42780 3660 42832
rect 9680 42780 9732 42832
rect 10140 42848 10192 42900
rect 10876 42891 10928 42900
rect 10876 42857 10885 42891
rect 10885 42857 10919 42891
rect 10919 42857 10928 42891
rect 10876 42848 10928 42857
rect 12900 42848 12952 42900
rect 14280 42848 14332 42900
rect 11336 42780 11388 42832
rect 12072 42780 12124 42832
rect 13452 42780 13504 42832
rect 14648 42780 14700 42832
rect 15108 42780 15160 42832
rect 1676 42687 1728 42696
rect 1676 42653 1685 42687
rect 1685 42653 1719 42687
rect 1719 42653 1728 42687
rect 1676 42644 1728 42653
rect 1952 42687 2004 42696
rect 1952 42653 1961 42687
rect 1961 42653 1995 42687
rect 1995 42653 2004 42687
rect 1952 42644 2004 42653
rect 2964 42644 3016 42696
rect 3332 42644 3384 42696
rect 3792 42712 3844 42764
rect 3884 42712 3936 42764
rect 4252 42712 4304 42764
rect 4344 42712 4396 42764
rect 4988 42712 5040 42764
rect 5356 42712 5408 42764
rect 6276 42712 6328 42764
rect 6460 42712 6512 42764
rect 8024 42755 8076 42764
rect 8024 42721 8033 42755
rect 8033 42721 8067 42755
rect 8067 42721 8076 42755
rect 8024 42712 8076 42721
rect 8300 42712 8352 42764
rect 5908 42644 5960 42696
rect 6920 42644 6972 42696
rect 1492 42551 1544 42560
rect 1492 42517 1501 42551
rect 1501 42517 1535 42551
rect 1535 42517 1544 42551
rect 1492 42508 1544 42517
rect 2688 42619 2740 42628
rect 2688 42585 2697 42619
rect 2697 42585 2731 42619
rect 2731 42585 2740 42619
rect 2688 42576 2740 42585
rect 3792 42576 3844 42628
rect 2964 42508 3016 42560
rect 3148 42508 3200 42560
rect 4252 42576 4304 42628
rect 4988 42619 5040 42628
rect 4988 42585 4997 42619
rect 4997 42585 5031 42619
rect 5031 42585 5040 42619
rect 4988 42576 5040 42585
rect 5816 42576 5868 42628
rect 6552 42576 6604 42628
rect 7012 42619 7064 42628
rect 7012 42585 7021 42619
rect 7021 42585 7055 42619
rect 7055 42585 7064 42619
rect 7012 42576 7064 42585
rect 8024 42576 8076 42628
rect 9496 42687 9548 42696
rect 9496 42653 9527 42687
rect 9527 42653 9548 42687
rect 9496 42644 9548 42653
rect 9956 42712 10008 42764
rect 10140 42644 10192 42696
rect 10324 42687 10376 42696
rect 10324 42653 10333 42687
rect 10333 42653 10367 42687
rect 10367 42653 10376 42687
rect 10324 42644 10376 42653
rect 12624 42712 12676 42764
rect 10876 42644 10928 42696
rect 11336 42687 11388 42696
rect 11336 42653 11345 42687
rect 11345 42653 11379 42687
rect 11379 42653 11388 42687
rect 11336 42644 11388 42653
rect 11888 42644 11940 42696
rect 12072 42687 12124 42696
rect 12072 42653 12081 42687
rect 12081 42653 12115 42687
rect 12115 42653 12124 42687
rect 12072 42644 12124 42653
rect 12532 42687 12584 42696
rect 12532 42653 12541 42687
rect 12541 42653 12575 42687
rect 12575 42653 12584 42687
rect 12532 42644 12584 42653
rect 12808 42687 12860 42696
rect 12808 42653 12817 42687
rect 12817 42653 12851 42687
rect 12851 42653 12860 42687
rect 12808 42644 12860 42653
rect 14924 42712 14976 42764
rect 13176 42687 13228 42696
rect 13176 42653 13185 42687
rect 13185 42653 13219 42687
rect 13219 42653 13228 42687
rect 13176 42644 13228 42653
rect 13636 42644 13688 42696
rect 15384 42687 15436 42696
rect 15384 42653 15393 42687
rect 15393 42653 15427 42687
rect 15427 42653 15436 42687
rect 15384 42644 15436 42653
rect 15476 42644 15528 42696
rect 9128 42551 9180 42560
rect 9128 42517 9137 42551
rect 9137 42517 9171 42551
rect 9171 42517 9180 42551
rect 9128 42508 9180 42517
rect 9680 42551 9732 42560
rect 9680 42517 9689 42551
rect 9689 42517 9723 42551
rect 9723 42517 9732 42551
rect 9680 42508 9732 42517
rect 10140 42551 10192 42560
rect 10140 42517 10149 42551
rect 10149 42517 10183 42551
rect 10183 42517 10192 42551
rect 10140 42508 10192 42517
rect 11152 42508 11204 42560
rect 11428 42508 11480 42560
rect 11520 42551 11572 42560
rect 11520 42517 11529 42551
rect 11529 42517 11563 42551
rect 11563 42517 11572 42551
rect 11520 42508 11572 42517
rect 11796 42551 11848 42560
rect 11796 42517 11805 42551
rect 11805 42517 11839 42551
rect 11839 42517 11848 42551
rect 11796 42508 11848 42517
rect 12256 42576 12308 42628
rect 12348 42551 12400 42560
rect 12348 42517 12357 42551
rect 12357 42517 12391 42551
rect 12391 42517 12400 42551
rect 12348 42508 12400 42517
rect 12624 42551 12676 42560
rect 12624 42517 12633 42551
rect 12633 42517 12667 42551
rect 12667 42517 12676 42551
rect 12624 42508 12676 42517
rect 16488 42891 16540 42900
rect 16488 42857 16497 42891
rect 16497 42857 16531 42891
rect 16531 42857 16540 42891
rect 16488 42848 16540 42857
rect 17960 42848 18012 42900
rect 19984 42848 20036 42900
rect 17500 42780 17552 42832
rect 19524 42780 19576 42832
rect 16764 42712 16816 42764
rect 17316 42712 17368 42764
rect 17868 42712 17920 42764
rect 19064 42712 19116 42764
rect 16212 42687 16264 42696
rect 16212 42653 16221 42687
rect 16221 42653 16255 42687
rect 16255 42653 16264 42687
rect 16212 42644 16264 42653
rect 16856 42644 16908 42696
rect 13544 42551 13596 42560
rect 13544 42517 13553 42551
rect 13553 42517 13587 42551
rect 13587 42517 13596 42551
rect 13544 42508 13596 42517
rect 14004 42508 14056 42560
rect 14648 42551 14700 42560
rect 14648 42517 14657 42551
rect 14657 42517 14691 42551
rect 14691 42517 14700 42551
rect 14648 42508 14700 42517
rect 14924 42551 14976 42560
rect 14924 42517 14933 42551
rect 14933 42517 14967 42551
rect 14967 42517 14976 42551
rect 14924 42508 14976 42517
rect 15016 42508 15068 42560
rect 15476 42551 15528 42560
rect 15476 42517 15485 42551
rect 15485 42517 15519 42551
rect 15519 42517 15528 42551
rect 15476 42508 15528 42517
rect 16396 42619 16448 42628
rect 16396 42585 16405 42619
rect 16405 42585 16439 42619
rect 16439 42585 16448 42619
rect 16396 42576 16448 42585
rect 16948 42619 17000 42628
rect 16948 42585 16957 42619
rect 16957 42585 16991 42619
rect 16991 42585 17000 42619
rect 16948 42576 17000 42585
rect 17500 42619 17552 42628
rect 17500 42585 17509 42619
rect 17509 42585 17543 42619
rect 17543 42585 17552 42619
rect 17500 42576 17552 42585
rect 18880 42576 18932 42628
rect 19892 42576 19944 42628
rect 16120 42508 16172 42560
rect 16212 42508 16264 42560
rect 17776 42508 17828 42560
rect 18328 42551 18380 42560
rect 18328 42517 18337 42551
rect 18337 42517 18371 42551
rect 18371 42517 18380 42551
rect 18328 42508 18380 42517
rect 18696 42508 18748 42560
rect 5894 42406 5946 42458
rect 5958 42406 6010 42458
rect 6022 42406 6074 42458
rect 6086 42406 6138 42458
rect 6150 42406 6202 42458
rect 10839 42406 10891 42458
rect 10903 42406 10955 42458
rect 10967 42406 11019 42458
rect 11031 42406 11083 42458
rect 11095 42406 11147 42458
rect 15784 42406 15836 42458
rect 15848 42406 15900 42458
rect 15912 42406 15964 42458
rect 15976 42406 16028 42458
rect 16040 42406 16092 42458
rect 20729 42406 20781 42458
rect 20793 42406 20845 42458
rect 20857 42406 20909 42458
rect 20921 42406 20973 42458
rect 20985 42406 21037 42458
rect 1492 42304 1544 42356
rect 2504 42304 2556 42356
rect 2596 42347 2648 42356
rect 2596 42313 2605 42347
rect 2605 42313 2639 42347
rect 2639 42313 2648 42347
rect 2596 42304 2648 42313
rect 4068 42304 4120 42356
rect 4804 42304 4856 42356
rect 5172 42304 5224 42356
rect 5724 42304 5776 42356
rect 3608 42236 3660 42288
rect 940 42168 992 42220
rect 3240 42168 3292 42220
rect 3332 42211 3384 42220
rect 3332 42177 3341 42211
rect 3341 42177 3375 42211
rect 3375 42177 3384 42211
rect 3332 42168 3384 42177
rect 4344 42236 4396 42288
rect 6828 42304 6880 42356
rect 7564 42304 7616 42356
rect 8024 42304 8076 42356
rect 8116 42304 8168 42356
rect 8944 42347 8996 42356
rect 8944 42313 8953 42347
rect 8953 42313 8987 42347
rect 8987 42313 8996 42347
rect 8944 42304 8996 42313
rect 1676 42100 1728 42152
rect 2872 42100 2924 42152
rect 4896 42211 4948 42220
rect 4896 42177 4905 42211
rect 4905 42177 4939 42211
rect 4939 42177 4948 42211
rect 4896 42168 4948 42177
rect 5540 42211 5592 42220
rect 5540 42177 5549 42211
rect 5549 42177 5583 42211
rect 5583 42177 5592 42211
rect 5540 42168 5592 42177
rect 848 42032 900 42084
rect 3700 42075 3752 42084
rect 3700 42041 3709 42075
rect 3709 42041 3743 42075
rect 3743 42041 3752 42075
rect 3700 42032 3752 42041
rect 4068 42100 4120 42152
rect 4528 42100 4580 42152
rect 3976 42032 4028 42084
rect 9588 42304 9640 42356
rect 9772 42236 9824 42288
rect 6276 42168 6328 42220
rect 7104 42211 7156 42220
rect 7104 42177 7113 42211
rect 7113 42177 7147 42211
rect 7147 42177 7156 42211
rect 7104 42168 7156 42177
rect 8208 42211 8260 42220
rect 8208 42177 8217 42211
rect 8217 42177 8251 42211
rect 8251 42177 8260 42211
rect 8208 42168 8260 42177
rect 8852 42211 8904 42220
rect 8852 42177 8861 42211
rect 8861 42177 8895 42211
rect 8895 42177 8904 42211
rect 8852 42168 8904 42177
rect 8944 42168 8996 42220
rect 6920 42100 6972 42152
rect 7748 42100 7800 42152
rect 9496 42168 9548 42220
rect 10048 42211 10100 42220
rect 10048 42177 10057 42211
rect 10057 42177 10091 42211
rect 10091 42177 10100 42211
rect 10048 42168 10100 42177
rect 10600 42211 10652 42220
rect 10600 42177 10609 42211
rect 10609 42177 10643 42211
rect 10643 42177 10652 42211
rect 10600 42168 10652 42177
rect 12348 42304 12400 42356
rect 13452 42304 13504 42356
rect 13544 42304 13596 42356
rect 11612 42236 11664 42288
rect 11336 42211 11388 42220
rect 11336 42177 11345 42211
rect 11345 42177 11379 42211
rect 11379 42177 11388 42211
rect 11336 42168 11388 42177
rect 12348 42211 12400 42220
rect 12348 42177 12357 42211
rect 12357 42177 12391 42211
rect 12391 42177 12400 42211
rect 12348 42168 12400 42177
rect 13728 42304 13780 42356
rect 14648 42304 14700 42356
rect 5172 41964 5224 42016
rect 7012 42032 7064 42084
rect 13636 42100 13688 42152
rect 14464 42211 14516 42220
rect 14464 42177 14473 42211
rect 14473 42177 14507 42211
rect 14507 42177 14516 42211
rect 14464 42168 14516 42177
rect 14648 42168 14700 42220
rect 15292 42304 15344 42356
rect 15476 42304 15528 42356
rect 16120 42304 16172 42356
rect 16212 42304 16264 42356
rect 14924 42168 14976 42220
rect 16488 42236 16540 42288
rect 18972 42304 19024 42356
rect 21180 42304 21232 42356
rect 16304 42168 16356 42220
rect 16580 42168 16632 42220
rect 17132 42211 17184 42220
rect 17132 42177 17141 42211
rect 17141 42177 17175 42211
rect 17175 42177 17184 42211
rect 17132 42168 17184 42177
rect 17316 42168 17368 42220
rect 18236 42279 18288 42288
rect 18236 42245 18245 42279
rect 18245 42245 18279 42279
rect 18279 42245 18288 42279
rect 18236 42236 18288 42245
rect 18604 42279 18656 42288
rect 18604 42245 18613 42279
rect 18613 42245 18647 42279
rect 18647 42245 18656 42279
rect 18604 42236 18656 42245
rect 10324 42032 10376 42084
rect 9496 42007 9548 42016
rect 9496 41973 9505 42007
rect 9505 41973 9539 42007
rect 9539 41973 9548 42007
rect 9496 41964 9548 41973
rect 9772 41964 9824 42016
rect 10416 42007 10468 42016
rect 10416 41973 10425 42007
rect 10425 41973 10459 42007
rect 10459 41973 10468 42007
rect 10416 41964 10468 41973
rect 17868 42100 17920 42152
rect 19616 42168 19668 42220
rect 20628 42168 20680 42220
rect 19156 42100 19208 42152
rect 12164 42007 12216 42016
rect 12164 41973 12173 42007
rect 12173 41973 12207 42007
rect 12207 41973 12216 42007
rect 12164 41964 12216 41973
rect 13176 42007 13228 42016
rect 13176 41973 13185 42007
rect 13185 41973 13219 42007
rect 13219 41973 13228 42007
rect 13176 41964 13228 41973
rect 13268 41964 13320 42016
rect 13912 42007 13964 42016
rect 13912 41973 13921 42007
rect 13921 41973 13955 42007
rect 13955 41973 13964 42007
rect 13912 41964 13964 41973
rect 14280 42007 14332 42016
rect 14280 41973 14289 42007
rect 14289 41973 14323 42007
rect 14323 41973 14332 42007
rect 14280 41964 14332 41973
rect 14372 41964 14424 42016
rect 14832 41964 14884 42016
rect 15292 41964 15344 42016
rect 15384 42007 15436 42016
rect 15384 41973 15393 42007
rect 15393 41973 15427 42007
rect 15427 41973 15436 42007
rect 15384 41964 15436 41973
rect 15476 41964 15528 42016
rect 15844 41964 15896 42016
rect 19340 42007 19392 42016
rect 19340 41973 19349 42007
rect 19349 41973 19383 42007
rect 19383 41973 19392 42007
rect 19340 41964 19392 41973
rect 19892 41964 19944 42016
rect 3422 41862 3474 41914
rect 3486 41862 3538 41914
rect 3550 41862 3602 41914
rect 3614 41862 3666 41914
rect 3678 41862 3730 41914
rect 8367 41862 8419 41914
rect 8431 41862 8483 41914
rect 8495 41862 8547 41914
rect 8559 41862 8611 41914
rect 8623 41862 8675 41914
rect 13312 41862 13364 41914
rect 13376 41862 13428 41914
rect 13440 41862 13492 41914
rect 13504 41862 13556 41914
rect 13568 41862 13620 41914
rect 18257 41862 18309 41914
rect 18321 41862 18373 41914
rect 18385 41862 18437 41914
rect 18449 41862 18501 41914
rect 18513 41862 18565 41914
rect 2136 41760 2188 41812
rect 2688 41760 2740 41812
rect 3056 41760 3108 41812
rect 3148 41803 3200 41812
rect 3148 41769 3157 41803
rect 3157 41769 3191 41803
rect 3191 41769 3200 41803
rect 3148 41760 3200 41769
rect 3240 41760 3292 41812
rect 2964 41692 3016 41744
rect 3976 41760 4028 41812
rect 4160 41803 4212 41812
rect 4160 41769 4169 41803
rect 4169 41769 4203 41803
rect 4203 41769 4212 41803
rect 4160 41760 4212 41769
rect 4252 41760 4304 41812
rect 5540 41760 5592 41812
rect 6644 41760 6696 41812
rect 7012 41760 7064 41812
rect 7104 41760 7156 41812
rect 8208 41760 8260 41812
rect 20 41624 72 41676
rect 5448 41692 5500 41744
rect 2504 41599 2556 41608
rect 2504 41565 2513 41599
rect 2513 41565 2547 41599
rect 2547 41565 2556 41599
rect 2504 41556 2556 41565
rect 2044 41488 2096 41540
rect 3056 41599 3108 41608
rect 3056 41565 3065 41599
rect 3065 41565 3099 41599
rect 3099 41565 3108 41599
rect 3056 41556 3108 41565
rect 3884 41556 3936 41608
rect 4712 41556 4764 41608
rect 5080 41556 5132 41608
rect 5172 41599 5224 41608
rect 5172 41565 5181 41599
rect 5181 41565 5215 41599
rect 5215 41565 5224 41599
rect 5172 41556 5224 41565
rect 5448 41599 5500 41608
rect 5448 41565 5457 41599
rect 5457 41565 5491 41599
rect 5491 41565 5500 41599
rect 5448 41556 5500 41565
rect 5540 41556 5592 41608
rect 480 41420 532 41472
rect 5172 41420 5224 41472
rect 5540 41463 5592 41472
rect 5540 41429 5549 41463
rect 5549 41429 5583 41463
rect 5583 41429 5592 41463
rect 5540 41420 5592 41429
rect 5632 41420 5684 41472
rect 7196 41692 7248 41744
rect 7196 41599 7248 41608
rect 7196 41565 7205 41599
rect 7205 41565 7239 41599
rect 7239 41565 7248 41599
rect 7196 41556 7248 41565
rect 7748 41599 7800 41608
rect 7748 41565 7757 41599
rect 7757 41565 7791 41599
rect 7791 41565 7800 41599
rect 7748 41556 7800 41565
rect 9496 41760 9548 41812
rect 8760 41692 8812 41744
rect 8760 41599 8812 41608
rect 8760 41565 8769 41599
rect 8769 41565 8803 41599
rect 8803 41565 8812 41599
rect 8760 41556 8812 41565
rect 9128 41599 9180 41608
rect 9128 41565 9137 41599
rect 9137 41565 9171 41599
rect 9171 41565 9180 41599
rect 9128 41556 9180 41565
rect 12624 41760 12676 41812
rect 14096 41760 14148 41812
rect 15016 41760 15068 41812
rect 12440 41692 12492 41744
rect 13820 41692 13872 41744
rect 13544 41556 13596 41608
rect 13636 41599 13688 41608
rect 13636 41565 13645 41599
rect 13645 41565 13679 41599
rect 13679 41565 13688 41599
rect 13636 41556 13688 41565
rect 14188 41692 14240 41744
rect 14924 41692 14976 41744
rect 18788 41760 18840 41812
rect 19432 41760 19484 41812
rect 15752 41692 15804 41744
rect 16580 41692 16632 41744
rect 17224 41692 17276 41744
rect 18236 41692 18288 41744
rect 9956 41488 10008 41540
rect 10232 41488 10284 41540
rect 11704 41488 11756 41540
rect 12348 41488 12400 41540
rect 12808 41488 12860 41540
rect 7012 41463 7064 41472
rect 7012 41429 7021 41463
rect 7021 41429 7055 41463
rect 7055 41429 7064 41463
rect 7012 41420 7064 41429
rect 14464 41420 14516 41472
rect 14832 41463 14884 41472
rect 14832 41429 14841 41463
rect 14841 41429 14875 41463
rect 14875 41429 14884 41463
rect 14832 41420 14884 41429
rect 15660 41556 15712 41608
rect 15936 41556 15988 41608
rect 16304 41556 16356 41608
rect 16396 41599 16448 41608
rect 16396 41565 16405 41599
rect 16405 41565 16439 41599
rect 16439 41565 16448 41599
rect 16396 41556 16448 41565
rect 16488 41556 16540 41608
rect 16764 41599 16816 41608
rect 16764 41565 16773 41599
rect 16773 41565 16807 41599
rect 16807 41565 16816 41599
rect 16764 41556 16816 41565
rect 16948 41556 17000 41608
rect 17224 41556 17276 41608
rect 17592 41599 17644 41608
rect 17592 41565 17601 41599
rect 17601 41565 17635 41599
rect 17635 41565 17644 41599
rect 17592 41556 17644 41565
rect 17684 41556 17736 41608
rect 18052 41556 18104 41608
rect 21272 41624 21324 41676
rect 20444 41556 20496 41608
rect 16028 41420 16080 41472
rect 18144 41531 18196 41540
rect 18144 41497 18153 41531
rect 18153 41497 18187 41531
rect 18187 41497 18196 41531
rect 18144 41488 18196 41497
rect 18788 41488 18840 41540
rect 19432 41531 19484 41540
rect 19432 41497 19441 41531
rect 19441 41497 19475 41531
rect 19475 41497 19484 41531
rect 19432 41488 19484 41497
rect 16856 41463 16908 41472
rect 16856 41429 16865 41463
rect 16865 41429 16899 41463
rect 16899 41429 16908 41463
rect 16856 41420 16908 41429
rect 17408 41463 17460 41472
rect 17408 41429 17417 41463
rect 17417 41429 17451 41463
rect 17451 41429 17460 41463
rect 17408 41420 17460 41429
rect 17960 41420 18012 41472
rect 19064 41420 19116 41472
rect 19340 41420 19392 41472
rect 20536 41531 20588 41540
rect 20536 41497 20545 41531
rect 20545 41497 20579 41531
rect 20579 41497 20588 41531
rect 20536 41488 20588 41497
rect 5894 41318 5946 41370
rect 5958 41318 6010 41370
rect 6022 41318 6074 41370
rect 6086 41318 6138 41370
rect 6150 41318 6202 41370
rect 10839 41318 10891 41370
rect 10903 41318 10955 41370
rect 10967 41318 11019 41370
rect 11031 41318 11083 41370
rect 11095 41318 11147 41370
rect 15784 41318 15836 41370
rect 15848 41318 15900 41370
rect 15912 41318 15964 41370
rect 15976 41318 16028 41370
rect 16040 41318 16092 41370
rect 20729 41318 20781 41370
rect 20793 41318 20845 41370
rect 20857 41318 20909 41370
rect 20921 41318 20973 41370
rect 20985 41318 21037 41370
rect 3332 41216 3384 41268
rect 3792 41216 3844 41268
rect 3976 41259 4028 41268
rect 3976 41225 3985 41259
rect 3985 41225 4019 41259
rect 4019 41225 4028 41259
rect 3976 41216 4028 41225
rect 4896 41216 4948 41268
rect 4988 41216 5040 41268
rect 5264 41216 5316 41268
rect 5816 41259 5868 41268
rect 5816 41225 5825 41259
rect 5825 41225 5859 41259
rect 5859 41225 5868 41259
rect 5816 41216 5868 41225
rect 6552 41259 6604 41268
rect 6552 41225 6561 41259
rect 6561 41225 6595 41259
rect 6595 41225 6604 41259
rect 6552 41216 6604 41225
rect 6736 41216 6788 41268
rect 7380 41216 7432 41268
rect 14372 41259 14424 41268
rect 14372 41225 14381 41259
rect 14381 41225 14415 41259
rect 14415 41225 14424 41259
rect 14372 41216 14424 41225
rect 14556 41216 14608 41268
rect 14648 41259 14700 41268
rect 14648 41225 14657 41259
rect 14657 41225 14691 41259
rect 14691 41225 14700 41259
rect 14648 41216 14700 41225
rect 14740 41216 14792 41268
rect 1952 41148 2004 41200
rect 2688 41148 2740 41200
rect 2780 41080 2832 41132
rect 3608 41123 3660 41132
rect 3608 41089 3617 41123
rect 3617 41089 3651 41123
rect 3651 41089 3660 41123
rect 3608 41080 3660 41089
rect 4068 41080 4120 41132
rect 4344 41080 4396 41132
rect 4436 41123 4488 41132
rect 4436 41089 4445 41123
rect 4445 41089 4479 41123
rect 4479 41089 4488 41123
rect 4436 41080 4488 41089
rect 4988 41123 5040 41132
rect 4988 41089 4997 41123
rect 4997 41089 5031 41123
rect 5031 41089 5040 41123
rect 4988 41080 5040 41089
rect 5080 41080 5132 41132
rect 5356 41012 5408 41064
rect 6920 41148 6972 41200
rect 15016 41216 15068 41268
rect 15200 41259 15252 41268
rect 15200 41225 15209 41259
rect 15209 41225 15243 41259
rect 15243 41225 15252 41259
rect 15200 41216 15252 41225
rect 15568 41216 15620 41268
rect 16396 41216 16448 41268
rect 16948 41216 17000 41268
rect 6276 41012 6328 41064
rect 2136 40876 2188 40928
rect 5724 40876 5776 40928
rect 7196 40944 7248 40996
rect 7932 41123 7984 41132
rect 7932 41089 7941 41123
rect 7941 41089 7975 41123
rect 7975 41089 7984 41123
rect 7932 41080 7984 41089
rect 8760 41012 8812 41064
rect 14556 41123 14608 41132
rect 14556 41089 14565 41123
rect 14565 41089 14599 41123
rect 14599 41089 14608 41123
rect 14556 41080 14608 41089
rect 16764 41148 16816 41200
rect 17224 41216 17276 41268
rect 17500 41216 17552 41268
rect 18236 41216 18288 41268
rect 19248 41216 19300 41268
rect 15384 41123 15436 41132
rect 15384 41089 15393 41123
rect 15393 41089 15427 41123
rect 15427 41089 15436 41123
rect 15384 41080 15436 41089
rect 15568 41080 15620 41132
rect 15476 41012 15528 41064
rect 16212 41080 16264 41132
rect 16304 41123 16356 41132
rect 16304 41089 16313 41123
rect 16313 41089 16347 41123
rect 16347 41089 16356 41123
rect 16304 41080 16356 41089
rect 16672 41080 16724 41132
rect 16856 41123 16908 41132
rect 16856 41089 16865 41123
rect 16865 41089 16899 41123
rect 16899 41089 16908 41123
rect 16856 41080 16908 41089
rect 16948 41080 17000 41132
rect 17408 41148 17460 41200
rect 17224 41123 17276 41132
rect 17224 41089 17233 41123
rect 17233 41089 17267 41123
rect 17267 41089 17276 41123
rect 17224 41080 17276 41089
rect 17500 41123 17552 41132
rect 17500 41089 17509 41123
rect 17509 41089 17543 41123
rect 17543 41089 17552 41123
rect 17500 41080 17552 41089
rect 12808 40944 12860 40996
rect 17040 41012 17092 41064
rect 18236 41123 18288 41132
rect 18236 41089 18245 41123
rect 18245 41089 18279 41123
rect 18279 41089 18288 41123
rect 18236 41080 18288 41089
rect 18972 41080 19024 41132
rect 19064 41123 19116 41132
rect 19064 41089 19073 41123
rect 19073 41089 19107 41123
rect 19107 41089 19116 41123
rect 19064 41080 19116 41089
rect 21088 41080 21140 41132
rect 16764 40944 16816 40996
rect 17592 40944 17644 40996
rect 14924 40876 14976 40928
rect 15384 40876 15436 40928
rect 16396 40876 16448 40928
rect 16488 40876 16540 40928
rect 17776 40944 17828 40996
rect 19156 41012 19208 41064
rect 17868 40876 17920 40928
rect 18052 40919 18104 40928
rect 18052 40885 18061 40919
rect 18061 40885 18095 40919
rect 18095 40885 18104 40919
rect 18052 40876 18104 40885
rect 20168 40876 20220 40928
rect 3422 40774 3474 40826
rect 3486 40774 3538 40826
rect 3550 40774 3602 40826
rect 3614 40774 3666 40826
rect 3678 40774 3730 40826
rect 8367 40774 8419 40826
rect 8431 40774 8483 40826
rect 8495 40774 8547 40826
rect 8559 40774 8611 40826
rect 8623 40774 8675 40826
rect 13312 40774 13364 40826
rect 13376 40774 13428 40826
rect 13440 40774 13492 40826
rect 13504 40774 13556 40826
rect 13568 40774 13620 40826
rect 18257 40774 18309 40826
rect 18321 40774 18373 40826
rect 18385 40774 18437 40826
rect 18449 40774 18501 40826
rect 18513 40774 18565 40826
rect 756 40536 808 40588
rect 5632 40672 5684 40724
rect 5264 40604 5316 40656
rect 13084 40672 13136 40724
rect 15200 40715 15252 40724
rect 15200 40681 15209 40715
rect 15209 40681 15243 40715
rect 15243 40681 15252 40715
rect 15200 40672 15252 40681
rect 15476 40715 15528 40724
rect 15476 40681 15485 40715
rect 15485 40681 15519 40715
rect 15519 40681 15528 40715
rect 15476 40672 15528 40681
rect 15660 40672 15712 40724
rect 16212 40715 16264 40724
rect 16212 40681 16221 40715
rect 16221 40681 16255 40715
rect 16255 40681 16264 40715
rect 16212 40672 16264 40681
rect 16764 40672 16816 40724
rect 17224 40672 17276 40724
rect 19432 40672 19484 40724
rect 19524 40715 19576 40724
rect 19524 40681 19533 40715
rect 19533 40681 19567 40715
rect 19567 40681 19576 40715
rect 19524 40672 19576 40681
rect 17040 40604 17092 40656
rect 4068 40536 4120 40588
rect 7564 40536 7616 40588
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 13544 40468 13596 40520
rect 13636 40468 13688 40520
rect 15384 40511 15436 40520
rect 15384 40477 15393 40511
rect 15393 40477 15427 40511
rect 15427 40477 15436 40511
rect 15384 40468 15436 40477
rect 15660 40511 15712 40520
rect 15660 40477 15669 40511
rect 15669 40477 15703 40511
rect 15703 40477 15712 40511
rect 15660 40468 15712 40477
rect 1952 40443 2004 40452
rect 1952 40409 1961 40443
rect 1961 40409 1995 40443
rect 1995 40409 2004 40443
rect 1952 40400 2004 40409
rect 2688 40443 2740 40452
rect 2688 40409 2697 40443
rect 2697 40409 2731 40443
rect 2731 40409 2740 40443
rect 2688 40400 2740 40409
rect 7656 40332 7708 40384
rect 12440 40332 12492 40384
rect 14924 40375 14976 40384
rect 14924 40341 14933 40375
rect 14933 40341 14967 40375
rect 14967 40341 14976 40375
rect 14924 40332 14976 40341
rect 15292 40400 15344 40452
rect 16120 40468 16172 40520
rect 16764 40468 16816 40520
rect 16488 40400 16540 40452
rect 17408 40468 17460 40520
rect 16212 40332 16264 40384
rect 16948 40332 17000 40384
rect 17040 40332 17092 40384
rect 17776 40511 17828 40520
rect 17776 40477 17785 40511
rect 17785 40477 17819 40511
rect 17819 40477 17828 40511
rect 17776 40468 17828 40477
rect 18144 40468 18196 40520
rect 17776 40332 17828 40384
rect 18420 40332 18472 40384
rect 19064 40511 19116 40520
rect 19064 40477 19073 40511
rect 19073 40477 19107 40511
rect 19107 40477 19116 40511
rect 19064 40468 19116 40477
rect 19432 40511 19484 40520
rect 19432 40477 19441 40511
rect 19441 40477 19475 40511
rect 19475 40477 19484 40511
rect 19432 40468 19484 40477
rect 19800 40536 19852 40588
rect 19984 40511 20036 40520
rect 19984 40477 19993 40511
rect 19993 40477 20027 40511
rect 20027 40477 20036 40511
rect 19984 40468 20036 40477
rect 20352 40400 20404 40452
rect 21272 40400 21324 40452
rect 19800 40375 19852 40384
rect 19800 40341 19809 40375
rect 19809 40341 19843 40375
rect 19843 40341 19852 40375
rect 19800 40332 19852 40341
rect 5894 40230 5946 40282
rect 5958 40230 6010 40282
rect 6022 40230 6074 40282
rect 6086 40230 6138 40282
rect 6150 40230 6202 40282
rect 10839 40230 10891 40282
rect 10903 40230 10955 40282
rect 10967 40230 11019 40282
rect 11031 40230 11083 40282
rect 11095 40230 11147 40282
rect 15784 40230 15836 40282
rect 15848 40230 15900 40282
rect 15912 40230 15964 40282
rect 15976 40230 16028 40282
rect 16040 40230 16092 40282
rect 20729 40230 20781 40282
rect 20793 40230 20845 40282
rect 20857 40230 20909 40282
rect 20921 40230 20973 40282
rect 20985 40230 21037 40282
rect 7656 40128 7708 40180
rect 1308 40060 1360 40112
rect 2688 40060 2740 40112
rect 1308 39924 1360 39976
rect 2044 39924 2096 39976
rect 3056 40035 3108 40044
rect 3056 40001 3065 40035
rect 3065 40001 3099 40035
rect 3099 40001 3108 40035
rect 3056 39992 3108 40001
rect 4896 39992 4948 40044
rect 4068 39924 4120 39976
rect 7840 40002 7892 40054
rect 15568 40128 15620 40180
rect 16120 40171 16172 40180
rect 16120 40137 16129 40171
rect 16129 40137 16163 40171
rect 16163 40137 16172 40171
rect 16120 40128 16172 40137
rect 16672 40128 16724 40180
rect 17316 40128 17368 40180
rect 17684 40128 17736 40180
rect 19064 40128 19116 40180
rect 19800 40128 19852 40180
rect 11336 39992 11388 40044
rect 16948 40060 17000 40112
rect 12808 39992 12860 40044
rect 14188 39992 14240 40044
rect 14648 40035 14700 40044
rect 14648 40001 14657 40035
rect 14657 40001 14691 40035
rect 14691 40001 14700 40035
rect 14648 39992 14700 40001
rect 18052 40060 18104 40112
rect 18236 40060 18288 40112
rect 20260 40128 20312 40180
rect 17592 40035 17644 40044
rect 17592 40001 17601 40035
rect 17601 40001 17635 40035
rect 17635 40001 17644 40035
rect 17592 39992 17644 40001
rect 17868 40035 17920 40044
rect 17868 40001 17877 40035
rect 17877 40001 17911 40035
rect 17911 40001 17920 40035
rect 17868 39992 17920 40001
rect 18328 39992 18380 40044
rect 18880 39992 18932 40044
rect 19248 39992 19300 40044
rect 19340 39992 19392 40044
rect 19892 39992 19944 40044
rect 20260 39992 20312 40044
rect 3792 39788 3844 39840
rect 11428 39924 11480 39976
rect 16488 39924 16540 39976
rect 16580 39924 16632 39976
rect 16672 39924 16724 39976
rect 18052 39856 18104 39908
rect 5448 39788 5500 39840
rect 5540 39831 5592 39840
rect 5540 39797 5549 39831
rect 5549 39797 5583 39831
rect 5583 39797 5592 39831
rect 5540 39788 5592 39797
rect 7564 39788 7616 39840
rect 7932 39788 7984 39840
rect 14924 39788 14976 39840
rect 18144 39788 18196 39840
rect 18696 39788 18748 39840
rect 18880 39831 18932 39840
rect 18880 39797 18889 39831
rect 18889 39797 18923 39831
rect 18923 39797 18932 39831
rect 18880 39788 18932 39797
rect 19064 39788 19116 39840
rect 19524 39831 19576 39840
rect 19524 39797 19533 39831
rect 19533 39797 19567 39831
rect 19567 39797 19576 39831
rect 19524 39788 19576 39797
rect 19800 39831 19852 39840
rect 19800 39797 19809 39831
rect 19809 39797 19843 39831
rect 19843 39797 19852 39831
rect 19800 39788 19852 39797
rect 20996 39788 21048 39840
rect 3422 39686 3474 39738
rect 3486 39686 3538 39738
rect 3550 39686 3602 39738
rect 3614 39686 3666 39738
rect 3678 39686 3730 39738
rect 8367 39686 8419 39738
rect 8431 39686 8483 39738
rect 8495 39686 8547 39738
rect 8559 39686 8611 39738
rect 8623 39686 8675 39738
rect 13312 39686 13364 39738
rect 13376 39686 13428 39738
rect 13440 39686 13492 39738
rect 13504 39686 13556 39738
rect 13568 39686 13620 39738
rect 18257 39686 18309 39738
rect 18321 39686 18373 39738
rect 18385 39686 18437 39738
rect 18449 39686 18501 39738
rect 18513 39686 18565 39738
rect 1400 39423 1452 39432
rect 1400 39389 1409 39423
rect 1409 39389 1443 39423
rect 1443 39389 1452 39423
rect 1400 39380 1452 39389
rect 2136 39380 2188 39432
rect 3792 39516 3844 39568
rect 4068 39423 4120 39432
rect 4068 39389 4075 39423
rect 4075 39389 4109 39423
rect 4109 39389 4120 39423
rect 4068 39380 4120 39389
rect 7564 39584 7616 39636
rect 13728 39584 13780 39636
rect 15660 39584 15712 39636
rect 7380 39559 7432 39568
rect 7380 39525 7389 39559
rect 7389 39525 7423 39559
rect 7423 39525 7432 39559
rect 7380 39516 7432 39525
rect 17592 39584 17644 39636
rect 17684 39584 17736 39636
rect 17868 39584 17920 39636
rect 17960 39584 18012 39636
rect 19340 39584 19392 39636
rect 19432 39584 19484 39636
rect 20168 39584 20220 39636
rect 16212 39559 16264 39568
rect 16212 39525 16221 39559
rect 16221 39525 16255 39559
rect 16255 39525 16264 39559
rect 16212 39516 16264 39525
rect 16580 39516 16632 39568
rect 18512 39516 18564 39568
rect 12624 39448 12676 39500
rect 17592 39448 17644 39500
rect 6644 39423 6696 39432
rect 6644 39389 6651 39423
rect 6651 39389 6685 39423
rect 6685 39389 6696 39423
rect 6644 39380 6696 39389
rect 11428 39380 11480 39432
rect 9588 39312 9640 39364
rect 15292 39380 15344 39432
rect 15476 39423 15528 39432
rect 15476 39389 15485 39423
rect 15485 39389 15519 39423
rect 15519 39389 15528 39423
rect 15476 39380 15528 39389
rect 16856 39423 16908 39432
rect 16856 39389 16865 39423
rect 16865 39389 16899 39423
rect 16899 39389 16908 39423
rect 16856 39380 16908 39389
rect 17132 39423 17184 39432
rect 17132 39389 17141 39423
rect 17141 39389 17175 39423
rect 17175 39389 17184 39423
rect 17132 39380 17184 39389
rect 17408 39423 17460 39432
rect 17408 39389 17417 39423
rect 17417 39389 17451 39423
rect 17451 39389 17460 39423
rect 17408 39380 17460 39389
rect 18236 39423 18288 39432
rect 18236 39389 18245 39423
rect 18245 39389 18279 39423
rect 18279 39389 18288 39423
rect 18236 39380 18288 39389
rect 18052 39312 18104 39364
rect 18144 39312 18196 39364
rect 18328 39312 18380 39364
rect 19248 39380 19300 39432
rect 19432 39380 19484 39432
rect 19708 39380 19760 39432
rect 3792 39244 3844 39296
rect 4712 39244 4764 39296
rect 5448 39244 5500 39296
rect 16856 39244 16908 39296
rect 17316 39244 17368 39296
rect 18788 39244 18840 39296
rect 18972 39244 19024 39296
rect 21272 39312 21324 39364
rect 19984 39244 20036 39296
rect 5894 39142 5946 39194
rect 5958 39142 6010 39194
rect 6022 39142 6074 39194
rect 6086 39142 6138 39194
rect 6150 39142 6202 39194
rect 10839 39142 10891 39194
rect 10903 39142 10955 39194
rect 10967 39142 11019 39194
rect 11031 39142 11083 39194
rect 11095 39142 11147 39194
rect 15784 39142 15836 39194
rect 15848 39142 15900 39194
rect 15912 39142 15964 39194
rect 15976 39142 16028 39194
rect 16040 39142 16092 39194
rect 20729 39142 20781 39194
rect 20793 39142 20845 39194
rect 20857 39142 20909 39194
rect 20921 39142 20973 39194
rect 20985 39142 21037 39194
rect 11244 39040 11296 39092
rect 14556 39040 14608 39092
rect 16396 39040 16448 39092
rect 1492 38904 1544 38956
rect 1952 38947 2004 38956
rect 1952 38913 1961 38947
rect 1961 38913 1995 38947
rect 1995 38913 2004 38947
rect 1952 38904 2004 38913
rect 4252 38972 4304 39024
rect 4620 38972 4672 39024
rect 4804 39015 4856 39024
rect 4804 38981 4813 39015
rect 4813 38981 4847 39015
rect 4847 38981 4856 39015
rect 4804 38972 4856 38981
rect 5540 38972 5592 39024
rect 17408 39040 17460 39092
rect 18236 39040 18288 39092
rect 18328 39040 18380 39092
rect 18972 39040 19024 39092
rect 5172 38904 5224 38956
rect 5632 38947 5684 38956
rect 5632 38913 5655 38947
rect 5655 38913 5684 38947
rect 5632 38904 5684 38913
rect 7932 38947 7984 38956
rect 7932 38913 7941 38947
rect 7941 38913 7975 38947
rect 7975 38913 7984 38947
rect 7932 38904 7984 38913
rect 12440 38904 12492 38956
rect 13084 38904 13136 38956
rect 15200 38904 15252 38956
rect 16856 38904 16908 38956
rect 17776 38972 17828 39024
rect 18052 38904 18104 38956
rect 18328 38904 18380 38956
rect 18420 38947 18472 38956
rect 18420 38913 18437 38947
rect 18437 38913 18471 38947
rect 18471 38913 18472 38947
rect 18420 38904 18472 38913
rect 19248 39040 19300 39092
rect 19616 39040 19668 39092
rect 19340 38904 19392 38956
rect 2320 38836 2372 38888
rect 3884 38836 3936 38888
rect 4712 38836 4764 38888
rect 6552 38836 6604 38888
rect 6920 38879 6972 38888
rect 6920 38845 6929 38879
rect 6929 38845 6963 38879
rect 6963 38845 6972 38879
rect 6920 38836 6972 38845
rect 7380 38879 7432 38888
rect 7380 38845 7389 38879
rect 7389 38845 7423 38879
rect 7423 38845 7432 38879
rect 7380 38836 7432 38845
rect 4068 38768 4120 38820
rect 7840 38836 7892 38888
rect 14096 38836 14148 38888
rect 14648 38836 14700 38888
rect 20628 39040 20680 39092
rect 20076 38972 20128 39024
rect 19892 38904 19944 38956
rect 18144 38768 18196 38820
rect 20352 38836 20404 38888
rect 18420 38768 18472 38820
rect 19524 38768 19576 38820
rect 4160 38700 4212 38752
rect 5816 38743 5868 38752
rect 5816 38709 5825 38743
rect 5825 38709 5859 38743
rect 5859 38709 5868 38743
rect 5816 38700 5868 38709
rect 13820 38700 13872 38752
rect 19708 38700 19760 38752
rect 20444 38743 20496 38752
rect 20444 38709 20453 38743
rect 20453 38709 20487 38743
rect 20487 38709 20496 38743
rect 20444 38700 20496 38709
rect 3422 38598 3474 38650
rect 3486 38598 3538 38650
rect 3550 38598 3602 38650
rect 3614 38598 3666 38650
rect 3678 38598 3730 38650
rect 8367 38598 8419 38650
rect 8431 38598 8483 38650
rect 8495 38598 8547 38650
rect 8559 38598 8611 38650
rect 8623 38598 8675 38650
rect 13312 38598 13364 38650
rect 13376 38598 13428 38650
rect 13440 38598 13492 38650
rect 13504 38598 13556 38650
rect 13568 38598 13620 38650
rect 18257 38598 18309 38650
rect 18321 38598 18373 38650
rect 18385 38598 18437 38650
rect 18449 38598 18501 38650
rect 18513 38598 18565 38650
rect 7288 38496 7340 38548
rect 9680 38428 9732 38480
rect 1584 38360 1636 38412
rect 2320 38403 2372 38412
rect 2320 38369 2329 38403
rect 2329 38369 2363 38403
rect 2363 38369 2372 38403
rect 2320 38360 2372 38369
rect 3792 38360 3844 38412
rect 5264 38360 5316 38412
rect 6276 38360 6328 38412
rect 10324 38360 10376 38412
rect 15200 38428 15252 38480
rect 1124 38292 1176 38344
rect 2688 38292 2740 38344
rect 4160 38292 4212 38344
rect 1676 38267 1728 38276
rect 1676 38233 1685 38267
rect 1685 38233 1719 38267
rect 1719 38233 1728 38267
rect 1676 38224 1728 38233
rect 4804 38292 4856 38344
rect 4896 38292 4948 38344
rect 5632 38292 5684 38344
rect 9772 38292 9824 38344
rect 10508 38335 10560 38344
rect 10508 38301 10517 38335
rect 10517 38301 10551 38335
rect 10551 38301 10560 38335
rect 10508 38292 10560 38301
rect 10784 38335 10836 38344
rect 10784 38301 10791 38335
rect 10791 38301 10825 38335
rect 10825 38301 10836 38335
rect 10784 38292 10836 38301
rect 4988 38224 5040 38276
rect 5172 38224 5224 38276
rect 9956 38224 10008 38276
rect 12256 38292 12308 38344
rect 13820 38292 13872 38344
rect 12164 38267 12216 38276
rect 12164 38233 12173 38267
rect 12173 38233 12207 38267
rect 12207 38233 12216 38267
rect 12164 38224 12216 38233
rect 12440 38224 12492 38276
rect 14096 38335 14148 38344
rect 14096 38301 14105 38335
rect 14105 38301 14139 38335
rect 14139 38301 14148 38335
rect 14096 38292 14148 38301
rect 16396 38496 16448 38548
rect 18328 38496 18380 38548
rect 19248 38496 19300 38548
rect 19432 38428 19484 38480
rect 19800 38496 19852 38548
rect 19984 38428 20036 38480
rect 3332 38199 3384 38208
rect 3332 38165 3341 38199
rect 3341 38165 3375 38199
rect 3375 38165 3384 38199
rect 3332 38156 3384 38165
rect 4160 38156 4212 38208
rect 4620 38156 4672 38208
rect 4896 38156 4948 38208
rect 5264 38199 5316 38208
rect 5264 38165 5273 38199
rect 5273 38165 5307 38199
rect 5307 38165 5316 38199
rect 5264 38156 5316 38165
rect 9128 38156 9180 38208
rect 10416 38156 10468 38208
rect 10508 38156 10560 38208
rect 10784 38156 10836 38208
rect 11520 38199 11572 38208
rect 11520 38165 11529 38199
rect 11529 38165 11563 38199
rect 11563 38165 11572 38199
rect 11520 38156 11572 38165
rect 13728 38199 13780 38208
rect 13728 38165 13737 38199
rect 13737 38165 13771 38199
rect 13771 38165 13780 38199
rect 13728 38156 13780 38165
rect 15016 38224 15068 38276
rect 17684 38335 17736 38344
rect 17684 38301 17693 38335
rect 17693 38301 17727 38335
rect 17727 38301 17736 38335
rect 17684 38292 17736 38301
rect 18144 38335 18196 38344
rect 18144 38301 18153 38335
rect 18153 38301 18187 38335
rect 18187 38301 18196 38335
rect 18144 38292 18196 38301
rect 18328 38292 18380 38344
rect 15476 38156 15528 38208
rect 15568 38199 15620 38208
rect 15568 38165 15577 38199
rect 15577 38165 15611 38199
rect 15611 38165 15620 38199
rect 15568 38156 15620 38165
rect 17776 38267 17828 38276
rect 17776 38233 17785 38267
rect 17785 38233 17819 38267
rect 17819 38233 17828 38267
rect 17776 38224 17828 38233
rect 18144 38156 18196 38208
rect 19432 38335 19484 38344
rect 19432 38301 19441 38335
rect 19441 38301 19475 38335
rect 19475 38301 19484 38335
rect 19432 38292 19484 38301
rect 19524 38335 19576 38344
rect 19524 38301 19533 38335
rect 19533 38301 19567 38335
rect 19567 38301 19576 38335
rect 19524 38292 19576 38301
rect 20076 38360 20128 38412
rect 18972 38156 19024 38208
rect 21272 38224 21324 38276
rect 19616 38199 19668 38208
rect 19616 38165 19625 38199
rect 19625 38165 19659 38199
rect 19659 38165 19668 38199
rect 19616 38156 19668 38165
rect 19984 38199 20036 38208
rect 19984 38165 19993 38199
rect 19993 38165 20027 38199
rect 20027 38165 20036 38199
rect 19984 38156 20036 38165
rect 5894 38054 5946 38106
rect 5958 38054 6010 38106
rect 6022 38054 6074 38106
rect 6086 38054 6138 38106
rect 6150 38054 6202 38106
rect 10839 38054 10891 38106
rect 10903 38054 10955 38106
rect 10967 38054 11019 38106
rect 11031 38054 11083 38106
rect 11095 38054 11147 38106
rect 15784 38054 15836 38106
rect 15848 38054 15900 38106
rect 15912 38054 15964 38106
rect 15976 38054 16028 38106
rect 16040 38054 16092 38106
rect 20729 38054 20781 38106
rect 20793 38054 20845 38106
rect 20857 38054 20909 38106
rect 20921 38054 20973 38106
rect 20985 38054 21037 38106
rect 3332 37884 3384 37936
rect 1860 37816 1912 37868
rect 2964 37816 3016 37868
rect 3792 37884 3844 37936
rect 4160 37884 4212 37936
rect 4528 37952 4580 38004
rect 6460 37952 6512 38004
rect 9680 37952 9732 38004
rect 9956 37995 10008 38004
rect 9956 37961 9965 37995
rect 9965 37961 9999 37995
rect 9999 37961 10008 37995
rect 9956 37952 10008 37961
rect 10324 37952 10376 38004
rect 10600 37952 10652 38004
rect 11520 37952 11572 38004
rect 6276 37884 6328 37936
rect 10232 37927 10284 37936
rect 10232 37893 10241 37927
rect 10241 37893 10275 37927
rect 10275 37893 10284 37927
rect 10232 37884 10284 37893
rect 13728 37952 13780 38004
rect 14372 37952 14424 38004
rect 15476 37952 15528 38004
rect 15568 37952 15620 38004
rect 2320 37748 2372 37800
rect 2780 37748 2832 37800
rect 4896 37816 4948 37868
rect 5540 37859 5592 37868
rect 5540 37825 5549 37859
rect 5549 37825 5583 37859
rect 5583 37825 5592 37859
rect 5540 37816 5592 37825
rect 6644 37816 6696 37868
rect 7380 37816 7432 37868
rect 10048 37816 10100 37868
rect 10600 37816 10652 37868
rect 10784 37816 10836 37868
rect 5356 37748 5408 37800
rect 5908 37748 5960 37800
rect 11888 37816 11940 37868
rect 11520 37791 11572 37800
rect 11520 37757 11529 37791
rect 11529 37757 11563 37791
rect 11563 37757 11572 37791
rect 11520 37748 11572 37757
rect 1400 37680 1452 37732
rect 4160 37655 4212 37664
rect 4160 37621 4169 37655
rect 4169 37621 4203 37655
rect 4203 37621 4212 37655
rect 4160 37612 4212 37621
rect 6368 37612 6420 37664
rect 6736 37612 6788 37664
rect 7472 37612 7524 37664
rect 9036 37680 9088 37732
rect 9588 37680 9640 37732
rect 7932 37612 7984 37664
rect 8760 37612 8812 37664
rect 9220 37612 9272 37664
rect 9496 37612 9548 37664
rect 12992 37612 13044 37664
rect 15108 37816 15160 37868
rect 15292 37859 15344 37868
rect 15292 37825 15301 37859
rect 15301 37825 15335 37859
rect 15335 37825 15344 37859
rect 15292 37816 15344 37825
rect 13912 37748 13964 37800
rect 17684 37995 17736 38004
rect 17684 37961 17693 37995
rect 17693 37961 17727 37995
rect 17727 37961 17736 37995
rect 17684 37952 17736 37961
rect 18144 37884 18196 37936
rect 19524 37952 19576 38004
rect 20260 37952 20312 38004
rect 19340 37884 19392 37936
rect 15844 37816 15896 37868
rect 17868 37816 17920 37868
rect 16488 37748 16540 37800
rect 16672 37791 16724 37800
rect 16672 37757 16681 37791
rect 16681 37757 16715 37791
rect 16715 37757 16724 37791
rect 16672 37748 16724 37757
rect 18972 37816 19024 37868
rect 19248 37816 19300 37868
rect 19524 37816 19576 37868
rect 19892 37748 19944 37800
rect 17776 37612 17828 37664
rect 19340 37612 19392 37664
rect 19800 37655 19852 37664
rect 19800 37621 19809 37655
rect 19809 37621 19843 37655
rect 19843 37621 19852 37655
rect 19800 37612 19852 37621
rect 19892 37612 19944 37664
rect 20168 37859 20220 37868
rect 20168 37825 20177 37859
rect 20177 37825 20211 37859
rect 20211 37825 20220 37859
rect 20168 37816 20220 37825
rect 20444 37655 20496 37664
rect 20444 37621 20453 37655
rect 20453 37621 20487 37655
rect 20487 37621 20496 37655
rect 20444 37612 20496 37621
rect 3422 37510 3474 37562
rect 3486 37510 3538 37562
rect 3550 37510 3602 37562
rect 3614 37510 3666 37562
rect 3678 37510 3730 37562
rect 8367 37510 8419 37562
rect 8431 37510 8483 37562
rect 8495 37510 8547 37562
rect 8559 37510 8611 37562
rect 8623 37510 8675 37562
rect 13312 37510 13364 37562
rect 13376 37510 13428 37562
rect 13440 37510 13492 37562
rect 13504 37510 13556 37562
rect 13568 37510 13620 37562
rect 18257 37510 18309 37562
rect 18321 37510 18373 37562
rect 18385 37510 18437 37562
rect 18449 37510 18501 37562
rect 18513 37510 18565 37562
rect 1032 37408 1084 37460
rect 1584 37272 1636 37324
rect 2780 37408 2832 37460
rect 4068 37408 4120 37460
rect 10600 37408 10652 37460
rect 3792 37340 3844 37392
rect 5264 37340 5316 37392
rect 9680 37340 9732 37392
rect 11520 37408 11572 37460
rect 14004 37408 14056 37460
rect 15108 37451 15160 37460
rect 15108 37417 15117 37451
rect 15117 37417 15151 37451
rect 15151 37417 15160 37451
rect 15108 37408 15160 37417
rect 18972 37408 19024 37460
rect 19156 37408 19208 37460
rect 17592 37340 17644 37392
rect 4068 37272 4120 37324
rect 5908 37315 5960 37324
rect 5908 37281 5917 37315
rect 5917 37281 5951 37315
rect 5951 37281 5960 37315
rect 5908 37272 5960 37281
rect 7472 37315 7524 37324
rect 7472 37281 7481 37315
rect 7481 37281 7515 37315
rect 7515 37281 7524 37315
rect 7472 37272 7524 37281
rect 12072 37272 12124 37324
rect 13636 37272 13688 37324
rect 2044 37204 2096 37256
rect 2688 37204 2740 37256
rect 1216 37136 1268 37188
rect 1308 37068 1360 37120
rect 4252 37204 4304 37256
rect 5264 37204 5316 37256
rect 5448 37136 5500 37188
rect 5540 37136 5592 37188
rect 6276 37136 6328 37188
rect 6368 37136 6420 37188
rect 6736 37136 6788 37188
rect 9036 37194 9088 37246
rect 9956 37204 10008 37256
rect 10784 37204 10836 37256
rect 9404 37136 9456 37188
rect 11244 37204 11296 37256
rect 13452 37136 13504 37188
rect 15568 37204 15620 37256
rect 16488 37204 16540 37256
rect 6920 37111 6972 37120
rect 6920 37077 6929 37111
rect 6929 37077 6963 37111
rect 6963 37077 6972 37111
rect 6920 37068 6972 37077
rect 8484 37111 8536 37120
rect 8484 37077 8493 37111
rect 8493 37077 8527 37111
rect 8527 37077 8536 37111
rect 8484 37068 8536 37077
rect 9036 37068 9088 37120
rect 11796 37068 11848 37120
rect 12072 37111 12124 37120
rect 12072 37077 12081 37111
rect 12081 37077 12115 37111
rect 12115 37077 12124 37111
rect 12072 37068 12124 37077
rect 19800 37340 19852 37392
rect 19340 37272 19392 37324
rect 21548 37340 21600 37392
rect 20260 37315 20312 37324
rect 20260 37281 20269 37315
rect 20269 37281 20303 37315
rect 20303 37281 20312 37315
rect 20260 37272 20312 37281
rect 21824 37272 21876 37324
rect 18696 37247 18748 37256
rect 18696 37213 18705 37247
rect 18705 37213 18739 37247
rect 18739 37213 18748 37247
rect 18696 37204 18748 37213
rect 18788 37204 18840 37256
rect 18972 37247 19024 37256
rect 18972 37213 18981 37247
rect 18981 37213 19015 37247
rect 19015 37213 19024 37247
rect 18972 37204 19024 37213
rect 20168 37204 20220 37256
rect 19708 37136 19760 37188
rect 19800 37179 19852 37188
rect 19800 37145 19809 37179
rect 19809 37145 19843 37179
rect 19843 37145 19852 37179
rect 19800 37136 19852 37145
rect 15844 37068 15896 37120
rect 17316 37068 17368 37120
rect 5894 36966 5946 37018
rect 5958 36966 6010 37018
rect 6022 36966 6074 37018
rect 6086 36966 6138 37018
rect 6150 36966 6202 37018
rect 10839 36966 10891 37018
rect 10903 36966 10955 37018
rect 10967 36966 11019 37018
rect 11031 36966 11083 37018
rect 11095 36966 11147 37018
rect 15784 36966 15836 37018
rect 15848 36966 15900 37018
rect 15912 36966 15964 37018
rect 15976 36966 16028 37018
rect 16040 36966 16092 37018
rect 20729 36966 20781 37018
rect 20793 36966 20845 37018
rect 20857 36966 20909 37018
rect 20921 36966 20973 37018
rect 20985 36966 21037 37018
rect 3056 36864 3108 36916
rect 664 36796 716 36848
rect 1768 36796 1820 36848
rect 6276 36864 6328 36916
rect 1492 36771 1544 36780
rect 1492 36737 1501 36771
rect 1501 36737 1535 36771
rect 1535 36737 1544 36771
rect 1492 36728 1544 36737
rect 1952 36771 2004 36780
rect 1952 36737 1961 36771
rect 1961 36737 1995 36771
rect 1995 36737 2004 36771
rect 1952 36728 2004 36737
rect 1216 36660 1268 36712
rect 3332 36660 3384 36712
rect 1308 36592 1360 36644
rect 6644 36796 6696 36848
rect 10416 36796 10468 36848
rect 13728 36796 13780 36848
rect 14004 36801 14056 36848
rect 4252 36771 4304 36780
rect 4252 36737 4261 36771
rect 4261 36737 4295 36771
rect 4295 36737 4304 36771
rect 4252 36728 4304 36737
rect 5356 36728 5408 36780
rect 5448 36728 5500 36780
rect 7472 36728 7524 36780
rect 8760 36771 8812 36780
rect 8760 36737 8769 36771
rect 8769 36737 8803 36771
rect 8803 36737 8812 36771
rect 8760 36728 8812 36737
rect 9036 36771 9088 36780
rect 9036 36737 9045 36771
rect 9045 36737 9079 36771
rect 9079 36737 9088 36771
rect 9036 36728 9088 36737
rect 9680 36728 9732 36780
rect 10048 36771 10100 36780
rect 10048 36737 10055 36771
rect 10055 36737 10089 36771
rect 10089 36737 10100 36771
rect 10048 36728 10100 36737
rect 11428 36728 11480 36780
rect 14004 36796 14029 36801
rect 14029 36796 14056 36801
rect 18696 36864 18748 36916
rect 18972 36864 19024 36916
rect 19156 36864 19208 36916
rect 19432 36864 19484 36916
rect 19248 36796 19300 36848
rect 2136 36524 2188 36576
rect 3240 36524 3292 36576
rect 5172 36660 5224 36712
rect 15384 36728 15436 36780
rect 15568 36728 15620 36780
rect 18144 36771 18196 36780
rect 18144 36737 18153 36771
rect 18153 36737 18187 36771
rect 18187 36737 18196 36771
rect 18144 36728 18196 36737
rect 18420 36771 18472 36780
rect 18420 36737 18429 36771
rect 18429 36737 18463 36771
rect 18463 36737 18472 36771
rect 18420 36728 18472 36737
rect 20168 36771 20220 36780
rect 20168 36737 20177 36771
rect 20177 36737 20211 36771
rect 20211 36737 20220 36771
rect 20168 36728 20220 36737
rect 7564 36660 7616 36712
rect 8024 36703 8076 36712
rect 8024 36669 8033 36703
rect 8033 36669 8067 36703
rect 8067 36669 8076 36703
rect 8024 36660 8076 36669
rect 8484 36703 8536 36712
rect 8484 36669 8493 36703
rect 8493 36669 8527 36703
rect 8527 36669 8536 36703
rect 8484 36660 8536 36669
rect 4160 36592 4212 36644
rect 7380 36592 7432 36644
rect 9772 36703 9824 36712
rect 7012 36524 7064 36576
rect 9036 36524 9088 36576
rect 9772 36669 9781 36703
rect 9781 36669 9815 36703
rect 9815 36669 9824 36703
rect 9772 36660 9824 36669
rect 9588 36524 9640 36576
rect 11336 36524 11388 36576
rect 13452 36660 13504 36712
rect 14740 36660 14792 36712
rect 16672 36660 16724 36712
rect 11796 36524 11848 36576
rect 12716 36524 12768 36576
rect 12900 36524 12952 36576
rect 13176 36524 13228 36576
rect 17040 36592 17092 36644
rect 14740 36567 14792 36576
rect 14740 36533 14749 36567
rect 14749 36533 14783 36567
rect 14783 36533 14792 36567
rect 14740 36524 14792 36533
rect 15200 36567 15252 36576
rect 15200 36533 15209 36567
rect 15209 36533 15243 36567
rect 15243 36533 15252 36567
rect 15200 36524 15252 36533
rect 15476 36524 15528 36576
rect 19892 36524 19944 36576
rect 21272 36524 21324 36576
rect 3422 36422 3474 36474
rect 3486 36422 3538 36474
rect 3550 36422 3602 36474
rect 3614 36422 3666 36474
rect 3678 36422 3730 36474
rect 8367 36422 8419 36474
rect 8431 36422 8483 36474
rect 8495 36422 8547 36474
rect 8559 36422 8611 36474
rect 8623 36422 8675 36474
rect 13312 36422 13364 36474
rect 13376 36422 13428 36474
rect 13440 36422 13492 36474
rect 13504 36422 13556 36474
rect 13568 36422 13620 36474
rect 18257 36422 18309 36474
rect 18321 36422 18373 36474
rect 18385 36422 18437 36474
rect 18449 36422 18501 36474
rect 18513 36422 18565 36474
rect 388 36320 440 36372
rect 2596 36320 2648 36372
rect 2872 36320 2924 36372
rect 6920 36320 6972 36372
rect 2228 36227 2280 36236
rect 2228 36193 2237 36227
rect 2237 36193 2271 36227
rect 2271 36193 2280 36227
rect 2228 36184 2280 36193
rect 4160 36252 4212 36304
rect 7472 36320 7524 36372
rect 3884 36184 3936 36236
rect 7564 36227 7616 36236
rect 7564 36193 7598 36227
rect 7598 36193 7616 36227
rect 7564 36184 7616 36193
rect 7932 36184 7984 36236
rect 756 36116 808 36168
rect 1032 36116 1084 36168
rect 1584 36159 1636 36168
rect 1584 36125 1593 36159
rect 1593 36125 1627 36159
rect 1627 36125 1636 36159
rect 1584 36116 1636 36125
rect 1768 36159 1820 36168
rect 1768 36125 1777 36159
rect 1777 36125 1811 36159
rect 1811 36125 1820 36159
rect 1768 36116 1820 36125
rect 2596 36159 2648 36168
rect 2596 36125 2630 36159
rect 2630 36125 2648 36159
rect 2596 36116 2648 36125
rect 2780 36159 2832 36168
rect 2780 36125 2789 36159
rect 2789 36125 2823 36159
rect 2823 36125 2832 36159
rect 2780 36116 2832 36125
rect 3976 36116 4028 36168
rect 4804 36116 4856 36168
rect 6552 36159 6604 36168
rect 6552 36125 6561 36159
rect 6561 36125 6595 36159
rect 6595 36125 6604 36159
rect 6552 36116 6604 36125
rect 6644 36116 6696 36168
rect 6920 36116 6972 36168
rect 7472 36159 7524 36168
rect 7472 36125 7481 36159
rect 7481 36125 7515 36159
rect 7515 36125 7524 36159
rect 7472 36116 7524 36125
rect 4620 36091 4672 36100
rect 4620 36057 4629 36091
rect 4629 36057 4663 36091
rect 4663 36057 4672 36091
rect 4620 36048 4672 36057
rect 4988 36091 5040 36100
rect 4988 36057 4997 36091
rect 4997 36057 5031 36091
rect 5031 36057 5040 36091
rect 4988 36048 5040 36057
rect 15292 36320 15344 36372
rect 15476 36320 15528 36372
rect 12348 36252 12400 36304
rect 13912 36252 13964 36304
rect 11244 36227 11296 36236
rect 11244 36193 11253 36227
rect 11253 36193 11287 36227
rect 11287 36193 11296 36227
rect 11244 36184 11296 36193
rect 14096 36227 14148 36236
rect 14096 36193 14105 36227
rect 14105 36193 14139 36227
rect 14139 36193 14148 36227
rect 14096 36184 14148 36193
rect 9036 36116 9088 36168
rect 9404 36116 9456 36168
rect 8760 36048 8812 36100
rect 11888 36116 11940 36168
rect 16672 36116 16724 36168
rect 18512 36320 18564 36372
rect 20168 36320 20220 36372
rect 18328 36252 18380 36304
rect 18972 36252 19024 36304
rect 20076 36252 20128 36304
rect 17408 36159 17460 36168
rect 17408 36125 17417 36159
rect 17417 36125 17451 36159
rect 17451 36125 17460 36159
rect 17408 36116 17460 36125
rect 15292 36048 15344 36100
rect 16212 36048 16264 36100
rect 18420 36116 18472 36168
rect 18972 36116 19024 36168
rect 19892 36116 19944 36168
rect 20536 36116 20588 36168
rect 2596 35980 2648 36032
rect 2872 35980 2924 36032
rect 3792 35980 3844 36032
rect 4160 35980 4212 36032
rect 4528 35980 4580 36032
rect 4896 35980 4948 36032
rect 6736 35980 6788 36032
rect 9956 35980 10008 36032
rect 10324 35980 10376 36032
rect 11428 35980 11480 36032
rect 11612 35980 11664 36032
rect 11888 35980 11940 36032
rect 13728 36023 13780 36032
rect 13728 35989 13737 36023
rect 13737 35989 13771 36023
rect 13771 35989 13780 36023
rect 13728 35980 13780 35989
rect 13820 35980 13872 36032
rect 15476 36023 15528 36032
rect 15476 35989 15485 36023
rect 15485 35989 15519 36023
rect 15519 35989 15528 36023
rect 15476 35980 15528 35989
rect 18880 36048 18932 36100
rect 19340 36048 19392 36100
rect 17224 35980 17276 36032
rect 17684 36023 17736 36032
rect 17684 35989 17693 36023
rect 17693 35989 17727 36023
rect 17727 35989 17736 36023
rect 17684 35980 17736 35989
rect 19524 35980 19576 36032
rect 5894 35878 5946 35930
rect 5958 35878 6010 35930
rect 6022 35878 6074 35930
rect 6086 35878 6138 35930
rect 6150 35878 6202 35930
rect 10839 35878 10891 35930
rect 10903 35878 10955 35930
rect 10967 35878 11019 35930
rect 11031 35878 11083 35930
rect 11095 35878 11147 35930
rect 15784 35878 15836 35930
rect 15848 35878 15900 35930
rect 15912 35878 15964 35930
rect 15976 35878 16028 35930
rect 16040 35878 16092 35930
rect 20729 35878 20781 35930
rect 20793 35878 20845 35930
rect 20857 35878 20909 35930
rect 20921 35878 20973 35930
rect 20985 35878 21037 35930
rect 2780 35776 2832 35828
rect 3884 35819 3936 35828
rect 3884 35785 3893 35819
rect 3893 35785 3927 35819
rect 3927 35785 3936 35819
rect 3884 35776 3936 35785
rect 4620 35776 4672 35828
rect 1400 35708 1452 35760
rect 1860 35708 1912 35760
rect 2320 35640 2372 35692
rect 2596 35640 2648 35692
rect 3148 35683 3200 35692
rect 3148 35649 3155 35683
rect 3155 35649 3189 35683
rect 3189 35649 3200 35683
rect 3148 35640 3200 35649
rect 5632 35708 5684 35760
rect 10140 35776 10192 35828
rect 10232 35776 10284 35828
rect 10784 35776 10836 35828
rect 4620 35683 4672 35692
rect 4620 35649 4627 35683
rect 4627 35649 4661 35683
rect 4661 35649 4672 35683
rect 4620 35640 4672 35649
rect 9772 35751 9824 35760
rect 9772 35717 9781 35751
rect 9781 35717 9815 35751
rect 9815 35717 9824 35751
rect 9772 35708 9824 35717
rect 9864 35708 9916 35760
rect 10140 35683 10192 35692
rect 10140 35649 10149 35683
rect 10149 35649 10183 35683
rect 10183 35649 10192 35683
rect 10140 35640 10192 35649
rect 10508 35751 10560 35760
rect 10508 35717 10517 35751
rect 10517 35717 10551 35751
rect 10551 35717 10560 35751
rect 10508 35708 10560 35717
rect 1400 35572 1452 35624
rect 4160 35572 4212 35624
rect 5724 35572 5776 35624
rect 6368 35572 6420 35624
rect 9588 35572 9640 35624
rect 10600 35572 10652 35624
rect 13728 35776 13780 35828
rect 15384 35819 15436 35828
rect 15384 35785 15393 35819
rect 15393 35785 15427 35819
rect 15427 35785 15436 35819
rect 15384 35776 15436 35785
rect 15476 35776 15528 35828
rect 17408 35776 17460 35828
rect 17684 35776 17736 35828
rect 18328 35776 18380 35828
rect 12716 35683 12768 35692
rect 12716 35649 12725 35683
rect 12725 35649 12759 35683
rect 12759 35649 12768 35683
rect 12716 35640 12768 35649
rect 15200 35708 15252 35760
rect 16212 35708 16264 35760
rect 17040 35683 17092 35692
rect 17040 35649 17049 35683
rect 17049 35649 17083 35683
rect 17083 35649 17092 35683
rect 17040 35640 17092 35649
rect 18512 35776 18564 35828
rect 19524 35776 19576 35828
rect 19616 35776 19668 35828
rect 17960 35640 18012 35692
rect 11612 35572 11664 35624
rect 11796 35572 11848 35624
rect 12072 35572 12124 35624
rect 10784 35504 10836 35556
rect 10876 35504 10928 35556
rect 3332 35436 3384 35488
rect 6736 35436 6788 35488
rect 14648 35572 14700 35624
rect 14740 35615 14792 35624
rect 14740 35581 14749 35615
rect 14749 35581 14783 35615
rect 14783 35581 14792 35615
rect 14740 35572 14792 35581
rect 13544 35504 13596 35556
rect 15200 35572 15252 35624
rect 17224 35572 17276 35624
rect 19156 35640 19208 35692
rect 19432 35640 19484 35692
rect 18696 35572 18748 35624
rect 19616 35683 19668 35692
rect 19616 35649 19625 35683
rect 19625 35649 19659 35683
rect 19659 35649 19668 35683
rect 19616 35640 19668 35649
rect 19984 35708 20036 35760
rect 20076 35683 20128 35692
rect 20076 35649 20085 35683
rect 20085 35649 20119 35683
rect 20119 35649 20128 35683
rect 20076 35640 20128 35649
rect 20536 35683 20588 35692
rect 20536 35649 20545 35683
rect 20545 35649 20579 35683
rect 20579 35649 20588 35683
rect 20536 35640 20588 35649
rect 20628 35572 20680 35624
rect 12808 35436 12860 35488
rect 13176 35436 13228 35488
rect 14372 35436 14424 35488
rect 16580 35436 16632 35488
rect 17132 35436 17184 35488
rect 17224 35479 17276 35488
rect 17224 35445 17233 35479
rect 17233 35445 17267 35479
rect 17267 35445 17276 35479
rect 17224 35436 17276 35445
rect 18144 35436 18196 35488
rect 19248 35504 19300 35556
rect 19892 35504 19944 35556
rect 19156 35479 19208 35488
rect 19156 35445 19165 35479
rect 19165 35445 19199 35479
rect 19199 35445 19208 35479
rect 19156 35436 19208 35445
rect 19708 35436 19760 35488
rect 19984 35436 20036 35488
rect 21364 35436 21416 35488
rect 3422 35334 3474 35386
rect 3486 35334 3538 35386
rect 3550 35334 3602 35386
rect 3614 35334 3666 35386
rect 3678 35334 3730 35386
rect 8367 35334 8419 35386
rect 8431 35334 8483 35386
rect 8495 35334 8547 35386
rect 8559 35334 8611 35386
rect 8623 35334 8675 35386
rect 13312 35334 13364 35386
rect 13376 35334 13428 35386
rect 13440 35334 13492 35386
rect 13504 35334 13556 35386
rect 13568 35334 13620 35386
rect 18257 35334 18309 35386
rect 18321 35334 18373 35386
rect 18385 35334 18437 35386
rect 18449 35334 18501 35386
rect 18513 35334 18565 35386
rect 2228 35232 2280 35284
rect 5080 35232 5132 35284
rect 2504 35164 2556 35216
rect 6460 35232 6512 35284
rect 7748 35232 7800 35284
rect 10324 35232 10376 35284
rect 10600 35232 10652 35284
rect 11428 35232 11480 35284
rect 11888 35232 11940 35284
rect 8760 35164 8812 35216
rect 9312 35164 9364 35216
rect 9496 35164 9548 35216
rect 1124 35096 1176 35148
rect 1400 35139 1452 35148
rect 1400 35105 1409 35139
rect 1409 35105 1443 35139
rect 1443 35105 1452 35139
rect 1400 35096 1452 35105
rect 1676 35071 1728 35080
rect 1676 35037 1683 35071
rect 1683 35037 1717 35071
rect 1717 35037 1728 35071
rect 3148 35096 3200 35148
rect 1676 35028 1728 35037
rect 2780 35071 2832 35080
rect 2780 35037 2789 35071
rect 2789 35037 2823 35071
rect 2823 35037 2832 35071
rect 2780 35028 2832 35037
rect 3792 35071 3844 35080
rect 3792 35037 3801 35071
rect 3801 35037 3835 35071
rect 3835 35037 3844 35071
rect 3792 35028 3844 35037
rect 4068 35003 4120 35012
rect 4068 34969 4077 35003
rect 4077 34969 4111 35003
rect 4111 34969 4120 35003
rect 4068 34960 4120 34969
rect 4712 34960 4764 35012
rect 2320 34892 2372 34944
rect 4620 34892 4672 34944
rect 5264 35028 5316 35080
rect 6736 35071 6788 35080
rect 6736 35037 6743 35071
rect 6743 35037 6777 35071
rect 6777 35037 6788 35071
rect 6736 35028 6788 35037
rect 7932 35028 7984 35080
rect 8760 35028 8812 35080
rect 9036 35028 9088 35080
rect 12072 35164 12124 35216
rect 12256 35232 12308 35284
rect 11244 35096 11296 35148
rect 11428 35096 11480 35148
rect 11796 35096 11848 35148
rect 13820 35232 13872 35284
rect 6920 34960 6972 35012
rect 7012 34960 7064 35012
rect 11612 35028 11664 35080
rect 12440 35071 12492 35080
rect 12440 35037 12449 35071
rect 12449 35037 12483 35071
rect 12483 35037 12492 35071
rect 12440 35028 12492 35037
rect 12532 35028 12584 35080
rect 12716 35071 12768 35080
rect 12716 35037 12725 35071
rect 12725 35037 12759 35071
rect 12759 35037 12768 35071
rect 12716 35028 12768 35037
rect 14004 35028 14056 35080
rect 14372 35071 14424 35080
rect 14372 35037 14381 35071
rect 14381 35037 14415 35071
rect 14415 35037 14424 35071
rect 14372 35028 14424 35037
rect 14556 35028 14608 35080
rect 15844 35207 15896 35216
rect 15844 35173 15853 35207
rect 15853 35173 15887 35207
rect 15887 35173 15896 35207
rect 15844 35164 15896 35173
rect 17040 35232 17092 35284
rect 18880 35275 18932 35284
rect 18880 35241 18889 35275
rect 18889 35241 18923 35275
rect 18923 35241 18932 35275
rect 18880 35232 18932 35241
rect 19432 35232 19484 35284
rect 20352 35232 20404 35284
rect 10324 34960 10376 35012
rect 5908 34892 5960 34944
rect 6828 34892 6880 34944
rect 7564 34892 7616 34944
rect 9772 34892 9824 34944
rect 9956 34892 10008 34944
rect 10876 34892 10928 34944
rect 11336 34892 11388 34944
rect 13820 34960 13872 35012
rect 14188 34960 14240 35012
rect 14372 34892 14424 34944
rect 15292 34892 15344 34944
rect 16488 35028 16540 35080
rect 17408 35028 17460 35080
rect 18696 35028 18748 35080
rect 19156 35028 19208 35080
rect 19432 35096 19484 35148
rect 20444 35096 20496 35148
rect 16212 34960 16264 35012
rect 18052 34960 18104 35012
rect 18144 34960 18196 35012
rect 16396 34892 16448 34944
rect 18512 34935 18564 34944
rect 18512 34901 18521 34935
rect 18521 34901 18555 34935
rect 18555 34901 18564 34935
rect 18512 34892 18564 34901
rect 18604 34892 18656 34944
rect 18972 34892 19024 34944
rect 21272 34892 21324 34944
rect 5894 34790 5946 34842
rect 5958 34790 6010 34842
rect 6022 34790 6074 34842
rect 6086 34790 6138 34842
rect 6150 34790 6202 34842
rect 10839 34790 10891 34842
rect 10903 34790 10955 34842
rect 10967 34790 11019 34842
rect 11031 34790 11083 34842
rect 11095 34790 11147 34842
rect 15784 34790 15836 34842
rect 15848 34790 15900 34842
rect 15912 34790 15964 34842
rect 15976 34790 16028 34842
rect 16040 34790 16092 34842
rect 20729 34790 20781 34842
rect 20793 34790 20845 34842
rect 20857 34790 20909 34842
rect 20921 34790 20973 34842
rect 20985 34790 21037 34842
rect 1768 34688 1820 34740
rect 1216 34552 1268 34604
rect 1952 34595 2004 34604
rect 1952 34561 1961 34595
rect 1961 34561 1995 34595
rect 1995 34561 2004 34595
rect 1952 34552 2004 34561
rect 2320 34552 2372 34604
rect 2596 34620 2648 34672
rect 3056 34620 3108 34672
rect 3424 34688 3476 34740
rect 5264 34688 5316 34740
rect 5448 34731 5500 34740
rect 5448 34697 5457 34731
rect 5457 34697 5491 34731
rect 5491 34697 5500 34731
rect 5448 34688 5500 34697
rect 6736 34688 6788 34740
rect 8024 34688 8076 34740
rect 8944 34688 8996 34740
rect 9128 34688 9180 34740
rect 3332 34552 3384 34604
rect 4620 34620 4672 34672
rect 7288 34620 7340 34672
rect 7380 34663 7432 34672
rect 7380 34629 7389 34663
rect 7389 34629 7423 34663
rect 7423 34629 7432 34663
rect 7380 34620 7432 34629
rect 8300 34620 8352 34672
rect 9956 34688 10008 34740
rect 10324 34688 10376 34740
rect 11704 34688 11756 34740
rect 12716 34688 12768 34740
rect 19340 34688 19392 34740
rect 20536 34688 20588 34740
rect 1768 34484 1820 34536
rect 2412 34484 2464 34536
rect 1492 34348 1544 34400
rect 3424 34348 3476 34400
rect 3884 34348 3936 34400
rect 4712 34595 4764 34604
rect 4712 34561 4719 34595
rect 4719 34561 4753 34595
rect 4753 34561 4764 34595
rect 4712 34552 4764 34561
rect 5264 34552 5316 34604
rect 7748 34552 7800 34604
rect 7840 34595 7892 34604
rect 7840 34561 7849 34595
rect 7849 34561 7883 34595
rect 7883 34561 7892 34595
rect 7840 34552 7892 34561
rect 11428 34620 11480 34672
rect 9864 34552 9916 34604
rect 12532 34620 12584 34672
rect 12164 34552 12216 34604
rect 18052 34620 18104 34672
rect 13820 34552 13872 34604
rect 14280 34552 14332 34604
rect 16672 34595 16724 34604
rect 16672 34561 16681 34595
rect 16681 34561 16715 34595
rect 16715 34561 16724 34595
rect 16672 34552 16724 34561
rect 16948 34595 17000 34604
rect 16948 34561 16982 34595
rect 16982 34561 17000 34595
rect 16948 34552 17000 34561
rect 18512 34620 18564 34672
rect 19524 34620 19576 34672
rect 5908 34484 5960 34536
rect 7564 34484 7616 34536
rect 8852 34527 8904 34536
rect 8852 34493 8861 34527
rect 8861 34493 8895 34527
rect 8895 34493 8904 34527
rect 8852 34484 8904 34493
rect 8944 34484 8996 34536
rect 9956 34484 10008 34536
rect 11060 34527 11112 34536
rect 11060 34493 11069 34527
rect 11069 34493 11103 34527
rect 11103 34493 11112 34527
rect 11060 34484 11112 34493
rect 15016 34484 15068 34536
rect 4896 34348 4948 34400
rect 9036 34416 9088 34468
rect 16580 34416 16632 34468
rect 19340 34595 19392 34604
rect 19340 34561 19349 34595
rect 19349 34561 19383 34595
rect 19383 34561 19392 34595
rect 19340 34552 19392 34561
rect 19432 34552 19484 34604
rect 19892 34595 19944 34604
rect 19892 34561 19901 34595
rect 19901 34561 19935 34595
rect 19935 34561 19944 34595
rect 19892 34552 19944 34561
rect 9312 34348 9364 34400
rect 10600 34391 10652 34400
rect 10600 34357 10609 34391
rect 10609 34357 10643 34391
rect 10643 34357 10652 34391
rect 10600 34348 10652 34357
rect 12256 34348 12308 34400
rect 12716 34348 12768 34400
rect 12992 34348 13044 34400
rect 14280 34348 14332 34400
rect 15016 34348 15068 34400
rect 17592 34348 17644 34400
rect 18696 34348 18748 34400
rect 20352 34348 20404 34400
rect 20444 34391 20496 34400
rect 20444 34357 20453 34391
rect 20453 34357 20487 34391
rect 20487 34357 20496 34391
rect 20444 34348 20496 34357
rect 3422 34246 3474 34298
rect 3486 34246 3538 34298
rect 3550 34246 3602 34298
rect 3614 34246 3666 34298
rect 3678 34246 3730 34298
rect 8367 34246 8419 34298
rect 8431 34246 8483 34298
rect 8495 34246 8547 34298
rect 8559 34246 8611 34298
rect 8623 34246 8675 34298
rect 13312 34246 13364 34298
rect 13376 34246 13428 34298
rect 13440 34246 13492 34298
rect 13504 34246 13556 34298
rect 13568 34246 13620 34298
rect 18257 34246 18309 34298
rect 18321 34246 18373 34298
rect 18385 34246 18437 34298
rect 18449 34246 18501 34298
rect 18513 34246 18565 34298
rect 2320 34051 2372 34060
rect 2320 34017 2329 34051
rect 2329 34017 2363 34051
rect 2363 34017 2372 34051
rect 2320 34008 2372 34017
rect 4436 34144 4488 34196
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 2044 33872 2096 33924
rect 3240 33940 3292 33992
rect 4252 33940 4304 33992
rect 4620 33940 4672 33992
rect 8576 34144 8628 34196
rect 8852 34144 8904 34196
rect 9312 34144 9364 34196
rect 6552 34076 6604 34128
rect 6828 34076 6880 34128
rect 7104 34076 7156 34128
rect 8760 34076 8812 34128
rect 9956 34144 10008 34196
rect 10140 34144 10192 34196
rect 10416 34144 10468 34196
rect 15384 34144 15436 34196
rect 16580 34144 16632 34196
rect 16856 34144 16908 34196
rect 17592 34187 17644 34196
rect 17592 34153 17601 34187
rect 17601 34153 17635 34187
rect 17635 34153 17644 34187
rect 17592 34144 17644 34153
rect 18512 34144 18564 34196
rect 19340 34144 19392 34196
rect 19524 34187 19576 34196
rect 19524 34153 19533 34187
rect 19533 34153 19567 34187
rect 19567 34153 19576 34187
rect 19524 34144 19576 34153
rect 19616 34144 19668 34196
rect 13820 34119 13872 34128
rect 13820 34085 13829 34119
rect 13829 34085 13863 34119
rect 13863 34085 13872 34119
rect 13820 34076 13872 34085
rect 4896 34008 4948 34060
rect 7472 34051 7524 34060
rect 7472 34017 7481 34051
rect 7481 34017 7515 34051
rect 7515 34017 7524 34051
rect 7472 34008 7524 34017
rect 7656 34008 7708 34060
rect 5264 33983 5316 33992
rect 5264 33949 5271 33983
rect 5271 33949 5305 33983
rect 5305 33949 5316 33983
rect 5264 33940 5316 33949
rect 6644 33940 6696 33992
rect 6736 33983 6788 33992
rect 6736 33949 6745 33983
rect 6745 33949 6779 33983
rect 6779 33949 6788 33983
rect 6736 33940 6788 33949
rect 7932 34008 7984 34060
rect 8116 34008 8168 34060
rect 8668 34008 8720 34060
rect 1308 33804 1360 33856
rect 3332 33847 3384 33856
rect 3332 33813 3341 33847
rect 3341 33813 3375 33847
rect 3375 33813 3384 33847
rect 3332 33804 3384 33813
rect 4160 33804 4212 33856
rect 4620 33804 4672 33856
rect 5540 33804 5592 33856
rect 8484 33804 8536 33856
rect 8760 33983 8812 33992
rect 8760 33949 8769 33983
rect 8769 33949 8803 33983
rect 8803 33949 8812 33983
rect 8760 33940 8812 33949
rect 9772 34008 9824 34060
rect 9404 33940 9456 33992
rect 10324 33940 10376 33992
rect 12532 34008 12584 34060
rect 13728 34008 13780 34060
rect 13912 34051 13964 34060
rect 13912 34017 13921 34051
rect 13921 34017 13955 34051
rect 13955 34017 13964 34051
rect 13912 34008 13964 34017
rect 8944 33804 8996 33856
rect 11244 33872 11296 33924
rect 9496 33804 9548 33856
rect 11612 33872 11664 33924
rect 12164 33872 12216 33924
rect 11796 33847 11848 33856
rect 11796 33813 11805 33847
rect 11805 33813 11839 33847
rect 11839 33813 11848 33847
rect 11796 33804 11848 33813
rect 12624 33804 12676 33856
rect 13176 33804 13228 33856
rect 14740 33940 14792 33992
rect 15660 33940 15712 33992
rect 16764 34008 16816 34060
rect 16948 33940 17000 33992
rect 18604 34008 18656 34060
rect 19156 34076 19208 34128
rect 13820 33872 13872 33924
rect 14556 33872 14608 33924
rect 16580 33872 16632 33924
rect 18236 33983 18288 33992
rect 18236 33949 18245 33983
rect 18245 33949 18279 33983
rect 18279 33949 18288 33983
rect 18236 33940 18288 33949
rect 18696 33940 18748 33992
rect 20076 34008 20128 34060
rect 18880 33940 18932 33992
rect 19432 33983 19484 33992
rect 19432 33949 19441 33983
rect 19441 33949 19475 33983
rect 19475 33949 19484 33983
rect 19432 33940 19484 33949
rect 19616 33983 19668 33992
rect 19616 33949 19625 33983
rect 19625 33949 19659 33983
rect 19659 33949 19668 33983
rect 19616 33940 19668 33949
rect 20168 33940 20220 33992
rect 14740 33804 14792 33856
rect 15200 33804 15252 33856
rect 17132 33804 17184 33856
rect 17592 33804 17644 33856
rect 19156 33804 19208 33856
rect 19800 33847 19852 33856
rect 19800 33813 19809 33847
rect 19809 33813 19843 33847
rect 19843 33813 19852 33847
rect 19800 33804 19852 33813
rect 21180 33804 21232 33856
rect 5894 33702 5946 33754
rect 5958 33702 6010 33754
rect 6022 33702 6074 33754
rect 6086 33702 6138 33754
rect 6150 33702 6202 33754
rect 10839 33702 10891 33754
rect 10903 33702 10955 33754
rect 10967 33702 11019 33754
rect 11031 33702 11083 33754
rect 11095 33702 11147 33754
rect 15784 33702 15836 33754
rect 15848 33702 15900 33754
rect 15912 33702 15964 33754
rect 15976 33702 16028 33754
rect 16040 33702 16092 33754
rect 20729 33702 20781 33754
rect 20793 33702 20845 33754
rect 20857 33702 20909 33754
rect 20921 33702 20973 33754
rect 20985 33702 21037 33754
rect 1676 33600 1728 33652
rect 3332 33600 3384 33652
rect 1860 33532 1912 33584
rect 3240 33532 3292 33584
rect 3700 33575 3752 33584
rect 3700 33541 3709 33575
rect 3709 33541 3743 33575
rect 3743 33541 3752 33575
rect 3700 33532 3752 33541
rect 3976 33575 4028 33584
rect 3976 33541 3985 33575
rect 3985 33541 4019 33575
rect 4019 33541 4028 33575
rect 3976 33532 4028 33541
rect 2780 33507 2832 33516
rect 2780 33473 2789 33507
rect 2789 33473 2823 33507
rect 2823 33473 2832 33507
rect 2780 33464 2832 33473
rect 7196 33600 7248 33652
rect 7656 33600 7708 33652
rect 7840 33600 7892 33652
rect 8760 33600 8812 33652
rect 4528 33532 4580 33584
rect 6276 33532 6328 33584
rect 4436 33507 4488 33516
rect 4436 33473 4445 33507
rect 4445 33473 4479 33507
rect 4479 33473 4488 33507
rect 4436 33464 4488 33473
rect 4988 33464 5040 33516
rect 6828 33532 6880 33584
rect 7564 33507 7616 33516
rect 7564 33473 7573 33507
rect 7573 33473 7607 33507
rect 7607 33473 7616 33507
rect 7564 33464 7616 33473
rect 8852 33507 8904 33516
rect 1308 33396 1360 33448
rect 3884 33396 3936 33448
rect 5264 33396 5316 33448
rect 7380 33396 7432 33448
rect 8024 33396 8076 33448
rect 8852 33473 8859 33507
rect 8859 33473 8893 33507
rect 8893 33473 8904 33507
rect 8852 33464 8904 33473
rect 8944 33464 8996 33516
rect 7104 33328 7156 33380
rect 2412 33303 2464 33312
rect 2412 33269 2421 33303
rect 2421 33269 2455 33303
rect 2455 33269 2464 33303
rect 2412 33260 2464 33269
rect 6736 33260 6788 33312
rect 7564 33260 7616 33312
rect 7656 33260 7708 33312
rect 11244 33464 11296 33516
rect 12072 33532 12124 33584
rect 13820 33532 13872 33584
rect 12992 33464 13044 33516
rect 14740 33600 14792 33652
rect 15016 33600 15068 33652
rect 16580 33600 16632 33652
rect 18236 33600 18288 33652
rect 18512 33600 18564 33652
rect 13912 33396 13964 33448
rect 15200 33507 15252 33516
rect 15200 33473 15209 33507
rect 15209 33473 15243 33507
rect 15243 33473 15252 33507
rect 15200 33464 15252 33473
rect 16120 33507 16172 33516
rect 16120 33473 16129 33507
rect 16129 33473 16163 33507
rect 16163 33473 16172 33507
rect 16120 33464 16172 33473
rect 8484 33260 8536 33312
rect 9496 33260 9548 33312
rect 12348 33260 12400 33312
rect 13176 33260 13228 33312
rect 14740 33396 14792 33448
rect 15016 33439 15068 33448
rect 15016 33405 15050 33439
rect 15050 33405 15068 33439
rect 15016 33396 15068 33405
rect 14372 33328 14424 33380
rect 19616 33600 19668 33652
rect 18972 33464 19024 33516
rect 19524 33464 19576 33516
rect 20260 33464 20312 33516
rect 19340 33260 19392 33312
rect 20444 33303 20496 33312
rect 20444 33269 20453 33303
rect 20453 33269 20487 33303
rect 20487 33269 20496 33303
rect 20444 33260 20496 33269
rect 3422 33158 3474 33210
rect 3486 33158 3538 33210
rect 3550 33158 3602 33210
rect 3614 33158 3666 33210
rect 3678 33158 3730 33210
rect 8367 33158 8419 33210
rect 8431 33158 8483 33210
rect 8495 33158 8547 33210
rect 8559 33158 8611 33210
rect 8623 33158 8675 33210
rect 13312 33158 13364 33210
rect 13376 33158 13428 33210
rect 13440 33158 13492 33210
rect 13504 33158 13556 33210
rect 13568 33158 13620 33210
rect 18257 33158 18309 33210
rect 18321 33158 18373 33210
rect 18385 33158 18437 33210
rect 18449 33158 18501 33210
rect 18513 33158 18565 33210
rect 1952 33056 2004 33108
rect 3056 33056 3108 33108
rect 4344 33056 4396 33108
rect 4988 33056 5040 33108
rect 5172 33056 5224 33108
rect 7564 33056 7616 33108
rect 7748 33056 7800 33108
rect 8208 33056 8260 33108
rect 9312 33056 9364 33108
rect 10508 33056 10560 33108
rect 6644 32988 6696 33040
rect 7288 32988 7340 33040
rect 8576 32988 8628 33040
rect 12440 33056 12492 33108
rect 12532 33056 12584 33108
rect 15384 33056 15436 33108
rect 16120 33056 16172 33108
rect 17224 33056 17276 33108
rect 18052 33056 18104 33108
rect 1308 32920 1360 32972
rect 756 32852 808 32904
rect 1492 32784 1544 32836
rect 2964 32920 3016 32972
rect 4804 32920 4856 32972
rect 5448 32920 5500 32972
rect 6920 32920 6972 32972
rect 7104 32920 7156 32972
rect 2228 32895 2280 32904
rect 2228 32861 2235 32895
rect 2235 32861 2269 32895
rect 2269 32861 2280 32895
rect 2228 32852 2280 32861
rect 2872 32852 2924 32904
rect 4068 32895 4120 32904
rect 4068 32861 4077 32895
rect 4077 32861 4111 32895
rect 4111 32861 4120 32895
rect 4068 32852 4120 32861
rect 2688 32784 2740 32836
rect 1216 32716 1268 32768
rect 3056 32716 3108 32768
rect 3332 32784 3384 32836
rect 3884 32784 3936 32836
rect 5540 32895 5592 32904
rect 5540 32861 5549 32895
rect 5549 32861 5583 32895
rect 5583 32861 5592 32895
rect 5540 32852 5592 32861
rect 6460 32852 6512 32904
rect 6644 32852 6696 32904
rect 7012 32852 7064 32904
rect 8852 32920 8904 32972
rect 5172 32759 5224 32768
rect 5172 32725 5181 32759
rect 5181 32725 5215 32759
rect 5215 32725 5224 32759
rect 5172 32716 5224 32725
rect 5632 32784 5684 32836
rect 6368 32784 6420 32836
rect 8116 32852 8168 32904
rect 11796 33031 11848 33040
rect 11796 32997 11805 33031
rect 11805 32997 11839 33031
rect 11839 32997 11848 33031
rect 11796 32988 11848 32997
rect 11704 32920 11756 32972
rect 12348 32963 12400 32972
rect 12348 32929 12357 32963
rect 12357 32929 12391 32963
rect 12391 32929 12400 32963
rect 12348 32920 12400 32929
rect 12532 32920 12584 32972
rect 8944 32784 8996 32836
rect 6736 32716 6788 32768
rect 6920 32716 6972 32768
rect 11152 32895 11204 32904
rect 11152 32861 11161 32895
rect 11161 32861 11195 32895
rect 11195 32861 11204 32895
rect 11152 32852 11204 32861
rect 9864 32716 9916 32768
rect 12164 32895 12216 32904
rect 12164 32861 12198 32895
rect 12198 32861 12216 32895
rect 14004 32920 14056 32972
rect 12164 32852 12216 32861
rect 15660 32895 15712 32904
rect 15660 32861 15669 32895
rect 15669 32861 15703 32895
rect 15703 32861 15712 32895
rect 15660 32852 15712 32861
rect 13820 32784 13872 32836
rect 17408 32852 17460 32904
rect 18604 32852 18656 32904
rect 19432 33056 19484 33108
rect 19708 33056 19760 33108
rect 21272 32988 21324 33040
rect 19340 32895 19392 32904
rect 19340 32861 19349 32895
rect 19349 32861 19383 32895
rect 19383 32861 19392 32895
rect 19340 32852 19392 32861
rect 18788 32784 18840 32836
rect 19616 32784 19668 32836
rect 19984 32852 20036 32904
rect 20076 32852 20128 32904
rect 20536 32827 20588 32836
rect 20536 32793 20545 32827
rect 20545 32793 20579 32827
rect 20579 32793 20588 32827
rect 20536 32784 20588 32793
rect 12440 32716 12492 32768
rect 12992 32716 13044 32768
rect 13728 32716 13780 32768
rect 14004 32716 14056 32768
rect 14556 32716 14608 32768
rect 14832 32716 14884 32768
rect 16212 32716 16264 32768
rect 16856 32716 16908 32768
rect 17316 32716 17368 32768
rect 19432 32716 19484 32768
rect 21640 32716 21692 32768
rect 5894 32614 5946 32666
rect 5958 32614 6010 32666
rect 6022 32614 6074 32666
rect 6086 32614 6138 32666
rect 6150 32614 6202 32666
rect 10839 32614 10891 32666
rect 10903 32614 10955 32666
rect 10967 32614 11019 32666
rect 11031 32614 11083 32666
rect 11095 32614 11147 32666
rect 15784 32614 15836 32666
rect 15848 32614 15900 32666
rect 15912 32614 15964 32666
rect 15976 32614 16028 32666
rect 16040 32614 16092 32666
rect 20729 32614 20781 32666
rect 20793 32614 20845 32666
rect 20857 32614 20909 32666
rect 20921 32614 20973 32666
rect 20985 32614 21037 32666
rect 1308 32512 1360 32564
rect 1860 32444 1912 32496
rect 1400 32419 1452 32428
rect 1400 32385 1409 32419
rect 1409 32385 1443 32419
rect 1443 32385 1452 32419
rect 1400 32376 1452 32385
rect 3056 32444 3108 32496
rect 3332 32487 3384 32496
rect 3332 32453 3341 32487
rect 3341 32453 3375 32487
rect 3375 32453 3384 32487
rect 3332 32444 3384 32453
rect 2780 32376 2832 32428
rect 2964 32419 3016 32428
rect 2964 32385 2973 32419
rect 2973 32385 3007 32419
rect 3007 32385 3016 32419
rect 2964 32376 3016 32385
rect 4068 32512 4120 32564
rect 5448 32444 5500 32496
rect 7472 32444 7524 32496
rect 3884 32376 3936 32428
rect 4344 32376 4396 32428
rect 4804 32376 4856 32428
rect 5540 32376 5592 32428
rect 6920 32376 6972 32428
rect 7104 32419 7156 32428
rect 7104 32385 7113 32419
rect 7113 32385 7147 32419
rect 7147 32385 7156 32419
rect 7104 32376 7156 32385
rect 7380 32419 7432 32428
rect 7380 32385 7387 32419
rect 7387 32385 7421 32419
rect 7421 32385 7432 32419
rect 7380 32376 7432 32385
rect 8024 32512 8076 32564
rect 9312 32512 9364 32564
rect 13820 32555 13872 32564
rect 13820 32521 13829 32555
rect 13829 32521 13863 32555
rect 13863 32521 13872 32555
rect 13820 32512 13872 32521
rect 9404 32444 9456 32496
rect 14280 32444 14332 32496
rect 16672 32512 16724 32564
rect 17132 32555 17184 32564
rect 17132 32521 17141 32555
rect 17141 32521 17175 32555
rect 17175 32521 17184 32555
rect 17132 32512 17184 32521
rect 19340 32512 19392 32564
rect 2412 32308 2464 32360
rect 2136 32240 2188 32292
rect 3516 32283 3568 32292
rect 3516 32249 3525 32283
rect 3525 32249 3559 32283
rect 3559 32249 3568 32283
rect 3516 32240 3568 32249
rect 8944 32308 8996 32360
rect 9680 32376 9732 32428
rect 10784 32376 10836 32428
rect 11612 32376 11664 32428
rect 13176 32376 13228 32428
rect 13820 32376 13872 32428
rect 4896 32172 4948 32224
rect 5356 32172 5408 32224
rect 5448 32215 5500 32224
rect 5448 32181 5457 32215
rect 5457 32181 5491 32215
rect 5491 32181 5500 32215
rect 5448 32172 5500 32181
rect 6552 32172 6604 32224
rect 9496 32172 9548 32224
rect 10232 32172 10284 32224
rect 10508 32215 10560 32224
rect 10508 32181 10517 32215
rect 10517 32181 10551 32215
rect 10551 32181 10560 32215
rect 10508 32172 10560 32181
rect 11060 32172 11112 32224
rect 11980 32172 12032 32224
rect 12164 32172 12216 32224
rect 14280 32351 14332 32360
rect 14280 32317 14289 32351
rect 14289 32317 14323 32351
rect 14323 32317 14332 32351
rect 14280 32308 14332 32317
rect 15292 32419 15344 32428
rect 15292 32385 15301 32419
rect 15301 32385 15335 32419
rect 15335 32385 15344 32419
rect 15292 32376 15344 32385
rect 15108 32351 15160 32360
rect 15108 32317 15142 32351
rect 15142 32317 15160 32351
rect 16212 32419 16264 32428
rect 16212 32385 16221 32419
rect 16221 32385 16255 32419
rect 16255 32385 16264 32419
rect 16212 32376 16264 32385
rect 16580 32376 16632 32428
rect 17960 32376 18012 32428
rect 18236 32376 18288 32428
rect 19524 32444 19576 32496
rect 15108 32308 15160 32317
rect 14556 32240 14608 32292
rect 14832 32240 14884 32292
rect 15752 32240 15804 32292
rect 16580 32240 16632 32292
rect 19892 32240 19944 32292
rect 13084 32172 13136 32224
rect 13176 32172 13228 32224
rect 14004 32172 14056 32224
rect 15844 32172 15896 32224
rect 15936 32215 15988 32224
rect 15936 32181 15945 32215
rect 15945 32181 15979 32215
rect 15979 32181 15988 32215
rect 15936 32172 15988 32181
rect 16396 32215 16448 32224
rect 16396 32181 16405 32215
rect 16405 32181 16439 32215
rect 16439 32181 16448 32215
rect 16396 32172 16448 32181
rect 18604 32172 18656 32224
rect 20168 32172 20220 32224
rect 3422 32070 3474 32122
rect 3486 32070 3538 32122
rect 3550 32070 3602 32122
rect 3614 32070 3666 32122
rect 3678 32070 3730 32122
rect 8367 32070 8419 32122
rect 8431 32070 8483 32122
rect 8495 32070 8547 32122
rect 8559 32070 8611 32122
rect 8623 32070 8675 32122
rect 13312 32070 13364 32122
rect 13376 32070 13428 32122
rect 13440 32070 13492 32122
rect 13504 32070 13556 32122
rect 13568 32070 13620 32122
rect 18257 32070 18309 32122
rect 18321 32070 18373 32122
rect 18385 32070 18437 32122
rect 18449 32070 18501 32122
rect 18513 32070 18565 32122
rect 1860 31968 1912 32020
rect 4068 31968 4120 32020
rect 6920 31968 6972 32020
rect 2596 31900 2648 31952
rect 1124 31832 1176 31884
rect 1860 31764 1912 31816
rect 2136 31696 2188 31748
rect 3056 31807 3108 31816
rect 3056 31773 3065 31807
rect 3065 31773 3099 31807
rect 3099 31773 3108 31807
rect 3056 31764 3108 31773
rect 4620 31807 4672 31816
rect 4620 31773 4629 31807
rect 4629 31773 4663 31807
rect 4663 31773 4672 31807
rect 4620 31764 4672 31773
rect 5448 31832 5500 31884
rect 6276 31832 6328 31884
rect 3608 31739 3660 31748
rect 3608 31705 3617 31739
rect 3617 31705 3651 31739
rect 3651 31705 3660 31739
rect 3608 31696 3660 31705
rect 3792 31739 3844 31748
rect 3792 31705 3801 31739
rect 3801 31705 3835 31739
rect 3835 31705 3844 31739
rect 3792 31696 3844 31705
rect 5172 31739 5224 31748
rect 5172 31705 5181 31739
rect 5181 31705 5215 31739
rect 5215 31705 5224 31739
rect 5172 31696 5224 31705
rect 1676 31628 1728 31680
rect 2228 31628 2280 31680
rect 2688 31628 2740 31680
rect 5356 31764 5408 31816
rect 5448 31739 5500 31748
rect 5448 31705 5457 31739
rect 5457 31705 5491 31739
rect 5491 31705 5500 31739
rect 5448 31696 5500 31705
rect 7104 31764 7156 31816
rect 13084 31968 13136 32020
rect 14188 31968 14240 32020
rect 14280 31968 14332 32020
rect 9312 31832 9364 31884
rect 14464 31900 14516 31952
rect 14740 31943 14792 31952
rect 14740 31909 14749 31943
rect 14749 31909 14783 31943
rect 14783 31909 14792 31943
rect 14740 31900 14792 31909
rect 15200 31968 15252 32020
rect 15660 31968 15712 32020
rect 17960 31900 18012 31952
rect 15108 31875 15160 31884
rect 15108 31841 15142 31875
rect 15142 31841 15160 31875
rect 15108 31832 15160 31841
rect 15476 31832 15528 31884
rect 15844 31832 15896 31884
rect 16856 31832 16908 31884
rect 6276 31739 6328 31748
rect 6276 31705 6285 31739
rect 6285 31705 6319 31739
rect 6319 31705 6328 31739
rect 6276 31696 6328 31705
rect 7380 31696 7432 31748
rect 5816 31628 5868 31680
rect 7840 31628 7892 31680
rect 8852 31696 8904 31748
rect 9404 31696 9456 31748
rect 10140 31764 10192 31816
rect 11612 31807 11664 31816
rect 11612 31773 11621 31807
rect 11621 31773 11655 31807
rect 11655 31773 11664 31807
rect 11612 31764 11664 31773
rect 12532 31764 12584 31816
rect 13912 31764 13964 31816
rect 11796 31628 11848 31680
rect 11980 31696 12032 31748
rect 18604 31968 18656 32020
rect 19708 31968 19760 32020
rect 19064 31832 19116 31884
rect 12440 31671 12492 31680
rect 12440 31637 12449 31671
rect 12449 31637 12483 31671
rect 12483 31637 12492 31671
rect 12440 31628 12492 31637
rect 13084 31628 13136 31680
rect 16856 31696 16908 31748
rect 17592 31696 17644 31748
rect 17868 31696 17920 31748
rect 18420 31696 18472 31748
rect 14924 31628 14976 31680
rect 15752 31628 15804 31680
rect 15936 31628 15988 31680
rect 16304 31628 16356 31680
rect 16580 31628 16632 31680
rect 18604 31628 18656 31680
rect 18788 31696 18840 31748
rect 19064 31696 19116 31748
rect 19340 31696 19392 31748
rect 20628 31764 20680 31816
rect 19616 31696 19668 31748
rect 21916 31696 21968 31748
rect 19984 31628 20036 31680
rect 20260 31671 20312 31680
rect 20260 31637 20269 31671
rect 20269 31637 20303 31671
rect 20303 31637 20312 31671
rect 20260 31628 20312 31637
rect 5894 31526 5946 31578
rect 5958 31526 6010 31578
rect 6022 31526 6074 31578
rect 6086 31526 6138 31578
rect 6150 31526 6202 31578
rect 10839 31526 10891 31578
rect 10903 31526 10955 31578
rect 10967 31526 11019 31578
rect 11031 31526 11083 31578
rect 11095 31526 11147 31578
rect 15784 31526 15836 31578
rect 15848 31526 15900 31578
rect 15912 31526 15964 31578
rect 15976 31526 16028 31578
rect 16040 31526 16092 31578
rect 20729 31526 20781 31578
rect 20793 31526 20845 31578
rect 20857 31526 20909 31578
rect 20921 31526 20973 31578
rect 20985 31526 21037 31578
rect 1584 31424 1636 31476
rect 1952 31288 2004 31340
rect 1584 31220 1636 31272
rect 572 31152 624 31204
rect 3056 31356 3108 31408
rect 5356 31424 5408 31476
rect 5540 31356 5592 31408
rect 2228 31288 2280 31340
rect 2412 31288 2464 31340
rect 3332 31288 3384 31340
rect 4804 31288 4856 31340
rect 5080 31288 5132 31340
rect 4896 31263 4948 31272
rect 4896 31229 4905 31263
rect 4905 31229 4939 31263
rect 4939 31229 4948 31263
rect 4896 31220 4948 31229
rect 7104 31288 7156 31340
rect 7656 31424 7708 31476
rect 10416 31424 10468 31476
rect 11796 31424 11848 31476
rect 12072 31424 12124 31476
rect 12164 31424 12216 31476
rect 12532 31467 12584 31476
rect 12532 31433 12541 31467
rect 12541 31433 12575 31467
rect 12575 31433 12584 31467
rect 12532 31424 12584 31433
rect 13820 31424 13872 31476
rect 8208 31288 8260 31340
rect 10048 31331 10100 31340
rect 10048 31297 10057 31331
rect 10057 31297 10091 31331
rect 10091 31297 10100 31331
rect 10048 31288 10100 31297
rect 10324 31331 10376 31340
rect 10324 31297 10333 31331
rect 10333 31297 10367 31331
rect 10367 31297 10376 31331
rect 10324 31288 10376 31297
rect 11152 31288 11204 31340
rect 12348 31356 12400 31408
rect 12440 31356 12492 31408
rect 15476 31424 15528 31476
rect 11796 31331 11848 31340
rect 11796 31297 11803 31331
rect 11803 31297 11837 31331
rect 11837 31297 11848 31331
rect 11796 31288 11848 31297
rect 12532 31288 12584 31340
rect 12716 31288 12768 31340
rect 2412 31084 2464 31136
rect 7104 31152 7156 31204
rect 3240 31084 3292 31136
rect 3608 31084 3660 31136
rect 5356 31084 5408 31136
rect 7196 31084 7248 31136
rect 7380 31084 7432 31136
rect 8208 31084 8260 31136
rect 9404 31220 9456 31272
rect 12992 31220 13044 31272
rect 13176 31220 13228 31272
rect 13820 31263 13872 31272
rect 13820 31229 13829 31263
rect 13829 31229 13863 31263
rect 13863 31229 13872 31263
rect 13820 31220 13872 31229
rect 14004 31220 14056 31272
rect 14924 31356 14976 31408
rect 18788 31424 18840 31476
rect 20260 31424 20312 31476
rect 20628 31424 20680 31476
rect 21824 31424 21876 31476
rect 16304 31288 16356 31340
rect 17592 31288 17644 31340
rect 9772 31195 9824 31204
rect 9772 31161 9781 31195
rect 9781 31161 9815 31195
rect 9815 31161 9824 31195
rect 9772 31152 9824 31161
rect 9864 31152 9916 31204
rect 16580 31220 16632 31272
rect 18236 31220 18288 31272
rect 18512 31288 18564 31340
rect 18696 31331 18748 31340
rect 18696 31297 18705 31331
rect 18705 31297 18739 31331
rect 18739 31297 18748 31331
rect 18696 31288 18748 31297
rect 18788 31220 18840 31272
rect 19248 31288 19300 31340
rect 19064 31220 19116 31272
rect 10508 31084 10560 31136
rect 14188 31084 14240 31136
rect 15568 31152 15620 31204
rect 16948 31152 17000 31204
rect 19248 31195 19300 31204
rect 19248 31161 19257 31195
rect 19257 31161 19291 31195
rect 19291 31161 19300 31195
rect 19248 31152 19300 31161
rect 19616 31331 19668 31340
rect 19616 31297 19625 31331
rect 19625 31297 19659 31331
rect 19659 31297 19668 31331
rect 19616 31288 19668 31297
rect 19800 31288 19852 31340
rect 19984 31263 20036 31272
rect 19984 31229 19993 31263
rect 19993 31229 20027 31263
rect 20027 31229 20036 31263
rect 19984 31220 20036 31229
rect 16764 31127 16816 31136
rect 16764 31093 16773 31127
rect 16773 31093 16807 31127
rect 16807 31093 16816 31127
rect 16764 31084 16816 31093
rect 18420 31084 18472 31136
rect 18696 31084 18748 31136
rect 19708 31084 19760 31136
rect 21732 31152 21784 31204
rect 20444 31127 20496 31136
rect 20444 31093 20453 31127
rect 20453 31093 20487 31127
rect 20487 31093 20496 31127
rect 20444 31084 20496 31093
rect 3422 30982 3474 31034
rect 3486 30982 3538 31034
rect 3550 30982 3602 31034
rect 3614 30982 3666 31034
rect 3678 30982 3730 31034
rect 8367 30982 8419 31034
rect 8431 30982 8483 31034
rect 8495 30982 8547 31034
rect 8559 30982 8611 31034
rect 8623 30982 8675 31034
rect 13312 30982 13364 31034
rect 13376 30982 13428 31034
rect 13440 30982 13492 31034
rect 13504 30982 13556 31034
rect 13568 30982 13620 31034
rect 18257 30982 18309 31034
rect 18321 30982 18373 31034
rect 18385 30982 18437 31034
rect 18449 30982 18501 31034
rect 18513 30982 18565 31034
rect 664 30880 716 30932
rect 4160 30880 4212 30932
rect 5632 30880 5684 30932
rect 8208 30880 8260 30932
rect 9404 30880 9456 30932
rect 10324 30880 10376 30932
rect 1860 30812 1912 30864
rect 1308 30608 1360 30660
rect 2596 30787 2648 30796
rect 2596 30753 2630 30787
rect 2630 30753 2648 30787
rect 2596 30744 2648 30753
rect 7840 30744 7892 30796
rect 2504 30719 2556 30728
rect 2504 30685 2513 30719
rect 2513 30685 2547 30719
rect 2547 30685 2556 30719
rect 2504 30676 2556 30685
rect 2780 30719 2832 30728
rect 2780 30685 2789 30719
rect 2789 30685 2823 30719
rect 2823 30685 2832 30719
rect 2780 30676 2832 30685
rect 3424 30676 3476 30728
rect 5080 30676 5132 30728
rect 5356 30676 5408 30728
rect 6736 30676 6788 30728
rect 8852 30812 8904 30864
rect 9312 30744 9364 30796
rect 11152 30880 11204 30932
rect 11244 30880 11296 30932
rect 8300 30676 8352 30728
rect 8484 30719 8536 30728
rect 8484 30685 8493 30719
rect 8493 30685 8527 30719
rect 8527 30685 8536 30719
rect 8484 30676 8536 30685
rect 3608 30540 3660 30592
rect 3792 30540 3844 30592
rect 5172 30540 5224 30592
rect 7196 30608 7248 30660
rect 7840 30608 7892 30660
rect 7932 30608 7984 30660
rect 9772 30676 9824 30728
rect 10048 30676 10100 30728
rect 10600 30676 10652 30728
rect 11888 30744 11940 30796
rect 12256 30744 12308 30796
rect 13360 30880 13412 30932
rect 13728 30880 13780 30932
rect 13820 30880 13872 30932
rect 15016 30880 15068 30932
rect 16212 30880 16264 30932
rect 16764 30880 16816 30932
rect 14740 30855 14792 30864
rect 14740 30821 14749 30855
rect 14749 30821 14783 30855
rect 14783 30821 14792 30855
rect 14740 30812 14792 30821
rect 15292 30787 15344 30796
rect 15292 30753 15301 30787
rect 15301 30753 15335 30787
rect 15335 30753 15344 30787
rect 15292 30744 15344 30753
rect 15660 30744 15712 30796
rect 16120 30744 16172 30796
rect 16580 30744 16632 30796
rect 11060 30719 11112 30728
rect 11060 30685 11069 30719
rect 11069 30685 11112 30719
rect 11060 30676 11112 30685
rect 12348 30676 12400 30728
rect 14188 30676 14240 30728
rect 11888 30608 11940 30660
rect 15016 30719 15068 30728
rect 15016 30685 15025 30719
rect 15025 30685 15059 30719
rect 15059 30685 15068 30719
rect 15016 30676 15068 30685
rect 15108 30719 15160 30728
rect 15108 30685 15142 30719
rect 15142 30685 15160 30719
rect 15108 30676 15160 30685
rect 16396 30719 16448 30728
rect 16396 30685 16405 30719
rect 16405 30685 16439 30719
rect 16439 30685 16448 30719
rect 16396 30676 16448 30685
rect 19248 30923 19300 30932
rect 19248 30889 19257 30923
rect 19257 30889 19291 30923
rect 19291 30889 19300 30923
rect 19248 30880 19300 30889
rect 17684 30744 17736 30796
rect 16304 30608 16356 30660
rect 17776 30719 17828 30728
rect 17776 30685 17785 30719
rect 17785 30685 17819 30719
rect 17819 30685 17828 30719
rect 17776 30676 17828 30685
rect 17960 30676 18012 30728
rect 18144 30719 18196 30728
rect 18144 30685 18153 30719
rect 18153 30685 18187 30719
rect 18187 30685 18196 30719
rect 18144 30676 18196 30685
rect 18788 30719 18840 30728
rect 18788 30685 18797 30719
rect 18797 30685 18831 30719
rect 18831 30685 18840 30719
rect 18788 30676 18840 30685
rect 18236 30608 18288 30660
rect 19524 30676 19576 30728
rect 19800 30676 19852 30728
rect 21272 30608 21324 30660
rect 7564 30540 7616 30592
rect 8116 30583 8168 30592
rect 8116 30549 8125 30583
rect 8125 30549 8159 30583
rect 8159 30549 8168 30583
rect 8116 30540 8168 30549
rect 8576 30583 8628 30592
rect 8576 30549 8585 30583
rect 8585 30549 8619 30583
rect 8619 30549 8628 30583
rect 8576 30540 8628 30549
rect 10416 30583 10468 30592
rect 10416 30549 10425 30583
rect 10425 30549 10459 30583
rect 10459 30549 10468 30583
rect 10416 30540 10468 30549
rect 10600 30540 10652 30592
rect 11336 30540 11388 30592
rect 11796 30583 11848 30592
rect 11796 30549 11805 30583
rect 11805 30549 11839 30583
rect 11839 30549 11848 30583
rect 11796 30540 11848 30549
rect 13084 30540 13136 30592
rect 16764 30540 16816 30592
rect 17316 30583 17368 30592
rect 17316 30549 17325 30583
rect 17325 30549 17359 30583
rect 17359 30549 17368 30583
rect 17316 30540 17368 30549
rect 17592 30583 17644 30592
rect 17592 30549 17601 30583
rect 17601 30549 17635 30583
rect 17635 30549 17644 30583
rect 17592 30540 17644 30549
rect 17684 30540 17736 30592
rect 19984 30540 20036 30592
rect 5894 30438 5946 30490
rect 5958 30438 6010 30490
rect 6022 30438 6074 30490
rect 6086 30438 6138 30490
rect 6150 30438 6202 30490
rect 10839 30438 10891 30490
rect 10903 30438 10955 30490
rect 10967 30438 11019 30490
rect 11031 30438 11083 30490
rect 11095 30438 11147 30490
rect 15784 30438 15836 30490
rect 15848 30438 15900 30490
rect 15912 30438 15964 30490
rect 15976 30438 16028 30490
rect 16040 30438 16092 30490
rect 20729 30438 20781 30490
rect 20793 30438 20845 30490
rect 20857 30438 20909 30490
rect 20921 30438 20973 30490
rect 20985 30438 21037 30490
rect 1400 30268 1452 30320
rect 756 30200 808 30252
rect 4804 30336 4856 30388
rect 2978 30243 3030 30252
rect 2978 30209 2991 30243
rect 2991 30209 3025 30243
rect 3025 30209 3030 30243
rect 2978 30200 3030 30209
rect 3976 30243 4028 30252
rect 3976 30209 3985 30243
rect 3985 30209 4019 30243
rect 4019 30209 4028 30243
rect 3976 30200 4028 30209
rect 4344 30200 4396 30252
rect 5172 30243 5224 30252
rect 5172 30209 5181 30243
rect 5181 30209 5215 30243
rect 5215 30209 5224 30243
rect 5172 30200 5224 30209
rect 2228 30175 2280 30184
rect 2228 30141 2237 30175
rect 2237 30141 2271 30175
rect 2271 30141 2280 30175
rect 2228 30132 2280 30141
rect 2596 30064 2648 30116
rect 2688 30107 2740 30116
rect 2688 30073 2697 30107
rect 2697 30073 2731 30107
rect 2731 30073 2740 30107
rect 2688 30064 2740 30073
rect 1400 29996 1452 30048
rect 1768 30039 1820 30048
rect 1768 30005 1777 30039
rect 1777 30005 1811 30039
rect 1811 30005 1820 30039
rect 1768 29996 1820 30005
rect 3222 30175 3274 30184
rect 3222 30141 3235 30175
rect 3235 30141 3269 30175
rect 3269 30141 3274 30175
rect 3222 30132 3274 30141
rect 4160 30175 4212 30184
rect 4160 30141 4169 30175
rect 4169 30141 4203 30175
rect 4203 30141 4212 30175
rect 4160 30132 4212 30141
rect 3976 30064 4028 30116
rect 4620 30107 4672 30116
rect 4620 30073 4629 30107
rect 4629 30073 4663 30107
rect 4663 30073 4672 30107
rect 4620 30064 4672 30073
rect 5356 30132 5408 30184
rect 7196 30336 7248 30388
rect 7656 30336 7708 30388
rect 8300 30336 8352 30388
rect 9588 30336 9640 30388
rect 11612 30336 11664 30388
rect 11980 30336 12032 30388
rect 14004 30336 14056 30388
rect 14648 30336 14700 30388
rect 16304 30379 16356 30388
rect 16304 30345 16313 30379
rect 16313 30345 16347 30379
rect 16347 30345 16356 30379
rect 16304 30336 16356 30345
rect 17132 30336 17184 30388
rect 17408 30336 17460 30388
rect 17592 30336 17644 30388
rect 17776 30336 17828 30388
rect 18788 30336 18840 30388
rect 19616 30336 19668 30388
rect 19708 30336 19760 30388
rect 20168 30336 20220 30388
rect 6920 30268 6972 30320
rect 7012 30268 7064 30320
rect 7564 30200 7616 30252
rect 9128 30268 9180 30320
rect 8668 30243 8720 30252
rect 8668 30209 8677 30243
rect 8677 30209 8711 30243
rect 8711 30209 8720 30243
rect 8668 30200 8720 30209
rect 11980 30200 12032 30252
rect 13360 30200 13412 30252
rect 14004 30243 14056 30252
rect 14004 30209 14038 30243
rect 14038 30209 14056 30243
rect 14004 30200 14056 30209
rect 15108 30200 15160 30252
rect 6644 30064 6696 30116
rect 8484 30132 8536 30184
rect 8576 30175 8628 30184
rect 8576 30141 8585 30175
rect 8585 30141 8619 30175
rect 8619 30141 8628 30175
rect 8576 30132 8628 30141
rect 13084 30132 13136 30184
rect 13176 30175 13228 30184
rect 13176 30141 13185 30175
rect 13185 30141 13219 30175
rect 13219 30141 13228 30175
rect 13176 30132 13228 30141
rect 13912 30175 13964 30184
rect 13912 30141 13921 30175
rect 13921 30141 13955 30175
rect 13955 30141 13964 30175
rect 13912 30132 13964 30141
rect 5080 29996 5132 30048
rect 5264 29996 5316 30048
rect 6552 29996 6604 30048
rect 13636 30107 13688 30116
rect 13636 30073 13645 30107
rect 13645 30073 13679 30107
rect 13679 30073 13688 30107
rect 13636 30064 13688 30073
rect 8116 29996 8168 30048
rect 8760 29996 8812 30048
rect 9680 30039 9732 30048
rect 9680 30005 9689 30039
rect 9689 30005 9723 30039
rect 9723 30005 9732 30039
rect 9680 29996 9732 30005
rect 10048 29996 10100 30048
rect 10876 29996 10928 30048
rect 14832 29996 14884 30048
rect 16672 30243 16724 30252
rect 16672 30209 16681 30243
rect 16681 30209 16715 30243
rect 16715 30209 16724 30243
rect 16672 30200 16724 30209
rect 17316 30200 17368 30252
rect 18144 30243 18196 30252
rect 18144 30209 18153 30243
rect 18153 30209 18187 30243
rect 18187 30209 18196 30243
rect 18144 30200 18196 30209
rect 18972 30243 19024 30252
rect 18972 30209 18981 30243
rect 18981 30209 19015 30243
rect 19015 30209 19024 30243
rect 18972 30200 19024 30209
rect 19616 30243 19668 30252
rect 19616 30209 19625 30243
rect 19625 30209 19659 30243
rect 19659 30209 19668 30243
rect 19616 30200 19668 30209
rect 19708 30243 19760 30252
rect 19708 30209 19717 30243
rect 19717 30209 19751 30243
rect 19751 30209 19760 30243
rect 19708 30200 19760 30209
rect 20076 30132 20128 30184
rect 18696 29996 18748 30048
rect 18880 29996 18932 30048
rect 20076 29996 20128 30048
rect 20352 29996 20404 30048
rect 20444 30039 20496 30048
rect 20444 30005 20453 30039
rect 20453 30005 20487 30039
rect 20487 30005 20496 30039
rect 20444 29996 20496 30005
rect 3422 29894 3474 29946
rect 3486 29894 3538 29946
rect 3550 29894 3602 29946
rect 3614 29894 3666 29946
rect 3678 29894 3730 29946
rect 8367 29894 8419 29946
rect 8431 29894 8483 29946
rect 8495 29894 8547 29946
rect 8559 29894 8611 29946
rect 8623 29894 8675 29946
rect 13312 29894 13364 29946
rect 13376 29894 13428 29946
rect 13440 29894 13492 29946
rect 13504 29894 13556 29946
rect 13568 29894 13620 29946
rect 18257 29894 18309 29946
rect 18321 29894 18373 29946
rect 18385 29894 18437 29946
rect 18449 29894 18501 29946
rect 18513 29894 18565 29946
rect 2228 29792 2280 29844
rect 1032 29724 1084 29776
rect 1492 29656 1544 29708
rect 1676 29656 1728 29708
rect 2688 29792 2740 29844
rect 4528 29792 4580 29844
rect 4620 29792 4672 29844
rect 6920 29792 6972 29844
rect 13636 29792 13688 29844
rect 3792 29699 3844 29708
rect 3792 29665 3801 29699
rect 3801 29665 3835 29699
rect 3835 29665 3844 29699
rect 3792 29656 3844 29665
rect 1492 29563 1544 29572
rect 1492 29529 1501 29563
rect 1501 29529 1535 29563
rect 1535 29529 1544 29563
rect 1492 29520 1544 29529
rect 1676 29563 1728 29572
rect 1676 29529 1685 29563
rect 1685 29529 1719 29563
rect 1719 29529 1728 29563
rect 1676 29520 1728 29529
rect 2780 29588 2832 29640
rect 3148 29588 3200 29640
rect 3332 29631 3384 29640
rect 3332 29597 3341 29631
rect 3341 29597 3375 29631
rect 3375 29597 3384 29631
rect 3332 29588 3384 29597
rect 2228 29520 2280 29572
rect 3240 29520 3292 29572
rect 3976 29588 4028 29640
rect 6736 29656 6788 29708
rect 7196 29656 7248 29708
rect 4160 29520 4212 29572
rect 5264 29588 5316 29640
rect 4528 29520 4580 29572
rect 5172 29520 5224 29572
rect 6276 29631 6328 29640
rect 6276 29597 6285 29631
rect 6285 29597 6319 29631
rect 6319 29597 6328 29631
rect 6276 29588 6328 29597
rect 1032 29452 1084 29504
rect 2596 29452 2648 29504
rect 3332 29452 3384 29504
rect 4804 29452 4856 29504
rect 7196 29495 7248 29504
rect 7196 29461 7205 29495
rect 7205 29461 7239 29495
rect 7239 29461 7248 29495
rect 7196 29452 7248 29461
rect 8944 29656 8996 29708
rect 10416 29656 10468 29708
rect 11704 29656 11756 29708
rect 13544 29724 13596 29776
rect 14556 29792 14608 29844
rect 8208 29588 8260 29640
rect 9312 29631 9364 29640
rect 9312 29597 9319 29631
rect 9319 29597 9353 29631
rect 9353 29597 9364 29631
rect 9312 29588 9364 29597
rect 10876 29631 10928 29640
rect 10876 29597 10885 29631
rect 10885 29597 10919 29631
rect 10919 29597 10928 29631
rect 10876 29588 10928 29597
rect 11796 29588 11848 29640
rect 15568 29656 15620 29708
rect 17132 29792 17184 29844
rect 18144 29792 18196 29844
rect 18972 29792 19024 29844
rect 17592 29724 17644 29776
rect 18604 29656 18656 29708
rect 13176 29588 13228 29640
rect 14556 29631 14608 29640
rect 7380 29520 7432 29572
rect 8300 29520 8352 29572
rect 11244 29520 11296 29572
rect 14556 29597 14563 29631
rect 14563 29597 14597 29631
rect 14597 29597 14608 29631
rect 14556 29588 14608 29597
rect 14648 29520 14700 29572
rect 16948 29588 17000 29640
rect 7656 29452 7708 29504
rect 9864 29452 9916 29504
rect 10048 29495 10100 29504
rect 10048 29461 10057 29495
rect 10057 29461 10091 29495
rect 10091 29461 10100 29495
rect 10048 29452 10100 29461
rect 11612 29452 11664 29504
rect 11704 29495 11756 29504
rect 11704 29461 11713 29495
rect 11713 29461 11747 29495
rect 11747 29461 11756 29495
rect 11704 29452 11756 29461
rect 12440 29452 12492 29504
rect 12716 29452 12768 29504
rect 14556 29452 14608 29504
rect 15016 29452 15068 29504
rect 15476 29452 15528 29504
rect 18604 29452 18656 29504
rect 19524 29724 19576 29776
rect 19892 29792 19944 29844
rect 21272 29520 21324 29572
rect 5894 29350 5946 29402
rect 5958 29350 6010 29402
rect 6022 29350 6074 29402
rect 6086 29350 6138 29402
rect 6150 29350 6202 29402
rect 10839 29350 10891 29402
rect 10903 29350 10955 29402
rect 10967 29350 11019 29402
rect 11031 29350 11083 29402
rect 11095 29350 11147 29402
rect 15784 29350 15836 29402
rect 15848 29350 15900 29402
rect 15912 29350 15964 29402
rect 15976 29350 16028 29402
rect 16040 29350 16092 29402
rect 20729 29350 20781 29402
rect 20793 29350 20845 29402
rect 20857 29350 20909 29402
rect 20921 29350 20973 29402
rect 20985 29350 21037 29402
rect 1308 29248 1360 29300
rect 3884 29248 3936 29300
rect 3976 29248 4028 29300
rect 4252 29248 4304 29300
rect 4436 29291 4488 29300
rect 4436 29257 4445 29291
rect 4445 29257 4479 29291
rect 4479 29257 4488 29291
rect 4436 29248 4488 29257
rect 4712 29291 4764 29300
rect 4712 29257 4721 29291
rect 4721 29257 4755 29291
rect 4755 29257 4764 29291
rect 4712 29248 4764 29257
rect 4988 29248 5040 29300
rect 1032 29112 1084 29164
rect 2044 29180 2096 29232
rect 2044 29078 2096 29130
rect 2596 29112 2648 29164
rect 2964 29180 3016 29232
rect 7656 29248 7708 29300
rect 8208 29248 8260 29300
rect 2872 29155 2924 29164
rect 2872 29121 2881 29155
rect 2881 29121 2915 29155
rect 2915 29121 2924 29155
rect 2872 29112 2924 29121
rect 4252 29155 4304 29164
rect 4252 29121 4261 29155
rect 4261 29121 4295 29155
rect 4295 29121 4304 29155
rect 4252 29112 4304 29121
rect 572 28908 624 28960
rect 2504 28908 2556 28960
rect 3792 29044 3844 29096
rect 5448 29180 5500 29232
rect 4804 29044 4856 29096
rect 3884 29019 3936 29028
rect 3884 28985 3893 29019
rect 3893 28985 3927 29019
rect 3927 28985 3936 29019
rect 3884 28976 3936 28985
rect 7104 29180 7156 29232
rect 7196 29180 7248 29232
rect 7380 29185 7432 29232
rect 7380 29180 7405 29185
rect 7405 29180 7432 29185
rect 7564 29180 7616 29232
rect 9220 29248 9272 29300
rect 9680 29248 9732 29300
rect 9864 29248 9916 29300
rect 10508 29248 10560 29300
rect 11704 29248 11756 29300
rect 12256 29248 12308 29300
rect 13176 29248 13228 29300
rect 14740 29248 14792 29300
rect 17592 29248 17644 29300
rect 9404 29223 9456 29232
rect 9404 29189 9413 29223
rect 9413 29189 9447 29223
rect 9447 29189 9456 29223
rect 9404 29180 9456 29189
rect 10692 29180 10744 29232
rect 11336 29180 11388 29232
rect 2872 28908 2924 28960
rect 4804 28908 4856 28960
rect 6920 28976 6972 29028
rect 7012 28976 7064 29028
rect 17316 29180 17368 29232
rect 18880 29248 18932 29300
rect 19616 29248 19668 29300
rect 14096 29112 14148 29164
rect 17776 29112 17828 29164
rect 18880 29155 18932 29164
rect 18880 29121 18889 29155
rect 18889 29121 18923 29155
rect 18923 29121 18932 29155
rect 18880 29112 18932 29121
rect 19156 29155 19208 29164
rect 19156 29121 19165 29155
rect 19165 29121 19199 29155
rect 19199 29121 19208 29155
rect 19156 29112 19208 29121
rect 20168 29223 20220 29232
rect 20168 29189 20177 29223
rect 20177 29189 20211 29223
rect 20211 29189 20220 29223
rect 20168 29180 20220 29189
rect 10416 29019 10468 29028
rect 10416 28985 10425 29019
rect 10425 28985 10459 29019
rect 10459 28985 10468 29019
rect 10416 28976 10468 28985
rect 12716 29044 12768 29096
rect 14556 29087 14608 29096
rect 12256 28976 12308 29028
rect 6736 28908 6788 28960
rect 7104 28908 7156 28960
rect 10324 28908 10376 28960
rect 11244 28908 11296 28960
rect 11612 28908 11664 28960
rect 14556 29053 14565 29087
rect 14565 29053 14599 29087
rect 14599 29053 14608 29087
rect 14556 29044 14608 29053
rect 19248 29044 19300 29096
rect 19892 29112 19944 29164
rect 19800 29044 19852 29096
rect 17868 28976 17920 29028
rect 19156 28976 19208 29028
rect 14188 28951 14240 28960
rect 14188 28917 14197 28951
rect 14197 28917 14231 28951
rect 14231 28917 14240 28951
rect 14188 28908 14240 28917
rect 15476 28908 15528 28960
rect 20444 29019 20496 29028
rect 20444 28985 20453 29019
rect 20453 28985 20487 29019
rect 20487 28985 20496 29019
rect 20444 28976 20496 28985
rect 19616 28951 19668 28960
rect 19616 28917 19625 28951
rect 19625 28917 19659 28951
rect 19659 28917 19668 28951
rect 19616 28908 19668 28917
rect 19800 28951 19852 28960
rect 19800 28917 19809 28951
rect 19809 28917 19843 28951
rect 19843 28917 19852 28951
rect 19800 28908 19852 28917
rect 3422 28806 3474 28858
rect 3486 28806 3538 28858
rect 3550 28806 3602 28858
rect 3614 28806 3666 28858
rect 3678 28806 3730 28858
rect 8367 28806 8419 28858
rect 8431 28806 8483 28858
rect 8495 28806 8547 28858
rect 8559 28806 8611 28858
rect 8623 28806 8675 28858
rect 13312 28806 13364 28858
rect 13376 28806 13428 28858
rect 13440 28806 13492 28858
rect 13504 28806 13556 28858
rect 13568 28806 13620 28858
rect 18257 28806 18309 28858
rect 18321 28806 18373 28858
rect 18385 28806 18437 28858
rect 18449 28806 18501 28858
rect 18513 28806 18565 28858
rect 1216 28568 1268 28620
rect 2596 28611 2648 28620
rect 2596 28577 2605 28611
rect 2605 28577 2639 28611
rect 2639 28577 2648 28611
rect 2596 28568 2648 28577
rect 4436 28704 4488 28756
rect 4896 28704 4948 28756
rect 5540 28636 5592 28688
rect 5724 28636 5776 28688
rect 6828 28704 6880 28756
rect 6920 28704 6972 28756
rect 7932 28636 7984 28688
rect 756 28500 808 28552
rect 3240 28543 3292 28552
rect 3240 28509 3249 28543
rect 3249 28509 3283 28543
rect 3283 28509 3292 28543
rect 3240 28500 3292 28509
rect 4620 28500 4672 28552
rect 5356 28500 5408 28552
rect 5448 28500 5500 28552
rect 5724 28543 5776 28552
rect 5724 28509 5733 28543
rect 5733 28509 5767 28543
rect 5767 28509 5776 28543
rect 5724 28500 5776 28509
rect 6460 28543 6512 28552
rect 6460 28509 6469 28543
rect 6469 28509 6503 28543
rect 6503 28509 6512 28543
rect 6460 28500 6512 28509
rect 6552 28543 6604 28552
rect 7104 28568 7156 28620
rect 8760 28704 8812 28756
rect 12900 28704 12952 28756
rect 13544 28704 13596 28756
rect 14188 28704 14240 28756
rect 14832 28568 14884 28620
rect 15476 28568 15528 28620
rect 18880 28704 18932 28756
rect 19248 28747 19300 28756
rect 19248 28713 19257 28747
rect 19257 28713 19291 28747
rect 19291 28713 19300 28747
rect 19248 28704 19300 28713
rect 19616 28704 19668 28756
rect 20076 28704 20128 28756
rect 19708 28636 19760 28688
rect 6552 28509 6586 28543
rect 6586 28509 6604 28543
rect 6552 28500 6604 28509
rect 8668 28500 8720 28552
rect 9588 28500 9640 28552
rect 10048 28500 10100 28552
rect 10324 28500 10376 28552
rect 11704 28500 11756 28552
rect 11888 28500 11940 28552
rect 12716 28500 12768 28552
rect 12992 28500 13044 28552
rect 13084 28500 13136 28552
rect 15200 28500 15252 28552
rect 1676 28475 1728 28484
rect 1676 28441 1685 28475
rect 1685 28441 1719 28475
rect 1719 28441 1728 28475
rect 1676 28432 1728 28441
rect 940 28364 992 28416
rect 2596 28364 2648 28416
rect 4988 28407 5040 28416
rect 4988 28373 4997 28407
rect 4997 28373 5031 28407
rect 5031 28373 5040 28407
rect 4988 28364 5040 28373
rect 8300 28364 8352 28416
rect 9404 28407 9456 28416
rect 9404 28373 9413 28407
rect 9413 28373 9447 28407
rect 9447 28373 9456 28407
rect 9404 28364 9456 28373
rect 14280 28432 14332 28484
rect 10508 28407 10560 28416
rect 10508 28373 10517 28407
rect 10517 28373 10551 28407
rect 10551 28373 10560 28407
rect 10508 28364 10560 28373
rect 10692 28407 10744 28416
rect 10692 28373 10701 28407
rect 10701 28373 10735 28407
rect 10735 28373 10744 28407
rect 10692 28364 10744 28373
rect 11612 28364 11664 28416
rect 11980 28364 12032 28416
rect 12716 28364 12768 28416
rect 14648 28364 14700 28416
rect 15016 28364 15068 28416
rect 15200 28364 15252 28416
rect 16672 28500 16724 28552
rect 16304 28475 16356 28484
rect 16304 28441 16327 28475
rect 16327 28441 16356 28475
rect 16304 28432 16356 28441
rect 19156 28432 19208 28484
rect 19984 28500 20036 28552
rect 18052 28364 18104 28416
rect 19984 28364 20036 28416
rect 20076 28364 20128 28416
rect 20444 28407 20496 28416
rect 20444 28373 20453 28407
rect 20453 28373 20487 28407
rect 20487 28373 20496 28407
rect 20444 28364 20496 28373
rect 5894 28262 5946 28314
rect 5958 28262 6010 28314
rect 6022 28262 6074 28314
rect 6086 28262 6138 28314
rect 6150 28262 6202 28314
rect 10839 28262 10891 28314
rect 10903 28262 10955 28314
rect 10967 28262 11019 28314
rect 11031 28262 11083 28314
rect 11095 28262 11147 28314
rect 15784 28262 15836 28314
rect 15848 28262 15900 28314
rect 15912 28262 15964 28314
rect 15976 28262 16028 28314
rect 16040 28262 16092 28314
rect 20729 28262 20781 28314
rect 20793 28262 20845 28314
rect 20857 28262 20909 28314
rect 20921 28262 20973 28314
rect 20985 28262 21037 28314
rect 1400 28160 1452 28212
rect 2044 28160 2096 28212
rect 2412 28160 2464 28212
rect 4252 28160 4304 28212
rect 5908 28160 5960 28212
rect 6552 28160 6604 28212
rect 8668 28160 8720 28212
rect 296 28092 348 28144
rect 1308 28092 1360 28144
rect 3976 28092 4028 28144
rect 5080 28092 5132 28144
rect 5356 28092 5408 28144
rect 8208 28092 8260 28144
rect 2044 28024 2096 28076
rect 3056 28024 3108 28076
rect 756 27956 808 28008
rect 1400 27999 1452 28008
rect 1400 27965 1409 27999
rect 1409 27965 1443 27999
rect 1443 27965 1452 27999
rect 1400 27956 1452 27965
rect 4804 28067 4856 28076
rect 4804 28033 4811 28067
rect 4811 28033 4845 28067
rect 4845 28033 4856 28067
rect 4804 28024 4856 28033
rect 3056 27931 3108 27940
rect 3056 27897 3065 27931
rect 3065 27897 3099 27931
rect 3099 27897 3108 27931
rect 3056 27888 3108 27897
rect 1032 27820 1084 27872
rect 2412 27863 2464 27872
rect 2412 27829 2421 27863
rect 2421 27829 2455 27863
rect 2455 27829 2464 27863
rect 2412 27820 2464 27829
rect 4528 27999 4580 28008
rect 4528 27965 4537 27999
rect 4537 27965 4571 27999
rect 4571 27965 4580 27999
rect 4528 27956 4580 27965
rect 9128 28024 9180 28076
rect 9404 28092 9456 28144
rect 10324 28092 10376 28144
rect 10784 28092 10836 28144
rect 10876 28092 10928 28144
rect 11612 28092 11664 28144
rect 11704 28092 11756 28144
rect 15292 28160 15344 28212
rect 17960 28160 18012 28212
rect 19432 28160 19484 28212
rect 19708 28160 19760 28212
rect 12716 28067 12768 28076
rect 12716 28033 12725 28067
rect 12725 28033 12759 28067
rect 12759 28033 12768 28067
rect 12716 28024 12768 28033
rect 7288 27956 7340 28008
rect 7656 27956 7708 28008
rect 8944 27999 8996 28008
rect 8944 27965 8953 27999
rect 8953 27965 8987 27999
rect 8987 27965 8996 27999
rect 8944 27956 8996 27965
rect 11612 27956 11664 28008
rect 11704 27999 11756 28008
rect 11704 27965 11713 27999
rect 11713 27965 11747 27999
rect 11747 27965 11756 27999
rect 11704 27956 11756 27965
rect 12256 27956 12308 28008
rect 12440 27999 12492 28008
rect 12440 27965 12449 27999
rect 12449 27965 12483 27999
rect 12483 27965 12492 27999
rect 12440 27956 12492 27965
rect 12900 27956 12952 28008
rect 14188 28024 14240 28076
rect 14280 28067 14332 28076
rect 14280 28033 14289 28067
rect 14289 28033 14323 28067
rect 14323 28033 14332 28067
rect 14280 28024 14332 28033
rect 15292 28067 15344 28076
rect 15292 28033 15326 28067
rect 15326 28033 15344 28067
rect 15292 28024 15344 28033
rect 16304 28024 16356 28076
rect 16856 28024 16908 28076
rect 18788 28097 18840 28144
rect 18788 28092 18813 28097
rect 18813 28092 18840 28097
rect 19064 28092 19116 28144
rect 19616 28092 19668 28144
rect 19800 28092 19852 28144
rect 18880 28024 18932 28076
rect 20628 28024 20680 28076
rect 4160 27863 4212 27872
rect 4160 27829 4169 27863
rect 4169 27829 4203 27863
rect 4203 27829 4212 27863
rect 4160 27820 4212 27829
rect 13176 27888 13228 27940
rect 14372 27956 14424 28008
rect 14648 27956 14700 28008
rect 15476 27999 15528 28008
rect 15476 27965 15485 27999
rect 15485 27965 15519 27999
rect 15519 27965 15528 27999
rect 15476 27956 15528 27965
rect 6828 27820 6880 27872
rect 7288 27820 7340 27872
rect 13084 27820 13136 27872
rect 13912 27820 13964 27872
rect 14464 27820 14516 27872
rect 17868 27956 17920 28008
rect 17132 27820 17184 27872
rect 17592 27820 17644 27872
rect 17776 27820 17828 27872
rect 20444 27863 20496 27872
rect 20444 27829 20453 27863
rect 20453 27829 20487 27863
rect 20487 27829 20496 27863
rect 20444 27820 20496 27829
rect 3422 27718 3474 27770
rect 3486 27718 3538 27770
rect 3550 27718 3602 27770
rect 3614 27718 3666 27770
rect 3678 27718 3730 27770
rect 8367 27718 8419 27770
rect 8431 27718 8483 27770
rect 8495 27718 8547 27770
rect 8559 27718 8611 27770
rect 8623 27718 8675 27770
rect 13312 27718 13364 27770
rect 13376 27718 13428 27770
rect 13440 27718 13492 27770
rect 13504 27718 13556 27770
rect 13568 27718 13620 27770
rect 18257 27718 18309 27770
rect 18321 27718 18373 27770
rect 18385 27718 18437 27770
rect 18449 27718 18501 27770
rect 18513 27718 18565 27770
rect 3056 27616 3108 27668
rect 1032 27548 1084 27600
rect 2412 27480 2464 27532
rect 2964 27480 3016 27532
rect 3700 27480 3752 27532
rect 4988 27480 5040 27532
rect 7840 27659 7892 27668
rect 7840 27625 7849 27659
rect 7849 27625 7883 27659
rect 7883 27625 7892 27659
rect 7840 27616 7892 27625
rect 8116 27480 8168 27532
rect 10324 27616 10376 27668
rect 11520 27616 11572 27668
rect 12256 27616 12308 27668
rect 13176 27616 13228 27668
rect 14188 27616 14240 27668
rect 15476 27616 15528 27668
rect 17776 27616 17828 27668
rect 10508 27548 10560 27600
rect 12716 27548 12768 27600
rect 18052 27548 18104 27600
rect 19892 27616 19944 27668
rect 21272 27616 21324 27668
rect 21824 27616 21876 27668
rect 13636 27480 13688 27532
rect 15476 27523 15528 27532
rect 15476 27489 15485 27523
rect 15485 27489 15519 27523
rect 15519 27489 15528 27523
rect 15476 27480 15528 27489
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 1124 27344 1176 27396
rect 4620 27412 4672 27464
rect 5080 27412 5132 27464
rect 1952 27344 2004 27396
rect 2228 27387 2280 27396
rect 2228 27353 2237 27387
rect 2237 27353 2271 27387
rect 2271 27353 2280 27387
rect 2228 27344 2280 27353
rect 2320 27344 2372 27396
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 5816 27412 5868 27464
rect 6368 27412 6420 27464
rect 6828 27455 6880 27464
rect 6828 27421 6837 27455
rect 6837 27421 6871 27455
rect 6871 27421 6880 27455
rect 6828 27412 6880 27421
rect 7104 27455 7156 27464
rect 7104 27421 7111 27455
rect 7111 27421 7145 27455
rect 7145 27421 7156 27455
rect 7104 27412 7156 27421
rect 8392 27455 8444 27464
rect 8392 27421 8401 27455
rect 8401 27421 8435 27455
rect 8435 27421 8444 27455
rect 8392 27412 8444 27421
rect 8668 27412 8720 27464
rect 9128 27412 9180 27464
rect 10784 27412 10836 27464
rect 11520 27412 11572 27464
rect 12072 27412 12124 27464
rect 12532 27412 12584 27464
rect 2964 27319 3016 27328
rect 2964 27285 2973 27319
rect 2973 27285 3007 27319
rect 3007 27285 3016 27319
rect 2964 27276 3016 27285
rect 4068 27276 4120 27328
rect 4436 27276 4488 27328
rect 4712 27276 4764 27328
rect 4896 27276 4948 27328
rect 5356 27276 5408 27328
rect 12256 27344 12308 27396
rect 8300 27276 8352 27328
rect 11980 27276 12032 27328
rect 12164 27276 12216 27328
rect 16948 27455 17000 27464
rect 16948 27421 16957 27455
rect 16957 27421 16991 27455
rect 16991 27421 17000 27455
rect 16948 27412 17000 27421
rect 16304 27344 16356 27396
rect 17592 27455 17644 27464
rect 17592 27421 17601 27455
rect 17601 27421 17635 27455
rect 17635 27421 17644 27455
rect 17592 27412 17644 27421
rect 14188 27276 14240 27328
rect 17040 27319 17092 27328
rect 17040 27285 17049 27319
rect 17049 27285 17083 27319
rect 17083 27285 17092 27319
rect 17040 27276 17092 27285
rect 17776 27276 17828 27328
rect 18052 27276 18104 27328
rect 18788 27455 18840 27464
rect 18788 27421 18797 27455
rect 18797 27421 18831 27455
rect 18831 27421 18840 27455
rect 18788 27412 18840 27421
rect 21272 27480 21324 27532
rect 19984 27412 20036 27464
rect 20536 27387 20588 27396
rect 20536 27353 20545 27387
rect 20545 27353 20579 27387
rect 20579 27353 20588 27387
rect 20536 27344 20588 27353
rect 5894 27174 5946 27226
rect 5958 27174 6010 27226
rect 6022 27174 6074 27226
rect 6086 27174 6138 27226
rect 6150 27174 6202 27226
rect 10839 27174 10891 27226
rect 10903 27174 10955 27226
rect 10967 27174 11019 27226
rect 11031 27174 11083 27226
rect 11095 27174 11147 27226
rect 15784 27174 15836 27226
rect 15848 27174 15900 27226
rect 15912 27174 15964 27226
rect 15976 27174 16028 27226
rect 16040 27174 16092 27226
rect 20729 27174 20781 27226
rect 20793 27174 20845 27226
rect 20857 27174 20909 27226
rect 20921 27174 20973 27226
rect 20985 27174 21037 27226
rect 2228 27072 2280 27124
rect 6736 27072 6788 27124
rect 1308 27004 1360 27056
rect 756 26936 808 26988
rect 2412 26936 2464 26988
rect 1216 26732 1268 26784
rect 3240 26979 3292 26988
rect 3240 26945 3249 26979
rect 3249 26945 3283 26979
rect 3283 26945 3292 26979
rect 3240 26936 3292 26945
rect 3608 27004 3660 27056
rect 4160 27004 4212 27056
rect 5448 27004 5500 27056
rect 6920 27004 6972 27056
rect 4804 26979 4856 26988
rect 4804 26945 4813 26979
rect 4813 26945 4847 26979
rect 4847 26945 4856 26979
rect 4804 26936 4856 26945
rect 5172 26979 5224 26988
rect 5172 26945 5195 26979
rect 5195 26945 5224 26979
rect 5172 26936 5224 26945
rect 5356 26936 5408 26988
rect 5816 26936 5868 26988
rect 8392 27072 8444 27124
rect 9956 27072 10008 27124
rect 10600 27072 10652 27124
rect 8116 27004 8168 27056
rect 8760 27004 8812 27056
rect 7564 26979 7616 26988
rect 7564 26945 7573 26979
rect 7573 26945 7607 26979
rect 7607 26945 7616 26979
rect 7564 26936 7616 26945
rect 7932 26979 7984 26988
rect 7932 26945 7941 26979
rect 7941 26945 7975 26979
rect 7975 26945 7984 26979
rect 7932 26936 7984 26945
rect 3056 26868 3108 26920
rect 3700 26868 3752 26920
rect 3884 26868 3936 26920
rect 7840 26868 7892 26920
rect 9404 26868 9456 26920
rect 10692 27004 10744 27056
rect 13820 27072 13872 27124
rect 13912 27072 13964 27124
rect 14096 27072 14148 27124
rect 16304 27072 16356 27124
rect 16948 27072 17000 27124
rect 12072 27004 12124 27056
rect 12716 27004 12768 27056
rect 13912 26979 13964 26988
rect 13912 26945 13921 26979
rect 13921 26945 13955 26979
rect 13955 26945 13964 26979
rect 13912 26936 13964 26945
rect 14188 26979 14240 26988
rect 14188 26945 14197 26979
rect 14197 26945 14231 26979
rect 14231 26945 14240 26979
rect 14188 26936 14240 26945
rect 15200 26936 15252 26988
rect 17040 27004 17092 27056
rect 18788 27072 18840 27124
rect 18972 27072 19024 27124
rect 19156 27115 19208 27124
rect 19156 27081 19165 27115
rect 19165 27081 19199 27115
rect 19199 27081 19208 27115
rect 19156 27072 19208 27081
rect 19340 27072 19392 27124
rect 19984 27072 20036 27124
rect 21548 27072 21600 27124
rect 17868 26936 17920 26988
rect 10968 26868 11020 26920
rect 3148 26843 3200 26852
rect 3148 26809 3157 26843
rect 3157 26809 3191 26843
rect 3191 26809 3200 26843
rect 3148 26800 3200 26809
rect 5356 26843 5408 26852
rect 5356 26809 5365 26843
rect 5365 26809 5399 26843
rect 5399 26809 5408 26843
rect 5356 26800 5408 26809
rect 4068 26732 4120 26784
rect 10508 26732 10560 26784
rect 10968 26732 11020 26784
rect 11060 26775 11112 26784
rect 11060 26741 11069 26775
rect 11069 26741 11103 26775
rect 11103 26741 11112 26775
rect 11060 26732 11112 26741
rect 12440 26868 12492 26920
rect 12256 26800 12308 26852
rect 12348 26732 12400 26784
rect 13636 26843 13688 26852
rect 13636 26809 13645 26843
rect 13645 26809 13679 26843
rect 13679 26809 13688 26843
rect 13636 26800 13688 26809
rect 14556 26732 14608 26784
rect 16948 26911 17000 26920
rect 16948 26877 16957 26911
rect 16957 26877 16991 26911
rect 16991 26877 17000 26911
rect 16948 26868 17000 26877
rect 18604 26911 18656 26920
rect 18604 26877 18613 26911
rect 18613 26877 18647 26911
rect 18647 26877 18656 26911
rect 18604 26868 18656 26877
rect 18788 26868 18840 26920
rect 15292 26732 15344 26784
rect 17040 26732 17092 26784
rect 17316 26732 17368 26784
rect 19064 26800 19116 26852
rect 21548 26868 21600 26920
rect 21916 26868 21968 26920
rect 17684 26732 17736 26784
rect 17868 26732 17920 26784
rect 19708 26732 19760 26784
rect 19892 26775 19944 26784
rect 19892 26741 19901 26775
rect 19901 26741 19935 26775
rect 19935 26741 19944 26775
rect 19892 26732 19944 26741
rect 20628 26732 20680 26784
rect 3422 26630 3474 26682
rect 3486 26630 3538 26682
rect 3550 26630 3602 26682
rect 3614 26630 3666 26682
rect 3678 26630 3730 26682
rect 8367 26630 8419 26682
rect 8431 26630 8483 26682
rect 8495 26630 8547 26682
rect 8559 26630 8611 26682
rect 8623 26630 8675 26682
rect 13312 26630 13364 26682
rect 13376 26630 13428 26682
rect 13440 26630 13492 26682
rect 13504 26630 13556 26682
rect 13568 26630 13620 26682
rect 18257 26630 18309 26682
rect 18321 26630 18373 26682
rect 18385 26630 18437 26682
rect 18449 26630 18501 26682
rect 18513 26630 18565 26682
rect 1308 26528 1360 26580
rect 3240 26528 3292 26580
rect 4804 26528 4856 26580
rect 4896 26528 4948 26580
rect 7104 26528 7156 26580
rect 7288 26528 7340 26580
rect 7564 26528 7616 26580
rect 9128 26528 9180 26580
rect 10140 26528 10192 26580
rect 13636 26571 13688 26580
rect 13636 26537 13645 26571
rect 13645 26537 13679 26571
rect 13679 26537 13688 26571
rect 13636 26528 13688 26537
rect 14832 26528 14884 26580
rect 17316 26528 17368 26580
rect 17868 26528 17920 26580
rect 18052 26528 18104 26580
rect 3056 26503 3108 26512
rect 3056 26469 3065 26503
rect 3065 26469 3099 26503
rect 3099 26469 3108 26503
rect 3056 26460 3108 26469
rect 3976 26460 4028 26512
rect 5448 26460 5500 26512
rect 7012 26460 7064 26512
rect 11980 26503 12032 26512
rect 11980 26469 11989 26503
rect 11989 26469 12023 26503
rect 12023 26469 12032 26503
rect 11980 26460 12032 26469
rect 1308 26324 1360 26376
rect 1768 26367 1820 26376
rect 1768 26333 1775 26367
rect 1775 26333 1809 26367
rect 1809 26333 1820 26367
rect 1768 26324 1820 26333
rect 3056 26324 3108 26376
rect 3148 26367 3200 26376
rect 3148 26333 3157 26367
rect 3157 26333 3191 26367
rect 3191 26333 3200 26367
rect 3148 26324 3200 26333
rect 6828 26392 6880 26444
rect 11060 26392 11112 26444
rect 16212 26392 16264 26444
rect 16580 26392 16632 26444
rect 4528 26367 4580 26376
rect 4528 26333 4537 26367
rect 4537 26333 4571 26367
rect 4571 26333 4580 26367
rect 4528 26324 4580 26333
rect 4712 26324 4764 26376
rect 8668 26324 8720 26376
rect 7564 26256 7616 26308
rect 8024 26256 8076 26308
rect 8116 26256 8168 26308
rect 10968 26367 11020 26376
rect 10968 26333 10977 26367
rect 10977 26333 11011 26367
rect 11011 26333 11020 26367
rect 10968 26324 11020 26333
rect 10324 26256 10376 26308
rect 10600 26256 10652 26308
rect 11796 26324 11848 26376
rect 12532 26324 12584 26376
rect 12900 26367 12952 26376
rect 1584 26188 1636 26240
rect 2044 26188 2096 26240
rect 2228 26188 2280 26240
rect 2504 26231 2556 26240
rect 2504 26197 2513 26231
rect 2513 26197 2547 26231
rect 2547 26197 2556 26231
rect 2504 26188 2556 26197
rect 2596 26188 2648 26240
rect 3516 26188 3568 26240
rect 3608 26188 3660 26240
rect 4988 26188 5040 26240
rect 5632 26188 5684 26240
rect 7012 26188 7064 26240
rect 9404 26188 9456 26240
rect 10048 26188 10100 26240
rect 11704 26256 11756 26308
rect 12900 26333 12907 26367
rect 12907 26333 12941 26367
rect 12941 26333 12952 26367
rect 12900 26324 12952 26333
rect 14556 26324 14608 26376
rect 15200 26324 15252 26376
rect 16764 26367 16816 26376
rect 16764 26333 16773 26367
rect 16773 26333 16807 26367
rect 16807 26333 16816 26367
rect 16764 26324 16816 26333
rect 16948 26367 17000 26376
rect 16948 26333 16957 26367
rect 16957 26333 16991 26367
rect 16991 26333 17000 26367
rect 16948 26324 17000 26333
rect 17040 26324 17092 26376
rect 17684 26367 17736 26376
rect 17684 26333 17693 26367
rect 17693 26333 17727 26367
rect 17727 26333 17736 26367
rect 17684 26324 17736 26333
rect 13084 26256 13136 26308
rect 14372 26256 14424 26308
rect 15016 26256 15068 26308
rect 16396 26256 16448 26308
rect 18144 26324 18196 26376
rect 18604 26528 18656 26580
rect 18788 26460 18840 26512
rect 19340 26460 19392 26512
rect 20076 26460 20128 26512
rect 20260 26460 20312 26512
rect 18512 26367 18564 26376
rect 18512 26333 18521 26367
rect 18521 26333 18555 26367
rect 18555 26333 18564 26367
rect 18512 26324 18564 26333
rect 18788 26367 18840 26376
rect 18788 26333 18797 26367
rect 18797 26333 18831 26367
rect 18831 26333 18840 26367
rect 18788 26324 18840 26333
rect 18880 26324 18932 26376
rect 20260 26367 20312 26376
rect 11612 26188 11664 26240
rect 11888 26188 11940 26240
rect 11980 26188 12032 26240
rect 12716 26188 12768 26240
rect 13176 26188 13228 26240
rect 15660 26188 15712 26240
rect 16488 26231 16540 26240
rect 16488 26197 16497 26231
rect 16497 26197 16531 26231
rect 16531 26197 16540 26231
rect 16488 26188 16540 26197
rect 20260 26333 20269 26367
rect 20269 26333 20303 26367
rect 20303 26333 20312 26367
rect 20260 26324 20312 26333
rect 21272 26324 21324 26376
rect 20076 26188 20128 26240
rect 20444 26188 20496 26240
rect 20536 26231 20588 26240
rect 20536 26197 20545 26231
rect 20545 26197 20579 26231
rect 20579 26197 20588 26231
rect 20536 26188 20588 26197
rect 20720 26188 20772 26240
rect 21916 26188 21968 26240
rect 388 26120 440 26172
rect 848 26120 900 26172
rect 5894 26086 5946 26138
rect 5958 26086 6010 26138
rect 6022 26086 6074 26138
rect 6086 26086 6138 26138
rect 6150 26086 6202 26138
rect 10839 26086 10891 26138
rect 10903 26086 10955 26138
rect 10967 26086 11019 26138
rect 11031 26086 11083 26138
rect 11095 26086 11147 26138
rect 15784 26086 15836 26138
rect 15848 26086 15900 26138
rect 15912 26086 15964 26138
rect 15976 26086 16028 26138
rect 16040 26086 16092 26138
rect 20729 26086 20781 26138
rect 20793 26086 20845 26138
rect 20857 26086 20909 26138
rect 20921 26086 20973 26138
rect 20985 26086 21037 26138
rect 1676 25984 1728 26036
rect 2320 25984 2372 26036
rect 2596 25984 2648 26036
rect 5172 25984 5224 26036
rect 5264 25984 5316 26036
rect 5540 25984 5592 26036
rect 5632 25984 5684 26036
rect 5816 25984 5868 26036
rect 6276 25984 6328 26036
rect 1952 25916 2004 25968
rect 2228 25959 2280 25968
rect 2228 25925 2237 25959
rect 2237 25925 2271 25959
rect 2271 25925 2280 25959
rect 2228 25916 2280 25925
rect 2872 25916 2924 25968
rect 756 25848 808 25900
rect 2504 25848 2556 25900
rect 3240 25848 3292 25900
rect 3700 25848 3752 25900
rect 4160 25916 4212 25968
rect 4528 25848 4580 25900
rect 5172 25891 5224 25900
rect 5172 25857 5179 25891
rect 5179 25857 5213 25891
rect 5213 25857 5224 25891
rect 5172 25848 5224 25857
rect 7104 25916 7156 25968
rect 7840 25984 7892 26036
rect 9220 25984 9272 26036
rect 9404 26027 9456 26036
rect 9404 25993 9413 26027
rect 9413 25993 9447 26027
rect 9447 25993 9456 26027
rect 9404 25984 9456 25993
rect 7932 25916 7984 25968
rect 8300 25916 8352 25968
rect 10048 25984 10100 26036
rect 11520 25984 11572 26036
rect 7748 25891 7800 25900
rect 7748 25857 7757 25891
rect 7757 25857 7800 25891
rect 3148 25687 3200 25696
rect 3148 25653 3157 25687
rect 3157 25653 3191 25687
rect 3191 25653 3200 25687
rect 3148 25644 3200 25653
rect 4804 25780 4856 25832
rect 7748 25848 7800 25857
rect 7012 25780 7064 25832
rect 7288 25780 7340 25832
rect 4528 25687 4580 25696
rect 4528 25653 4537 25687
rect 4537 25653 4571 25687
rect 4571 25653 4580 25687
rect 4528 25644 4580 25653
rect 5172 25644 5224 25696
rect 5816 25644 5868 25696
rect 7012 25687 7064 25696
rect 7012 25653 7021 25687
rect 7021 25653 7055 25687
rect 7055 25653 7064 25687
rect 7012 25644 7064 25653
rect 8208 25644 8260 25696
rect 10140 25959 10192 25968
rect 10140 25925 10149 25959
rect 10149 25925 10183 25959
rect 10183 25925 10192 25959
rect 10140 25916 10192 25925
rect 11244 25916 11296 25968
rect 12348 25984 12400 26036
rect 12900 25984 12952 26036
rect 12164 25916 12216 25968
rect 10692 25848 10744 25900
rect 12532 25848 12584 25900
rect 13728 25916 13780 25968
rect 14740 25984 14792 26036
rect 15016 25984 15068 26036
rect 15108 25916 15160 25968
rect 15476 25916 15528 25968
rect 16212 25984 16264 26036
rect 16764 25984 16816 26036
rect 18788 25984 18840 26036
rect 16856 25852 16908 25904
rect 18696 25891 18748 25900
rect 18696 25857 18730 25891
rect 18730 25857 18748 25891
rect 12716 25755 12768 25764
rect 12716 25721 12725 25755
rect 12725 25721 12759 25755
rect 12759 25721 12768 25755
rect 13360 25780 13412 25832
rect 12716 25712 12768 25721
rect 9220 25644 9272 25696
rect 10600 25644 10652 25696
rect 10692 25687 10744 25696
rect 10692 25653 10701 25687
rect 10701 25653 10735 25687
rect 10735 25653 10744 25687
rect 10692 25644 10744 25653
rect 11796 25644 11848 25696
rect 12164 25644 12216 25696
rect 18696 25848 18748 25857
rect 13728 25823 13780 25832
rect 13728 25789 13737 25823
rect 13737 25789 13771 25823
rect 13771 25789 13780 25823
rect 13728 25780 13780 25789
rect 14648 25780 14700 25832
rect 15108 25780 15160 25832
rect 15292 25780 15344 25832
rect 15568 25780 15620 25832
rect 16396 25780 16448 25832
rect 18144 25780 18196 25832
rect 13728 25644 13780 25696
rect 17776 25712 17828 25764
rect 14740 25687 14792 25696
rect 14740 25653 14749 25687
rect 14749 25653 14783 25687
rect 14783 25653 14792 25687
rect 14740 25644 14792 25653
rect 16764 25644 16816 25696
rect 20444 25687 20496 25696
rect 20444 25653 20453 25687
rect 20453 25653 20487 25687
rect 20487 25653 20496 25687
rect 20444 25644 20496 25653
rect 3422 25542 3474 25594
rect 3486 25542 3538 25594
rect 3550 25542 3602 25594
rect 3614 25542 3666 25594
rect 3678 25542 3730 25594
rect 8367 25542 8419 25594
rect 8431 25542 8483 25594
rect 8495 25542 8547 25594
rect 8559 25542 8611 25594
rect 8623 25542 8675 25594
rect 13312 25542 13364 25594
rect 13376 25542 13428 25594
rect 13440 25542 13492 25594
rect 13504 25542 13556 25594
rect 13568 25542 13620 25594
rect 18257 25542 18309 25594
rect 18321 25542 18373 25594
rect 18385 25542 18437 25594
rect 18449 25542 18501 25594
rect 18513 25542 18565 25594
rect 2228 25440 2280 25492
rect 5816 25440 5868 25492
rect 2504 25372 2556 25424
rect 3240 25372 3292 25424
rect 1308 25304 1360 25356
rect 3976 25304 4028 25356
rect 6920 25440 6972 25492
rect 7012 25440 7064 25492
rect 7288 25372 7340 25424
rect 7380 25372 7432 25424
rect 7012 25304 7064 25356
rect 664 25236 716 25288
rect 1768 25279 1820 25288
rect 1768 25245 1777 25279
rect 1777 25245 1811 25279
rect 1811 25245 1820 25279
rect 1768 25236 1820 25245
rect 2136 25236 2188 25288
rect 2412 25236 2464 25288
rect 4712 25279 4764 25288
rect 1308 25168 1360 25220
rect 4712 25245 4721 25279
rect 4721 25245 4755 25279
rect 4755 25245 4764 25279
rect 4712 25236 4764 25245
rect 5632 25279 5684 25288
rect 5632 25245 5641 25279
rect 5641 25245 5675 25279
rect 5675 25245 5684 25279
rect 5632 25236 5684 25245
rect 5724 25236 5776 25288
rect 6736 25236 6788 25288
rect 6828 25279 6880 25288
rect 6828 25245 6837 25279
rect 6837 25245 6871 25279
rect 6871 25245 6880 25279
rect 6828 25236 6880 25245
rect 2596 25100 2648 25152
rect 4252 25211 4304 25220
rect 4252 25177 4261 25211
rect 4261 25177 4295 25211
rect 4295 25177 4304 25211
rect 4252 25168 4304 25177
rect 4620 25168 4672 25220
rect 4804 25168 4856 25220
rect 7840 25372 7892 25424
rect 8208 25440 8260 25492
rect 9036 25440 9088 25492
rect 10048 25304 10100 25356
rect 11428 25304 11480 25356
rect 8576 25236 8628 25288
rect 8208 25168 8260 25220
rect 8760 25211 8812 25220
rect 8760 25177 8769 25211
rect 8769 25177 8803 25211
rect 8803 25177 8812 25211
rect 8760 25168 8812 25177
rect 9220 25249 9272 25288
rect 9220 25236 9245 25249
rect 9245 25236 9272 25249
rect 4068 25100 4120 25152
rect 5080 25143 5132 25152
rect 5080 25109 5089 25143
rect 5089 25109 5123 25143
rect 5123 25109 5132 25143
rect 5080 25100 5132 25109
rect 5264 25143 5316 25152
rect 5264 25109 5273 25143
rect 5273 25109 5307 25143
rect 5307 25109 5316 25143
rect 5264 25100 5316 25109
rect 5448 25100 5500 25152
rect 7472 25143 7524 25152
rect 7472 25109 7481 25143
rect 7481 25109 7515 25143
rect 7515 25109 7524 25143
rect 7472 25100 7524 25109
rect 9036 25100 9088 25152
rect 9220 25100 9272 25152
rect 10784 25236 10836 25288
rect 11244 25168 11296 25220
rect 12164 25483 12216 25492
rect 12164 25449 12173 25483
rect 12173 25449 12207 25483
rect 12207 25449 12216 25483
rect 12164 25440 12216 25449
rect 12532 25440 12584 25492
rect 13360 25440 13412 25492
rect 13912 25440 13964 25492
rect 16396 25440 16448 25492
rect 16948 25440 17000 25492
rect 17224 25440 17276 25492
rect 19064 25440 19116 25492
rect 20260 25483 20312 25492
rect 20260 25449 20269 25483
rect 20269 25449 20303 25483
rect 20303 25449 20312 25483
rect 20260 25440 20312 25449
rect 14096 25372 14148 25424
rect 16212 25372 16264 25424
rect 17040 25372 17092 25424
rect 18972 25372 19024 25424
rect 12072 25279 12124 25288
rect 12072 25245 12081 25279
rect 12081 25245 12115 25279
rect 12115 25245 12124 25279
rect 12072 25236 12124 25245
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 15292 25304 15344 25356
rect 12624 25279 12676 25288
rect 12624 25245 12633 25279
rect 12633 25245 12667 25279
rect 12667 25245 12676 25279
rect 12624 25236 12676 25245
rect 13268 25236 13320 25288
rect 13728 25236 13780 25288
rect 13912 25236 13964 25288
rect 16580 25304 16632 25356
rect 16856 25304 16908 25356
rect 17132 25304 17184 25356
rect 16488 25236 16540 25288
rect 17132 25168 17184 25220
rect 19524 25279 19576 25288
rect 19524 25245 19531 25279
rect 19531 25245 19565 25279
rect 19565 25245 19576 25279
rect 19524 25236 19576 25245
rect 9404 25100 9456 25152
rect 9956 25143 10008 25152
rect 9956 25109 9965 25143
rect 9965 25109 9999 25143
rect 9999 25109 10008 25143
rect 9956 25100 10008 25109
rect 10140 25100 10192 25152
rect 10600 25100 10652 25152
rect 14096 25100 14148 25152
rect 14280 25100 14332 25152
rect 14832 25100 14884 25152
rect 15292 25100 15344 25152
rect 15568 25100 15620 25152
rect 16580 25100 16632 25152
rect 17868 25100 17920 25152
rect 19340 25100 19392 25152
rect 5894 24998 5946 25050
rect 5958 24998 6010 25050
rect 6022 24998 6074 25050
rect 6086 24998 6138 25050
rect 6150 24998 6202 25050
rect 10839 24998 10891 25050
rect 10903 24998 10955 25050
rect 10967 24998 11019 25050
rect 11031 24998 11083 25050
rect 11095 24998 11147 25050
rect 15784 24998 15836 25050
rect 15848 24998 15900 25050
rect 15912 24998 15964 25050
rect 15976 24998 16028 25050
rect 16040 24998 16092 25050
rect 20729 24998 20781 25050
rect 20793 24998 20845 25050
rect 20857 24998 20909 25050
rect 20921 24998 20973 25050
rect 20985 24998 21037 25050
rect 1768 24896 1820 24948
rect 2688 24828 2740 24880
rect 3976 24939 4028 24948
rect 3976 24905 3985 24939
rect 3985 24905 4019 24939
rect 4019 24905 4028 24939
rect 3976 24896 4028 24905
rect 4160 24896 4212 24948
rect 4712 24896 4764 24948
rect 6184 24896 6236 24948
rect 6368 24896 6420 24948
rect 7472 24896 7524 24948
rect 7932 24939 7984 24948
rect 7932 24905 7941 24939
rect 7941 24905 7975 24939
rect 7975 24905 7984 24939
rect 7932 24896 7984 24905
rect 1216 24760 1268 24812
rect 6828 24828 6880 24880
rect 3240 24803 3292 24812
rect 3240 24769 3249 24803
rect 3249 24769 3292 24803
rect 1400 24735 1452 24744
rect 1400 24701 1409 24735
rect 1409 24701 1443 24735
rect 1443 24701 1452 24735
rect 1400 24692 1452 24701
rect 3240 24760 3292 24769
rect 4160 24760 4212 24812
rect 4712 24760 4764 24812
rect 4804 24803 4856 24812
rect 4804 24769 4813 24803
rect 4813 24769 4847 24803
rect 4847 24769 4856 24803
rect 4804 24760 4856 24769
rect 4896 24803 4948 24812
rect 4896 24769 4905 24803
rect 4905 24769 4939 24803
rect 4939 24769 4948 24803
rect 4896 24760 4948 24769
rect 5264 24803 5316 24812
rect 5264 24769 5273 24803
rect 5273 24769 5307 24803
rect 5307 24769 5316 24803
rect 5264 24760 5316 24769
rect 5448 24760 5500 24812
rect 1308 24624 1360 24676
rect 2872 24692 2924 24744
rect 4528 24692 4580 24744
rect 5908 24760 5960 24812
rect 6736 24760 6788 24812
rect 8944 24828 8996 24880
rect 9404 24896 9456 24948
rect 9680 24896 9732 24948
rect 10416 24896 10468 24948
rect 10600 24896 10652 24948
rect 11428 24896 11480 24948
rect 10508 24828 10560 24880
rect 11888 24828 11940 24880
rect 12256 24896 12308 24948
rect 8484 24803 8536 24812
rect 8484 24769 8491 24803
rect 8491 24769 8525 24803
rect 8525 24769 8536 24803
rect 8484 24760 8536 24769
rect 9404 24760 9456 24812
rect 10324 24760 10376 24812
rect 10784 24760 10836 24812
rect 12900 24760 12952 24812
rect 13176 24760 13228 24812
rect 13636 24803 13688 24812
rect 13636 24769 13645 24803
rect 13645 24769 13679 24803
rect 13679 24769 13688 24803
rect 13636 24760 13688 24769
rect 13728 24803 13780 24812
rect 13728 24769 13737 24803
rect 13737 24769 13771 24803
rect 13771 24769 13780 24803
rect 13728 24760 13780 24769
rect 6000 24692 6052 24744
rect 2504 24667 2556 24676
rect 2504 24633 2513 24667
rect 2513 24633 2547 24667
rect 2547 24633 2556 24667
rect 2504 24624 2556 24633
rect 2688 24556 2740 24608
rect 3976 24556 4028 24608
rect 9496 24692 9548 24744
rect 10324 24624 10376 24676
rect 11796 24735 11848 24744
rect 11796 24701 11805 24735
rect 11805 24701 11839 24735
rect 11839 24701 11848 24735
rect 11796 24692 11848 24701
rect 17868 24896 17920 24948
rect 18604 24828 18656 24880
rect 14832 24760 14884 24812
rect 16580 24760 16632 24812
rect 13360 24624 13412 24676
rect 14280 24692 14332 24744
rect 12808 24599 12860 24608
rect 12808 24565 12817 24599
rect 12817 24565 12851 24599
rect 12851 24565 12860 24599
rect 12808 24556 12860 24565
rect 12992 24556 13044 24608
rect 13912 24556 13964 24608
rect 16120 24624 16172 24676
rect 16856 24735 16908 24744
rect 16856 24701 16865 24735
rect 16865 24701 16899 24735
rect 16899 24701 16908 24735
rect 16856 24692 16908 24701
rect 17684 24692 17736 24744
rect 18144 24692 18196 24744
rect 19616 24692 19668 24744
rect 15292 24556 15344 24608
rect 15568 24599 15620 24608
rect 15568 24565 15577 24599
rect 15577 24565 15611 24599
rect 15611 24565 15620 24599
rect 15568 24556 15620 24565
rect 17868 24599 17920 24608
rect 17868 24565 17877 24599
rect 17877 24565 17911 24599
rect 17911 24565 17920 24599
rect 17868 24556 17920 24565
rect 18604 24556 18656 24608
rect 19432 24556 19484 24608
rect 20260 24599 20312 24608
rect 20260 24565 20269 24599
rect 20269 24565 20303 24599
rect 20303 24565 20312 24599
rect 20260 24556 20312 24565
rect 3422 24454 3474 24506
rect 3486 24454 3538 24506
rect 3550 24454 3602 24506
rect 3614 24454 3666 24506
rect 3678 24454 3730 24506
rect 8367 24454 8419 24506
rect 8431 24454 8483 24506
rect 8495 24454 8547 24506
rect 8559 24454 8611 24506
rect 8623 24454 8675 24506
rect 13312 24454 13364 24506
rect 13376 24454 13428 24506
rect 13440 24454 13492 24506
rect 13504 24454 13556 24506
rect 13568 24454 13620 24506
rect 18257 24454 18309 24506
rect 18321 24454 18373 24506
rect 18385 24454 18437 24506
rect 18449 24454 18501 24506
rect 18513 24454 18565 24506
rect 4068 24352 4120 24404
rect 848 24216 900 24268
rect 1492 24259 1544 24268
rect 1492 24225 1501 24259
rect 1501 24225 1535 24259
rect 1535 24225 1544 24259
rect 1492 24216 1544 24225
rect 2964 24216 3016 24268
rect 4620 24352 4672 24404
rect 4896 24352 4948 24404
rect 5724 24352 5776 24404
rect 5816 24352 5868 24404
rect 6000 24352 6052 24404
rect 4712 24284 4764 24336
rect 5264 24259 5316 24268
rect 5264 24225 5273 24259
rect 5273 24225 5307 24259
rect 5307 24225 5316 24259
rect 5264 24216 5316 24225
rect 7104 24395 7156 24404
rect 7104 24361 7113 24395
rect 7113 24361 7147 24395
rect 7147 24361 7156 24395
rect 7104 24352 7156 24361
rect 7196 24352 7248 24404
rect 8760 24352 8812 24404
rect 8944 24352 8996 24404
rect 9496 24352 9548 24404
rect 10784 24395 10836 24404
rect 10784 24361 10793 24395
rect 10793 24361 10827 24395
rect 10827 24361 10836 24395
rect 10784 24352 10836 24361
rect 7012 24284 7064 24336
rect 6828 24216 6880 24268
rect 2228 24148 2280 24200
rect 1308 24080 1360 24132
rect 3700 24148 3752 24200
rect 4620 24148 4672 24200
rect 5080 24148 5132 24200
rect 5448 24191 5500 24200
rect 5448 24157 5457 24191
rect 5457 24157 5491 24191
rect 5491 24157 5500 24191
rect 5448 24148 5500 24157
rect 6184 24191 6236 24200
rect 6184 24157 6193 24191
rect 6193 24157 6227 24191
rect 6227 24157 6236 24191
rect 6184 24148 6236 24157
rect 10508 24216 10560 24268
rect 3240 24080 3292 24132
rect 4160 24080 4212 24132
rect 8208 24148 8260 24200
rect 8300 24148 8352 24200
rect 9772 24191 9824 24200
rect 9772 24157 9781 24191
rect 9781 24157 9815 24191
rect 9815 24157 9824 24191
rect 9772 24148 9824 24157
rect 10324 24148 10376 24200
rect 2412 24012 2464 24064
rect 2964 24012 3016 24064
rect 4068 24012 4120 24064
rect 5080 24012 5132 24064
rect 7840 24080 7892 24132
rect 9956 24080 10008 24132
rect 10140 24080 10192 24132
rect 10508 24080 10560 24132
rect 10784 24216 10836 24268
rect 11428 24259 11480 24268
rect 11428 24225 11437 24259
rect 11437 24225 11471 24259
rect 11471 24225 11480 24259
rect 11428 24216 11480 24225
rect 12072 24259 12124 24268
rect 12072 24225 12081 24259
rect 12081 24225 12115 24259
rect 12115 24225 12124 24259
rect 12072 24216 12124 24225
rect 12808 24216 12860 24268
rect 13544 24352 13596 24404
rect 15568 24352 15620 24404
rect 7564 24012 7616 24064
rect 9496 24055 9548 24064
rect 9496 24021 9505 24055
rect 9505 24021 9539 24055
rect 9539 24021 9548 24055
rect 9496 24012 9548 24021
rect 10876 24012 10928 24064
rect 11428 24012 11480 24064
rect 12348 24191 12400 24200
rect 12348 24157 12357 24191
rect 12357 24157 12391 24191
rect 12391 24157 12400 24191
rect 12348 24148 12400 24157
rect 13636 24148 13688 24200
rect 13728 24148 13780 24200
rect 13912 24148 13964 24200
rect 14096 24216 14148 24268
rect 14556 24191 14608 24200
rect 14556 24157 14565 24191
rect 14565 24157 14599 24191
rect 14599 24157 14608 24191
rect 14556 24148 14608 24157
rect 14740 24148 14792 24200
rect 17684 24352 17736 24404
rect 18236 24352 18288 24404
rect 13912 24012 13964 24064
rect 14096 24012 14148 24064
rect 17868 24191 17920 24200
rect 17868 24157 17877 24191
rect 17877 24157 17911 24191
rect 17911 24157 17920 24191
rect 17868 24148 17920 24157
rect 18972 24284 19024 24336
rect 20352 24148 20404 24200
rect 20628 24148 20680 24200
rect 15660 24012 15712 24064
rect 19616 24080 19668 24132
rect 18604 24012 18656 24064
rect 20260 24055 20312 24064
rect 20260 24021 20269 24055
rect 20269 24021 20303 24055
rect 20303 24021 20312 24055
rect 20260 24012 20312 24021
rect 5894 23910 5946 23962
rect 5958 23910 6010 23962
rect 6022 23910 6074 23962
rect 6086 23910 6138 23962
rect 6150 23910 6202 23962
rect 10839 23910 10891 23962
rect 10903 23910 10955 23962
rect 10967 23910 11019 23962
rect 11031 23910 11083 23962
rect 11095 23910 11147 23962
rect 15784 23910 15836 23962
rect 15848 23910 15900 23962
rect 15912 23910 15964 23962
rect 15976 23910 16028 23962
rect 16040 23910 16092 23962
rect 20729 23910 20781 23962
rect 20793 23910 20845 23962
rect 20857 23910 20909 23962
rect 20921 23910 20973 23962
rect 20985 23910 21037 23962
rect 2964 23808 3016 23860
rect 3240 23851 3292 23860
rect 3240 23817 3249 23851
rect 3249 23817 3283 23851
rect 3283 23817 3292 23851
rect 3240 23808 3292 23817
rect 3700 23808 3752 23860
rect 2136 23783 2188 23792
rect 2136 23749 2145 23783
rect 2145 23749 2179 23783
rect 2179 23749 2188 23783
rect 2136 23740 2188 23749
rect 9496 23851 9548 23860
rect 9496 23817 9505 23851
rect 9505 23817 9539 23851
rect 9539 23817 9548 23851
rect 9496 23808 9548 23817
rect 9772 23783 9824 23792
rect 756 23672 808 23724
rect 1676 23715 1728 23724
rect 1676 23681 1685 23715
rect 1685 23681 1719 23715
rect 1719 23681 1728 23715
rect 1676 23672 1728 23681
rect 2688 23672 2740 23724
rect 2780 23672 2832 23724
rect 5080 23672 5132 23724
rect 5172 23715 5224 23724
rect 5172 23681 5179 23715
rect 5179 23681 5213 23715
rect 5213 23681 5224 23715
rect 5172 23672 5224 23681
rect 2412 23604 2464 23656
rect 3792 23604 3844 23656
rect 1860 23579 1912 23588
rect 1860 23545 1869 23579
rect 1869 23545 1903 23579
rect 1903 23545 1912 23579
rect 1860 23536 1912 23545
rect 3884 23468 3936 23520
rect 5172 23468 5224 23520
rect 6276 23672 6328 23724
rect 7564 23715 7616 23724
rect 7564 23681 7573 23715
rect 7573 23681 7607 23715
rect 7607 23681 7616 23715
rect 7564 23672 7616 23681
rect 9772 23749 9777 23783
rect 9777 23749 9811 23783
rect 9811 23749 9824 23783
rect 9772 23740 9824 23749
rect 9956 23740 10008 23792
rect 11244 23808 11296 23860
rect 11428 23740 11480 23792
rect 12992 23808 13044 23860
rect 13176 23808 13228 23860
rect 14188 23808 14240 23860
rect 14556 23808 14608 23860
rect 15016 23808 15068 23860
rect 16120 23808 16172 23860
rect 17868 23808 17920 23860
rect 19432 23808 19484 23860
rect 13820 23672 13872 23724
rect 14832 23672 14884 23724
rect 17132 23740 17184 23792
rect 19340 23715 19392 23724
rect 19340 23681 19349 23715
rect 19349 23681 19383 23715
rect 19383 23681 19392 23715
rect 19340 23672 19392 23681
rect 20260 23808 20312 23860
rect 6460 23604 6512 23656
rect 6644 23604 6696 23656
rect 7104 23604 7156 23656
rect 7472 23604 7524 23656
rect 10048 23604 10100 23656
rect 11428 23604 11480 23656
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 12532 23647 12584 23656
rect 12532 23613 12566 23647
rect 12566 23613 12584 23647
rect 12532 23604 12584 23613
rect 18696 23604 18748 23656
rect 6828 23536 6880 23588
rect 11244 23536 11296 23588
rect 11888 23536 11940 23588
rect 6368 23468 6420 23520
rect 8208 23511 8260 23520
rect 8208 23477 8217 23511
rect 8217 23477 8251 23511
rect 8251 23477 8260 23511
rect 8208 23468 8260 23477
rect 10784 23511 10836 23520
rect 10784 23477 10793 23511
rect 10793 23477 10827 23511
rect 10827 23477 10836 23511
rect 10784 23468 10836 23477
rect 11152 23468 11204 23520
rect 11796 23468 11848 23520
rect 12072 23468 12124 23520
rect 13176 23536 13228 23588
rect 19340 23536 19392 23588
rect 20076 23536 20128 23588
rect 12440 23468 12492 23520
rect 14280 23468 14332 23520
rect 15200 23511 15252 23520
rect 15200 23477 15209 23511
rect 15209 23477 15243 23511
rect 15243 23477 15252 23511
rect 15200 23468 15252 23477
rect 15660 23468 15712 23520
rect 19064 23511 19116 23520
rect 19064 23477 19073 23511
rect 19073 23477 19107 23511
rect 19107 23477 19116 23511
rect 19064 23468 19116 23477
rect 20444 23511 20496 23520
rect 20444 23477 20453 23511
rect 20453 23477 20487 23511
rect 20487 23477 20496 23511
rect 20444 23468 20496 23477
rect 3422 23366 3474 23418
rect 3486 23366 3538 23418
rect 3550 23366 3602 23418
rect 3614 23366 3666 23418
rect 3678 23366 3730 23418
rect 8367 23366 8419 23418
rect 8431 23366 8483 23418
rect 8495 23366 8547 23418
rect 8559 23366 8611 23418
rect 8623 23366 8675 23418
rect 13312 23366 13364 23418
rect 13376 23366 13428 23418
rect 13440 23366 13492 23418
rect 13504 23366 13556 23418
rect 13568 23366 13620 23418
rect 18257 23366 18309 23418
rect 18321 23366 18373 23418
rect 18385 23366 18437 23418
rect 18449 23366 18501 23418
rect 18513 23366 18565 23418
rect 2320 23264 2372 23316
rect 2688 23264 2740 23316
rect 1952 23196 2004 23248
rect 3700 23128 3752 23180
rect 5356 23264 5408 23316
rect 5264 23196 5316 23248
rect 6000 23196 6052 23248
rect 5356 23128 5408 23180
rect 5632 23128 5684 23180
rect 756 23060 808 23112
rect 940 22992 992 23044
rect 2688 23060 2740 23112
rect 4068 23103 4120 23112
rect 4068 23069 4075 23103
rect 4075 23069 4109 23103
rect 4109 23069 4120 23103
rect 4068 23060 4120 23069
rect 2504 22992 2556 23044
rect 6828 23196 6880 23248
rect 6460 23171 6512 23180
rect 6460 23137 6469 23171
rect 6469 23137 6503 23171
rect 6503 23137 6512 23171
rect 6460 23128 6512 23137
rect 6736 23128 6788 23180
rect 7472 23171 7524 23180
rect 7472 23137 7506 23171
rect 7506 23137 7524 23171
rect 7472 23128 7524 23137
rect 7656 23171 7708 23180
rect 7656 23137 7665 23171
rect 7665 23137 7699 23171
rect 7699 23137 7708 23171
rect 7656 23128 7708 23137
rect 8208 23264 8260 23316
rect 8208 23128 8260 23180
rect 6552 23060 6604 23112
rect 6828 23060 6880 23112
rect 9036 23264 9088 23316
rect 9496 23264 9548 23316
rect 9956 23264 10008 23316
rect 11520 23264 11572 23316
rect 8668 23196 8720 23248
rect 9220 23196 9272 23248
rect 12072 23264 12124 23316
rect 13912 23264 13964 23316
rect 13728 23196 13780 23248
rect 15200 23264 15252 23316
rect 16120 23264 16172 23316
rect 18052 23264 18104 23316
rect 18696 23264 18748 23316
rect 19064 23264 19116 23316
rect 1584 22924 1636 22976
rect 1952 22924 2004 22976
rect 2320 22924 2372 22976
rect 9496 23060 9548 23112
rect 9036 22992 9088 23044
rect 12900 23060 12952 23112
rect 13084 23060 13136 23112
rect 13912 23128 13964 23180
rect 16212 23196 16264 23248
rect 18880 23196 18932 23248
rect 15200 23128 15252 23180
rect 15384 23171 15436 23180
rect 15384 23137 15393 23171
rect 15393 23137 15427 23171
rect 15427 23137 15436 23171
rect 15384 23128 15436 23137
rect 13820 23060 13872 23112
rect 10508 22992 10560 23044
rect 11152 22992 11204 23044
rect 11888 22992 11940 23044
rect 14832 23060 14884 23112
rect 15660 23103 15712 23112
rect 15660 23069 15669 23103
rect 15669 23069 15703 23103
rect 15703 23069 15712 23103
rect 15660 23060 15712 23069
rect 4068 22924 4120 22976
rect 5172 22924 5224 22976
rect 5448 22924 5500 22976
rect 8760 22924 8812 22976
rect 9312 22924 9364 22976
rect 15200 22924 15252 22976
rect 17684 23128 17736 23180
rect 17960 23128 18012 23180
rect 19892 23264 19944 23316
rect 20076 23264 20128 23316
rect 21640 23264 21692 23316
rect 19156 23196 19208 23248
rect 19708 23196 19760 23248
rect 20260 23196 20312 23248
rect 18604 23060 18656 23112
rect 19892 23128 19944 23180
rect 18696 22924 18748 22976
rect 19708 23103 19760 23112
rect 19708 23069 19717 23103
rect 19717 23069 19751 23103
rect 19751 23069 19760 23103
rect 19708 23060 19760 23069
rect 20076 22992 20128 23044
rect 20260 22992 20312 23044
rect 21272 22992 21324 23044
rect 20444 22924 20496 22976
rect 5894 22822 5946 22874
rect 5958 22822 6010 22874
rect 6022 22822 6074 22874
rect 6086 22822 6138 22874
rect 6150 22822 6202 22874
rect 10839 22822 10891 22874
rect 10903 22822 10955 22874
rect 10967 22822 11019 22874
rect 11031 22822 11083 22874
rect 11095 22822 11147 22874
rect 15784 22822 15836 22874
rect 15848 22822 15900 22874
rect 15912 22822 15964 22874
rect 15976 22822 16028 22874
rect 16040 22822 16092 22874
rect 20729 22822 20781 22874
rect 20793 22822 20845 22874
rect 20857 22822 20909 22874
rect 20921 22822 20973 22874
rect 20985 22822 21037 22874
rect 1032 22720 1084 22772
rect 1676 22720 1728 22772
rect 112 22652 164 22704
rect 1308 22652 1360 22704
rect 2320 22695 2372 22704
rect 2320 22661 2329 22695
rect 2329 22661 2363 22695
rect 2363 22661 2372 22695
rect 2320 22652 2372 22661
rect 3148 22695 3200 22704
rect 3148 22661 3157 22695
rect 3157 22661 3191 22695
rect 3191 22661 3200 22695
rect 3148 22652 3200 22661
rect 3332 22763 3384 22772
rect 3332 22729 3341 22763
rect 3341 22729 3375 22763
rect 3375 22729 3384 22763
rect 3332 22720 3384 22729
rect 3976 22720 4028 22772
rect 4344 22720 4396 22772
rect 4620 22720 4672 22772
rect 7564 22720 7616 22772
rect 8852 22720 8904 22772
rect 9036 22720 9088 22772
rect 9220 22720 9272 22772
rect 9404 22720 9456 22772
rect 9588 22720 9640 22772
rect 9772 22720 9824 22772
rect 10232 22720 10284 22772
rect 10508 22720 10560 22772
rect 13820 22720 13872 22772
rect 15568 22720 15620 22772
rect 4436 22695 4488 22704
rect 4436 22661 4445 22695
rect 4445 22661 4479 22695
rect 4479 22661 4488 22695
rect 4436 22652 4488 22661
rect 5172 22652 5224 22704
rect 756 22584 808 22636
rect 2412 22627 2464 22636
rect 2412 22593 2421 22627
rect 2421 22593 2455 22627
rect 2455 22593 2464 22627
rect 2412 22584 2464 22593
rect 2780 22627 2832 22636
rect 2780 22593 2789 22627
rect 2789 22593 2823 22627
rect 2823 22593 2832 22627
rect 2780 22584 2832 22593
rect 3608 22584 3660 22636
rect 3976 22627 4028 22636
rect 3976 22593 3985 22627
rect 3985 22593 4019 22627
rect 4019 22593 4028 22627
rect 3976 22584 4028 22593
rect 4068 22627 4120 22636
rect 4068 22593 4077 22627
rect 4077 22593 4111 22627
rect 4111 22593 4120 22627
rect 4068 22584 4120 22593
rect 4988 22584 5040 22636
rect 5908 22584 5960 22636
rect 6000 22584 6052 22636
rect 6828 22584 6880 22636
rect 9588 22627 9640 22636
rect 9588 22593 9597 22627
rect 9597 22593 9631 22627
rect 9631 22593 9640 22627
rect 9588 22584 9640 22593
rect 10140 22652 10192 22704
rect 2504 22516 2556 22568
rect 3884 22516 3936 22568
rect 4804 22516 4856 22568
rect 7196 22516 7248 22568
rect 7840 22516 7892 22568
rect 9220 22448 9272 22500
rect 9496 22516 9548 22568
rect 10324 22627 10376 22636
rect 10324 22593 10331 22627
rect 10331 22593 10365 22627
rect 10365 22593 10376 22627
rect 10324 22584 10376 22593
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 5080 22380 5132 22432
rect 6920 22380 6972 22432
rect 7196 22380 7248 22432
rect 8024 22380 8076 22432
rect 8852 22380 8904 22432
rect 11336 22584 11388 22636
rect 12256 22584 12308 22636
rect 13084 22584 13136 22636
rect 13912 22584 13964 22636
rect 16764 22652 16816 22704
rect 17224 22652 17276 22704
rect 16488 22584 16540 22636
rect 19708 22720 19760 22772
rect 19892 22720 19944 22772
rect 18512 22584 18564 22636
rect 18696 22695 18748 22704
rect 18696 22661 18730 22695
rect 18730 22661 18748 22695
rect 18696 22652 18748 22661
rect 20444 22652 20496 22704
rect 11152 22516 11204 22568
rect 12256 22448 12308 22500
rect 15108 22491 15160 22500
rect 15108 22457 15117 22491
rect 15117 22457 15151 22491
rect 15151 22457 15160 22491
rect 15108 22448 15160 22457
rect 10508 22380 10560 22432
rect 11060 22423 11112 22432
rect 11060 22389 11069 22423
rect 11069 22389 11103 22423
rect 11103 22389 11112 22423
rect 11060 22380 11112 22389
rect 11428 22380 11480 22432
rect 14188 22380 14240 22432
rect 14648 22380 14700 22432
rect 15568 22516 15620 22568
rect 18144 22448 18196 22500
rect 19064 22380 19116 22432
rect 20444 22423 20496 22432
rect 20444 22389 20453 22423
rect 20453 22389 20487 22423
rect 20487 22389 20496 22423
rect 20444 22380 20496 22389
rect 3422 22278 3474 22330
rect 3486 22278 3538 22330
rect 3550 22278 3602 22330
rect 3614 22278 3666 22330
rect 3678 22278 3730 22330
rect 8367 22278 8419 22330
rect 8431 22278 8483 22330
rect 8495 22278 8547 22330
rect 8559 22278 8611 22330
rect 8623 22278 8675 22330
rect 13312 22278 13364 22330
rect 13376 22278 13428 22330
rect 13440 22278 13492 22330
rect 13504 22278 13556 22330
rect 13568 22278 13620 22330
rect 18257 22278 18309 22330
rect 18321 22278 18373 22330
rect 18385 22278 18437 22330
rect 18449 22278 18501 22330
rect 18513 22278 18565 22330
rect 2780 22176 2832 22228
rect 3976 22176 4028 22228
rect 6368 22176 6420 22228
rect 7840 22176 7892 22228
rect 9588 22176 9640 22228
rect 1952 22040 2004 22092
rect 2780 22040 2832 22092
rect 4160 22108 4212 22160
rect 6000 22151 6052 22160
rect 6000 22117 6009 22151
rect 6009 22117 6043 22151
rect 6043 22117 6052 22151
rect 6000 22108 6052 22117
rect 14740 22176 14792 22228
rect 15108 22176 15160 22228
rect 12256 22108 12308 22160
rect 13268 22108 13320 22160
rect 848 21972 900 22024
rect 1032 21836 1084 21888
rect 5540 22040 5592 22092
rect 5908 22040 5960 22092
rect 9312 22040 9364 22092
rect 3424 22015 3476 22024
rect 3424 21981 3433 22015
rect 3433 21981 3467 22015
rect 3467 21981 3476 22015
rect 3424 21972 3476 21981
rect 3976 21972 4028 22024
rect 4436 21972 4488 22024
rect 4988 22015 5040 22024
rect 4988 21981 4997 22015
rect 4997 21981 5031 22015
rect 5031 21981 5040 22015
rect 4988 21972 5040 21981
rect 6184 21972 6236 22024
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 8760 21972 8812 22024
rect 9220 22015 9272 22024
rect 9220 21981 9229 22015
rect 9229 21981 9263 22015
rect 9263 21981 9272 22015
rect 9220 21972 9272 21981
rect 9772 21972 9824 22024
rect 10508 21972 10560 22024
rect 11152 21972 11204 22024
rect 11428 22015 11480 22024
rect 11428 21981 11451 22015
rect 11451 21981 11480 22015
rect 11428 21972 11480 21981
rect 12072 21972 12124 22024
rect 12256 21972 12308 22024
rect 2412 21836 2464 21888
rect 3608 21879 3660 21888
rect 3608 21845 3617 21879
rect 3617 21845 3651 21879
rect 3651 21845 3660 21879
rect 3608 21836 3660 21845
rect 4712 21879 4764 21888
rect 4712 21845 4721 21879
rect 4721 21845 4755 21879
rect 4755 21845 4764 21879
rect 4712 21836 4764 21845
rect 4988 21836 5040 21888
rect 5632 21836 5684 21888
rect 6184 21836 6236 21888
rect 10140 21904 10192 21956
rect 10232 21904 10284 21956
rect 13912 21972 13964 22024
rect 12532 21904 12584 21956
rect 15016 21972 15068 22024
rect 16948 22176 17000 22228
rect 18604 22176 18656 22228
rect 20260 22219 20312 22228
rect 20260 22185 20269 22219
rect 20269 22185 20303 22219
rect 20303 22185 20312 22219
rect 20260 22176 20312 22185
rect 18420 22108 18472 22160
rect 18696 22108 18748 22160
rect 19156 22108 19208 22160
rect 18328 22040 18380 22092
rect 18972 22040 19024 22092
rect 16396 21904 16448 21956
rect 16764 22015 16816 22024
rect 16764 21981 16773 22015
rect 16773 21981 16807 22015
rect 16807 21981 16816 22015
rect 16764 21972 16816 21981
rect 18144 21972 18196 22024
rect 14832 21836 14884 21888
rect 15292 21836 15344 21888
rect 16304 21836 16356 21888
rect 18420 21972 18472 22024
rect 19064 22015 19116 22024
rect 19064 21981 19073 22015
rect 19073 21981 19107 22015
rect 19107 21981 19116 22015
rect 19064 21972 19116 21981
rect 21548 21972 21600 22024
rect 18972 21904 19024 21956
rect 19708 21904 19760 21956
rect 18328 21879 18380 21888
rect 18328 21845 18337 21879
rect 18337 21845 18371 21879
rect 18371 21845 18380 21879
rect 18328 21836 18380 21845
rect 19248 21836 19300 21888
rect 5894 21734 5946 21786
rect 5958 21734 6010 21786
rect 6022 21734 6074 21786
rect 6086 21734 6138 21786
rect 6150 21734 6202 21786
rect 10839 21734 10891 21786
rect 10903 21734 10955 21786
rect 10967 21734 11019 21786
rect 11031 21734 11083 21786
rect 11095 21734 11147 21786
rect 15784 21734 15836 21786
rect 15848 21734 15900 21786
rect 15912 21734 15964 21786
rect 15976 21734 16028 21786
rect 16040 21734 16092 21786
rect 20729 21734 20781 21786
rect 20793 21734 20845 21786
rect 20857 21734 20909 21786
rect 20921 21734 20973 21786
rect 20985 21734 21037 21786
rect 1584 21632 1636 21684
rect 2044 21632 2096 21684
rect 2504 21675 2556 21684
rect 2504 21641 2513 21675
rect 2513 21641 2547 21675
rect 2547 21641 2556 21675
rect 2504 21632 2556 21641
rect 1952 21564 2004 21616
rect 1676 21496 1728 21548
rect 2412 21496 2464 21548
rect 3884 21564 3936 21616
rect 4896 21632 4948 21684
rect 5540 21632 5592 21684
rect 7656 21632 7708 21684
rect 3240 21496 3292 21548
rect 3792 21496 3844 21548
rect 4160 21496 4212 21548
rect 4436 21496 4488 21548
rect 5080 21564 5132 21616
rect 5448 21496 5500 21548
rect 7748 21564 7800 21616
rect 10416 21632 10468 21684
rect 11428 21632 11480 21684
rect 6736 21496 6788 21548
rect 8208 21564 8260 21616
rect 9036 21564 9088 21616
rect 12992 21632 13044 21684
rect 13820 21632 13872 21684
rect 16764 21632 16816 21684
rect 17224 21632 17276 21684
rect 18328 21632 18380 21684
rect 21272 21632 21324 21684
rect 8852 21496 8904 21548
rect 9496 21496 9548 21548
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 13084 21539 13136 21548
rect 13084 21505 13118 21539
rect 13118 21505 13136 21539
rect 13084 21496 13136 21505
rect 13268 21539 13320 21548
rect 13268 21505 13277 21539
rect 13277 21505 13311 21539
rect 13311 21505 13320 21539
rect 13268 21496 13320 21505
rect 14188 21539 14240 21548
rect 14188 21505 14197 21539
rect 14197 21505 14231 21539
rect 14231 21505 14240 21539
rect 14188 21496 14240 21505
rect 15016 21539 15068 21548
rect 18880 21564 18932 21616
rect 15016 21505 15050 21539
rect 15050 21505 15068 21539
rect 15016 21496 15068 21505
rect 2320 21428 2372 21480
rect 2504 21428 2556 21480
rect 20 21360 72 21412
rect 1216 21360 1268 21412
rect 388 21292 440 21344
rect 1032 21292 1084 21344
rect 1952 21292 2004 21344
rect 3332 21292 3384 21344
rect 4620 21292 4672 21344
rect 8208 21428 8260 21480
rect 9404 21428 9456 21480
rect 9956 21428 10008 21480
rect 10048 21471 10100 21480
rect 10048 21437 10057 21471
rect 10057 21437 10091 21471
rect 10091 21437 10100 21471
rect 10048 21428 10100 21437
rect 9312 21403 9364 21412
rect 9312 21369 9321 21403
rect 9321 21369 9355 21403
rect 9355 21369 9364 21403
rect 9312 21360 9364 21369
rect 7288 21292 7340 21344
rect 7380 21335 7432 21344
rect 7380 21301 7389 21335
rect 7389 21301 7423 21335
rect 7423 21301 7432 21335
rect 7380 21292 7432 21301
rect 9956 21292 10008 21344
rect 11980 21428 12032 21480
rect 12992 21471 13044 21480
rect 12992 21437 13001 21471
rect 13001 21437 13035 21471
rect 13035 21437 13044 21471
rect 12992 21428 13044 21437
rect 12072 21360 12124 21412
rect 12716 21403 12768 21412
rect 12716 21369 12725 21403
rect 12725 21369 12759 21403
rect 12759 21369 12768 21403
rect 12716 21360 12768 21369
rect 11796 21292 11848 21344
rect 12440 21292 12492 21344
rect 15384 21428 15436 21480
rect 13728 21292 13780 21344
rect 14464 21292 14516 21344
rect 14924 21292 14976 21344
rect 15936 21335 15988 21344
rect 15936 21301 15945 21335
rect 15945 21301 15979 21335
rect 15979 21301 15988 21335
rect 15936 21292 15988 21301
rect 19248 21539 19300 21548
rect 19248 21505 19257 21539
rect 19257 21505 19291 21539
rect 19291 21505 19300 21539
rect 19248 21496 19300 21505
rect 20168 21607 20220 21616
rect 20168 21573 20177 21607
rect 20177 21573 20211 21607
rect 20211 21573 20220 21607
rect 20168 21564 20220 21573
rect 20536 21496 20588 21548
rect 19340 21428 19392 21480
rect 20444 21428 20496 21480
rect 18144 21292 18196 21344
rect 19248 21292 19300 21344
rect 19340 21335 19392 21344
rect 19340 21301 19349 21335
rect 19349 21301 19383 21335
rect 19383 21301 19392 21335
rect 19340 21292 19392 21301
rect 19892 21335 19944 21344
rect 19892 21301 19901 21335
rect 19901 21301 19935 21335
rect 19935 21301 19944 21335
rect 19892 21292 19944 21301
rect 3422 21190 3474 21242
rect 3486 21190 3538 21242
rect 3550 21190 3602 21242
rect 3614 21190 3666 21242
rect 3678 21190 3730 21242
rect 8367 21190 8419 21242
rect 8431 21190 8483 21242
rect 8495 21190 8547 21242
rect 8559 21190 8611 21242
rect 8623 21190 8675 21242
rect 13312 21190 13364 21242
rect 13376 21190 13428 21242
rect 13440 21190 13492 21242
rect 13504 21190 13556 21242
rect 13568 21190 13620 21242
rect 18257 21190 18309 21242
rect 18321 21190 18373 21242
rect 18385 21190 18437 21242
rect 18449 21190 18501 21242
rect 18513 21190 18565 21242
rect 3700 21020 3752 21072
rect 7380 21088 7432 21140
rect 8208 21088 8260 21140
rect 9036 21088 9088 21140
rect 11336 21088 11388 21140
rect 12440 21088 12492 21140
rect 12992 21088 13044 21140
rect 15936 21088 15988 21140
rect 17040 21088 17092 21140
rect 3424 20884 3476 20936
rect 3608 20884 3660 20936
rect 296 20816 348 20868
rect 1124 20816 1176 20868
rect 2228 20859 2280 20868
rect 2228 20825 2237 20859
rect 2237 20825 2271 20859
rect 2271 20825 2280 20859
rect 2228 20816 2280 20825
rect 2504 20816 2556 20868
rect 3056 20816 3108 20868
rect 4896 20884 4948 20936
rect 5172 20884 5224 20936
rect 5816 20884 5868 20936
rect 5908 20884 5960 20936
rect 10508 21020 10560 21072
rect 10600 20952 10652 21004
rect 11428 20952 11480 21004
rect 11520 20995 11572 21004
rect 11520 20961 11529 20995
rect 11529 20961 11563 20995
rect 11563 20961 11572 20995
rect 11520 20952 11572 20961
rect 13544 21020 13596 21072
rect 14648 21020 14700 21072
rect 2872 20748 2924 20800
rect 4252 20816 4304 20868
rect 4988 20816 5040 20868
rect 4068 20748 4120 20800
rect 6368 20816 6420 20868
rect 7288 20816 7340 20868
rect 8668 20884 8720 20936
rect 8760 20816 8812 20868
rect 9036 20816 9088 20868
rect 11060 20927 11112 20936
rect 11060 20893 11069 20927
rect 11069 20893 11103 20927
rect 11103 20893 11112 20927
rect 11060 20884 11112 20893
rect 11796 20927 11848 20936
rect 11796 20893 11823 20927
rect 11823 20893 11848 20927
rect 11796 20884 11848 20893
rect 12072 20927 12124 20936
rect 12072 20893 12081 20927
rect 12081 20893 12115 20927
rect 12115 20893 12124 20927
rect 12072 20884 12124 20893
rect 13544 20884 13596 20936
rect 8024 20748 8076 20800
rect 8208 20748 8260 20800
rect 10968 20748 11020 20800
rect 12164 20748 12216 20800
rect 12624 20748 12676 20800
rect 13084 20748 13136 20800
rect 13820 20748 13872 20800
rect 14096 20927 14148 20936
rect 14096 20893 14105 20927
rect 14105 20893 14139 20927
rect 14139 20893 14148 20927
rect 14096 20884 14148 20893
rect 14188 20816 14240 20868
rect 18420 21088 18472 21140
rect 19708 21088 19760 21140
rect 19892 21020 19944 21072
rect 14464 20884 14516 20936
rect 15016 20927 15068 20936
rect 15016 20893 15025 20927
rect 15025 20893 15059 20927
rect 15059 20893 15068 20927
rect 15016 20884 15068 20893
rect 15292 20927 15344 20936
rect 15292 20893 15301 20927
rect 15301 20893 15335 20927
rect 15335 20893 15344 20927
rect 15292 20884 15344 20893
rect 15016 20748 15068 20800
rect 16120 20748 16172 20800
rect 16396 20927 16448 20936
rect 16396 20893 16405 20927
rect 16405 20893 16439 20927
rect 16439 20893 16448 20927
rect 16396 20884 16448 20893
rect 19340 20952 19392 21004
rect 20352 20952 20404 21004
rect 21732 20952 21784 21004
rect 18880 20927 18932 20936
rect 18880 20893 18889 20927
rect 18889 20893 18923 20927
rect 18923 20893 18932 20927
rect 18880 20884 18932 20893
rect 18972 20884 19024 20936
rect 19432 20927 19484 20936
rect 19432 20893 19441 20927
rect 19441 20893 19475 20927
rect 19475 20893 19484 20927
rect 19432 20884 19484 20893
rect 19984 20927 20036 20936
rect 19984 20893 19993 20927
rect 19993 20893 20027 20927
rect 20027 20893 20036 20927
rect 19984 20884 20036 20893
rect 16488 20859 16540 20868
rect 16488 20825 16497 20859
rect 16497 20825 16531 20859
rect 16531 20825 16540 20859
rect 16488 20816 16540 20825
rect 16580 20859 16632 20868
rect 16580 20825 16589 20859
rect 16589 20825 16623 20859
rect 16623 20825 16632 20859
rect 16580 20816 16632 20825
rect 19340 20816 19392 20868
rect 21272 20816 21324 20868
rect 17132 20748 17184 20800
rect 17500 20748 17552 20800
rect 19708 20748 19760 20800
rect 21548 20748 21600 20800
rect 5894 20646 5946 20698
rect 5958 20646 6010 20698
rect 6022 20646 6074 20698
rect 6086 20646 6138 20698
rect 6150 20646 6202 20698
rect 10839 20646 10891 20698
rect 10903 20646 10955 20698
rect 10967 20646 11019 20698
rect 11031 20646 11083 20698
rect 11095 20646 11147 20698
rect 15784 20646 15836 20698
rect 15848 20646 15900 20698
rect 15912 20646 15964 20698
rect 15976 20646 16028 20698
rect 16040 20646 16092 20698
rect 20729 20646 20781 20698
rect 20793 20646 20845 20698
rect 20857 20646 20909 20698
rect 20921 20646 20973 20698
rect 20985 20646 21037 20698
rect 1584 20544 1636 20596
rect 1860 20544 1912 20596
rect 2228 20544 2280 20596
rect 3608 20544 3660 20596
rect 1860 20451 1912 20460
rect 1860 20417 1867 20451
rect 1867 20417 1901 20451
rect 1901 20417 1912 20451
rect 1860 20408 1912 20417
rect 3884 20476 3936 20528
rect 4620 20476 4672 20528
rect 6736 20544 6788 20596
rect 8300 20544 8352 20596
rect 11612 20544 11664 20596
rect 3516 20408 3568 20460
rect 4712 20408 4764 20460
rect 8944 20476 8996 20528
rect 10876 20476 10928 20528
rect 11796 20476 11848 20528
rect 12716 20587 12768 20596
rect 12716 20553 12725 20587
rect 12725 20553 12759 20587
rect 12759 20553 12768 20587
rect 12716 20544 12768 20553
rect 13084 20544 13136 20596
rect 14464 20544 14516 20596
rect 15292 20544 15344 20596
rect 16120 20544 16172 20596
rect 16396 20544 16448 20596
rect 16580 20544 16632 20596
rect 16856 20544 16908 20596
rect 17776 20544 17828 20596
rect 18788 20544 18840 20596
rect 7380 20451 7432 20460
rect 7380 20417 7387 20451
rect 7387 20417 7421 20451
rect 7421 20417 7432 20451
rect 7380 20408 7432 20417
rect 7472 20408 7524 20460
rect 7840 20408 7892 20460
rect 8760 20408 8812 20460
rect 10784 20408 10836 20460
rect 12072 20408 12124 20460
rect 16028 20476 16080 20528
rect 2320 20204 2372 20256
rect 6736 20340 6788 20392
rect 4436 20272 4488 20324
rect 5816 20272 5868 20324
rect 4068 20204 4120 20256
rect 8208 20340 8260 20392
rect 10600 20340 10652 20392
rect 8208 20204 8260 20256
rect 8668 20204 8720 20256
rect 8852 20247 8904 20256
rect 8852 20213 8861 20247
rect 8861 20213 8895 20247
rect 8895 20213 8904 20247
rect 8852 20204 8904 20213
rect 9956 20247 10008 20256
rect 9956 20213 9965 20247
rect 9965 20213 9999 20247
rect 9999 20213 10008 20247
rect 9956 20204 10008 20213
rect 13176 20340 13228 20392
rect 12164 20204 12216 20256
rect 12532 20204 12584 20256
rect 13084 20204 13136 20256
rect 14096 20408 14148 20460
rect 14464 20408 14516 20460
rect 14924 20451 14976 20460
rect 14924 20417 14931 20451
rect 14931 20417 14965 20451
rect 14965 20417 14976 20451
rect 14924 20408 14976 20417
rect 17500 20408 17552 20460
rect 18420 20408 18472 20460
rect 19340 20408 19392 20460
rect 20076 20451 20128 20460
rect 14096 20272 14148 20324
rect 16672 20383 16724 20392
rect 16672 20349 16681 20383
rect 16681 20349 16715 20383
rect 16715 20349 16724 20383
rect 16672 20340 16724 20349
rect 16580 20204 16632 20256
rect 17960 20204 18012 20256
rect 18880 20204 18932 20256
rect 20076 20417 20085 20451
rect 20085 20417 20119 20451
rect 20119 20417 20128 20451
rect 20076 20408 20128 20417
rect 19708 20340 19760 20392
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 19984 20204 20036 20213
rect 20260 20247 20312 20256
rect 20260 20213 20269 20247
rect 20269 20213 20303 20247
rect 20303 20213 20312 20247
rect 20260 20204 20312 20213
rect 204 20068 256 20120
rect 3422 20102 3474 20154
rect 3486 20102 3538 20154
rect 3550 20102 3602 20154
rect 3614 20102 3666 20154
rect 3678 20102 3730 20154
rect 8367 20102 8419 20154
rect 8431 20102 8483 20154
rect 8495 20102 8547 20154
rect 8559 20102 8611 20154
rect 8623 20102 8675 20154
rect 13312 20102 13364 20154
rect 13376 20102 13428 20154
rect 13440 20102 13492 20154
rect 13504 20102 13556 20154
rect 13568 20102 13620 20154
rect 18257 20102 18309 20154
rect 18321 20102 18373 20154
rect 18385 20102 18437 20154
rect 18449 20102 18501 20154
rect 18513 20102 18565 20154
rect 3700 20000 3752 20052
rect 1400 19907 1452 19916
rect 1400 19873 1409 19907
rect 1409 19873 1443 19907
rect 1443 19873 1452 19907
rect 1400 19864 1452 19873
rect 1676 19907 1728 19916
rect 1676 19873 1685 19907
rect 1685 19873 1719 19907
rect 1719 19873 1728 19907
rect 1676 19864 1728 19873
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 4068 19864 4120 19916
rect 5172 19864 5224 19916
rect 7472 20000 7524 20052
rect 6736 19932 6788 19984
rect 2688 19796 2740 19848
rect 3240 19728 3292 19780
rect 3332 19703 3384 19712
rect 3332 19669 3341 19703
rect 3341 19669 3375 19703
rect 3375 19669 3384 19703
rect 3332 19660 3384 19669
rect 3700 19660 3752 19712
rect 3884 19660 3936 19712
rect 4252 19728 4304 19780
rect 5724 19796 5776 19848
rect 6368 19796 6420 19848
rect 8576 19932 8628 19984
rect 8852 19932 8904 19984
rect 8668 19864 8720 19916
rect 11520 20000 11572 20052
rect 12256 20000 12308 20052
rect 13176 20000 13228 20052
rect 14096 20000 14148 20052
rect 11520 19864 11572 19916
rect 15384 19864 15436 19916
rect 16396 20000 16448 20052
rect 16856 20000 16908 20052
rect 17776 20000 17828 20052
rect 18972 20000 19024 20052
rect 16396 19864 16448 19916
rect 16764 19864 16816 19916
rect 8208 19796 8260 19848
rect 4620 19660 4672 19712
rect 4896 19660 4948 19712
rect 5632 19660 5684 19712
rect 8852 19660 8904 19712
rect 9128 19839 9180 19848
rect 9128 19805 9137 19839
rect 9137 19805 9171 19839
rect 9171 19805 9180 19839
rect 9128 19796 9180 19805
rect 9496 19839 9548 19848
rect 9496 19805 9503 19839
rect 9503 19805 9537 19839
rect 9537 19805 9548 19839
rect 9496 19796 9548 19805
rect 10048 19796 10100 19848
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 10784 19796 10836 19848
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 14096 19839 14148 19848
rect 14096 19805 14105 19839
rect 14105 19805 14139 19839
rect 14139 19805 14148 19839
rect 14096 19796 14148 19805
rect 14372 19839 14424 19848
rect 14372 19805 14379 19839
rect 14379 19805 14413 19839
rect 14413 19805 14424 19839
rect 14372 19796 14424 19805
rect 18144 19864 18196 19916
rect 10048 19660 10100 19712
rect 10232 19703 10284 19712
rect 10232 19669 10241 19703
rect 10241 19669 10275 19703
rect 10275 19669 10284 19703
rect 10232 19660 10284 19669
rect 10600 19660 10652 19712
rect 11980 19660 12032 19712
rect 12164 19660 12216 19712
rect 12992 19703 13044 19712
rect 12992 19669 13001 19703
rect 13001 19669 13035 19703
rect 13035 19669 13044 19703
rect 12992 19660 13044 19669
rect 14832 19728 14884 19780
rect 19984 20000 20036 20052
rect 20076 20000 20128 20052
rect 14372 19660 14424 19712
rect 14648 19660 14700 19712
rect 15660 19660 15712 19712
rect 16212 19660 16264 19712
rect 19340 19728 19392 19780
rect 17592 19703 17644 19712
rect 17592 19669 17601 19703
rect 17601 19669 17635 19703
rect 17635 19669 17644 19703
rect 17592 19660 17644 19669
rect 18420 19660 18472 19712
rect 19064 19660 19116 19712
rect 19524 19660 19576 19712
rect 20996 19660 21048 19712
rect 5894 19558 5946 19610
rect 5958 19558 6010 19610
rect 6022 19558 6074 19610
rect 6086 19558 6138 19610
rect 6150 19558 6202 19610
rect 10839 19558 10891 19610
rect 10903 19558 10955 19610
rect 10967 19558 11019 19610
rect 11031 19558 11083 19610
rect 11095 19558 11147 19610
rect 15784 19558 15836 19610
rect 15848 19558 15900 19610
rect 15912 19558 15964 19610
rect 15976 19558 16028 19610
rect 16040 19558 16092 19610
rect 20729 19558 20781 19610
rect 20793 19558 20845 19610
rect 20857 19558 20909 19610
rect 20921 19558 20973 19610
rect 20985 19558 21037 19610
rect 3240 19456 3292 19508
rect 3332 19456 3384 19508
rect 756 19388 808 19440
rect 2136 19388 2188 19440
rect 4344 19456 4396 19508
rect 7288 19456 7340 19508
rect 3700 19388 3752 19440
rect 4620 19431 4672 19440
rect 4620 19397 4629 19431
rect 4629 19397 4663 19431
rect 4663 19397 4672 19431
rect 4620 19388 4672 19397
rect 5264 19388 5316 19440
rect 8944 19456 8996 19508
rect 9128 19456 9180 19508
rect 4252 19363 4304 19372
rect 4252 19329 4261 19363
rect 4261 19329 4295 19363
rect 4295 19329 4304 19363
rect 4252 19320 4304 19329
rect 4712 19320 4764 19372
rect 5632 19320 5684 19372
rect 7656 19363 7708 19372
rect 7656 19329 7665 19363
rect 7665 19329 7699 19363
rect 7699 19329 7708 19363
rect 7656 19320 7708 19329
rect 9680 19388 9732 19440
rect 10232 19456 10284 19508
rect 11888 19456 11940 19508
rect 13544 19456 13596 19508
rect 14372 19456 14424 19508
rect 15108 19456 15160 19508
rect 15660 19456 15712 19508
rect 17868 19456 17920 19508
rect 13084 19388 13136 19440
rect 13360 19388 13412 19440
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 8668 19363 8720 19372
rect 8668 19329 8702 19363
rect 8702 19329 8720 19363
rect 8668 19320 8720 19329
rect 8852 19363 8904 19372
rect 8852 19329 8861 19363
rect 8861 19329 8895 19363
rect 8895 19329 8904 19363
rect 8852 19320 8904 19329
rect 10508 19363 10560 19372
rect 10508 19329 10517 19363
rect 10517 19329 10551 19363
rect 10551 19329 10560 19363
rect 10508 19320 10560 19329
rect 11152 19320 11204 19372
rect 12532 19363 12584 19372
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 14004 19320 14056 19372
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 17224 19363 17276 19372
rect 17224 19329 17231 19363
rect 17231 19329 17265 19363
rect 17265 19329 17276 19363
rect 17224 19320 17276 19329
rect 17592 19320 17644 19372
rect 18420 19456 18472 19508
rect 20260 19456 20312 19508
rect 19984 19388 20036 19440
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 20260 19363 20312 19372
rect 20260 19329 20269 19363
rect 20269 19329 20303 19363
rect 20303 19329 20312 19363
rect 20260 19320 20312 19329
rect 1308 19116 1360 19168
rect 8300 19295 8352 19304
rect 8300 19261 8309 19295
rect 8309 19261 8343 19295
rect 8343 19261 8352 19295
rect 8300 19252 8352 19261
rect 9956 19252 10008 19304
rect 12992 19252 13044 19304
rect 14648 19252 14700 19304
rect 15016 19252 15068 19304
rect 15108 19295 15160 19304
rect 15108 19261 15117 19295
rect 15117 19261 15151 19295
rect 15151 19261 15160 19295
rect 15108 19252 15160 19261
rect 4804 19227 4856 19236
rect 4804 19193 4813 19227
rect 4813 19193 4847 19227
rect 4847 19193 4856 19227
rect 4804 19184 4856 19193
rect 4896 19184 4948 19236
rect 2044 19116 2096 19168
rect 2320 19116 2372 19168
rect 2780 19116 2832 19168
rect 3424 19116 3476 19168
rect 5264 19116 5316 19168
rect 6828 19184 6880 19236
rect 8116 19184 8168 19236
rect 11060 19227 11112 19236
rect 11060 19193 11069 19227
rect 11069 19193 11103 19227
rect 11103 19193 11112 19227
rect 11060 19184 11112 19193
rect 16120 19184 16172 19236
rect 7564 19116 7616 19168
rect 7932 19116 7984 19168
rect 9404 19116 9456 19168
rect 9496 19159 9548 19168
rect 9496 19125 9505 19159
rect 9505 19125 9539 19159
rect 9539 19125 9548 19159
rect 9496 19116 9548 19125
rect 15016 19116 15068 19168
rect 15476 19116 15528 19168
rect 15844 19116 15896 19168
rect 19340 19252 19392 19304
rect 20352 19252 20404 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 18144 19184 18196 19236
rect 19156 19116 19208 19168
rect 19248 19116 19300 19168
rect 20076 19159 20128 19168
rect 20076 19125 20085 19159
rect 20085 19125 20119 19159
rect 20119 19125 20128 19159
rect 20076 19116 20128 19125
rect 20352 19159 20404 19168
rect 20352 19125 20361 19159
rect 20361 19125 20395 19159
rect 20395 19125 20404 19159
rect 20352 19116 20404 19125
rect 3422 19014 3474 19066
rect 3486 19014 3538 19066
rect 3550 19014 3602 19066
rect 3614 19014 3666 19066
rect 3678 19014 3730 19066
rect 8367 19014 8419 19066
rect 8431 19014 8483 19066
rect 8495 19014 8547 19066
rect 8559 19014 8611 19066
rect 8623 19014 8675 19066
rect 13312 19014 13364 19066
rect 13376 19014 13428 19066
rect 13440 19014 13492 19066
rect 13504 19014 13556 19066
rect 13568 19014 13620 19066
rect 18257 19014 18309 19066
rect 18321 19014 18373 19066
rect 18385 19014 18437 19066
rect 18449 19014 18501 19066
rect 18513 19014 18565 19066
rect 3056 18912 3108 18964
rect 4344 18912 4396 18964
rect 5172 18912 5224 18964
rect 6552 18912 6604 18964
rect 6736 18912 6788 18964
rect 7564 18912 7616 18964
rect 8300 18912 8352 18964
rect 12532 18912 12584 18964
rect 1584 18844 1636 18896
rect 1768 18844 1820 18896
rect 1216 18776 1268 18828
rect 756 18708 808 18760
rect 1216 18640 1268 18692
rect 2688 18751 2740 18760
rect 2688 18717 2697 18751
rect 2697 18717 2731 18751
rect 2731 18717 2740 18751
rect 2688 18708 2740 18717
rect 3700 18776 3752 18828
rect 4896 18776 4948 18828
rect 9680 18776 9732 18828
rect 11520 18776 11572 18828
rect 3056 18708 3108 18760
rect 3332 18708 3384 18760
rect 4436 18708 4488 18760
rect 6460 18708 6512 18760
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 7288 18708 7340 18760
rect 7380 18708 7432 18760
rect 1860 18683 1912 18692
rect 1860 18649 1869 18683
rect 1869 18649 1903 18683
rect 1903 18649 1912 18683
rect 1860 18640 1912 18649
rect 2044 18683 2096 18692
rect 2044 18649 2053 18683
rect 2053 18649 2087 18683
rect 2087 18649 2096 18683
rect 2044 18640 2096 18649
rect 5172 18640 5224 18692
rect 12072 18708 12124 18760
rect 12532 18751 12584 18760
rect 12532 18717 12539 18751
rect 12539 18717 12573 18751
rect 12573 18717 12584 18751
rect 12532 18708 12584 18717
rect 9772 18640 9824 18692
rect 10048 18683 10100 18692
rect 10048 18649 10057 18683
rect 10057 18649 10091 18683
rect 10091 18649 10100 18683
rect 10048 18640 10100 18649
rect 10232 18640 10284 18692
rect 10416 18683 10468 18692
rect 10416 18649 10425 18683
rect 10425 18649 10459 18683
rect 10459 18649 10468 18683
rect 10416 18640 10468 18649
rect 10508 18640 10560 18692
rect 11060 18640 11112 18692
rect 14280 18776 14332 18828
rect 14924 18819 14976 18828
rect 14924 18785 14933 18819
rect 14933 18785 14967 18819
rect 14967 18785 14976 18819
rect 14924 18776 14976 18785
rect 15568 18819 15620 18828
rect 15568 18785 15577 18819
rect 15577 18785 15611 18819
rect 15611 18785 15620 18819
rect 15568 18776 15620 18785
rect 20352 18912 20404 18964
rect 21548 18844 21600 18896
rect 21272 18776 21324 18828
rect 13820 18708 13872 18760
rect 15844 18751 15896 18760
rect 15844 18717 15853 18751
rect 15853 18717 15887 18751
rect 15887 18717 15896 18751
rect 15844 18708 15896 18717
rect 14924 18640 14976 18692
rect 2780 18572 2832 18624
rect 3148 18572 3200 18624
rect 5448 18572 5500 18624
rect 7656 18572 7708 18624
rect 8208 18572 8260 18624
rect 9220 18572 9272 18624
rect 11152 18615 11204 18624
rect 11152 18581 11161 18615
rect 11161 18581 11195 18615
rect 11195 18581 11204 18615
rect 11152 18572 11204 18581
rect 11336 18615 11388 18624
rect 11336 18581 11345 18615
rect 11345 18581 11379 18615
rect 11379 18581 11388 18615
rect 11336 18572 11388 18581
rect 12072 18572 12124 18624
rect 12900 18572 12952 18624
rect 14096 18572 14148 18624
rect 16948 18640 17000 18692
rect 20168 18751 20220 18760
rect 20168 18717 20177 18751
rect 20177 18717 20211 18751
rect 20211 18717 20220 18751
rect 20168 18708 20220 18717
rect 16764 18615 16816 18624
rect 16764 18581 16773 18615
rect 16773 18581 16807 18615
rect 16807 18581 16816 18615
rect 16764 18572 16816 18581
rect 18696 18572 18748 18624
rect 21640 18640 21692 18692
rect 5894 18470 5946 18522
rect 5958 18470 6010 18522
rect 6022 18470 6074 18522
rect 6086 18470 6138 18522
rect 6150 18470 6202 18522
rect 10839 18470 10891 18522
rect 10903 18470 10955 18522
rect 10967 18470 11019 18522
rect 11031 18470 11083 18522
rect 11095 18470 11147 18522
rect 15784 18470 15836 18522
rect 15848 18470 15900 18522
rect 15912 18470 15964 18522
rect 15976 18470 16028 18522
rect 16040 18470 16092 18522
rect 20729 18470 20781 18522
rect 20793 18470 20845 18522
rect 20857 18470 20909 18522
rect 20921 18470 20973 18522
rect 20985 18470 21037 18522
rect 1308 18368 1360 18420
rect 3148 18368 3200 18420
rect 4344 18368 4396 18420
rect 5080 18368 5132 18420
rect 7840 18368 7892 18420
rect 9496 18368 9548 18420
rect 756 18300 808 18352
rect 1952 18300 2004 18352
rect 3056 18300 3108 18352
rect 3240 18300 3292 18352
rect 3976 18300 4028 18352
rect 4620 18343 4672 18352
rect 4620 18309 4629 18343
rect 4629 18309 4663 18343
rect 4663 18309 4672 18343
rect 9680 18411 9732 18420
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 10416 18368 10468 18420
rect 4620 18300 4672 18309
rect 3608 18232 3660 18284
rect 3792 18275 3844 18284
rect 3792 18241 3801 18275
rect 3801 18241 3835 18275
rect 3835 18241 3844 18275
rect 3792 18232 3844 18241
rect 3884 18275 3936 18284
rect 3884 18241 3893 18275
rect 3893 18241 3927 18275
rect 3927 18241 3936 18275
rect 3884 18232 3936 18241
rect 4252 18275 4304 18284
rect 4252 18241 4261 18275
rect 4261 18241 4295 18275
rect 4295 18241 4304 18275
rect 4252 18232 4304 18241
rect 4896 18232 4948 18284
rect 5080 18232 5132 18284
rect 7472 18232 7524 18284
rect 8300 18232 8352 18284
rect 1952 18028 2004 18080
rect 2320 18028 2372 18080
rect 2688 18028 2740 18080
rect 11796 18300 11848 18352
rect 12072 18300 12124 18352
rect 12440 18300 12492 18352
rect 12900 18300 12952 18352
rect 13820 18300 13872 18352
rect 14280 18300 14332 18352
rect 15108 18368 15160 18420
rect 15384 18368 15436 18420
rect 16856 18368 16908 18420
rect 19616 18368 19668 18420
rect 18696 18343 18748 18352
rect 18696 18309 18708 18343
rect 18708 18309 18748 18343
rect 18696 18300 18748 18309
rect 19156 18300 19208 18352
rect 9588 18232 9640 18284
rect 9956 18164 10008 18216
rect 9496 18096 9548 18148
rect 7656 18028 7708 18080
rect 9956 18028 10008 18080
rect 10508 18028 10560 18080
rect 10784 18028 10836 18080
rect 15384 18232 15436 18284
rect 16212 18232 16264 18284
rect 17960 18232 18012 18284
rect 11520 18164 11572 18216
rect 12440 18164 12492 18216
rect 12900 18164 12952 18216
rect 13544 18164 13596 18216
rect 14096 18164 14148 18216
rect 15108 18164 15160 18216
rect 17316 18164 17368 18216
rect 12624 18028 12676 18080
rect 16396 18028 16448 18080
rect 20996 18028 21048 18080
rect 3422 17926 3474 17978
rect 3486 17926 3538 17978
rect 3550 17926 3602 17978
rect 3614 17926 3666 17978
rect 3678 17926 3730 17978
rect 8367 17926 8419 17978
rect 8431 17926 8483 17978
rect 8495 17926 8547 17978
rect 8559 17926 8611 17978
rect 8623 17926 8675 17978
rect 13312 17926 13364 17978
rect 13376 17926 13428 17978
rect 13440 17926 13492 17978
rect 13504 17926 13556 17978
rect 13568 17926 13620 17978
rect 18257 17926 18309 17978
rect 18321 17926 18373 17978
rect 18385 17926 18437 17978
rect 18449 17926 18501 17978
rect 18513 17926 18565 17978
rect 1676 17824 1728 17876
rect 1308 17756 1360 17808
rect 2228 17824 2280 17876
rect 2688 17867 2740 17876
rect 2688 17833 2697 17867
rect 2697 17833 2731 17867
rect 2731 17833 2740 17867
rect 2688 17824 2740 17833
rect 1860 17756 1912 17808
rect 848 17688 900 17740
rect 1584 17688 1636 17740
rect 2228 17688 2280 17740
rect 2412 17688 2464 17740
rect 7104 17824 7156 17876
rect 7472 17824 7524 17876
rect 6828 17731 6880 17740
rect 6828 17697 6837 17731
rect 6837 17697 6871 17731
rect 6871 17697 6880 17731
rect 6828 17688 6880 17697
rect 6920 17688 6972 17740
rect 8852 17688 8904 17740
rect 11520 17688 11572 17740
rect 13728 17824 13780 17876
rect 14556 17756 14608 17808
rect 15568 17824 15620 17876
rect 16580 17824 16632 17876
rect 19248 17824 19300 17876
rect 20260 17867 20312 17876
rect 20260 17833 20269 17867
rect 20269 17833 20303 17867
rect 20303 17833 20312 17867
rect 20260 17824 20312 17833
rect 14096 17688 14148 17740
rect 1492 17663 1544 17672
rect 1492 17629 1501 17663
rect 1501 17629 1535 17663
rect 1535 17629 1544 17663
rect 1492 17620 1544 17629
rect 1492 17484 1544 17536
rect 2136 17527 2188 17536
rect 2136 17493 2145 17527
rect 2145 17493 2179 17527
rect 2179 17493 2188 17527
rect 2136 17484 2188 17493
rect 3148 17620 3200 17672
rect 3332 17620 3384 17672
rect 3516 17663 3568 17672
rect 3516 17629 3525 17663
rect 3525 17629 3559 17663
rect 3559 17629 3568 17663
rect 3516 17620 3568 17629
rect 4436 17620 4488 17672
rect 4896 17620 4948 17672
rect 6552 17620 6604 17672
rect 7104 17663 7156 17672
rect 7104 17629 7113 17663
rect 7113 17629 7147 17663
rect 7147 17629 7156 17663
rect 7104 17620 7156 17629
rect 7390 17663 7442 17672
rect 7390 17629 7399 17663
rect 7399 17629 7433 17663
rect 7433 17629 7442 17663
rect 7390 17620 7442 17629
rect 9680 17620 9732 17672
rect 10232 17620 10284 17672
rect 12072 17620 12124 17672
rect 3608 17552 3660 17604
rect 5080 17595 5132 17604
rect 5080 17561 5089 17595
rect 5089 17561 5123 17595
rect 5123 17561 5132 17595
rect 5080 17552 5132 17561
rect 5724 17552 5776 17604
rect 9404 17552 9456 17604
rect 10048 17552 10100 17604
rect 10508 17595 10560 17604
rect 10508 17561 10517 17595
rect 10517 17561 10551 17595
rect 10551 17561 10560 17595
rect 10508 17552 10560 17561
rect 10784 17552 10836 17604
rect 10968 17552 11020 17604
rect 11704 17552 11756 17604
rect 13176 17620 13228 17672
rect 13728 17620 13780 17672
rect 13820 17620 13872 17672
rect 14372 17620 14424 17672
rect 16396 17663 16448 17672
rect 3976 17527 4028 17536
rect 3976 17493 3985 17527
rect 3985 17493 4019 17527
rect 4019 17493 4028 17527
rect 3976 17484 4028 17493
rect 5172 17484 5224 17536
rect 5356 17484 5408 17536
rect 5448 17484 5500 17536
rect 5908 17484 5960 17536
rect 7196 17484 7248 17536
rect 8024 17527 8076 17536
rect 8024 17493 8033 17527
rect 8033 17493 8067 17527
rect 8067 17493 8076 17527
rect 8024 17484 8076 17493
rect 10600 17484 10652 17536
rect 11244 17527 11296 17536
rect 11244 17493 11253 17527
rect 11253 17493 11287 17527
rect 11287 17493 11296 17527
rect 11244 17484 11296 17493
rect 12256 17484 12308 17536
rect 14464 17552 14516 17604
rect 14832 17552 14884 17604
rect 16396 17629 16403 17663
rect 16403 17629 16437 17663
rect 16437 17629 16448 17663
rect 16396 17620 16448 17629
rect 16672 17552 16724 17604
rect 18052 17552 18104 17604
rect 13084 17484 13136 17536
rect 14004 17484 14056 17536
rect 15200 17484 15252 17536
rect 15292 17484 15344 17536
rect 19156 17620 19208 17672
rect 19616 17620 19668 17672
rect 20536 17620 20588 17672
rect 20260 17484 20312 17536
rect 5894 17382 5946 17434
rect 5958 17382 6010 17434
rect 6022 17382 6074 17434
rect 6086 17382 6138 17434
rect 6150 17382 6202 17434
rect 10839 17382 10891 17434
rect 10903 17382 10955 17434
rect 10967 17382 11019 17434
rect 11031 17382 11083 17434
rect 11095 17382 11147 17434
rect 15784 17382 15836 17434
rect 15848 17382 15900 17434
rect 15912 17382 15964 17434
rect 15976 17382 16028 17434
rect 16040 17382 16092 17434
rect 20729 17382 20781 17434
rect 20793 17382 20845 17434
rect 20857 17382 20909 17434
rect 20921 17382 20973 17434
rect 20985 17382 21037 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 1952 17280 2004 17332
rect 2320 17217 2372 17264
rect 1952 17144 2004 17196
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 2320 17212 2345 17217
rect 2345 17212 2372 17217
rect 3608 17280 3660 17332
rect 3884 17280 3936 17332
rect 6828 17280 6880 17332
rect 7380 17280 7432 17332
rect 4160 17212 4212 17264
rect 4528 17212 4580 17264
rect 4896 17212 4948 17264
rect 4252 17144 4304 17196
rect 5632 17144 5684 17196
rect 2872 17076 2924 17128
rect 3056 17076 3108 17128
rect 4528 17076 4580 17128
rect 4896 17119 4948 17128
rect 4896 17085 4905 17119
rect 4905 17085 4939 17119
rect 4939 17085 4948 17119
rect 4896 17076 4948 17085
rect 6000 17212 6052 17264
rect 8024 17280 8076 17332
rect 8852 17323 8904 17332
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 9772 17280 9824 17332
rect 10416 17280 10468 17332
rect 5908 17144 5960 17196
rect 9956 17212 10008 17264
rect 2964 17008 3016 17060
rect 3424 17008 3476 17060
rect 2780 16940 2832 16992
rect 6000 16940 6052 16992
rect 7564 17076 7616 17128
rect 7288 16940 7340 16992
rect 8760 16940 8812 16992
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 10600 17144 10652 17196
rect 10784 17144 10836 17196
rect 11244 17144 11296 17196
rect 12072 17212 12124 17264
rect 13084 17187 13136 17196
rect 13084 17153 13093 17187
rect 13093 17153 13127 17187
rect 13127 17153 13136 17187
rect 13084 17144 13136 17153
rect 9220 17076 9272 17128
rect 9312 16940 9364 16992
rect 10600 16940 10652 16992
rect 12072 16940 12124 16992
rect 13912 17144 13964 17196
rect 14464 17280 14516 17332
rect 15476 17280 15528 17332
rect 15752 17280 15804 17332
rect 17500 17280 17552 17332
rect 19708 17280 19760 17332
rect 14832 17187 14884 17196
rect 14832 17153 14866 17187
rect 14866 17153 14884 17187
rect 14832 17144 14884 17153
rect 14188 17076 14240 17128
rect 12992 16940 13044 16992
rect 13176 16940 13228 16992
rect 14096 17008 14148 17060
rect 15200 17076 15252 17128
rect 15384 17076 15436 17128
rect 17776 17212 17828 17264
rect 19616 17212 19668 17264
rect 21272 17280 21324 17332
rect 17960 17144 18012 17196
rect 18052 17144 18104 17196
rect 18788 17144 18840 17196
rect 19984 17144 20036 17196
rect 16672 17119 16724 17128
rect 16672 17085 16681 17119
rect 16681 17085 16715 17119
rect 16715 17085 16724 17119
rect 16672 17076 16724 17085
rect 14832 16940 14884 16992
rect 15108 16940 15160 16992
rect 15476 16940 15528 16992
rect 16212 16940 16264 16992
rect 17868 16940 17920 16992
rect 18052 16940 18104 16992
rect 19800 16940 19852 16992
rect 20904 16940 20956 16992
rect 3422 16838 3474 16890
rect 3486 16838 3538 16890
rect 3550 16838 3602 16890
rect 3614 16838 3666 16890
rect 3678 16838 3730 16890
rect 8367 16838 8419 16890
rect 8431 16838 8483 16890
rect 8495 16838 8547 16890
rect 8559 16838 8611 16890
rect 8623 16838 8675 16890
rect 13312 16838 13364 16890
rect 13376 16838 13428 16890
rect 13440 16838 13492 16890
rect 13504 16838 13556 16890
rect 13568 16838 13620 16890
rect 18257 16838 18309 16890
rect 18321 16838 18373 16890
rect 18385 16838 18437 16890
rect 18449 16838 18501 16890
rect 18513 16838 18565 16890
rect 1768 16779 1820 16788
rect 1768 16745 1777 16779
rect 1777 16745 1811 16779
rect 1811 16745 1820 16779
rect 1768 16736 1820 16745
rect 1124 16668 1176 16720
rect 2688 16736 2740 16788
rect 3332 16779 3384 16788
rect 3332 16745 3341 16779
rect 3341 16745 3375 16779
rect 3375 16745 3384 16779
rect 3332 16736 3384 16745
rect 3056 16668 3108 16720
rect 2044 16600 2096 16652
rect 2964 16532 3016 16584
rect 3792 16532 3844 16584
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 204 16464 256 16516
rect 664 16464 716 16516
rect 3056 16464 3108 16516
rect 3332 16464 3384 16516
rect 5356 16711 5408 16720
rect 5356 16677 5365 16711
rect 5365 16677 5399 16711
rect 5399 16677 5408 16711
rect 5356 16668 5408 16677
rect 6644 16736 6696 16788
rect 6828 16736 6880 16788
rect 7012 16736 7064 16788
rect 9956 16736 10008 16788
rect 11336 16736 11388 16788
rect 2320 16396 2372 16448
rect 4896 16464 4948 16516
rect 7104 16600 7156 16652
rect 7380 16600 7432 16652
rect 5080 16532 5132 16584
rect 5540 16532 5592 16584
rect 7748 16575 7800 16584
rect 7748 16541 7755 16575
rect 7755 16541 7789 16575
rect 7789 16541 7800 16575
rect 7748 16532 7800 16541
rect 10140 16600 10192 16652
rect 11336 16600 11388 16652
rect 10416 16532 10468 16584
rect 14096 16736 14148 16788
rect 14188 16736 14240 16788
rect 16212 16736 16264 16788
rect 11428 16532 11480 16584
rect 11796 16532 11848 16584
rect 5356 16464 5408 16516
rect 7012 16464 7064 16516
rect 7564 16464 7616 16516
rect 8944 16464 8996 16516
rect 9864 16464 9916 16516
rect 10048 16464 10100 16516
rect 10232 16507 10284 16516
rect 10232 16473 10241 16507
rect 10241 16473 10275 16507
rect 10275 16473 10284 16507
rect 10232 16464 10284 16473
rect 5816 16396 5868 16448
rect 6184 16396 6236 16448
rect 6368 16396 6420 16448
rect 6552 16396 6604 16448
rect 9772 16396 9824 16448
rect 10784 16464 10836 16516
rect 12164 16464 12216 16516
rect 11244 16396 11296 16448
rect 11336 16396 11388 16448
rect 11428 16396 11480 16448
rect 13176 16532 13228 16584
rect 13728 16532 13780 16584
rect 12992 16464 13044 16516
rect 15108 16575 15160 16584
rect 15108 16541 15117 16575
rect 15117 16541 15151 16575
rect 15151 16541 15160 16575
rect 15752 16600 15804 16652
rect 16028 16643 16080 16652
rect 16028 16609 16037 16643
rect 16037 16609 16071 16643
rect 16071 16609 16080 16643
rect 16028 16600 16080 16609
rect 15108 16532 15160 16541
rect 15394 16575 15446 16584
rect 15394 16541 15403 16575
rect 15403 16541 15437 16575
rect 15437 16541 15446 16575
rect 15394 16532 15446 16541
rect 17500 16736 17552 16788
rect 17960 16736 18012 16788
rect 17960 16600 18012 16652
rect 18696 16600 18748 16652
rect 19616 16668 19668 16720
rect 16580 16464 16632 16516
rect 18420 16575 18472 16584
rect 18420 16541 18429 16575
rect 18429 16541 18463 16575
rect 18463 16541 18472 16575
rect 18420 16532 18472 16541
rect 18788 16532 18840 16584
rect 20444 16643 20496 16652
rect 20444 16609 20453 16643
rect 20453 16609 20487 16643
rect 20487 16609 20496 16643
rect 20444 16600 20496 16609
rect 19708 16575 19760 16584
rect 19708 16541 19717 16575
rect 19717 16541 19751 16575
rect 19751 16541 19760 16575
rect 19708 16532 19760 16541
rect 17684 16396 17736 16448
rect 18052 16396 18104 16448
rect 18512 16439 18564 16448
rect 18512 16405 18521 16439
rect 18521 16405 18555 16439
rect 18555 16405 18564 16439
rect 18512 16396 18564 16405
rect 18880 16396 18932 16448
rect 21088 16396 21140 16448
rect 5894 16294 5946 16346
rect 5958 16294 6010 16346
rect 6022 16294 6074 16346
rect 6086 16294 6138 16346
rect 6150 16294 6202 16346
rect 10839 16294 10891 16346
rect 10903 16294 10955 16346
rect 10967 16294 11019 16346
rect 11031 16294 11083 16346
rect 11095 16294 11147 16346
rect 15784 16294 15836 16346
rect 15848 16294 15900 16346
rect 15912 16294 15964 16346
rect 15976 16294 16028 16346
rect 16040 16294 16092 16346
rect 20729 16294 20781 16346
rect 20793 16294 20845 16346
rect 20857 16294 20909 16346
rect 20921 16294 20973 16346
rect 20985 16294 21037 16346
rect 1584 16235 1636 16244
rect 1584 16201 1593 16235
rect 1593 16201 1627 16235
rect 1627 16201 1636 16235
rect 1584 16192 1636 16201
rect 1952 16192 2004 16244
rect 3148 16192 3200 16244
rect 1676 16124 1728 16176
rect 2228 16124 2280 16176
rect 3424 16124 3476 16176
rect 1952 16056 2004 16108
rect 2504 16056 2556 16108
rect 2780 16056 2832 16108
rect 3148 16075 3155 16108
rect 3155 16075 3189 16108
rect 3189 16075 3200 16108
rect 3148 16056 3200 16075
rect 2136 15895 2188 15904
rect 2136 15861 2145 15895
rect 2145 15861 2179 15895
rect 2179 15861 2188 15895
rect 2136 15852 2188 15861
rect 3792 15852 3844 15904
rect 3884 15895 3936 15904
rect 3884 15861 3893 15895
rect 3893 15861 3927 15895
rect 3927 15861 3936 15895
rect 3884 15852 3936 15861
rect 6460 16192 6512 16244
rect 7380 16192 7432 16244
rect 7656 16192 7708 16244
rect 8116 16192 8168 16244
rect 4620 16056 4672 16108
rect 5264 16099 5316 16108
rect 5264 16065 5298 16099
rect 5298 16065 5316 16099
rect 5264 16056 5316 16065
rect 4344 15988 4396 16040
rect 4712 15920 4764 15972
rect 4528 15852 4580 15904
rect 7472 16099 7524 16108
rect 7472 16065 7506 16099
rect 7506 16065 7524 16099
rect 7472 16056 7524 16065
rect 7656 16099 7708 16108
rect 7656 16065 7665 16099
rect 7665 16065 7699 16099
rect 7699 16065 7708 16099
rect 7656 16056 7708 16065
rect 10048 16192 10100 16244
rect 14004 16192 14056 16244
rect 9772 16099 9824 16108
rect 9772 16065 9806 16099
rect 9806 16065 9824 16099
rect 9772 16056 9824 16065
rect 11704 16056 11756 16108
rect 12440 16056 12492 16108
rect 6000 15988 6052 16040
rect 6460 16031 6512 16040
rect 6460 15997 6469 16031
rect 6469 15997 6503 16031
rect 6503 15997 6512 16031
rect 6460 15988 6512 15997
rect 6552 15988 6604 16040
rect 6736 15988 6788 16040
rect 7196 15988 7248 16040
rect 7012 15920 7064 15972
rect 9404 15963 9456 15972
rect 9404 15929 9413 15963
rect 9413 15929 9447 15963
rect 9447 15929 9456 15963
rect 9404 15920 9456 15929
rect 6184 15852 6236 15904
rect 8760 15852 8812 15904
rect 10140 15988 10192 16040
rect 9864 15852 9916 15904
rect 10048 15852 10100 15904
rect 11796 15988 11848 16040
rect 14740 16192 14792 16244
rect 15200 16192 15252 16244
rect 18052 16192 18104 16244
rect 18420 16192 18472 16244
rect 18512 16192 18564 16244
rect 19708 16235 19760 16244
rect 19708 16201 19717 16235
rect 19717 16201 19751 16235
rect 19751 16201 19760 16235
rect 19708 16192 19760 16201
rect 15016 16099 15068 16108
rect 15016 16065 15025 16099
rect 15025 16065 15059 16099
rect 15059 16065 15068 16099
rect 15016 16056 15068 16065
rect 15292 16099 15344 16108
rect 15292 16065 15301 16099
rect 15301 16065 15335 16099
rect 15335 16065 15344 16099
rect 15292 16056 15344 16065
rect 14280 16031 14332 16040
rect 14280 15997 14289 16031
rect 14289 15997 14323 16031
rect 14323 15997 14332 16031
rect 14280 15988 14332 15997
rect 13820 15852 13872 15904
rect 14096 15920 14148 15972
rect 15660 15988 15712 16040
rect 16212 15988 16264 16040
rect 16948 16124 17000 16176
rect 16672 16056 16724 16108
rect 14740 15963 14792 15972
rect 14740 15929 14749 15963
rect 14749 15929 14783 15963
rect 14783 15929 14792 15963
rect 14740 15920 14792 15929
rect 18696 16031 18748 16040
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 16948 15852 17000 15904
rect 20444 15895 20496 15904
rect 20444 15861 20453 15895
rect 20453 15861 20487 15895
rect 20487 15861 20496 15895
rect 20444 15852 20496 15861
rect 3422 15750 3474 15802
rect 3486 15750 3538 15802
rect 3550 15750 3602 15802
rect 3614 15750 3666 15802
rect 3678 15750 3730 15802
rect 8367 15750 8419 15802
rect 8431 15750 8483 15802
rect 8495 15750 8547 15802
rect 8559 15750 8611 15802
rect 8623 15750 8675 15802
rect 13312 15750 13364 15802
rect 13376 15750 13428 15802
rect 13440 15750 13492 15802
rect 13504 15750 13556 15802
rect 13568 15750 13620 15802
rect 18257 15750 18309 15802
rect 18321 15750 18373 15802
rect 18385 15750 18437 15802
rect 18449 15750 18501 15802
rect 18513 15750 18565 15802
rect 1492 15691 1544 15700
rect 1492 15657 1501 15691
rect 1501 15657 1535 15691
rect 1535 15657 1544 15691
rect 1492 15648 1544 15657
rect 1676 15648 1728 15700
rect 2044 15487 2096 15496
rect 2044 15453 2051 15487
rect 2051 15453 2085 15487
rect 2085 15453 2096 15487
rect 2044 15444 2096 15453
rect 2136 15444 2188 15496
rect 2780 15444 2832 15496
rect 3148 15444 3200 15496
rect 6184 15648 6236 15700
rect 7564 15648 7616 15700
rect 4528 15580 4580 15632
rect 9956 15648 10008 15700
rect 10140 15648 10192 15700
rect 10508 15648 10560 15700
rect 11796 15580 11848 15632
rect 13912 15580 13964 15632
rect 15200 15648 15252 15700
rect 15384 15648 15436 15700
rect 19616 15691 19668 15700
rect 19616 15657 19625 15691
rect 19625 15657 19659 15691
rect 19659 15657 19668 15691
rect 19616 15648 19668 15657
rect 19708 15648 19760 15700
rect 19800 15648 19852 15700
rect 8944 15512 8996 15564
rect 2688 15308 2740 15360
rect 2872 15308 2924 15360
rect 3792 15351 3844 15360
rect 3792 15317 3801 15351
rect 3801 15317 3835 15351
rect 3835 15317 3844 15351
rect 3792 15308 3844 15317
rect 3884 15308 3936 15360
rect 5448 15444 5500 15496
rect 5816 15444 5868 15496
rect 6276 15444 6328 15496
rect 7472 15487 7524 15496
rect 7472 15453 7481 15487
rect 7481 15453 7515 15487
rect 7515 15453 7524 15487
rect 7472 15444 7524 15453
rect 7748 15487 7800 15496
rect 7748 15453 7755 15487
rect 7755 15453 7789 15487
rect 7789 15453 7800 15487
rect 7748 15444 7800 15453
rect 8668 15376 8720 15428
rect 9312 15487 9364 15496
rect 9312 15453 9319 15487
rect 9319 15453 9353 15487
rect 9353 15453 9364 15487
rect 9312 15444 9364 15453
rect 10140 15512 10192 15564
rect 9588 15376 9640 15428
rect 13176 15512 13228 15564
rect 11520 15444 11572 15496
rect 12440 15444 12492 15496
rect 14556 15580 14608 15632
rect 19524 15580 19576 15632
rect 15016 15555 15068 15564
rect 15016 15521 15025 15555
rect 15025 15521 15059 15555
rect 15059 15521 15068 15555
rect 15016 15512 15068 15521
rect 15200 15512 15252 15564
rect 15660 15512 15712 15564
rect 13912 15444 13964 15496
rect 14096 15487 14148 15496
rect 14096 15453 14105 15487
rect 14105 15453 14139 15487
rect 14139 15453 14148 15487
rect 14096 15444 14148 15453
rect 14464 15444 14516 15496
rect 15292 15487 15344 15496
rect 15292 15453 15301 15487
rect 15301 15453 15335 15487
rect 15335 15453 15344 15487
rect 15292 15444 15344 15453
rect 17316 15512 17368 15564
rect 19340 15512 19392 15564
rect 5448 15308 5500 15360
rect 6644 15308 6696 15360
rect 7564 15308 7616 15360
rect 7932 15308 7984 15360
rect 11244 15308 11296 15360
rect 16212 15444 16264 15496
rect 17408 15444 17460 15496
rect 16580 15376 16632 15428
rect 18696 15487 18748 15496
rect 18696 15453 18705 15487
rect 18705 15453 18739 15487
rect 18739 15453 18748 15487
rect 18696 15444 18748 15453
rect 19064 15487 19116 15496
rect 19064 15453 19073 15487
rect 19073 15453 19107 15487
rect 19107 15453 19116 15487
rect 19064 15444 19116 15453
rect 19248 15487 19300 15496
rect 19248 15453 19257 15487
rect 19257 15453 19291 15487
rect 19291 15453 19300 15487
rect 19248 15444 19300 15453
rect 19156 15376 19208 15428
rect 16948 15308 17000 15360
rect 18604 15308 18656 15360
rect 18788 15308 18840 15360
rect 19340 15351 19392 15360
rect 19340 15317 19349 15351
rect 19349 15317 19383 15351
rect 19383 15317 19392 15351
rect 19340 15308 19392 15317
rect 19984 15308 20036 15360
rect 21272 15376 21324 15428
rect 5894 15206 5946 15258
rect 5958 15206 6010 15258
rect 6022 15206 6074 15258
rect 6086 15206 6138 15258
rect 6150 15206 6202 15258
rect 10839 15206 10891 15258
rect 10903 15206 10955 15258
rect 10967 15206 11019 15258
rect 11031 15206 11083 15258
rect 11095 15206 11147 15258
rect 15784 15206 15836 15258
rect 15848 15206 15900 15258
rect 15912 15206 15964 15258
rect 15976 15206 16028 15258
rect 16040 15206 16092 15258
rect 20729 15206 20781 15258
rect 20793 15206 20845 15258
rect 20857 15206 20909 15258
rect 20921 15206 20973 15258
rect 20985 15206 21037 15258
rect 848 15104 900 15156
rect 1952 15104 2004 15156
rect 2228 15104 2280 15156
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 2044 14968 2096 15020
rect 2688 15036 2740 15088
rect 2964 15036 3016 15088
rect 3884 15036 3936 15088
rect 4068 15036 4120 15088
rect 4252 15036 4304 15088
rect 4528 14968 4580 15020
rect 5080 14968 5132 15020
rect 7288 15011 7340 15020
rect 7288 14977 7297 15011
rect 7297 14977 7331 15011
rect 7331 14977 7340 15011
rect 7288 14968 7340 14977
rect 8300 14968 8352 15020
rect 11336 15104 11388 15156
rect 11704 15104 11756 15156
rect 12072 15104 12124 15156
rect 12256 15104 12308 15156
rect 12624 15104 12676 15156
rect 14740 15104 14792 15156
rect 16120 15104 16172 15156
rect 16488 15104 16540 15156
rect 16580 15104 16632 15156
rect 20536 15104 20588 15156
rect 10968 15036 11020 15088
rect 11060 15036 11112 15088
rect 11520 15036 11572 15088
rect 13820 15036 13872 15088
rect 15660 15036 15712 15088
rect 11796 14968 11848 15020
rect 11980 14968 12032 15020
rect 12164 14968 12216 15020
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 14004 14968 14056 14977
rect 17684 15036 17736 15088
rect 2964 14900 3016 14952
rect 480 14764 532 14816
rect 1124 14764 1176 14816
rect 3148 14807 3200 14816
rect 3148 14773 3157 14807
rect 3157 14773 3191 14807
rect 3191 14773 3200 14807
rect 3148 14764 3200 14773
rect 4252 14900 4304 14952
rect 4712 14900 4764 14952
rect 6552 14943 6604 14952
rect 6552 14909 6561 14943
rect 6561 14909 6595 14943
rect 6595 14909 6604 14943
rect 6552 14900 6604 14909
rect 6644 14900 6696 14952
rect 7380 14943 7432 14952
rect 7380 14909 7414 14943
rect 7414 14909 7432 14943
rect 7380 14900 7432 14909
rect 6460 14832 6512 14884
rect 6920 14832 6972 14884
rect 8576 14832 8628 14884
rect 10968 14900 11020 14952
rect 11612 14900 11664 14952
rect 9128 14764 9180 14816
rect 9864 14832 9916 14884
rect 12440 14900 12492 14952
rect 12624 14900 12676 14952
rect 13268 14943 13320 14952
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 13636 14900 13688 14952
rect 13820 14900 13872 14952
rect 17500 14968 17552 15020
rect 18144 15011 18196 15020
rect 18144 14977 18153 15011
rect 18153 14977 18187 15011
rect 18187 14977 18196 15011
rect 18144 14968 18196 14977
rect 19432 15036 19484 15088
rect 18512 14968 18564 15020
rect 18696 15011 18748 15020
rect 18696 14977 18719 15011
rect 18719 14977 18748 15011
rect 18696 14968 18748 14977
rect 11612 14764 11664 14816
rect 11704 14764 11756 14816
rect 14832 14764 14884 14816
rect 15200 14764 15252 14816
rect 15660 14764 15712 14816
rect 15936 14807 15988 14816
rect 15936 14773 15945 14807
rect 15945 14773 15979 14807
rect 15979 14773 15988 14807
rect 15936 14764 15988 14773
rect 16120 14764 16172 14816
rect 18052 14807 18104 14816
rect 18052 14773 18061 14807
rect 18061 14773 18095 14807
rect 18095 14773 18104 14807
rect 18052 14764 18104 14773
rect 18604 14764 18656 14816
rect 19064 14764 19116 14816
rect 20076 14832 20128 14884
rect 19708 14764 19760 14816
rect 20444 14807 20496 14816
rect 20444 14773 20453 14807
rect 20453 14773 20487 14807
rect 20487 14773 20496 14807
rect 20444 14764 20496 14773
rect 3422 14662 3474 14714
rect 3486 14662 3538 14714
rect 3550 14662 3602 14714
rect 3614 14662 3666 14714
rect 3678 14662 3730 14714
rect 8367 14662 8419 14714
rect 8431 14662 8483 14714
rect 8495 14662 8547 14714
rect 8559 14662 8611 14714
rect 8623 14662 8675 14714
rect 13312 14662 13364 14714
rect 13376 14662 13428 14714
rect 13440 14662 13492 14714
rect 13504 14662 13556 14714
rect 13568 14662 13620 14714
rect 18257 14662 18309 14714
rect 18321 14662 18373 14714
rect 18385 14662 18437 14714
rect 18449 14662 18501 14714
rect 18513 14662 18565 14714
rect 664 14560 716 14612
rect 3148 14492 3200 14544
rect 664 14424 716 14476
rect 1308 14424 1360 14476
rect 2044 14424 2096 14476
rect 3700 14424 3752 14476
rect 4068 14424 4120 14476
rect 4712 14467 4764 14476
rect 4712 14433 4721 14467
rect 4721 14433 4755 14467
rect 4755 14433 4764 14467
rect 4712 14424 4764 14433
rect 4804 14467 4856 14476
rect 4804 14433 4838 14467
rect 4838 14433 4856 14467
rect 5448 14560 5500 14612
rect 11704 14560 11756 14612
rect 13636 14560 13688 14612
rect 14924 14560 14976 14612
rect 15936 14560 15988 14612
rect 9404 14492 9456 14544
rect 9864 14492 9916 14544
rect 4804 14424 4856 14433
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 2596 14399 2648 14408
rect 2596 14365 2603 14399
rect 2603 14365 2637 14399
rect 2637 14365 2648 14399
rect 2596 14356 2648 14365
rect 3148 14356 3200 14408
rect 2228 14220 2280 14272
rect 2504 14220 2556 14272
rect 5816 14356 5868 14408
rect 6920 14356 6972 14408
rect 6184 14288 6236 14340
rect 4344 14220 4396 14272
rect 4528 14220 4580 14272
rect 6276 14220 6328 14272
rect 7196 14356 7248 14408
rect 7288 14356 7340 14408
rect 7472 14399 7524 14408
rect 7472 14365 7481 14399
rect 7481 14365 7515 14399
rect 7515 14365 7524 14399
rect 7472 14356 7524 14365
rect 7748 14399 7800 14408
rect 7748 14365 7755 14399
rect 7755 14365 7789 14399
rect 7789 14365 7800 14399
rect 7748 14356 7800 14365
rect 10324 14467 10376 14476
rect 10324 14433 10358 14467
rect 10358 14433 10376 14467
rect 10324 14424 10376 14433
rect 11612 14424 11664 14476
rect 14004 14424 14056 14476
rect 16856 14467 16908 14476
rect 16856 14433 16865 14467
rect 16865 14433 16899 14467
rect 16899 14433 16908 14467
rect 16856 14424 16908 14433
rect 18604 14560 18656 14612
rect 19248 14560 19300 14612
rect 8668 14356 8720 14408
rect 9680 14356 9732 14408
rect 10508 14399 10560 14408
rect 10508 14365 10517 14399
rect 10517 14365 10551 14399
rect 10551 14365 10560 14399
rect 10508 14356 10560 14365
rect 11244 14356 11296 14408
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 14372 14399 14424 14408
rect 14372 14365 14379 14399
rect 14379 14365 14413 14399
rect 14413 14365 14424 14399
rect 14372 14356 14424 14365
rect 14740 14356 14792 14408
rect 15016 14356 15068 14408
rect 15384 14356 15436 14408
rect 12440 14288 12492 14340
rect 12624 14288 12676 14340
rect 16488 14356 16540 14408
rect 7472 14220 7524 14272
rect 11980 14220 12032 14272
rect 12992 14220 13044 14272
rect 16212 14288 16264 14340
rect 16580 14288 16632 14340
rect 14740 14220 14792 14272
rect 18144 14356 18196 14408
rect 18696 14492 18748 14544
rect 21916 14560 21968 14612
rect 18788 14424 18840 14476
rect 18972 14424 19024 14476
rect 19248 14467 19300 14476
rect 19248 14433 19257 14467
rect 19257 14433 19291 14467
rect 19291 14433 19300 14467
rect 19248 14424 19300 14433
rect 17408 14220 17460 14272
rect 17684 14220 17736 14272
rect 19432 14220 19484 14272
rect 19616 14220 19668 14272
rect 20168 14220 20220 14272
rect 5894 14118 5946 14170
rect 5958 14118 6010 14170
rect 6022 14118 6074 14170
rect 6086 14118 6138 14170
rect 6150 14118 6202 14170
rect 10839 14118 10891 14170
rect 10903 14118 10955 14170
rect 10967 14118 11019 14170
rect 11031 14118 11083 14170
rect 11095 14118 11147 14170
rect 15784 14118 15836 14170
rect 15848 14118 15900 14170
rect 15912 14118 15964 14170
rect 15976 14118 16028 14170
rect 16040 14118 16092 14170
rect 20729 14118 20781 14170
rect 20793 14118 20845 14170
rect 20857 14118 20909 14170
rect 20921 14118 20973 14170
rect 20985 14118 21037 14170
rect 1952 14059 2004 14068
rect 1952 14025 1961 14059
rect 1961 14025 1995 14059
rect 1995 14025 2004 14059
rect 1952 14016 2004 14025
rect 3056 14016 3108 14068
rect 1768 13948 1820 14000
rect 4068 13948 4120 14000
rect 3332 13923 3384 13932
rect 3332 13889 3366 13923
rect 3366 13889 3384 13923
rect 3332 13880 3384 13889
rect 3516 13923 3568 13932
rect 3516 13889 3525 13923
rect 3525 13889 3559 13923
rect 3559 13889 3568 13923
rect 3516 13880 3568 13889
rect 4160 13880 4212 13932
rect 4436 13923 4488 13932
rect 4436 13889 4445 13923
rect 4445 13889 4479 13923
rect 4479 13889 4488 13923
rect 4436 13880 4488 13889
rect 112 13812 164 13864
rect 2228 13812 2280 13864
rect 2504 13855 2556 13864
rect 2504 13821 2513 13855
rect 2513 13821 2547 13855
rect 2547 13821 2556 13855
rect 2504 13812 2556 13821
rect 2872 13812 2924 13864
rect 5080 13880 5132 13932
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 7288 13923 7340 13932
rect 7288 13889 7297 13923
rect 7297 13889 7331 13923
rect 7331 13889 7340 13923
rect 7288 13880 7340 13889
rect 7380 13923 7432 13932
rect 7380 13889 7414 13923
rect 7414 13889 7432 13923
rect 7380 13880 7432 13889
rect 1952 13676 2004 13728
rect 2320 13676 2372 13728
rect 3700 13676 3752 13728
rect 4068 13744 4120 13796
rect 4712 13744 4764 13796
rect 3976 13676 4028 13728
rect 4436 13676 4488 13728
rect 4804 13676 4856 13728
rect 6092 13812 6144 13864
rect 5816 13744 5868 13796
rect 5632 13676 5684 13728
rect 8208 13719 8260 13728
rect 8208 13685 8217 13719
rect 8217 13685 8251 13719
rect 8251 13685 8260 13719
rect 8208 13676 8260 13685
rect 8852 14016 8904 14068
rect 10232 14016 10284 14068
rect 10600 14016 10652 14068
rect 11428 14016 11480 14068
rect 13176 14016 13228 14068
rect 15660 14016 15712 14068
rect 9036 13948 9088 14000
rect 9496 13948 9548 14000
rect 12532 13948 12584 14000
rect 9036 13812 9088 13864
rect 9864 13880 9916 13932
rect 10600 13880 10652 13932
rect 12900 13948 12952 14000
rect 13820 13948 13872 14000
rect 14188 13948 14240 14000
rect 15200 13880 15252 13932
rect 15660 13880 15712 13932
rect 16212 13923 16264 13932
rect 16212 13889 16221 13923
rect 16221 13889 16255 13923
rect 16255 13889 16264 13923
rect 16212 13880 16264 13889
rect 18052 13948 18104 14000
rect 18696 13948 18748 14000
rect 8668 13744 8720 13796
rect 8852 13744 8904 13796
rect 9128 13744 9180 13796
rect 9404 13744 9456 13796
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 10876 13812 10928 13864
rect 12256 13812 12308 13864
rect 10140 13787 10192 13796
rect 10140 13753 10149 13787
rect 10149 13753 10183 13787
rect 10183 13753 10192 13787
rect 10140 13744 10192 13753
rect 11428 13676 11480 13728
rect 14004 13855 14056 13864
rect 14004 13821 14013 13855
rect 14013 13821 14047 13855
rect 14047 13821 14056 13855
rect 14004 13812 14056 13821
rect 15292 13812 15344 13864
rect 15384 13812 15436 13864
rect 17500 13880 17552 13932
rect 15568 13744 15620 13796
rect 15752 13744 15804 13796
rect 16212 13744 16264 13796
rect 16396 13676 16448 13728
rect 18144 13812 18196 13864
rect 18604 13923 18656 13932
rect 18604 13889 18613 13923
rect 18613 13889 18647 13923
rect 18647 13889 18656 13923
rect 18604 13880 18656 13889
rect 18972 13923 19024 13932
rect 18972 13889 18981 13923
rect 18981 13889 19015 13923
rect 19015 13889 19024 13923
rect 18972 13880 19024 13889
rect 19524 13855 19576 13864
rect 19524 13821 19533 13855
rect 19533 13821 19567 13855
rect 19567 13821 19576 13855
rect 19524 13812 19576 13821
rect 20168 14016 20220 14068
rect 21272 14016 21324 14068
rect 20168 13923 20220 13932
rect 20168 13889 20177 13923
rect 20177 13889 20211 13923
rect 20211 13889 20220 13923
rect 20168 13880 20220 13889
rect 19064 13744 19116 13796
rect 19340 13744 19392 13796
rect 17316 13676 17368 13728
rect 17592 13676 17644 13728
rect 18236 13676 18288 13728
rect 18604 13676 18656 13728
rect 3422 13574 3474 13626
rect 3486 13574 3538 13626
rect 3550 13574 3602 13626
rect 3614 13574 3666 13626
rect 3678 13574 3730 13626
rect 8367 13574 8419 13626
rect 8431 13574 8483 13626
rect 8495 13574 8547 13626
rect 8559 13574 8611 13626
rect 8623 13574 8675 13626
rect 13312 13574 13364 13626
rect 13376 13574 13428 13626
rect 13440 13574 13492 13626
rect 13504 13574 13556 13626
rect 13568 13574 13620 13626
rect 18257 13574 18309 13626
rect 18321 13574 18373 13626
rect 18385 13574 18437 13626
rect 18449 13574 18501 13626
rect 18513 13574 18565 13626
rect 1584 13515 1636 13524
rect 1584 13481 1593 13515
rect 1593 13481 1627 13515
rect 1627 13481 1636 13515
rect 1584 13472 1636 13481
rect 3332 13472 3384 13524
rect 3976 13515 4028 13524
rect 3976 13481 3985 13515
rect 3985 13481 4019 13515
rect 4019 13481 4028 13515
rect 3976 13472 4028 13481
rect 3700 13404 3752 13456
rect 204 13268 256 13320
rect 1584 13268 1636 13320
rect 8208 13472 8260 13524
rect 9588 13472 9640 13524
rect 6460 13404 6512 13456
rect 6644 13447 6696 13456
rect 6644 13413 6653 13447
rect 6653 13413 6687 13447
rect 6687 13413 6696 13447
rect 6644 13404 6696 13413
rect 9220 13404 9272 13456
rect 9404 13404 9456 13456
rect 10416 13472 10468 13524
rect 11612 13472 11664 13524
rect 14096 13472 14148 13524
rect 15292 13472 15344 13524
rect 1860 13200 1912 13252
rect 2228 13200 2280 13252
rect 4528 13311 4580 13320
rect 4528 13277 4537 13311
rect 4537 13277 4571 13311
rect 4571 13277 4580 13311
rect 4528 13268 4580 13277
rect 4804 13268 4856 13320
rect 4988 13268 5040 13320
rect 5356 13268 5408 13320
rect 6092 13336 6144 13388
rect 6368 13336 6420 13388
rect 14188 13404 14240 13456
rect 3148 13200 3200 13252
rect 4436 13200 4488 13252
rect 3608 13132 3660 13184
rect 4344 13175 4396 13184
rect 4344 13141 4353 13175
rect 4353 13141 4387 13175
rect 4387 13141 4396 13175
rect 4344 13132 4396 13141
rect 5080 13132 5132 13184
rect 6920 13311 6972 13320
rect 6920 13277 6929 13311
rect 6929 13277 6963 13311
rect 6963 13277 6972 13311
rect 6920 13268 6972 13277
rect 6552 13132 6604 13184
rect 7012 13132 7064 13184
rect 7840 13268 7892 13320
rect 9128 13268 9180 13320
rect 9680 13268 9732 13320
rect 11520 13336 11572 13388
rect 11888 13336 11940 13388
rect 14556 13404 14608 13456
rect 14740 13447 14792 13456
rect 14740 13413 14749 13447
rect 14749 13413 14783 13447
rect 14783 13413 14792 13447
rect 14740 13404 14792 13413
rect 14648 13336 14700 13388
rect 17408 13472 17460 13524
rect 18144 13472 18196 13524
rect 18972 13472 19024 13524
rect 19708 13472 19760 13524
rect 19248 13379 19300 13388
rect 19248 13345 19257 13379
rect 19257 13345 19291 13379
rect 19291 13345 19300 13379
rect 19248 13336 19300 13345
rect 9404 13200 9456 13252
rect 10784 13268 10836 13320
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 12164 13268 12216 13320
rect 12532 13268 12584 13320
rect 12716 13200 12768 13252
rect 14188 13268 14240 13320
rect 15016 13311 15068 13320
rect 15016 13277 15025 13311
rect 15025 13277 15059 13311
rect 15059 13277 15068 13311
rect 15016 13268 15068 13277
rect 16212 13268 16264 13320
rect 16672 13268 16724 13320
rect 13084 13200 13136 13252
rect 15936 13243 15988 13252
rect 15936 13209 15945 13243
rect 15945 13209 15979 13243
rect 15979 13209 15988 13243
rect 15936 13200 15988 13209
rect 16488 13200 16540 13252
rect 17040 13200 17092 13252
rect 17868 13200 17920 13252
rect 7840 13175 7892 13184
rect 7840 13141 7849 13175
rect 7849 13141 7883 13175
rect 7883 13141 7892 13175
rect 7840 13132 7892 13141
rect 8208 13132 8260 13184
rect 11980 13132 12032 13184
rect 12992 13132 13044 13184
rect 13912 13132 13964 13184
rect 18420 13132 18472 13184
rect 18604 13132 18656 13184
rect 5894 13030 5946 13082
rect 5958 13030 6010 13082
rect 6022 13030 6074 13082
rect 6086 13030 6138 13082
rect 6150 13030 6202 13082
rect 10839 13030 10891 13082
rect 10903 13030 10955 13082
rect 10967 13030 11019 13082
rect 11031 13030 11083 13082
rect 11095 13030 11147 13082
rect 15784 13030 15836 13082
rect 15848 13030 15900 13082
rect 15912 13030 15964 13082
rect 15976 13030 16028 13082
rect 16040 13030 16092 13082
rect 20729 13030 20781 13082
rect 20793 13030 20845 13082
rect 20857 13030 20909 13082
rect 20921 13030 20973 13082
rect 20985 13030 21037 13082
rect 1676 12928 1728 12980
rect 4344 12928 4396 12980
rect 3792 12860 3844 12912
rect 6736 12928 6788 12980
rect 7564 12928 7616 12980
rect 7840 12928 7892 12980
rect 8300 12971 8352 12980
rect 8300 12937 8309 12971
rect 8309 12937 8343 12971
rect 8343 12937 8352 12971
rect 8300 12928 8352 12937
rect 8668 12928 8720 12980
rect 2872 12792 2924 12844
rect 3240 12835 3292 12844
rect 3240 12801 3247 12835
rect 3247 12801 3281 12835
rect 3281 12801 3292 12835
rect 3240 12792 3292 12801
rect 3608 12792 3660 12844
rect 3700 12792 3752 12844
rect 2320 12724 2372 12776
rect 2964 12767 3016 12776
rect 2964 12733 2973 12767
rect 2973 12733 3007 12767
rect 3007 12733 3016 12767
rect 2964 12724 3016 12733
rect 4068 12724 4120 12776
rect 4988 12860 5040 12912
rect 7472 12792 7524 12844
rect 8116 12792 8168 12844
rect 9312 12860 9364 12912
rect 10508 12928 10560 12980
rect 11888 12928 11940 12980
rect 13728 12928 13780 12980
rect 11980 12860 12032 12912
rect 12164 12860 12216 12912
rect 13084 12860 13136 12912
rect 11704 12792 11756 12844
rect 12440 12835 12492 12844
rect 12440 12801 12449 12835
rect 12449 12801 12483 12835
rect 12483 12801 12492 12835
rect 12440 12792 12492 12801
rect 12992 12792 13044 12844
rect 14280 12860 14332 12912
rect 18052 12928 18104 12980
rect 18144 12928 18196 12980
rect 20168 12928 20220 12980
rect 21272 12928 21324 12980
rect 14004 12792 14056 12844
rect 14648 12792 14700 12844
rect 15292 12835 15344 12844
rect 15292 12801 15326 12835
rect 15326 12801 15344 12835
rect 15292 12792 15344 12801
rect 16396 12792 16448 12844
rect 16948 12835 17000 12844
rect 16948 12801 16955 12835
rect 16955 12801 16989 12835
rect 16989 12801 17000 12835
rect 16948 12792 17000 12801
rect 4804 12724 4856 12776
rect 2044 12631 2096 12640
rect 2044 12597 2053 12631
rect 2053 12597 2087 12631
rect 2087 12597 2096 12631
rect 2044 12588 2096 12597
rect 2596 12631 2648 12640
rect 2596 12597 2605 12631
rect 2605 12597 2639 12631
rect 2639 12597 2648 12631
rect 2596 12588 2648 12597
rect 2688 12588 2740 12640
rect 5632 12656 5684 12708
rect 5816 12588 5868 12640
rect 6368 12699 6420 12708
rect 6368 12665 6377 12699
rect 6377 12665 6411 12699
rect 6411 12665 6420 12699
rect 6368 12656 6420 12665
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 7380 12588 7432 12640
rect 12532 12724 12584 12776
rect 13176 12724 13228 12776
rect 10140 12588 10192 12640
rect 11888 12588 11940 12640
rect 14648 12588 14700 12640
rect 15016 12724 15068 12776
rect 15568 12588 15620 12640
rect 16212 12724 16264 12776
rect 19432 12860 19484 12912
rect 18604 12835 18656 12844
rect 18604 12801 18613 12835
rect 18613 12801 18647 12835
rect 18647 12801 18656 12835
rect 18604 12792 18656 12801
rect 18788 12792 18840 12844
rect 18328 12767 18380 12776
rect 18328 12733 18337 12767
rect 18337 12733 18371 12767
rect 18371 12733 18380 12767
rect 18328 12724 18380 12733
rect 18420 12724 18472 12776
rect 21364 12724 21416 12776
rect 16120 12699 16172 12708
rect 16120 12665 16129 12699
rect 16129 12665 16163 12699
rect 16163 12665 16172 12699
rect 16120 12656 16172 12665
rect 18144 12631 18196 12640
rect 18144 12597 18153 12631
rect 18153 12597 18187 12631
rect 18187 12597 18196 12631
rect 18144 12588 18196 12597
rect 18604 12588 18656 12640
rect 19524 12656 19576 12708
rect 19984 12656 20036 12708
rect 21272 12656 21324 12708
rect 19340 12631 19392 12640
rect 19340 12597 19349 12631
rect 19349 12597 19383 12631
rect 19383 12597 19392 12631
rect 19340 12588 19392 12597
rect 19892 12631 19944 12640
rect 19892 12597 19901 12631
rect 19901 12597 19935 12631
rect 19935 12597 19944 12631
rect 19892 12588 19944 12597
rect 3422 12486 3474 12538
rect 3486 12486 3538 12538
rect 3550 12486 3602 12538
rect 3614 12486 3666 12538
rect 3678 12486 3730 12538
rect 8367 12486 8419 12538
rect 8431 12486 8483 12538
rect 8495 12486 8547 12538
rect 8559 12486 8611 12538
rect 8623 12486 8675 12538
rect 13312 12486 13364 12538
rect 13376 12486 13428 12538
rect 13440 12486 13492 12538
rect 13504 12486 13556 12538
rect 13568 12486 13620 12538
rect 18257 12486 18309 12538
rect 18321 12486 18373 12538
rect 18385 12486 18437 12538
rect 18449 12486 18501 12538
rect 18513 12486 18565 12538
rect 940 12384 992 12436
rect 4160 12427 4212 12436
rect 4160 12393 4169 12427
rect 4169 12393 4203 12427
rect 4203 12393 4212 12427
rect 4160 12384 4212 12393
rect 4528 12384 4580 12436
rect 5172 12384 5224 12436
rect 5724 12384 5776 12436
rect 6368 12316 6420 12368
rect 6828 12316 6880 12368
rect 2320 12291 2372 12300
rect 2320 12257 2329 12291
rect 2329 12257 2363 12291
rect 2363 12257 2372 12291
rect 2320 12248 2372 12257
rect 4436 12248 4488 12300
rect 1584 12180 1636 12232
rect 20 12112 72 12164
rect 2320 12112 2372 12164
rect 2412 12112 2464 12164
rect 3608 12180 3660 12232
rect 3976 12180 4028 12232
rect 5172 12248 5224 12300
rect 5816 12291 5868 12300
rect 5816 12257 5825 12291
rect 5825 12257 5859 12291
rect 5859 12257 5868 12291
rect 5816 12248 5868 12257
rect 5540 12223 5592 12232
rect 5540 12189 5549 12223
rect 5549 12189 5583 12223
rect 5583 12189 5592 12223
rect 5540 12180 5592 12189
rect 5724 12180 5776 12232
rect 8208 12384 8260 12436
rect 9404 12384 9456 12436
rect 9588 12384 9640 12436
rect 8668 12316 8720 12368
rect 7380 12248 7432 12300
rect 8208 12248 8260 12300
rect 9220 12248 9272 12300
rect 11244 12384 11296 12436
rect 13912 12384 13964 12436
rect 14464 12384 14516 12436
rect 9864 12316 9916 12368
rect 14004 12316 14056 12368
rect 14648 12316 14700 12368
rect 18144 12384 18196 12436
rect 19064 12384 19116 12436
rect 18236 12316 18288 12368
rect 19156 12316 19208 12368
rect 19248 12316 19300 12368
rect 19984 12316 20036 12368
rect 10048 12291 10100 12300
rect 10048 12257 10057 12291
rect 10057 12257 10091 12291
rect 10091 12257 10100 12291
rect 10048 12248 10100 12257
rect 10140 12248 10192 12300
rect 10416 12291 10468 12300
rect 10416 12257 10450 12291
rect 10450 12257 10468 12291
rect 10416 12248 10468 12257
rect 12624 12248 12676 12300
rect 8300 12180 8352 12232
rect 8576 12180 8628 12232
rect 8852 12180 8904 12232
rect 2964 12044 3016 12096
rect 9312 12112 9364 12164
rect 4436 12044 4488 12096
rect 6552 12087 6604 12096
rect 6552 12053 6561 12087
rect 6561 12053 6595 12087
rect 6595 12053 6604 12087
rect 6552 12044 6604 12053
rect 6828 12087 6880 12096
rect 6828 12053 6837 12087
rect 6837 12053 6871 12087
rect 6871 12053 6880 12087
rect 6828 12044 6880 12053
rect 7104 12044 7156 12096
rect 7380 12044 7432 12096
rect 10600 12223 10652 12232
rect 10600 12189 10609 12223
rect 10609 12189 10643 12223
rect 10643 12189 10652 12223
rect 10600 12180 10652 12189
rect 12164 12223 12216 12232
rect 12164 12189 12173 12223
rect 12173 12189 12207 12223
rect 12207 12189 12216 12223
rect 12164 12180 12216 12189
rect 13084 12180 13136 12232
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 14096 12248 14148 12300
rect 14188 12223 14240 12232
rect 14188 12189 14197 12223
rect 14197 12189 14231 12223
rect 14231 12189 14240 12223
rect 14188 12180 14240 12189
rect 9864 12044 9916 12096
rect 10416 12044 10468 12096
rect 11244 12087 11296 12096
rect 11244 12053 11253 12087
rect 11253 12053 11287 12087
rect 11287 12053 11296 12087
rect 11244 12044 11296 12053
rect 11980 12044 12032 12096
rect 12256 12155 12308 12164
rect 12256 12121 12265 12155
rect 12265 12121 12299 12155
rect 12299 12121 12308 12155
rect 12256 12112 12308 12121
rect 13636 12112 13688 12164
rect 15292 12248 15344 12300
rect 17316 12248 17368 12300
rect 14556 12180 14608 12232
rect 16028 12180 16080 12232
rect 15936 12112 15988 12164
rect 16856 12180 16908 12232
rect 16764 12112 16816 12164
rect 16948 12112 17000 12164
rect 18052 12180 18104 12232
rect 18604 12180 18656 12232
rect 19708 12180 19760 12232
rect 12992 12087 13044 12096
rect 12992 12053 13001 12087
rect 13001 12053 13035 12087
rect 13035 12053 13044 12087
rect 12992 12044 13044 12053
rect 13084 12044 13136 12096
rect 18328 12044 18380 12096
rect 18512 12044 18564 12096
rect 18880 12044 18932 12096
rect 19248 12044 19300 12096
rect 20260 12223 20312 12232
rect 20260 12189 20269 12223
rect 20269 12189 20303 12223
rect 20303 12189 20312 12223
rect 20260 12180 20312 12189
rect 5894 11942 5946 11994
rect 5958 11942 6010 11994
rect 6022 11942 6074 11994
rect 6086 11942 6138 11994
rect 6150 11942 6202 11994
rect 10839 11942 10891 11994
rect 10903 11942 10955 11994
rect 10967 11942 11019 11994
rect 11031 11942 11083 11994
rect 11095 11942 11147 11994
rect 15784 11942 15836 11994
rect 15848 11942 15900 11994
rect 15912 11942 15964 11994
rect 15976 11942 16028 11994
rect 16040 11942 16092 11994
rect 20729 11942 20781 11994
rect 20793 11942 20845 11994
rect 20857 11942 20909 11994
rect 20921 11942 20973 11994
rect 20985 11942 21037 11994
rect 848 11840 900 11892
rect 3884 11840 3936 11892
rect 4896 11840 4948 11892
rect 1032 11772 1084 11824
rect 2596 11772 2648 11824
rect 2872 11772 2924 11824
rect 1952 11704 2004 11756
rect 2320 11747 2372 11756
rect 2320 11713 2329 11747
rect 2329 11713 2372 11747
rect 2320 11704 2372 11713
rect 3240 11704 3292 11756
rect 2044 11679 2096 11688
rect 2044 11645 2053 11679
rect 2053 11645 2087 11679
rect 2087 11645 2096 11679
rect 2044 11636 2096 11645
rect 3332 11636 3384 11688
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 4528 11704 4580 11756
rect 4160 11636 4212 11688
rect 3516 11568 3568 11620
rect 3884 11568 3936 11620
rect 4068 11611 4120 11620
rect 4068 11577 4077 11611
rect 4077 11577 4111 11611
rect 4111 11577 4120 11611
rect 4068 11568 4120 11577
rect 5356 11840 5408 11892
rect 5540 11883 5592 11892
rect 5540 11849 5549 11883
rect 5549 11849 5583 11883
rect 5583 11849 5592 11883
rect 5540 11840 5592 11849
rect 5632 11840 5684 11892
rect 6828 11840 6880 11892
rect 7012 11840 7064 11892
rect 10232 11840 10284 11892
rect 10692 11840 10744 11892
rect 12256 11840 12308 11892
rect 15384 11840 15436 11892
rect 15568 11840 15620 11892
rect 8668 11772 8720 11824
rect 5356 11704 5408 11756
rect 5540 11704 5592 11756
rect 6092 11704 6144 11756
rect 6184 11704 6236 11756
rect 7380 11747 7432 11756
rect 7380 11713 7414 11747
rect 7414 11713 7432 11747
rect 8852 11815 8904 11824
rect 8852 11781 8861 11815
rect 8861 11781 8895 11815
rect 8895 11781 8904 11815
rect 8852 11772 8904 11781
rect 9404 11772 9456 11824
rect 12164 11772 12216 11824
rect 7380 11704 7432 11713
rect 9036 11704 9088 11756
rect 9220 11747 9272 11756
rect 9220 11713 9229 11747
rect 9229 11713 9263 11747
rect 9263 11713 9272 11747
rect 9220 11704 9272 11713
rect 11612 11704 11664 11756
rect 11888 11704 11940 11756
rect 12256 11704 12308 11756
rect 12900 11772 12952 11824
rect 13268 11704 13320 11756
rect 13728 11747 13780 11756
rect 13728 11713 13737 11747
rect 13737 11713 13771 11747
rect 13771 11713 13780 11747
rect 13728 11704 13780 11713
rect 16304 11772 16356 11824
rect 14096 11704 14148 11756
rect 5724 11636 5776 11688
rect 6368 11679 6420 11688
rect 6368 11645 6377 11679
rect 6377 11645 6411 11679
rect 6411 11645 6420 11679
rect 6368 11636 6420 11645
rect 5448 11568 5500 11620
rect 5816 11568 5868 11620
rect 5908 11568 5960 11620
rect 6276 11568 6328 11620
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 7748 11636 7800 11688
rect 6828 11568 6880 11620
rect 6920 11568 6972 11620
rect 7104 11568 7156 11620
rect 2136 11500 2188 11552
rect 3148 11500 3200 11552
rect 3240 11500 3292 11552
rect 5632 11500 5684 11552
rect 11428 11636 11480 11688
rect 10232 11500 10284 11552
rect 12716 11500 12768 11552
rect 13820 11500 13872 11552
rect 14832 11704 14884 11756
rect 15476 11704 15528 11756
rect 18788 11840 18840 11892
rect 20536 11840 20588 11892
rect 16672 11704 16724 11756
rect 19800 11772 19852 11824
rect 16856 11704 16908 11756
rect 17500 11704 17552 11756
rect 15108 11679 15160 11688
rect 15108 11645 15117 11679
rect 15117 11645 15151 11679
rect 15151 11645 15160 11679
rect 15108 11636 15160 11645
rect 18236 11747 18288 11756
rect 18236 11713 18245 11747
rect 18245 11713 18279 11747
rect 18279 11713 18288 11747
rect 18236 11704 18288 11713
rect 18328 11747 18380 11756
rect 18328 11713 18337 11747
rect 18337 11713 18371 11747
rect 18371 11713 18380 11747
rect 18328 11704 18380 11713
rect 18512 11679 18564 11688
rect 18512 11645 18521 11679
rect 18521 11645 18555 11679
rect 18555 11645 18564 11679
rect 18512 11636 18564 11645
rect 14464 11500 14516 11552
rect 17500 11500 17552 11552
rect 18144 11543 18196 11552
rect 18144 11509 18153 11543
rect 18153 11509 18187 11543
rect 18187 11509 18196 11543
rect 18144 11500 18196 11509
rect 21272 11500 21324 11552
rect 20 11364 72 11416
rect 572 11364 624 11416
rect 3422 11398 3474 11450
rect 3486 11398 3538 11450
rect 3550 11398 3602 11450
rect 3614 11398 3666 11450
rect 3678 11398 3730 11450
rect 8367 11398 8419 11450
rect 8431 11398 8483 11450
rect 8495 11398 8547 11450
rect 8559 11398 8611 11450
rect 8623 11398 8675 11450
rect 13312 11398 13364 11450
rect 13376 11398 13428 11450
rect 13440 11398 13492 11450
rect 13504 11398 13556 11450
rect 13568 11398 13620 11450
rect 18257 11398 18309 11450
rect 18321 11398 18373 11450
rect 18385 11398 18437 11450
rect 18449 11398 18501 11450
rect 18513 11398 18565 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 480 11228 532 11280
rect 3240 11296 3292 11348
rect 4068 11296 4120 11348
rect 4528 11296 4580 11348
rect 4712 11296 4764 11348
rect 2136 11228 2188 11280
rect 3516 11228 3568 11280
rect 6644 11296 6696 11348
rect 9864 11296 9916 11348
rect 11336 11296 11388 11348
rect 12256 11296 12308 11348
rect 12440 11296 12492 11348
rect 13728 11296 13780 11348
rect 15292 11296 15344 11348
rect 2044 11160 2096 11212
rect 2320 11203 2372 11212
rect 2320 11169 2329 11203
rect 2329 11169 2363 11203
rect 2363 11169 2372 11203
rect 2320 11160 2372 11169
rect 3976 11203 4028 11212
rect 3976 11169 3985 11203
rect 3985 11169 4019 11203
rect 4019 11169 4028 11203
rect 3976 11160 4028 11169
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 4712 11203 4764 11212
rect 4712 11169 4721 11203
rect 4721 11169 4755 11203
rect 4755 11169 4764 11203
rect 4712 11160 4764 11169
rect 5172 11160 5224 11212
rect 2504 11092 2556 11144
rect 2964 11092 3016 11144
rect 3332 11092 3384 11144
rect 3608 11024 3660 11076
rect 2044 10999 2096 11008
rect 2044 10965 2053 10999
rect 2053 10965 2087 10999
rect 2087 10965 2096 10999
rect 2044 10956 2096 10965
rect 2136 10956 2188 11008
rect 2412 10956 2464 11008
rect 3240 10956 3292 11008
rect 6552 11228 6604 11280
rect 6920 11228 6972 11280
rect 7380 11228 7432 11280
rect 7472 11228 7524 11280
rect 4988 11135 5040 11144
rect 4988 11101 4997 11135
rect 4997 11101 5031 11135
rect 5031 11101 5040 11135
rect 4988 11092 5040 11101
rect 5558 11092 5610 11144
rect 4620 10956 4672 11008
rect 6644 11092 6696 11144
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 8116 11092 8168 11144
rect 10692 11228 10744 11280
rect 12072 11228 12124 11280
rect 9588 11160 9640 11212
rect 11520 11160 11572 11212
rect 13084 11228 13136 11280
rect 14096 11228 14148 11280
rect 14832 11228 14884 11280
rect 15016 11228 15068 11280
rect 17132 11339 17184 11348
rect 17132 11305 17141 11339
rect 17141 11305 17175 11339
rect 17175 11305 17184 11339
rect 17132 11296 17184 11305
rect 18052 11296 18104 11348
rect 18696 11339 18748 11348
rect 18696 11305 18705 11339
rect 18705 11305 18739 11339
rect 18739 11305 18748 11339
rect 18696 11296 18748 11305
rect 20076 11296 20128 11348
rect 18788 11228 18840 11280
rect 9220 11092 9272 11144
rect 9404 11092 9456 11144
rect 8392 11024 8444 11076
rect 11060 11092 11112 11144
rect 11336 11092 11388 11144
rect 11612 11092 11664 11144
rect 13912 11092 13964 11144
rect 14372 11135 14424 11144
rect 5816 10956 5868 11008
rect 5908 10956 5960 11008
rect 6000 10956 6052 11008
rect 6368 10956 6420 11008
rect 8024 10956 8076 11008
rect 8300 10956 8352 11008
rect 9404 10956 9456 11008
rect 9496 10999 9548 11008
rect 9496 10965 9505 10999
rect 9505 10965 9539 10999
rect 9539 10965 9548 10999
rect 9496 10956 9548 10965
rect 10232 11024 10284 11076
rect 10508 11024 10560 11076
rect 14372 11101 14379 11135
rect 14379 11101 14413 11135
rect 14413 11101 14424 11135
rect 14372 11092 14424 11101
rect 15660 11092 15712 11144
rect 16764 11092 16816 11144
rect 17500 11092 17552 11144
rect 19156 11160 19208 11212
rect 11796 10956 11848 11008
rect 12256 10956 12308 11008
rect 12992 10956 13044 11008
rect 15568 11024 15620 11076
rect 16120 11024 16172 11076
rect 13912 10956 13964 11008
rect 14924 10956 14976 11008
rect 15108 10956 15160 11008
rect 16212 10956 16264 11008
rect 17224 11024 17276 11076
rect 17408 11024 17460 11076
rect 18880 11135 18932 11144
rect 18880 11101 18889 11135
rect 18889 11101 18923 11135
rect 18923 11101 18932 11135
rect 18880 11092 18932 11101
rect 17776 11024 17828 11076
rect 18604 11024 18656 11076
rect 18788 11024 18840 11076
rect 19616 11024 19668 11076
rect 20076 11024 20128 11076
rect 17684 10956 17736 11008
rect 5894 10854 5946 10906
rect 5958 10854 6010 10906
rect 6022 10854 6074 10906
rect 6086 10854 6138 10906
rect 6150 10854 6202 10906
rect 10839 10854 10891 10906
rect 10903 10854 10955 10906
rect 10967 10854 11019 10906
rect 11031 10854 11083 10906
rect 11095 10854 11147 10906
rect 15784 10854 15836 10906
rect 15848 10854 15900 10906
rect 15912 10854 15964 10906
rect 15976 10854 16028 10906
rect 16040 10854 16092 10906
rect 20729 10854 20781 10906
rect 20793 10854 20845 10906
rect 20857 10854 20909 10906
rect 20921 10854 20973 10906
rect 20985 10854 21037 10906
rect 1032 10752 1084 10804
rect 1400 10752 1452 10804
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 20 10684 72 10736
rect 2504 10752 2556 10804
rect 4436 10752 4488 10804
rect 4988 10752 5040 10804
rect 5172 10752 5224 10804
rect 5264 10752 5316 10804
rect 6920 10752 6972 10804
rect 7012 10752 7064 10804
rect 8852 10752 8904 10804
rect 10048 10752 10100 10804
rect 10140 10752 10192 10804
rect 10416 10752 10468 10804
rect 10600 10752 10652 10804
rect 11152 10752 11204 10804
rect 12348 10752 12400 10804
rect 12532 10795 12584 10804
rect 12532 10761 12541 10795
rect 12541 10761 12575 10795
rect 12575 10761 12584 10795
rect 12532 10752 12584 10761
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 2228 10684 2280 10736
rect 2872 10684 2924 10736
rect 4252 10684 4304 10736
rect 4344 10684 4396 10736
rect 4896 10684 4948 10736
rect 2780 10616 2832 10668
rect 3148 10616 3200 10668
rect 6000 10684 6052 10736
rect 3516 10591 3568 10600
rect 3516 10557 3525 10591
rect 3525 10557 3559 10591
rect 3559 10557 3568 10591
rect 3516 10548 3568 10557
rect 4804 10548 4856 10600
rect 3608 10412 3660 10464
rect 5908 10616 5960 10668
rect 5816 10548 5868 10600
rect 6368 10616 6420 10668
rect 6644 10616 6696 10668
rect 6184 10548 6236 10600
rect 8116 10684 8168 10736
rect 8392 10689 8444 10736
rect 7472 10616 7524 10668
rect 8392 10684 8417 10689
rect 8417 10684 8444 10689
rect 9312 10684 9364 10736
rect 14924 10752 14976 10804
rect 16304 10752 16356 10804
rect 16396 10752 16448 10804
rect 13176 10684 13228 10736
rect 15384 10684 15436 10736
rect 15936 10684 15988 10736
rect 8024 10548 8076 10600
rect 9864 10616 9916 10668
rect 12440 10616 12492 10668
rect 5172 10412 5224 10464
rect 6000 10412 6052 10464
rect 7472 10412 7524 10464
rect 9312 10548 9364 10600
rect 8576 10412 8628 10464
rect 11520 10591 11572 10600
rect 11520 10557 11529 10591
rect 11529 10557 11563 10591
rect 11563 10557 11572 10591
rect 11520 10548 11572 10557
rect 12900 10548 12952 10600
rect 13176 10591 13228 10600
rect 13176 10557 13185 10591
rect 13185 10557 13219 10591
rect 13219 10557 13228 10591
rect 13176 10548 13228 10557
rect 10324 10480 10376 10532
rect 10968 10480 11020 10532
rect 9772 10412 9824 10464
rect 13912 10659 13964 10668
rect 13912 10625 13921 10659
rect 13921 10625 13955 10659
rect 13955 10625 13964 10659
rect 13912 10616 13964 10625
rect 14004 10659 14056 10668
rect 14004 10625 14038 10659
rect 14038 10625 14056 10659
rect 14004 10616 14056 10625
rect 15108 10616 15160 10668
rect 15200 10635 15207 10668
rect 15207 10635 15241 10668
rect 15241 10635 15252 10668
rect 15200 10616 15252 10635
rect 16120 10616 16172 10668
rect 18880 10752 18932 10804
rect 16580 10616 16632 10668
rect 17132 10684 17184 10736
rect 19248 10684 19300 10736
rect 17040 10616 17092 10668
rect 18696 10616 18748 10668
rect 20260 10659 20312 10668
rect 20260 10625 20269 10659
rect 20269 10625 20303 10659
rect 20303 10625 20312 10659
rect 20260 10616 20312 10625
rect 13728 10548 13780 10600
rect 16028 10548 16080 10600
rect 14832 10412 14884 10464
rect 15844 10480 15896 10532
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 17408 10480 17460 10532
rect 19616 10591 19668 10600
rect 19616 10557 19625 10591
rect 19625 10557 19659 10591
rect 19659 10557 19668 10591
rect 19616 10548 19668 10557
rect 19800 10480 19852 10532
rect 17776 10412 17828 10464
rect 3422 10310 3474 10362
rect 3486 10310 3538 10362
rect 3550 10310 3602 10362
rect 3614 10310 3666 10362
rect 3678 10310 3730 10362
rect 8367 10310 8419 10362
rect 8431 10310 8483 10362
rect 8495 10310 8547 10362
rect 8559 10310 8611 10362
rect 8623 10310 8675 10362
rect 13312 10310 13364 10362
rect 13376 10310 13428 10362
rect 13440 10310 13492 10362
rect 13504 10310 13556 10362
rect 13568 10310 13620 10362
rect 18257 10310 18309 10362
rect 18321 10310 18373 10362
rect 18385 10310 18437 10362
rect 18449 10310 18501 10362
rect 18513 10310 18565 10362
rect 1492 10208 1544 10260
rect 3332 10208 3384 10260
rect 3424 10208 3476 10260
rect 3056 10140 3108 10192
rect 4160 10251 4212 10260
rect 4160 10217 4169 10251
rect 4169 10217 4203 10251
rect 4203 10217 4212 10251
rect 4160 10208 4212 10217
rect 4712 10208 4764 10260
rect 4804 10208 4856 10260
rect 1492 10072 1544 10124
rect 2964 10072 3016 10124
rect 3516 10072 3568 10124
rect 1308 10004 1360 10056
rect 2872 10004 2924 10056
rect 3884 10072 3936 10124
rect 5448 10140 5500 10192
rect 2596 9936 2648 9988
rect 4436 10004 4488 10056
rect 4620 10004 4672 10056
rect 5080 10004 5132 10056
rect 6828 10208 6880 10260
rect 6000 10072 6052 10124
rect 7196 10208 7248 10260
rect 7288 10140 7340 10192
rect 5632 10004 5684 10056
rect 7012 10004 7064 10056
rect 2228 9868 2280 9920
rect 2872 9911 2924 9920
rect 2872 9877 2881 9911
rect 2881 9877 2915 9911
rect 2915 9877 2924 9911
rect 2872 9868 2924 9877
rect 2964 9868 3016 9920
rect 4068 9868 4120 9920
rect 7196 9936 7248 9988
rect 4344 9911 4396 9920
rect 4344 9877 4353 9911
rect 4353 9877 4387 9911
rect 4387 9877 4396 9911
rect 4344 9868 4396 9877
rect 4620 9868 4672 9920
rect 5080 9868 5132 9920
rect 5448 9868 5500 9920
rect 6184 9868 6236 9920
rect 6736 9868 6788 9920
rect 9312 10208 9364 10260
rect 9772 10208 9824 10260
rect 9404 10140 9456 10192
rect 8208 10072 8260 10124
rect 8760 10072 8812 10124
rect 9588 10115 9640 10124
rect 9588 10081 9597 10115
rect 9597 10081 9631 10115
rect 9631 10081 9640 10115
rect 9588 10072 9640 10081
rect 7564 9868 7616 9920
rect 8116 10004 8168 10056
rect 9956 10072 10008 10124
rect 12624 10208 12676 10260
rect 13912 10208 13964 10260
rect 14464 10208 14516 10260
rect 14556 10140 14608 10192
rect 15844 10208 15896 10260
rect 10508 10115 10560 10124
rect 10508 10081 10517 10115
rect 10517 10081 10551 10115
rect 10551 10081 10560 10115
rect 10508 10072 10560 10081
rect 10600 10115 10652 10124
rect 10600 10081 10634 10115
rect 10634 10081 10652 10115
rect 10600 10072 10652 10081
rect 10968 10072 11020 10124
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 12900 10072 12952 10124
rect 13176 10072 13228 10124
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 15108 10115 15160 10124
rect 15108 10081 15142 10115
rect 15142 10081 15160 10115
rect 15108 10072 15160 10081
rect 16764 10140 16816 10192
rect 18696 10208 18748 10260
rect 18788 10251 18840 10260
rect 18788 10217 18797 10251
rect 18797 10217 18831 10251
rect 18831 10217 18840 10251
rect 18788 10208 18840 10217
rect 18880 10208 18932 10260
rect 17224 10072 17276 10124
rect 17408 10115 17460 10124
rect 17408 10081 17417 10115
rect 17417 10081 17451 10115
rect 17451 10081 17460 10115
rect 17408 10072 17460 10081
rect 18788 10072 18840 10124
rect 19156 10072 19208 10124
rect 8300 10004 8352 10056
rect 8576 10004 8628 10056
rect 9680 10004 9732 10056
rect 9772 10047 9824 10056
rect 9772 10013 9781 10047
rect 9781 10013 9815 10047
rect 9815 10013 9824 10047
rect 9772 10004 9824 10013
rect 10784 10047 10836 10056
rect 10784 10013 10793 10047
rect 10793 10013 10827 10047
rect 10827 10013 10836 10047
rect 10784 10004 10836 10013
rect 11796 10047 11848 10056
rect 11796 10013 11803 10047
rect 11803 10013 11837 10047
rect 11837 10013 11848 10047
rect 11796 10004 11848 10013
rect 12348 10004 12400 10056
rect 14004 10004 14056 10056
rect 14188 10004 14240 10056
rect 8392 9868 8444 9920
rect 9404 9868 9456 9920
rect 12532 9936 12584 9988
rect 14464 10004 14516 10056
rect 15936 10004 15988 10056
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17736 10047
rect 17684 10004 17736 10013
rect 17776 10004 17828 10056
rect 18144 10004 18196 10056
rect 9772 9868 9824 9920
rect 10048 9868 10100 9920
rect 16120 9868 16172 9920
rect 19708 9936 19760 9988
rect 16396 9868 16448 9920
rect 5894 9766 5946 9818
rect 5958 9766 6010 9818
rect 6022 9766 6074 9818
rect 6086 9766 6138 9818
rect 6150 9766 6202 9818
rect 10839 9766 10891 9818
rect 10903 9766 10955 9818
rect 10967 9766 11019 9818
rect 11031 9766 11083 9818
rect 11095 9766 11147 9818
rect 15784 9766 15836 9818
rect 15848 9766 15900 9818
rect 15912 9766 15964 9818
rect 15976 9766 16028 9818
rect 16040 9766 16092 9818
rect 20729 9766 20781 9818
rect 20793 9766 20845 9818
rect 20857 9766 20909 9818
rect 20921 9766 20973 9818
rect 20985 9766 21037 9818
rect 1768 9707 1820 9716
rect 1768 9673 1777 9707
rect 1777 9673 1811 9707
rect 1811 9673 1820 9707
rect 1768 9664 1820 9673
rect 2412 9596 2464 9648
rect 112 9528 164 9580
rect 2780 9664 2832 9716
rect 3240 9664 3292 9716
rect 3332 9664 3384 9716
rect 5356 9664 5408 9716
rect 6552 9664 6604 9716
rect 6828 9664 6880 9716
rect 7748 9707 7800 9716
rect 7748 9673 7757 9707
rect 7757 9673 7791 9707
rect 7791 9673 7800 9707
rect 7748 9664 7800 9673
rect 4160 9596 4212 9648
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 3516 9528 3568 9580
rect 2780 9460 2832 9512
rect 4160 9460 4212 9512
rect 4712 9460 4764 9512
rect 4896 9460 4948 9512
rect 5264 9537 5291 9546
rect 5291 9537 5316 9546
rect 5264 9494 5316 9537
rect 5448 9518 5500 9570
rect 6368 9528 6420 9580
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 7288 9596 7340 9648
rect 5540 9503 5592 9512
rect 5540 9469 5549 9503
rect 5549 9469 5583 9503
rect 5583 9469 5592 9503
rect 5540 9460 5592 9469
rect 5908 9460 5960 9512
rect 7748 9528 7800 9580
rect 8392 9664 8444 9716
rect 9312 9596 9364 9648
rect 8484 9528 8536 9580
rect 9588 9596 9640 9648
rect 10416 9571 10468 9580
rect 10416 9537 10425 9571
rect 10425 9537 10459 9571
rect 10459 9537 10468 9571
rect 10416 9528 10468 9537
rect 10600 9528 10652 9580
rect 11704 9664 11756 9716
rect 12348 9664 12400 9716
rect 14924 9528 14976 9580
rect 15660 9528 15712 9580
rect 16028 9528 16080 9580
rect 16304 9664 16356 9716
rect 3056 9435 3108 9444
rect 3056 9401 3065 9435
rect 3065 9401 3099 9435
rect 3099 9401 3108 9435
rect 3056 9392 3108 9401
rect 4988 9435 5040 9444
rect 4988 9401 4997 9435
rect 4997 9401 5031 9435
rect 5031 9401 5040 9435
rect 4988 9392 5040 9401
rect 4620 9324 4672 9376
rect 4896 9324 4948 9376
rect 6276 9324 6328 9376
rect 6736 9324 6788 9376
rect 7840 9324 7892 9376
rect 9404 9460 9456 9512
rect 9772 9460 9824 9512
rect 9312 9392 9364 9444
rect 8392 9324 8444 9376
rect 11520 9460 11572 9512
rect 12624 9460 12676 9512
rect 13176 9460 13228 9512
rect 11336 9367 11388 9376
rect 11336 9333 11345 9367
rect 11345 9333 11379 9367
rect 11379 9333 11388 9367
rect 11336 9324 11388 9333
rect 11796 9324 11848 9376
rect 13912 9392 13964 9444
rect 14188 9460 14240 9512
rect 14556 9460 14608 9512
rect 16120 9460 16172 9512
rect 16304 9571 16356 9580
rect 16304 9537 16313 9571
rect 16313 9537 16347 9571
rect 16347 9537 16356 9571
rect 16304 9528 16356 9537
rect 17224 9664 17276 9716
rect 18604 9664 18656 9716
rect 18880 9664 18932 9716
rect 19064 9664 19116 9716
rect 16672 9596 16724 9648
rect 17868 9596 17920 9648
rect 19524 9596 19576 9648
rect 16672 9503 16724 9512
rect 16672 9469 16681 9503
rect 16681 9469 16715 9503
rect 16715 9469 16724 9503
rect 16672 9460 16724 9469
rect 14280 9392 14332 9444
rect 14464 9435 14516 9444
rect 14464 9401 14473 9435
rect 14473 9401 14507 9435
rect 14507 9401 14516 9435
rect 14464 9392 14516 9401
rect 18512 9528 18564 9580
rect 19062 9571 19114 9580
rect 19062 9537 19073 9571
rect 19073 9537 19114 9571
rect 19062 9528 19114 9537
rect 21916 9528 21968 9580
rect 18696 9460 18748 9512
rect 18788 9503 18840 9512
rect 18788 9469 18797 9503
rect 18797 9469 18831 9503
rect 18831 9469 18840 9503
rect 18788 9460 18840 9469
rect 12716 9367 12768 9376
rect 12716 9333 12725 9367
rect 12725 9333 12759 9367
rect 12759 9333 12768 9367
rect 12716 9324 12768 9333
rect 12808 9324 12860 9376
rect 15476 9324 15528 9376
rect 16580 9324 16632 9376
rect 19524 9392 19576 9444
rect 18144 9324 18196 9376
rect 20076 9324 20128 9376
rect 3422 9222 3474 9274
rect 3486 9222 3538 9274
rect 3550 9222 3602 9274
rect 3614 9222 3666 9274
rect 3678 9222 3730 9274
rect 8367 9222 8419 9274
rect 8431 9222 8483 9274
rect 8495 9222 8547 9274
rect 8559 9222 8611 9274
rect 8623 9222 8675 9274
rect 13312 9222 13364 9274
rect 13376 9222 13428 9274
rect 13440 9222 13492 9274
rect 13504 9222 13556 9274
rect 13568 9222 13620 9274
rect 18257 9222 18309 9274
rect 18321 9222 18373 9274
rect 18385 9222 18437 9274
rect 18449 9222 18501 9274
rect 18513 9222 18565 9274
rect 1768 9163 1820 9172
rect 1768 9129 1777 9163
rect 1777 9129 1811 9163
rect 1811 9129 1820 9163
rect 1768 9120 1820 9129
rect 2320 9120 2372 9172
rect 4252 9120 4304 9172
rect 5172 9120 5224 9172
rect 5558 9120 5610 9172
rect 6368 9120 6420 9172
rect 6552 9120 6604 9172
rect 12532 9120 12584 9172
rect 13728 9120 13780 9172
rect 14464 9120 14516 9172
rect 2044 8916 2096 8968
rect 2228 8916 2280 8968
rect 3148 8916 3200 8968
rect 3516 8984 3568 9036
rect 6920 9095 6972 9104
rect 6920 9061 6929 9095
rect 6929 9061 6963 9095
rect 6963 9061 6972 9095
rect 6920 9052 6972 9061
rect 9956 9052 10008 9104
rect 10140 9052 10192 9104
rect 4344 8916 4396 8968
rect 4252 8848 4304 8900
rect 5080 8916 5132 8968
rect 6092 8984 6144 9036
rect 6552 8984 6604 9036
rect 5816 8916 5868 8968
rect 6368 8916 6420 8968
rect 7214 8959 7266 8968
rect 6000 8848 6052 8900
rect 7214 8925 7239 8959
rect 7239 8925 7266 8959
rect 7214 8916 7266 8925
rect 8208 8984 8260 9036
rect 9680 8984 9732 9036
rect 9772 8984 9824 9036
rect 12716 9052 12768 9104
rect 14832 9052 14884 9104
rect 15384 9052 15436 9104
rect 10600 8984 10652 9036
rect 10784 8984 10836 9036
rect 11428 8984 11480 9036
rect 11980 9027 12032 9036
rect 11980 8993 11989 9027
rect 11989 8993 12023 9027
rect 12023 8993 12032 9027
rect 11980 8984 12032 8993
rect 8484 8916 8536 8968
rect 2504 8780 2556 8832
rect 3148 8780 3200 8832
rect 3700 8780 3752 8832
rect 5264 8780 5316 8832
rect 6920 8780 6972 8832
rect 7380 8780 7432 8832
rect 9404 8848 9456 8900
rect 9864 8848 9916 8900
rect 10416 8916 10468 8968
rect 10968 8959 11020 8968
rect 10968 8925 10977 8959
rect 10977 8925 11011 8959
rect 11011 8925 11020 8959
rect 10968 8916 11020 8925
rect 11244 8959 11296 8968
rect 11244 8925 11253 8959
rect 11253 8925 11287 8959
rect 11287 8925 11296 8959
rect 11244 8916 11296 8925
rect 11888 8916 11940 8968
rect 12256 8984 12308 9036
rect 12900 9027 12952 9036
rect 12900 8993 12909 9027
rect 12909 8993 12943 9027
rect 12943 8993 12952 9027
rect 12900 8984 12952 8993
rect 15568 9120 15620 9172
rect 16212 9120 16264 9172
rect 17132 9120 17184 9172
rect 12992 8959 13044 8968
rect 12992 8925 13026 8959
rect 13026 8925 13044 8959
rect 12992 8916 13044 8925
rect 13176 8959 13228 8968
rect 13176 8925 13185 8959
rect 13185 8925 13219 8959
rect 13219 8925 13228 8959
rect 13176 8916 13228 8925
rect 14372 8959 14424 8968
rect 13728 8848 13780 8900
rect 14372 8925 14379 8959
rect 14379 8925 14413 8959
rect 14413 8925 14424 8959
rect 14372 8916 14424 8925
rect 15200 8916 15252 8968
rect 8392 8780 8444 8832
rect 9588 8780 9640 8832
rect 10416 8780 10468 8832
rect 10876 8780 10928 8832
rect 10968 8780 11020 8832
rect 12624 8780 12676 8832
rect 13268 8780 13320 8832
rect 13912 8780 13964 8832
rect 16120 8916 16172 8968
rect 16396 8916 16448 8968
rect 16580 8916 16632 8968
rect 15936 8848 15988 8900
rect 17960 8916 18012 8968
rect 18052 8916 18104 8968
rect 18788 8916 18840 8968
rect 17316 8848 17368 8900
rect 17776 8848 17828 8900
rect 16028 8780 16080 8832
rect 18328 8848 18380 8900
rect 18696 8891 18748 8900
rect 18696 8857 18705 8891
rect 18705 8857 18739 8891
rect 18739 8857 18748 8891
rect 18696 8848 18748 8857
rect 18512 8780 18564 8832
rect 20352 9120 20404 9172
rect 20076 9052 20128 9104
rect 19248 9027 19300 9036
rect 19248 8993 19257 9027
rect 19257 8993 19291 9027
rect 19291 8993 19300 9027
rect 19248 8984 19300 8993
rect 19524 8959 19576 8968
rect 19524 8925 19531 8959
rect 19531 8925 19565 8959
rect 19565 8925 19576 8959
rect 19524 8916 19576 8925
rect 19616 8780 19668 8832
rect 5894 8678 5946 8730
rect 5958 8678 6010 8730
rect 6022 8678 6074 8730
rect 6086 8678 6138 8730
rect 6150 8678 6202 8730
rect 10839 8678 10891 8730
rect 10903 8678 10955 8730
rect 10967 8678 11019 8730
rect 11031 8678 11083 8730
rect 11095 8678 11147 8730
rect 15784 8678 15836 8730
rect 15848 8678 15900 8730
rect 15912 8678 15964 8730
rect 15976 8678 16028 8730
rect 16040 8678 16092 8730
rect 20729 8678 20781 8730
rect 20793 8678 20845 8730
rect 20857 8678 20909 8730
rect 20921 8678 20973 8730
rect 20985 8678 21037 8730
rect 1492 8576 1544 8628
rect 1860 8576 1912 8628
rect 2964 8576 3016 8628
rect 3148 8576 3200 8628
rect 4712 8576 4764 8628
rect 4988 8576 5040 8628
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 2504 8508 2556 8560
rect 3424 8483 3476 8492
rect 3424 8449 3433 8483
rect 3433 8449 3467 8483
rect 3467 8449 3476 8483
rect 3424 8440 3476 8449
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 1860 8372 1912 8424
rect 2872 8372 2924 8424
rect 4068 8372 4120 8424
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 5724 8440 5776 8492
rect 5908 8440 5960 8492
rect 8760 8576 8812 8628
rect 9404 8576 9456 8628
rect 9496 8576 9548 8628
rect 6092 8508 6144 8560
rect 7748 8508 7800 8560
rect 7840 8508 7892 8560
rect 8300 8551 8352 8560
rect 8300 8517 8331 8551
rect 8331 8517 8352 8551
rect 8300 8508 8352 8517
rect 8484 8508 8536 8560
rect 8576 8440 8628 8492
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 10416 8576 10468 8628
rect 10692 8576 10744 8628
rect 11060 8576 11112 8628
rect 15108 8576 15160 8628
rect 10324 8508 10376 8560
rect 11428 8508 11480 8560
rect 15476 8576 15528 8628
rect 16212 8576 16264 8628
rect 16672 8576 16724 8628
rect 12072 8440 12124 8492
rect 12164 8440 12216 8492
rect 12624 8440 12676 8492
rect 13544 8440 13596 8492
rect 572 8304 624 8356
rect 1032 8236 1084 8288
rect 2504 8236 2556 8288
rect 2872 8236 2924 8288
rect 6184 8372 6236 8424
rect 4344 8279 4396 8288
rect 4344 8245 4353 8279
rect 4353 8245 4387 8279
rect 4387 8245 4396 8279
rect 4344 8236 4396 8245
rect 4528 8236 4580 8288
rect 9312 8372 9364 8424
rect 5172 8236 5224 8288
rect 7748 8236 7800 8288
rect 9588 8279 9640 8288
rect 9588 8245 9597 8279
rect 9597 8245 9631 8279
rect 9631 8245 9640 8279
rect 9588 8236 9640 8245
rect 9772 8236 9824 8288
rect 10692 8372 10744 8424
rect 11612 8372 11664 8424
rect 11152 8304 11204 8356
rect 11888 8304 11940 8356
rect 12072 8304 12124 8356
rect 12992 8372 13044 8424
rect 13176 8372 13228 8424
rect 13820 8440 13872 8492
rect 14372 8440 14424 8492
rect 15200 8440 15252 8492
rect 13636 8304 13688 8356
rect 13452 8236 13504 8288
rect 15476 8440 15528 8492
rect 15844 8508 15896 8560
rect 16120 8508 16172 8560
rect 17224 8576 17276 8628
rect 17408 8576 17460 8628
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 16764 8440 16816 8492
rect 17592 8508 17644 8560
rect 17868 8508 17920 8560
rect 19432 8551 19484 8560
rect 15844 8372 15896 8424
rect 17132 8372 17184 8424
rect 17408 8372 17460 8424
rect 17776 8483 17828 8492
rect 17776 8449 17785 8483
rect 17785 8449 17819 8483
rect 17819 8449 17828 8483
rect 17776 8440 17828 8449
rect 18604 8440 18656 8492
rect 19432 8517 19466 8551
rect 19466 8517 19484 8551
rect 19432 8508 19484 8517
rect 19708 8508 19760 8560
rect 18512 8372 18564 8424
rect 15660 8236 15712 8288
rect 17132 8236 17184 8288
rect 17408 8236 17460 8288
rect 17684 8236 17736 8288
rect 18788 8347 18840 8356
rect 18788 8313 18797 8347
rect 18797 8313 18831 8347
rect 18831 8313 18840 8347
rect 18788 8304 18840 8313
rect 18144 8236 18196 8288
rect 19524 8236 19576 8288
rect 3422 8134 3474 8186
rect 3486 8134 3538 8186
rect 3550 8134 3602 8186
rect 3614 8134 3666 8186
rect 3678 8134 3730 8186
rect 8367 8134 8419 8186
rect 8431 8134 8483 8186
rect 8495 8134 8547 8186
rect 8559 8134 8611 8186
rect 8623 8134 8675 8186
rect 13312 8134 13364 8186
rect 13376 8134 13428 8186
rect 13440 8134 13492 8186
rect 13504 8134 13556 8186
rect 13568 8134 13620 8186
rect 18257 8134 18309 8186
rect 18321 8134 18373 8186
rect 18385 8134 18437 8186
rect 18449 8134 18501 8186
rect 18513 8134 18565 8186
rect 1952 8032 2004 8084
rect 1400 7896 1452 7948
rect 2044 7828 2096 7880
rect 4160 8032 4212 8084
rect 5172 8032 5224 8084
rect 3516 7964 3568 8016
rect 3884 7964 3936 8016
rect 4252 7896 4304 7948
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 6184 8032 6236 8084
rect 6552 8032 6604 8084
rect 5816 7896 5868 7948
rect 6092 7939 6144 7948
rect 6092 7905 6101 7939
rect 6101 7905 6135 7939
rect 6135 7905 6144 7939
rect 6092 7896 6144 7905
rect 8300 8032 8352 8084
rect 9220 8032 9272 8084
rect 9680 8032 9732 8084
rect 9956 8032 10008 8084
rect 10784 8032 10836 8084
rect 11244 8032 11296 8084
rect 13912 8032 13964 8084
rect 1400 7760 1452 7812
rect 1860 7760 1912 7812
rect 3240 7828 3292 7880
rect 3516 7760 3568 7812
rect 4896 7828 4948 7880
rect 5540 7828 5592 7880
rect 5632 7828 5684 7880
rect 2872 7692 2924 7744
rect 3332 7692 3384 7744
rect 4068 7692 4120 7744
rect 4896 7692 4948 7744
rect 6000 7760 6052 7812
rect 7012 7828 7064 7880
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7800 7871
rect 7748 7828 7800 7837
rect 8116 7862 8168 7914
rect 9772 7896 9824 7948
rect 11520 7896 11572 7948
rect 11888 7896 11940 7948
rect 12440 7896 12492 7948
rect 12716 8007 12768 8016
rect 12716 7973 12725 8007
rect 12725 7973 12759 8007
rect 12759 7973 12768 8007
rect 12716 7964 12768 7973
rect 15844 8032 15896 8084
rect 16120 8032 16172 8084
rect 16672 8032 16724 8084
rect 16764 8032 16816 8084
rect 12808 7896 12860 7948
rect 13820 7896 13872 7948
rect 8300 7828 8352 7880
rect 9312 7828 9364 7880
rect 7840 7760 7892 7812
rect 7932 7760 7984 7812
rect 8116 7760 8168 7812
rect 10692 7828 10744 7880
rect 12164 7828 12216 7880
rect 5908 7692 5960 7744
rect 7012 7692 7064 7744
rect 7472 7692 7524 7744
rect 7656 7692 7708 7744
rect 9680 7760 9732 7812
rect 9220 7692 9272 7744
rect 11796 7760 11848 7812
rect 12992 7871 13044 7880
rect 12992 7837 13001 7871
rect 13001 7837 13035 7871
rect 13035 7837 13044 7871
rect 12992 7828 13044 7837
rect 14740 7828 14792 7880
rect 15016 7896 15068 7948
rect 15476 7871 15528 7880
rect 15476 7837 15485 7871
rect 15485 7837 15519 7871
rect 15519 7837 15528 7871
rect 15476 7828 15528 7837
rect 15936 7828 15988 7880
rect 16488 7939 16540 7948
rect 16488 7905 16497 7939
rect 16497 7905 16531 7939
rect 16531 7905 16540 7939
rect 16488 7896 16540 7905
rect 18880 8007 18932 8016
rect 18880 7973 18889 8007
rect 18889 7973 18923 8007
rect 18923 7973 18932 8007
rect 18880 7964 18932 7973
rect 19892 7964 19944 8016
rect 17592 7896 17644 7948
rect 17684 7828 17736 7880
rect 18236 7828 18288 7880
rect 19524 7896 19576 7948
rect 19616 7871 19668 7880
rect 19616 7837 19625 7871
rect 19625 7837 19659 7871
rect 19659 7837 19668 7871
rect 19616 7828 19668 7837
rect 19892 7828 19944 7880
rect 11060 7692 11112 7744
rect 11980 7692 12032 7744
rect 14004 7692 14056 7744
rect 15660 7735 15712 7744
rect 15660 7701 15669 7735
rect 15669 7701 15703 7735
rect 15703 7701 15712 7735
rect 15660 7692 15712 7701
rect 15752 7692 15804 7744
rect 16304 7692 16356 7744
rect 16672 7692 16724 7744
rect 17776 7692 17828 7744
rect 18052 7692 18104 7744
rect 18788 7692 18840 7744
rect 19340 7692 19392 7744
rect 19616 7692 19668 7744
rect 296 7556 348 7608
rect 664 7556 716 7608
rect 5894 7590 5946 7642
rect 5958 7590 6010 7642
rect 6022 7590 6074 7642
rect 6086 7590 6138 7642
rect 6150 7590 6202 7642
rect 10839 7590 10891 7642
rect 10903 7590 10955 7642
rect 10967 7590 11019 7642
rect 11031 7590 11083 7642
rect 11095 7590 11147 7642
rect 15784 7590 15836 7642
rect 15848 7590 15900 7642
rect 15912 7590 15964 7642
rect 15976 7590 16028 7642
rect 16040 7590 16092 7642
rect 20729 7590 20781 7642
rect 20793 7590 20845 7642
rect 20857 7590 20909 7642
rect 20921 7590 20973 7642
rect 20985 7590 21037 7642
rect 21364 7624 21416 7676
rect 756 7488 808 7540
rect 1124 7488 1176 7540
rect 2596 7488 2648 7540
rect 3056 7488 3108 7540
rect 3148 7488 3200 7540
rect 4344 7488 4396 7540
rect 2228 7420 2280 7472
rect 4528 7420 4580 7472
rect 1860 7352 1912 7404
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4160 7352 4212 7404
rect 5264 7395 5316 7404
rect 5264 7361 5273 7395
rect 5273 7361 5307 7395
rect 5307 7361 5316 7395
rect 5264 7352 5316 7361
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 6184 7352 6236 7404
rect 6460 7352 6512 7404
rect 7012 7488 7064 7540
rect 7104 7352 7156 7404
rect 7840 7488 7892 7540
rect 8208 7420 8260 7472
rect 10600 7488 10652 7540
rect 12624 7488 12676 7540
rect 14004 7420 14056 7472
rect 14188 7420 14240 7472
rect 7840 7352 7892 7404
rect 1124 7284 1176 7336
rect 2872 7284 2924 7336
rect 3976 7284 4028 7336
rect 4252 7284 4304 7336
rect 4896 7284 4948 7336
rect 6092 7284 6144 7336
rect 7932 7284 7984 7336
rect 9036 7395 9088 7404
rect 9036 7361 9070 7395
rect 9070 7361 9088 7395
rect 9036 7352 9088 7361
rect 9220 7395 9272 7404
rect 9220 7361 9229 7395
rect 9229 7361 9263 7395
rect 9263 7361 9272 7395
rect 9220 7352 9272 7361
rect 11520 7352 11572 7404
rect 11704 7395 11756 7404
rect 11704 7361 11713 7395
rect 11713 7361 11747 7395
rect 11747 7361 11756 7395
rect 11704 7352 11756 7361
rect 11888 7352 11940 7404
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 12808 7395 12860 7404
rect 12808 7361 12842 7395
rect 12842 7361 12860 7395
rect 12808 7352 12860 7361
rect 12992 7395 13044 7404
rect 12992 7361 13001 7395
rect 13001 7361 13035 7395
rect 13035 7361 13044 7395
rect 12992 7352 13044 7361
rect 14556 7420 14608 7472
rect 14464 7352 14516 7404
rect 15752 7420 15804 7472
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 16212 7488 16264 7540
rect 16764 7420 16816 7472
rect 17132 7420 17184 7472
rect 17224 7420 17276 7472
rect 17684 7531 17736 7540
rect 17684 7497 17693 7531
rect 17693 7497 17727 7531
rect 17727 7497 17736 7531
rect 17684 7488 17736 7497
rect 19524 7488 19576 7540
rect 20260 7488 20312 7540
rect 20536 7488 20588 7540
rect 2780 7216 2832 7268
rect 4712 7216 4764 7268
rect 4988 7259 5040 7268
rect 4988 7225 4997 7259
rect 4997 7225 5031 7259
rect 5031 7225 5040 7259
rect 4988 7216 5040 7225
rect 7104 7216 7156 7268
rect 9772 7284 9824 7336
rect 10968 7284 11020 7336
rect 11612 7284 11664 7336
rect 1768 7148 1820 7200
rect 3700 7148 3752 7200
rect 3884 7148 3936 7200
rect 5264 7148 5316 7200
rect 5724 7148 5776 7200
rect 6368 7191 6420 7200
rect 6368 7157 6377 7191
rect 6377 7157 6411 7191
rect 6411 7157 6420 7191
rect 6368 7148 6420 7157
rect 8208 7148 8260 7200
rect 9036 7148 9088 7200
rect 11152 7216 11204 7268
rect 15476 7327 15528 7336
rect 12440 7259 12492 7268
rect 12440 7225 12449 7259
rect 12449 7225 12483 7259
rect 12483 7225 12492 7259
rect 12440 7216 12492 7225
rect 9864 7191 9916 7200
rect 9864 7157 9873 7191
rect 9873 7157 9907 7191
rect 9907 7157 9916 7191
rect 9864 7148 9916 7157
rect 10784 7148 10836 7200
rect 11520 7148 11572 7200
rect 11612 7148 11664 7200
rect 13636 7191 13688 7200
rect 13636 7157 13645 7191
rect 13645 7157 13679 7191
rect 13679 7157 13688 7191
rect 13636 7148 13688 7157
rect 13912 7259 13964 7268
rect 13912 7225 13921 7259
rect 13921 7225 13955 7259
rect 13955 7225 13964 7259
rect 13912 7216 13964 7225
rect 14004 7216 14056 7268
rect 15476 7293 15485 7327
rect 15485 7293 15519 7327
rect 15519 7293 15528 7327
rect 15476 7284 15528 7293
rect 16304 7395 16356 7404
rect 16304 7361 16313 7395
rect 16313 7361 16347 7395
rect 16347 7361 16356 7395
rect 16304 7352 16356 7361
rect 16856 7352 16908 7404
rect 16948 7395 17000 7404
rect 16948 7361 16955 7395
rect 16955 7361 16989 7395
rect 16989 7361 17000 7395
rect 16948 7352 17000 7361
rect 16488 7284 16540 7336
rect 16672 7327 16724 7336
rect 16672 7293 16681 7327
rect 16681 7293 16715 7327
rect 16715 7293 16724 7327
rect 16672 7284 16724 7293
rect 15384 7216 15436 7268
rect 15752 7216 15804 7268
rect 18052 7420 18104 7472
rect 17960 7352 18012 7404
rect 18236 7352 18288 7404
rect 18972 7352 19024 7404
rect 19708 7352 19760 7404
rect 19892 7420 19944 7472
rect 21456 7420 21508 7472
rect 18052 7216 18104 7268
rect 16212 7148 16264 7200
rect 16396 7148 16448 7200
rect 3422 7046 3474 7098
rect 3486 7046 3538 7098
rect 3550 7046 3602 7098
rect 3614 7046 3666 7098
rect 3678 7046 3730 7098
rect 8367 7046 8419 7098
rect 8431 7046 8483 7098
rect 8495 7046 8547 7098
rect 8559 7046 8611 7098
rect 8623 7046 8675 7098
rect 13312 7046 13364 7098
rect 13376 7046 13428 7098
rect 13440 7046 13492 7098
rect 13504 7046 13556 7098
rect 13568 7046 13620 7098
rect 18257 7046 18309 7098
rect 18321 7046 18373 7098
rect 18385 7046 18437 7098
rect 18449 7046 18501 7098
rect 18513 7046 18565 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 1584 6944 1636 6996
rect 2044 6944 2096 6996
rect 1124 6808 1176 6860
rect 2228 6808 2280 6860
rect 3056 6808 3108 6860
rect 5540 6944 5592 6996
rect 6920 6944 6972 6996
rect 6368 6876 6420 6928
rect 4344 6808 4396 6860
rect 5632 6808 5684 6860
rect 480 6740 532 6792
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2648 6783
rect 2596 6740 2648 6749
rect 1768 6604 1820 6656
rect 3056 6604 3108 6656
rect 3792 6604 3844 6656
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4896 6783 4948 6792
rect 4896 6749 4903 6783
rect 4903 6749 4937 6783
rect 4937 6749 4948 6783
rect 4896 6740 4948 6749
rect 5264 6740 5316 6792
rect 5816 6740 5868 6792
rect 6000 6740 6052 6792
rect 6184 6783 6236 6792
rect 6184 6749 6193 6783
rect 6193 6749 6227 6783
rect 6227 6749 6236 6783
rect 6184 6740 6236 6749
rect 6368 6740 6420 6792
rect 6828 6808 6880 6860
rect 6920 6851 6972 6860
rect 6920 6817 6929 6851
rect 6929 6817 6963 6851
rect 6963 6817 6972 6851
rect 6920 6808 6972 6817
rect 7840 6944 7892 6996
rect 9312 6944 9364 6996
rect 9404 6944 9456 6996
rect 7932 6876 7984 6928
rect 9772 6876 9824 6928
rect 8484 6808 8536 6860
rect 9956 6808 10008 6860
rect 10508 6808 10560 6860
rect 10692 6808 10744 6860
rect 11814 6876 11866 6928
rect 12164 6944 12216 6996
rect 12348 6944 12400 6996
rect 12992 6944 13044 6996
rect 14556 6944 14608 6996
rect 14648 6944 14700 6996
rect 13912 6876 13964 6928
rect 14096 6876 14148 6928
rect 7288 6783 7340 6792
rect 7288 6749 7322 6783
rect 7322 6749 7340 6783
rect 7288 6740 7340 6749
rect 7472 6783 7524 6792
rect 7472 6749 7481 6783
rect 7481 6749 7515 6783
rect 7515 6749 7524 6783
rect 7472 6740 7524 6749
rect 9220 6783 9272 6792
rect 9220 6749 9229 6783
rect 9229 6749 9263 6783
rect 9263 6749 9272 6783
rect 9220 6740 9272 6749
rect 11060 6783 11112 6792
rect 11060 6749 11069 6783
rect 11069 6749 11103 6783
rect 11103 6749 11112 6783
rect 11060 6740 11112 6749
rect 11152 6783 11204 6792
rect 11152 6749 11186 6783
rect 11186 6749 11204 6783
rect 11152 6740 11204 6749
rect 11336 6783 11388 6792
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 5264 6604 5316 6656
rect 5908 6604 5960 6656
rect 6460 6672 6512 6724
rect 9496 6672 9548 6724
rect 13360 6808 13412 6860
rect 15384 6808 15436 6860
rect 15660 6851 15712 6860
rect 15660 6817 15669 6851
rect 15669 6817 15703 6851
rect 15703 6817 15712 6851
rect 15660 6808 15712 6817
rect 16672 6808 16724 6860
rect 18604 6944 18656 6996
rect 19248 6944 19300 6996
rect 20076 6919 20128 6928
rect 20076 6885 20085 6919
rect 20085 6885 20119 6919
rect 20119 6885 20128 6919
rect 20076 6876 20128 6885
rect 12072 6783 12124 6792
rect 12072 6749 12081 6783
rect 12081 6749 12115 6783
rect 12115 6749 12124 6783
rect 12072 6740 12124 6749
rect 12716 6740 12768 6792
rect 13268 6740 13320 6792
rect 13636 6740 13688 6792
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14004 6740 14056 6792
rect 14924 6740 14976 6792
rect 15476 6740 15528 6792
rect 12624 6672 12676 6724
rect 17040 6740 17092 6792
rect 18052 6740 18104 6792
rect 18420 6740 18472 6792
rect 18604 6740 18656 6792
rect 18880 6740 18932 6792
rect 6828 6604 6880 6656
rect 9680 6604 9732 6656
rect 9864 6604 9916 6656
rect 10048 6604 10100 6656
rect 10508 6604 10560 6656
rect 14004 6604 14056 6656
rect 15200 6604 15252 6656
rect 15660 6604 15712 6656
rect 17776 6604 17828 6656
rect 18144 6647 18196 6656
rect 18144 6613 18153 6647
rect 18153 6613 18187 6647
rect 18187 6613 18196 6647
rect 18144 6604 18196 6613
rect 18604 6647 18656 6656
rect 18604 6613 18613 6647
rect 18613 6613 18647 6647
rect 18647 6613 18656 6647
rect 18604 6604 18656 6613
rect 18696 6604 18748 6656
rect 18880 6647 18932 6656
rect 18880 6613 18889 6647
rect 18889 6613 18923 6647
rect 18923 6613 18932 6647
rect 18880 6604 18932 6613
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 19892 6604 19944 6656
rect 20536 6604 20588 6656
rect 20996 6604 21048 6656
rect 5894 6502 5946 6554
rect 5958 6502 6010 6554
rect 6022 6502 6074 6554
rect 6086 6502 6138 6554
rect 6150 6502 6202 6554
rect 10839 6502 10891 6554
rect 10903 6502 10955 6554
rect 10967 6502 11019 6554
rect 11031 6502 11083 6554
rect 11095 6502 11147 6554
rect 15784 6502 15836 6554
rect 15848 6502 15900 6554
rect 15912 6502 15964 6554
rect 15976 6502 16028 6554
rect 16040 6502 16092 6554
rect 20729 6502 20781 6554
rect 20793 6502 20845 6554
rect 20857 6502 20909 6554
rect 20921 6502 20973 6554
rect 20985 6502 21037 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2320 6443 2372 6452
rect 2320 6409 2329 6443
rect 2329 6409 2363 6443
rect 2363 6409 2372 6443
rect 2320 6400 2372 6409
rect 2136 6332 2188 6384
rect 112 6264 164 6316
rect 2044 6307 2096 6316
rect 2044 6273 2053 6307
rect 2053 6273 2087 6307
rect 2087 6273 2096 6307
rect 2044 6264 2096 6273
rect 3884 6400 3936 6452
rect 4528 6400 4580 6452
rect 4988 6400 5040 6452
rect 5632 6400 5684 6452
rect 4344 6332 4396 6384
rect 3792 6307 3844 6316
rect 3792 6273 3801 6307
rect 3801 6273 3835 6307
rect 3835 6273 3844 6307
rect 3792 6264 3844 6273
rect 4712 6264 4764 6316
rect 5172 6264 5224 6316
rect 5632 6264 5684 6316
rect 5816 6264 5868 6316
rect 6092 6307 6144 6316
rect 6092 6273 6101 6307
rect 6101 6273 6135 6307
rect 6135 6273 6144 6307
rect 6092 6264 6144 6273
rect 2872 6196 2924 6248
rect 6276 6400 6328 6452
rect 8208 6443 8260 6452
rect 8208 6409 8217 6443
rect 8217 6409 8251 6443
rect 8251 6409 8260 6443
rect 8208 6400 8260 6409
rect 8484 6400 8536 6452
rect 7288 6332 7340 6384
rect 9220 6332 9272 6384
rect 9312 6332 9364 6384
rect 9864 6443 9916 6452
rect 9864 6409 9873 6443
rect 9873 6409 9907 6443
rect 9907 6409 9916 6443
rect 9864 6400 9916 6409
rect 10140 6400 10192 6452
rect 11796 6400 11848 6452
rect 12072 6400 12124 6452
rect 12348 6400 12400 6452
rect 12716 6400 12768 6452
rect 14464 6400 14516 6452
rect 14740 6400 14792 6452
rect 15752 6400 15804 6452
rect 15844 6443 15896 6452
rect 15844 6409 15853 6443
rect 15853 6409 15887 6443
rect 15887 6409 15896 6443
rect 15844 6400 15896 6409
rect 3056 6128 3108 6180
rect 3240 6171 3292 6180
rect 3240 6137 3249 6171
rect 3249 6137 3283 6171
rect 3283 6137 3292 6171
rect 3240 6128 3292 6137
rect 2596 6060 2648 6112
rect 3332 6060 3384 6112
rect 7104 6128 7156 6180
rect 5908 6103 5960 6112
rect 5908 6069 5917 6103
rect 5917 6069 5951 6103
rect 5951 6069 5960 6103
rect 5908 6060 5960 6069
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 9404 6196 9456 6248
rect 10232 6307 10284 6316
rect 10232 6273 10241 6307
rect 10241 6273 10275 6307
rect 10275 6273 10284 6307
rect 10232 6264 10284 6273
rect 11060 6307 11112 6316
rect 11060 6273 11069 6307
rect 11069 6273 11103 6307
rect 11103 6273 11112 6307
rect 11060 6264 11112 6273
rect 11152 6307 11204 6316
rect 11152 6273 11161 6307
rect 11161 6273 11195 6307
rect 11195 6273 11204 6307
rect 11152 6264 11204 6273
rect 11796 6307 11848 6316
rect 9956 6196 10008 6248
rect 11796 6273 11803 6307
rect 11803 6273 11837 6307
rect 11837 6273 11848 6307
rect 11796 6264 11848 6273
rect 11428 6196 11480 6248
rect 12348 6264 12400 6316
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13412 6307
rect 13360 6264 13412 6273
rect 13728 6332 13780 6384
rect 15108 6332 15160 6384
rect 14188 6264 14240 6316
rect 14740 6307 14792 6316
rect 14740 6273 14774 6307
rect 14774 6273 14792 6307
rect 14740 6264 14792 6273
rect 15200 6264 15252 6316
rect 12532 6128 12584 6180
rect 7564 6060 7616 6112
rect 10140 6060 10192 6112
rect 10600 6060 10652 6112
rect 12440 6060 12492 6112
rect 12624 6060 12676 6112
rect 12992 6060 13044 6112
rect 13751 6128 13803 6180
rect 15844 6264 15896 6316
rect 16028 6400 16080 6452
rect 16304 6400 16356 6452
rect 16028 6264 16080 6316
rect 16212 6264 16264 6316
rect 18052 6332 18104 6384
rect 18144 6332 18196 6384
rect 18236 6332 18288 6384
rect 18512 6332 18564 6384
rect 16580 6264 16632 6316
rect 16672 6264 16724 6316
rect 17132 6307 17184 6316
rect 17132 6273 17139 6307
rect 17139 6273 17173 6307
rect 17173 6273 17184 6307
rect 17132 6264 17184 6273
rect 17684 6264 17736 6316
rect 18696 6264 18748 6316
rect 16396 6239 16448 6248
rect 16396 6205 16405 6239
rect 16405 6205 16439 6239
rect 16439 6205 16448 6239
rect 16396 6196 16448 6205
rect 16764 6128 16816 6180
rect 14004 6060 14056 6112
rect 14464 6060 14516 6112
rect 15384 6060 15436 6112
rect 15568 6060 15620 6112
rect 16580 6060 16632 6112
rect 17868 6196 17920 6248
rect 18144 6196 18196 6248
rect 19616 6400 19668 6452
rect 19708 6264 19760 6316
rect 20352 6307 20404 6316
rect 20352 6273 20361 6307
rect 20361 6273 20395 6307
rect 20395 6273 20404 6307
rect 20352 6264 20404 6273
rect 17684 6128 17736 6180
rect 18880 6239 18932 6248
rect 18880 6205 18889 6239
rect 18889 6205 18923 6239
rect 18923 6205 18932 6239
rect 18880 6196 18932 6205
rect 18420 6171 18472 6180
rect 18420 6137 18429 6171
rect 18429 6137 18463 6171
rect 18463 6137 18472 6171
rect 18420 6128 18472 6137
rect 19892 6060 19944 6112
rect 20444 6103 20496 6112
rect 20444 6069 20453 6103
rect 20453 6069 20487 6103
rect 20487 6069 20496 6103
rect 20444 6060 20496 6069
rect 3422 5958 3474 6010
rect 3486 5958 3538 6010
rect 3550 5958 3602 6010
rect 3614 5958 3666 6010
rect 3678 5958 3730 6010
rect 8367 5958 8419 6010
rect 8431 5958 8483 6010
rect 8495 5958 8547 6010
rect 8559 5958 8611 6010
rect 8623 5958 8675 6010
rect 13312 5958 13364 6010
rect 13376 5958 13428 6010
rect 13440 5958 13492 6010
rect 13504 5958 13556 6010
rect 13568 5958 13620 6010
rect 18257 5958 18309 6010
rect 18321 5958 18373 6010
rect 18385 5958 18437 6010
rect 18449 5958 18501 6010
rect 18513 5958 18565 6010
rect 1124 5720 1176 5772
rect 2780 5856 2832 5908
rect 3240 5856 3292 5908
rect 3976 5899 4028 5908
rect 3976 5865 3985 5899
rect 3985 5865 4019 5899
rect 4019 5865 4028 5899
rect 3976 5856 4028 5865
rect 1676 5584 1728 5636
rect 2412 5652 2464 5704
rect 4160 5720 4212 5772
rect 4436 5652 4488 5704
rect 6828 5856 6880 5908
rect 6920 5856 6972 5908
rect 5816 5720 5868 5772
rect 3884 5627 3936 5636
rect 3884 5593 3893 5627
rect 3893 5593 3927 5627
rect 3927 5593 3936 5627
rect 3884 5584 3936 5593
rect 5540 5652 5592 5704
rect 5080 5584 5132 5636
rect 7196 5788 7248 5840
rect 8392 5720 8444 5772
rect 9220 5856 9272 5908
rect 9956 5899 10008 5908
rect 9956 5865 9965 5899
rect 9965 5865 9999 5899
rect 9999 5865 10008 5899
rect 9956 5856 10008 5865
rect 11336 5899 11388 5908
rect 11336 5865 11345 5899
rect 11345 5865 11379 5899
rect 11379 5865 11388 5899
rect 11336 5856 11388 5865
rect 12256 5856 12308 5908
rect 9220 5665 9272 5704
rect 6368 5584 6420 5636
rect 8760 5584 8812 5636
rect 9220 5652 9245 5665
rect 9245 5652 9272 5665
rect 9772 5788 9824 5840
rect 12716 5856 12768 5908
rect 12164 5720 12216 5772
rect 2504 5516 2556 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 4068 5516 4120 5568
rect 5540 5516 5592 5568
rect 7104 5516 7156 5568
rect 9772 5652 9824 5704
rect 11796 5652 11848 5704
rect 12440 5652 12492 5704
rect 10232 5584 10284 5636
rect 13084 5788 13136 5840
rect 14004 5788 14056 5840
rect 15384 5856 15436 5908
rect 18788 5856 18840 5908
rect 20076 5856 20128 5908
rect 13728 5763 13780 5772
rect 13728 5729 13737 5763
rect 13737 5729 13771 5763
rect 13771 5729 13780 5763
rect 13728 5720 13780 5729
rect 12900 5652 12952 5704
rect 13912 5720 13964 5772
rect 15568 5788 15620 5840
rect 15752 5788 15804 5840
rect 17132 5788 17184 5840
rect 15476 5720 15528 5772
rect 14372 5695 14424 5704
rect 14372 5661 14379 5695
rect 14379 5661 14413 5695
rect 14413 5661 14424 5695
rect 14372 5652 14424 5661
rect 10048 5516 10100 5568
rect 10784 5516 10836 5568
rect 12992 5516 13044 5568
rect 13636 5584 13688 5636
rect 13452 5516 13504 5568
rect 13728 5516 13780 5568
rect 13912 5627 13964 5636
rect 13912 5593 13921 5627
rect 13921 5593 13955 5627
rect 13955 5593 13964 5627
rect 13912 5584 13964 5593
rect 14096 5584 14148 5636
rect 15384 5652 15436 5704
rect 14832 5584 14884 5636
rect 16212 5652 16264 5704
rect 16488 5652 16540 5704
rect 18144 5720 18196 5772
rect 17960 5652 18012 5704
rect 18788 5652 18840 5704
rect 20168 5652 20220 5704
rect 14648 5516 14700 5568
rect 15200 5516 15252 5568
rect 15384 5516 15436 5568
rect 16120 5584 16172 5636
rect 16672 5584 16724 5636
rect 17868 5584 17920 5636
rect 19616 5584 19668 5636
rect 19800 5584 19852 5636
rect 16856 5516 16908 5568
rect 16948 5516 17000 5568
rect 5894 5414 5946 5466
rect 5958 5414 6010 5466
rect 6022 5414 6074 5466
rect 6086 5414 6138 5466
rect 6150 5414 6202 5466
rect 10839 5414 10891 5466
rect 10903 5414 10955 5466
rect 10967 5414 11019 5466
rect 11031 5414 11083 5466
rect 11095 5414 11147 5466
rect 15784 5414 15836 5466
rect 15848 5414 15900 5466
rect 15912 5414 15964 5466
rect 15976 5414 16028 5466
rect 16040 5414 16092 5466
rect 20729 5414 20781 5466
rect 20793 5414 20845 5466
rect 20857 5414 20909 5466
rect 20921 5414 20973 5466
rect 20985 5414 21037 5466
rect 1308 5312 1360 5364
rect 3884 5312 3936 5364
rect 3976 5312 4028 5364
rect 5448 5312 5500 5364
rect 6276 5312 6328 5364
rect 6736 5312 6788 5364
rect 7012 5312 7064 5364
rect 7840 5355 7892 5364
rect 7840 5321 7849 5355
rect 7849 5321 7883 5355
rect 7883 5321 7892 5355
rect 7840 5312 7892 5321
rect 7932 5312 7984 5364
rect 9220 5312 9272 5364
rect 9404 5355 9456 5364
rect 9404 5321 9413 5355
rect 9413 5321 9447 5355
rect 9447 5321 9456 5355
rect 9404 5312 9456 5321
rect 10048 5312 10100 5364
rect 10692 5312 10744 5364
rect 11244 5312 11296 5364
rect 11704 5312 11756 5364
rect 11796 5355 11848 5364
rect 11796 5321 11805 5355
rect 11805 5321 11839 5355
rect 11839 5321 11848 5355
rect 11796 5312 11848 5321
rect 12256 5312 12308 5364
rect 13360 5312 13412 5364
rect 1952 5176 2004 5228
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 2136 5176 2188 5185
rect 2320 5176 2372 5228
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2596 5176 2648 5228
rect 3378 5176 3430 5228
rect 4436 5176 4488 5228
rect 4528 5219 4580 5228
rect 4528 5185 4537 5219
rect 4537 5185 4571 5219
rect 4571 5185 4580 5219
rect 4528 5176 4580 5185
rect 5356 5219 5408 5228
rect 5356 5185 5390 5219
rect 5390 5185 5408 5219
rect 5356 5176 5408 5185
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 6828 5219 6880 5228
rect 6828 5185 6837 5219
rect 6837 5185 6871 5219
rect 6871 5185 6880 5219
rect 6828 5176 6880 5185
rect 7196 5176 7248 5228
rect 7380 5176 7432 5228
rect 7656 5287 7708 5296
rect 7656 5253 7665 5287
rect 7665 5253 7699 5287
rect 7699 5253 7708 5287
rect 7656 5244 7708 5253
rect 10324 5244 10376 5296
rect 8392 5219 8444 5228
rect 8392 5185 8401 5219
rect 8401 5185 8435 5219
rect 8435 5185 8444 5219
rect 8392 5176 8444 5185
rect 8668 5219 8720 5228
rect 8668 5185 8675 5219
rect 8675 5185 8709 5219
rect 8709 5185 8720 5219
rect 8668 5176 8720 5185
rect 9036 5176 9088 5228
rect 9220 5176 9272 5228
rect 2780 5108 2832 5160
rect 2228 5040 2280 5092
rect 2596 5040 2648 5092
rect 4160 5108 4212 5160
rect 6368 5108 6420 5160
rect 10968 5108 11020 5160
rect 11520 5108 11572 5160
rect 3976 5040 4028 5092
rect 2780 4972 2832 5024
rect 10692 5040 10744 5092
rect 12164 5244 12216 5296
rect 13636 5312 13688 5364
rect 13728 5312 13780 5364
rect 14188 5312 14240 5364
rect 14740 5312 14792 5364
rect 14924 5312 14976 5364
rect 15108 5312 15160 5364
rect 15384 5312 15436 5364
rect 15752 5312 15804 5364
rect 16212 5312 16264 5364
rect 12716 5176 12768 5228
rect 14280 5244 14332 5296
rect 15016 5244 15068 5296
rect 13084 5219 13136 5228
rect 13084 5185 13093 5219
rect 13093 5185 13127 5219
rect 13127 5185 13136 5219
rect 13084 5176 13136 5185
rect 13268 5176 13320 5228
rect 13360 5176 13412 5228
rect 12532 5108 12584 5160
rect 12716 5040 12768 5092
rect 13084 5040 13136 5092
rect 13636 5176 13688 5228
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 14924 5176 14976 5228
rect 15476 5219 15528 5228
rect 15476 5185 15485 5219
rect 15485 5185 15519 5219
rect 15519 5185 15528 5219
rect 15476 5176 15528 5185
rect 15200 5108 15252 5160
rect 13544 5040 13596 5092
rect 15108 5083 15160 5092
rect 15108 5049 15117 5083
rect 15117 5049 15151 5083
rect 15151 5049 15160 5083
rect 15108 5040 15160 5049
rect 15384 5040 15436 5092
rect 16764 5244 16816 5296
rect 17592 5312 17644 5364
rect 17684 5312 17736 5364
rect 19984 5312 20036 5364
rect 16304 5176 16356 5228
rect 16488 5176 16540 5228
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17500 5176 17552 5228
rect 17684 5219 17736 5228
rect 17684 5185 17693 5219
rect 17693 5185 17727 5219
rect 17727 5185 17736 5219
rect 17684 5176 17736 5185
rect 18788 5176 18840 5228
rect 18880 5176 18932 5228
rect 19432 5219 19484 5228
rect 19432 5185 19466 5219
rect 19466 5185 19484 5219
rect 19432 5176 19484 5185
rect 20444 5176 20496 5228
rect 16120 5040 16172 5092
rect 18604 5108 18656 5160
rect 5356 4972 5408 5024
rect 9864 4972 9916 5024
rect 13452 4972 13504 5024
rect 13728 4972 13780 5024
rect 14372 4972 14424 5024
rect 14464 4972 14516 5024
rect 16488 4972 16540 5024
rect 16764 4972 16816 5024
rect 18696 5083 18748 5092
rect 18696 5049 18705 5083
rect 18705 5049 18739 5083
rect 18739 5049 18748 5083
rect 18696 5040 18748 5049
rect 18788 4972 18840 5024
rect 3422 4870 3474 4922
rect 3486 4870 3538 4922
rect 3550 4870 3602 4922
rect 3614 4870 3666 4922
rect 3678 4870 3730 4922
rect 8367 4870 8419 4922
rect 8431 4870 8483 4922
rect 8495 4870 8547 4922
rect 8559 4870 8611 4922
rect 8623 4870 8675 4922
rect 13312 4870 13364 4922
rect 13376 4870 13428 4922
rect 13440 4870 13492 4922
rect 13504 4870 13556 4922
rect 13568 4870 13620 4922
rect 18257 4870 18309 4922
rect 18321 4870 18373 4922
rect 18385 4870 18437 4922
rect 18449 4870 18501 4922
rect 18513 4870 18565 4922
rect 1216 4768 1268 4820
rect 2044 4768 2096 4820
rect 572 4564 624 4616
rect 1768 4564 1820 4616
rect 2688 4768 2740 4820
rect 3332 4811 3384 4820
rect 3332 4777 3341 4811
rect 3341 4777 3375 4811
rect 3375 4777 3384 4811
rect 3332 4768 3384 4777
rect 3516 4768 3568 4820
rect 3976 4768 4028 4820
rect 3056 4700 3108 4752
rect 4988 4768 5040 4820
rect 3332 4632 3384 4684
rect 6368 4811 6420 4820
rect 6368 4777 6377 4811
rect 6377 4777 6411 4811
rect 6411 4777 6420 4811
rect 6368 4768 6420 4777
rect 7104 4768 7156 4820
rect 7196 4768 7248 4820
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 10508 4768 10560 4820
rect 10876 4768 10928 4820
rect 7564 4700 7616 4752
rect 9496 4700 9548 4752
rect 10416 4700 10468 4752
rect 6736 4675 6788 4684
rect 6736 4641 6745 4675
rect 6745 4641 6779 4675
rect 6779 4641 6788 4675
rect 6736 4632 6788 4641
rect 10048 4632 10100 4684
rect 11428 4768 11480 4820
rect 11612 4768 11664 4820
rect 13084 4768 13136 4820
rect 2504 4564 2556 4616
rect 3608 4564 3660 4616
rect 4068 4564 4120 4616
rect 4528 4564 4580 4616
rect 1952 4496 2004 4548
rect 4344 4496 4396 4548
rect 4436 4539 4488 4548
rect 4436 4505 4445 4539
rect 4445 4505 4479 4539
rect 4479 4505 4488 4539
rect 4436 4496 4488 4505
rect 10784 4632 10836 4684
rect 11152 4632 11204 4684
rect 11428 4632 11480 4684
rect 11888 4632 11940 4684
rect 12256 4632 12308 4684
rect 5448 4496 5500 4548
rect 6736 4496 6788 4548
rect 10692 4564 10744 4616
rect 10968 4564 11020 4616
rect 11980 4607 12032 4616
rect 11980 4573 11989 4607
rect 11989 4573 12023 4607
rect 12023 4573 12032 4607
rect 11980 4564 12032 4573
rect 12624 4632 12676 4684
rect 12992 4700 13044 4752
rect 13820 4811 13872 4820
rect 13820 4777 13829 4811
rect 13829 4777 13863 4811
rect 13863 4777 13872 4811
rect 13820 4768 13872 4777
rect 14096 4768 14148 4820
rect 13268 4700 13320 4752
rect 13176 4632 13228 4684
rect 13452 4632 13504 4684
rect 14556 4700 14608 4752
rect 15292 4768 15344 4820
rect 15200 4700 15252 4752
rect 14648 4632 14700 4684
rect 15568 4768 15620 4820
rect 15660 4768 15712 4820
rect 18788 4768 18840 4820
rect 17316 4700 17368 4752
rect 17776 4700 17828 4752
rect 19800 4700 19852 4752
rect 20076 4743 20128 4752
rect 20076 4709 20085 4743
rect 20085 4709 20119 4743
rect 20119 4709 20128 4743
rect 20076 4700 20128 4709
rect 6828 4428 6880 4480
rect 10048 4428 10100 4480
rect 11888 4428 11940 4480
rect 12440 4496 12492 4548
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13544 4564 13596 4616
rect 12164 4428 12216 4480
rect 14004 4496 14056 4548
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 14740 4607 14792 4616
rect 14740 4573 14749 4607
rect 14749 4573 14783 4607
rect 14783 4573 14792 4607
rect 14740 4564 14792 4573
rect 14832 4564 14884 4616
rect 15108 4641 15117 4650
rect 15117 4641 15151 4650
rect 15151 4641 15160 4650
rect 15108 4598 15160 4641
rect 16672 4632 16724 4684
rect 16948 4632 17000 4684
rect 18144 4632 18196 4684
rect 20444 4632 20496 4684
rect 16580 4564 16632 4616
rect 12992 4428 13044 4480
rect 14188 4428 14240 4480
rect 14464 4428 14516 4480
rect 14924 4496 14976 4548
rect 15752 4496 15804 4548
rect 17132 4496 17184 4548
rect 18236 4564 18288 4616
rect 19248 4607 19300 4616
rect 19248 4573 19257 4607
rect 19257 4573 19291 4607
rect 19291 4573 19300 4607
rect 19248 4564 19300 4573
rect 19616 4607 19668 4616
rect 19616 4573 19625 4607
rect 19625 4573 19659 4607
rect 19659 4573 19668 4607
rect 19616 4564 19668 4573
rect 17776 4496 17828 4548
rect 16488 4428 16540 4480
rect 16764 4471 16816 4480
rect 16764 4437 16773 4471
rect 16773 4437 16807 4471
rect 16807 4437 16816 4471
rect 16764 4428 16816 4437
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 17224 4428 17276 4480
rect 19064 4496 19116 4548
rect 19432 4496 19484 4548
rect 18788 4428 18840 4480
rect 21456 4428 21508 4480
rect 5894 4326 5946 4378
rect 5958 4326 6010 4378
rect 6022 4326 6074 4378
rect 6086 4326 6138 4378
rect 6150 4326 6202 4378
rect 10839 4326 10891 4378
rect 10903 4326 10955 4378
rect 10967 4326 11019 4378
rect 11031 4326 11083 4378
rect 11095 4326 11147 4378
rect 15784 4326 15836 4378
rect 15848 4326 15900 4378
rect 15912 4326 15964 4378
rect 15976 4326 16028 4378
rect 16040 4326 16092 4378
rect 20729 4326 20781 4378
rect 20793 4326 20845 4378
rect 20857 4326 20909 4378
rect 20921 4326 20973 4378
rect 20985 4326 21037 4378
rect 5356 4224 5408 4276
rect 10232 4224 10284 4276
rect 10416 4224 10468 4276
rect 10600 4224 10652 4276
rect 11152 4224 11204 4276
rect 11704 4224 11756 4276
rect 13360 4224 13412 4276
rect 13728 4224 13780 4276
rect 14096 4224 14148 4276
rect 5816 4156 5868 4208
rect 7288 4156 7340 4208
rect 10140 4156 10192 4208
rect 2320 4063 2372 4072
rect 2320 4029 2329 4063
rect 2329 4029 2363 4063
rect 2363 4029 2372 4063
rect 2320 4020 2372 4029
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 2688 4020 2740 4072
rect 2872 4020 2924 4072
rect 3424 4088 3476 4140
rect 3884 4020 3936 4072
rect 2228 3952 2280 4004
rect 2780 3952 2832 4004
rect 2964 3995 3016 4004
rect 2964 3961 2973 3995
rect 2973 3961 3007 3995
rect 3007 3961 3016 3995
rect 2964 3952 3016 3961
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 8760 4088 8812 4140
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 10600 4131 10652 4140
rect 10600 4097 10609 4131
rect 10609 4097 10643 4131
rect 10643 4097 10652 4131
rect 10600 4088 10652 4097
rect 5816 4020 5868 4072
rect 7472 4020 7524 4072
rect 11336 4131 11388 4140
rect 11336 4097 11345 4131
rect 11345 4097 11379 4131
rect 11379 4097 11388 4131
rect 11336 4088 11388 4097
rect 11520 4088 11572 4140
rect 11704 4088 11756 4140
rect 12072 4131 12124 4140
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12072 4088 12124 4097
rect 12348 4131 12400 4140
rect 12348 4097 12357 4131
rect 12357 4097 12391 4131
rect 12391 4097 12400 4131
rect 12348 4088 12400 4097
rect 13544 4156 13596 4208
rect 10600 3952 10652 4004
rect 11796 3952 11848 4004
rect 12532 4020 12584 4072
rect 5080 3884 5132 3936
rect 5632 3884 5684 3936
rect 6736 3884 6788 3936
rect 9036 3884 9088 3936
rect 9220 3927 9272 3936
rect 9220 3893 9229 3927
rect 9229 3893 9263 3927
rect 9263 3893 9272 3927
rect 9220 3884 9272 3893
rect 10048 3927 10100 3936
rect 10048 3893 10057 3927
rect 10057 3893 10091 3927
rect 10091 3893 10100 3927
rect 10048 3884 10100 3893
rect 10692 3927 10744 3936
rect 10692 3893 10701 3927
rect 10701 3893 10735 3927
rect 10735 3893 10744 3927
rect 10692 3884 10744 3893
rect 11336 3884 11388 3936
rect 11612 3884 11664 3936
rect 11888 3927 11940 3936
rect 11888 3893 11897 3927
rect 11897 3893 11931 3927
rect 11931 3893 11940 3927
rect 11888 3884 11940 3893
rect 12348 3952 12400 4004
rect 13084 4088 13136 4140
rect 13820 4156 13872 4208
rect 12992 4020 13044 4072
rect 13360 4020 13412 4072
rect 13176 3952 13228 4004
rect 14832 4156 14884 4208
rect 14924 4156 14976 4208
rect 15660 4156 15712 4208
rect 15844 4224 15896 4276
rect 16396 4224 16448 4276
rect 17224 4224 17276 4276
rect 13820 4020 13872 4072
rect 16120 4088 16172 4140
rect 16856 4199 16908 4208
rect 16856 4165 16865 4199
rect 16865 4165 16899 4199
rect 16899 4165 16908 4199
rect 16856 4156 16908 4165
rect 19156 4224 19208 4276
rect 19892 4267 19944 4276
rect 19892 4233 19901 4267
rect 19901 4233 19935 4267
rect 19935 4233 19944 4267
rect 19892 4224 19944 4233
rect 20444 4267 20496 4276
rect 20444 4233 20453 4267
rect 20453 4233 20487 4267
rect 20487 4233 20496 4267
rect 20444 4224 20496 4233
rect 16396 4088 16448 4140
rect 17500 4156 17552 4208
rect 17316 4088 17368 4140
rect 17408 4131 17460 4140
rect 17408 4097 17415 4131
rect 17415 4097 17449 4131
rect 17449 4097 17460 4131
rect 17408 4088 17460 4097
rect 13912 3952 13964 4004
rect 14004 3952 14056 4004
rect 15660 4020 15712 4072
rect 16028 4020 16080 4072
rect 18880 4156 18932 4208
rect 19064 4156 19116 4208
rect 18604 4088 18656 4140
rect 19708 4088 19760 4140
rect 17960 4020 18012 4072
rect 18144 4020 18196 4072
rect 21180 4020 21232 4072
rect 14464 3884 14516 3936
rect 15200 3884 15252 3936
rect 16948 3927 17000 3936
rect 16948 3893 16957 3927
rect 16957 3893 16991 3927
rect 16991 3893 17000 3927
rect 16948 3884 17000 3893
rect 17960 3884 18012 3936
rect 19156 3884 19208 3936
rect 3422 3782 3474 3834
rect 3486 3782 3538 3834
rect 3550 3782 3602 3834
rect 3614 3782 3666 3834
rect 3678 3782 3730 3834
rect 8367 3782 8419 3834
rect 8431 3782 8483 3834
rect 8495 3782 8547 3834
rect 8559 3782 8611 3834
rect 8623 3782 8675 3834
rect 13312 3782 13364 3834
rect 13376 3782 13428 3834
rect 13440 3782 13492 3834
rect 13504 3782 13556 3834
rect 13568 3782 13620 3834
rect 18257 3782 18309 3834
rect 18321 3782 18373 3834
rect 18385 3782 18437 3834
rect 18449 3782 18501 3834
rect 18513 3782 18565 3834
rect 2596 3723 2648 3732
rect 2596 3689 2605 3723
rect 2605 3689 2639 3723
rect 2639 3689 2648 3723
rect 2596 3680 2648 3689
rect 3148 3723 3200 3732
rect 3148 3689 3157 3723
rect 3157 3689 3191 3723
rect 3191 3689 3200 3723
rect 3148 3680 3200 3689
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 4344 3723 4396 3732
rect 4344 3689 4353 3723
rect 4353 3689 4387 3723
rect 4387 3689 4396 3723
rect 4344 3680 4396 3689
rect 4436 3680 4488 3732
rect 6368 3680 6420 3732
rect 7748 3680 7800 3732
rect 7840 3680 7892 3732
rect 9772 3680 9824 3732
rect 9864 3680 9916 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 11428 3680 11480 3732
rect 11520 3680 11572 3732
rect 12256 3680 12308 3732
rect 1768 3476 1820 3528
rect 5448 3612 5500 3664
rect 7196 3612 7248 3664
rect 11152 3612 11204 3664
rect 4528 3519 4580 3528
rect 4528 3485 4537 3519
rect 4537 3485 4571 3519
rect 4571 3485 4580 3519
rect 4528 3476 4580 3485
rect 3332 3408 3384 3460
rect 3976 3408 4028 3460
rect 1676 3340 1728 3392
rect 5724 3476 5776 3528
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 7012 3519 7064 3528
rect 7012 3485 7021 3519
rect 7021 3485 7055 3519
rect 7055 3485 7064 3519
rect 7012 3476 7064 3485
rect 7104 3476 7156 3528
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 9128 3519 9180 3528
rect 9128 3485 9137 3519
rect 9137 3485 9171 3519
rect 9171 3485 9180 3519
rect 9128 3476 9180 3485
rect 9404 3476 9456 3528
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 11060 3544 11112 3596
rect 5448 3408 5500 3460
rect 5356 3340 5408 3392
rect 6276 3340 6328 3392
rect 6828 3383 6880 3392
rect 6828 3349 6837 3383
rect 6837 3349 6871 3383
rect 6871 3349 6880 3383
rect 6828 3340 6880 3349
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 12164 3612 12216 3664
rect 12440 3612 12492 3664
rect 12900 3612 12952 3664
rect 13820 3612 13872 3664
rect 7748 3383 7800 3392
rect 7748 3349 7757 3383
rect 7757 3349 7791 3383
rect 7791 3349 7800 3383
rect 7748 3340 7800 3349
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 9404 3340 9456 3392
rect 10324 3340 10376 3392
rect 10600 3340 10652 3392
rect 11796 3476 11848 3528
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 12256 3519 12308 3528
rect 12256 3485 12265 3519
rect 12265 3485 12299 3519
rect 12299 3485 12308 3519
rect 12256 3476 12308 3485
rect 12532 3519 12584 3528
rect 12532 3485 12541 3519
rect 12541 3485 12575 3519
rect 12575 3485 12584 3519
rect 12532 3476 12584 3485
rect 12716 3544 12768 3596
rect 18696 3680 18748 3732
rect 19340 3680 19392 3732
rect 14096 3612 14148 3664
rect 14924 3612 14976 3664
rect 15384 3612 15436 3664
rect 16212 3612 16264 3664
rect 17224 3612 17276 3664
rect 13820 3476 13872 3528
rect 14832 3544 14884 3596
rect 15200 3544 15252 3596
rect 18144 3612 18196 3664
rect 12256 3340 12308 3392
rect 14832 3408 14884 3460
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 20168 3587 20220 3596
rect 20168 3553 20177 3587
rect 20177 3553 20211 3587
rect 20211 3553 20220 3587
rect 20168 3544 20220 3553
rect 15844 3476 15896 3528
rect 16304 3476 16356 3528
rect 12624 3340 12676 3392
rect 12808 3340 12860 3392
rect 12992 3340 13044 3392
rect 13358 3340 13410 3392
rect 13636 3340 13688 3392
rect 15384 3340 15436 3392
rect 16120 3340 16172 3392
rect 16856 3408 16908 3460
rect 17316 3408 17368 3460
rect 17960 3476 18012 3528
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 18328 3476 18380 3528
rect 19064 3476 19116 3528
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 18972 3408 19024 3460
rect 21272 3340 21324 3392
rect 5894 3238 5946 3290
rect 5958 3238 6010 3290
rect 6022 3238 6074 3290
rect 6086 3238 6138 3290
rect 6150 3238 6202 3290
rect 10839 3238 10891 3290
rect 10903 3238 10955 3290
rect 10967 3238 11019 3290
rect 11031 3238 11083 3290
rect 11095 3238 11147 3290
rect 15784 3238 15836 3290
rect 15848 3238 15900 3290
rect 15912 3238 15964 3290
rect 15976 3238 16028 3290
rect 16040 3238 16092 3290
rect 20729 3238 20781 3290
rect 20793 3238 20845 3290
rect 20857 3238 20909 3290
rect 20921 3238 20973 3290
rect 20985 3238 21037 3290
rect 1584 3179 1636 3188
rect 1584 3145 1593 3179
rect 1593 3145 1627 3179
rect 1627 3145 1636 3179
rect 1584 3136 1636 3145
rect 3056 3136 3108 3188
rect 3884 3136 3936 3188
rect 4160 3136 4212 3188
rect 7380 3136 7432 3188
rect 8300 3136 8352 3188
rect 2780 3068 2832 3120
rect 1768 3000 1820 3052
rect 3240 3068 3292 3120
rect 5540 3068 5592 3120
rect 3056 3000 3108 3052
rect 5724 3000 5776 3052
rect 6644 3043 6696 3052
rect 6644 3009 6653 3043
rect 6653 3009 6687 3043
rect 6687 3009 6696 3043
rect 6644 3000 6696 3009
rect 8392 3068 8444 3120
rect 4620 2932 4672 2984
rect 5816 2932 5868 2984
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 7932 3000 7984 3052
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8024 3000 8076 3009
rect 8300 3043 8352 3052
rect 8300 3009 8309 3043
rect 8309 3009 8343 3043
rect 8343 3009 8352 3043
rect 8300 3000 8352 3009
rect 8576 3043 8628 3052
rect 8576 3009 8585 3043
rect 8585 3009 8619 3043
rect 8619 3009 8628 3043
rect 8576 3000 8628 3009
rect 8852 3043 8904 3052
rect 8852 3009 8861 3043
rect 8861 3009 8895 3043
rect 8895 3009 8904 3043
rect 8852 3000 8904 3009
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 6552 2864 6604 2916
rect 7380 2864 7432 2916
rect 664 2796 716 2848
rect 3056 2796 3108 2848
rect 4896 2796 4948 2848
rect 5632 2796 5684 2848
rect 6644 2796 6696 2848
rect 6736 2839 6788 2848
rect 6736 2805 6745 2839
rect 6745 2805 6779 2839
rect 6779 2805 6788 2839
rect 6736 2796 6788 2805
rect 9220 2932 9272 2984
rect 10968 3136 11020 3188
rect 12716 3136 12768 3188
rect 12808 3136 12860 3188
rect 13360 3136 13412 3188
rect 9680 3043 9732 3052
rect 9680 3009 9689 3043
rect 9689 3009 9723 3043
rect 9723 3009 9732 3043
rect 9680 3000 9732 3009
rect 9956 3043 10008 3052
rect 9956 3009 9965 3043
rect 9965 3009 9999 3043
rect 9999 3009 10008 3043
rect 9956 3000 10008 3009
rect 10232 3000 10284 3052
rect 10784 3043 10836 3052
rect 10784 3009 10793 3043
rect 10793 3009 10827 3043
rect 10827 3009 10836 3043
rect 10784 3000 10836 3009
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11152 3043 11204 3052
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11704 3000 11756 3052
rect 10416 2932 10468 2984
rect 7564 2839 7616 2848
rect 7564 2805 7573 2839
rect 7573 2805 7607 2839
rect 7607 2805 7616 2839
rect 7564 2796 7616 2805
rect 7840 2839 7892 2848
rect 7840 2805 7849 2839
rect 7849 2805 7883 2839
rect 7883 2805 7892 2839
rect 7840 2796 7892 2805
rect 8116 2839 8168 2848
rect 8116 2805 8125 2839
rect 8125 2805 8159 2839
rect 8159 2805 8168 2839
rect 8116 2796 8168 2805
rect 8392 2839 8444 2848
rect 8392 2805 8401 2839
rect 8401 2805 8435 2839
rect 8435 2805 8444 2839
rect 8392 2796 8444 2805
rect 10048 2864 10100 2916
rect 11612 2932 11664 2984
rect 11888 3043 11940 3052
rect 11888 3009 11923 3043
rect 11923 3009 11940 3043
rect 11888 3000 11940 3009
rect 12072 3000 12124 3052
rect 12440 3000 12492 3052
rect 12808 3000 12860 3052
rect 13084 3000 13136 3052
rect 13912 3136 13964 3188
rect 14280 3136 14332 3188
rect 14372 3136 14424 3188
rect 14648 3136 14700 3188
rect 14832 3068 14884 3120
rect 15200 3136 15252 3188
rect 16764 3136 16816 3188
rect 16948 3136 17000 3188
rect 17316 3136 17368 3188
rect 17776 3136 17828 3188
rect 18236 3179 18288 3188
rect 18236 3145 18245 3179
rect 18245 3145 18279 3179
rect 18279 3145 18288 3179
rect 18236 3136 18288 3145
rect 18788 3136 18840 3188
rect 21824 3136 21876 3188
rect 15108 3068 15160 3120
rect 11888 2864 11940 2916
rect 12164 2864 12216 2916
rect 13728 2932 13780 2984
rect 12992 2864 13044 2916
rect 13360 2864 13412 2916
rect 14363 3000 14415 3052
rect 14004 2932 14056 2984
rect 14648 3043 14700 3052
rect 14648 3009 14657 3043
rect 14657 3009 14691 3043
rect 14691 3009 14700 3043
rect 14648 3000 14700 3009
rect 15476 3068 15528 3120
rect 16304 3111 16356 3120
rect 16304 3077 16313 3111
rect 16313 3077 16347 3111
rect 16347 3077 16356 3111
rect 16304 3068 16356 3077
rect 18328 3068 18380 3120
rect 18604 3068 18656 3120
rect 19524 3068 19576 3120
rect 16488 3043 16540 3052
rect 16488 3009 16497 3043
rect 16497 3009 16531 3043
rect 16531 3009 16540 3043
rect 16488 3000 16540 3009
rect 16580 3000 16632 3052
rect 17408 3000 17460 3052
rect 18788 3000 18840 3052
rect 14924 2975 14976 2984
rect 14924 2941 14933 2975
rect 14933 2941 14967 2975
rect 14967 2941 14976 2975
rect 14924 2932 14976 2941
rect 15292 2932 15344 2984
rect 15844 2932 15896 2984
rect 16672 2932 16724 2984
rect 8944 2839 8996 2848
rect 8944 2805 8953 2839
rect 8953 2805 8987 2839
rect 8987 2805 8996 2839
rect 8944 2796 8996 2805
rect 9220 2839 9272 2848
rect 9220 2805 9229 2839
rect 9229 2805 9263 2839
rect 9263 2805 9272 2839
rect 9220 2796 9272 2805
rect 9680 2796 9732 2848
rect 9772 2839 9824 2848
rect 9772 2805 9781 2839
rect 9781 2805 9815 2839
rect 9815 2805 9824 2839
rect 9772 2796 9824 2805
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 10692 2796 10744 2848
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 11428 2796 11480 2848
rect 13176 2796 13228 2848
rect 13820 2796 13872 2848
rect 13912 2839 13964 2848
rect 13912 2805 13921 2839
rect 13921 2805 13955 2839
rect 13955 2805 13964 2839
rect 13912 2796 13964 2805
rect 14280 2839 14332 2848
rect 14280 2805 14289 2839
rect 14289 2805 14323 2839
rect 14323 2805 14332 2839
rect 14280 2796 14332 2805
rect 15936 2864 15988 2916
rect 15292 2839 15344 2848
rect 15292 2805 15301 2839
rect 15301 2805 15335 2839
rect 15335 2805 15344 2839
rect 15292 2796 15344 2805
rect 15476 2796 15528 2848
rect 16120 2796 16172 2848
rect 16856 2796 16908 2848
rect 17224 2796 17276 2848
rect 3422 2694 3474 2746
rect 3486 2694 3538 2746
rect 3550 2694 3602 2746
rect 3614 2694 3666 2746
rect 3678 2694 3730 2746
rect 8367 2694 8419 2746
rect 8431 2694 8483 2746
rect 8495 2694 8547 2746
rect 8559 2694 8611 2746
rect 8623 2694 8675 2746
rect 13312 2694 13364 2746
rect 13376 2694 13428 2746
rect 13440 2694 13492 2746
rect 13504 2694 13556 2746
rect 13568 2694 13620 2746
rect 18257 2694 18309 2746
rect 18321 2694 18373 2746
rect 18385 2694 18437 2746
rect 18449 2694 18501 2746
rect 18513 2694 18565 2746
rect 1676 2635 1728 2644
rect 1676 2601 1685 2635
rect 1685 2601 1719 2635
rect 1719 2601 1728 2635
rect 1676 2592 1728 2601
rect 2964 2592 3016 2644
rect 3792 2592 3844 2644
rect 4436 2592 4488 2644
rect 5172 2592 5224 2644
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 6460 2592 6512 2644
rect 7012 2635 7064 2644
rect 7012 2601 7021 2635
rect 7021 2601 7055 2635
rect 7055 2601 7064 2635
rect 7012 2592 7064 2601
rect 7472 2592 7524 2644
rect 8392 2592 8444 2644
rect 9036 2592 9088 2644
rect 11428 2592 11480 2644
rect 11520 2592 11572 2644
rect 6276 2524 6328 2576
rect 1768 2456 1820 2508
rect 4068 2456 4120 2508
rect 3424 2431 3476 2440
rect 3424 2397 3433 2431
rect 3433 2397 3467 2431
rect 3467 2397 3476 2431
rect 3424 2388 3476 2397
rect 3792 2431 3844 2440
rect 3792 2397 3801 2431
rect 3801 2397 3835 2431
rect 3835 2397 3844 2431
rect 3792 2388 3844 2397
rect 4528 2431 4580 2440
rect 4528 2397 4537 2431
rect 4537 2397 4571 2431
rect 4571 2397 4580 2431
rect 4528 2388 4580 2397
rect 2964 2320 3016 2372
rect 4068 2320 4120 2372
rect 5632 2388 5684 2440
rect 6368 2388 6420 2440
rect 6644 2388 6696 2440
rect 7288 2388 7340 2440
rect 9312 2524 9364 2576
rect 11704 2524 11756 2576
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 5540 2363 5592 2372
rect 5540 2329 5549 2363
rect 5549 2329 5583 2363
rect 5583 2329 5592 2363
rect 5540 2320 5592 2329
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 5908 2252 5960 2304
rect 6276 2320 6328 2372
rect 9128 2388 9180 2440
rect 9496 2431 9548 2440
rect 9496 2397 9505 2431
rect 9505 2397 9539 2431
rect 9539 2397 9548 2431
rect 9496 2388 9548 2397
rect 10140 2431 10192 2440
rect 10140 2397 10149 2431
rect 10149 2397 10183 2431
rect 10183 2397 10192 2431
rect 10140 2388 10192 2397
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 11152 2388 11204 2440
rect 11244 2388 11296 2440
rect 11428 2431 11480 2440
rect 11428 2397 11437 2431
rect 11437 2397 11471 2431
rect 11471 2397 11480 2431
rect 11428 2388 11480 2397
rect 6184 2252 6236 2304
rect 8576 2252 8628 2304
rect 8944 2252 8996 2304
rect 9036 2295 9088 2304
rect 9036 2261 9045 2295
rect 9045 2261 9079 2295
rect 9079 2261 9088 2295
rect 9036 2252 9088 2261
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 9496 2252 9548 2304
rect 9864 2252 9916 2304
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 11244 2252 11296 2304
rect 11428 2252 11480 2304
rect 11612 2295 11664 2304
rect 11612 2261 11621 2295
rect 11621 2261 11655 2295
rect 11655 2261 11664 2295
rect 11612 2252 11664 2261
rect 12256 2431 12308 2440
rect 12256 2397 12265 2431
rect 12265 2397 12299 2431
rect 12299 2397 12308 2431
rect 12256 2388 12308 2397
rect 12532 2431 12584 2440
rect 12532 2397 12541 2431
rect 12541 2397 12575 2431
rect 12575 2397 12584 2431
rect 12532 2388 12584 2397
rect 12624 2388 12676 2440
rect 12900 2388 12952 2440
rect 13360 2388 13412 2440
rect 13912 2456 13964 2508
rect 14372 2524 14424 2576
rect 14648 2524 14700 2576
rect 13636 2388 13688 2440
rect 14188 2388 14240 2440
rect 11796 2320 11848 2372
rect 11980 2252 12032 2304
rect 12072 2295 12124 2304
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 14372 2320 14424 2372
rect 12440 2252 12492 2304
rect 12992 2295 13044 2304
rect 12992 2261 13001 2295
rect 13001 2261 13035 2295
rect 13035 2261 13044 2295
rect 12992 2252 13044 2261
rect 13728 2252 13780 2304
rect 14464 2252 14516 2304
rect 14832 2388 14884 2440
rect 16396 2635 16448 2644
rect 16396 2601 16405 2635
rect 16405 2601 16439 2635
rect 16439 2601 16448 2635
rect 16396 2592 16448 2601
rect 16580 2592 16632 2644
rect 20076 2592 20128 2644
rect 16488 2524 16540 2576
rect 19248 2524 19300 2576
rect 15660 2320 15712 2372
rect 15844 2320 15896 2372
rect 15936 2320 15988 2372
rect 17224 2456 17276 2508
rect 17500 2499 17552 2508
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17500 2456 17552 2465
rect 18696 2456 18748 2508
rect 16488 2388 16540 2440
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 19156 2320 19208 2372
rect 20260 2388 20312 2440
rect 14740 2252 14792 2304
rect 14924 2252 14976 2304
rect 16488 2252 16540 2304
rect 17040 2252 17092 2304
rect 17224 2252 17276 2304
rect 19248 2252 19300 2304
rect 19984 2295 20036 2304
rect 19984 2261 19993 2295
rect 19993 2261 20027 2295
rect 20027 2261 20036 2295
rect 19984 2252 20036 2261
rect 20352 2295 20404 2304
rect 20352 2261 20361 2295
rect 20361 2261 20395 2295
rect 20395 2261 20404 2295
rect 20352 2252 20404 2261
rect 5894 2150 5946 2202
rect 5958 2150 6010 2202
rect 6022 2150 6074 2202
rect 6086 2150 6138 2202
rect 6150 2150 6202 2202
rect 10839 2150 10891 2202
rect 10903 2150 10955 2202
rect 10967 2150 11019 2202
rect 11031 2150 11083 2202
rect 11095 2150 11147 2202
rect 15784 2150 15836 2202
rect 15848 2150 15900 2202
rect 15912 2150 15964 2202
rect 15976 2150 16028 2202
rect 16040 2150 16092 2202
rect 20729 2150 20781 2202
rect 20793 2150 20845 2202
rect 20857 2150 20909 2202
rect 20921 2150 20973 2202
rect 20985 2150 21037 2202
rect 1400 2048 1452 2100
rect 1308 1980 1360 2032
rect 4160 2048 4212 2100
rect 2412 2023 2464 2032
rect 2412 1989 2421 2023
rect 2421 1989 2455 2023
rect 2455 1989 2464 2023
rect 2412 1980 2464 1989
rect 2596 2023 2648 2032
rect 2596 1989 2605 2023
rect 2605 1989 2639 2023
rect 2639 1989 2648 2023
rect 2596 1980 2648 1989
rect 3240 1955 3292 1964
rect 3240 1921 3249 1955
rect 3249 1921 3283 1955
rect 3283 1921 3292 1955
rect 3240 1912 3292 1921
rect 756 1844 808 1896
rect 2780 1844 2832 1896
rect 3976 1955 4028 1964
rect 3976 1921 3985 1955
rect 3985 1921 4019 1955
rect 4019 1921 4028 1955
rect 3976 1912 4028 1921
rect 4160 1912 4212 1964
rect 4896 2048 4948 2100
rect 6552 2048 6604 2100
rect 6828 2048 6880 2100
rect 7012 2091 7064 2100
rect 7012 2057 7021 2091
rect 7021 2057 7055 2091
rect 7055 2057 7064 2091
rect 7012 2048 7064 2057
rect 7840 2048 7892 2100
rect 4988 1955 5040 1964
rect 4988 1921 4997 1955
rect 4997 1921 5031 1955
rect 5031 1921 5040 1955
rect 4988 1912 5040 1921
rect 5540 1912 5592 1964
rect 8116 1980 8168 2032
rect 8484 1980 8536 2032
rect 8576 1980 8628 2032
rect 9312 2048 9364 2100
rect 9956 2048 10008 2100
rect 11336 1980 11388 2032
rect 13544 1980 13596 2032
rect 14464 2048 14516 2100
rect 15292 2048 15344 2100
rect 16212 2048 16264 2100
rect 16396 2048 16448 2100
rect 16580 2048 16632 2100
rect 4712 1887 4764 1896
rect 4712 1853 4721 1887
rect 4721 1853 4755 1887
rect 4755 1853 4764 1887
rect 4712 1844 4764 1853
rect 5172 1844 5224 1896
rect 6276 1776 6328 1828
rect 4528 1708 4580 1760
rect 6000 1708 6052 1760
rect 6920 1912 6972 1964
rect 7564 1912 7616 1964
rect 7748 1912 7800 1964
rect 8208 1912 8260 1964
rect 9312 1955 9364 1964
rect 9312 1921 9321 1955
rect 9321 1921 9355 1955
rect 9355 1921 9364 1955
rect 9312 1912 9364 1921
rect 9588 1912 9640 1964
rect 7472 1776 7524 1828
rect 6920 1708 6972 1760
rect 7840 1776 7892 1828
rect 8852 1776 8904 1828
rect 9680 1776 9732 1828
rect 11888 1912 11940 1964
rect 12624 1912 12676 1964
rect 14280 1980 14332 2032
rect 14372 1980 14424 2032
rect 14924 1980 14976 2032
rect 11152 1844 11204 1896
rect 12440 1844 12492 1896
rect 12900 1844 12952 1896
rect 10876 1776 10928 1828
rect 7656 1708 7708 1760
rect 8116 1751 8168 1760
rect 8116 1717 8125 1751
rect 8125 1717 8159 1751
rect 8159 1717 8168 1751
rect 8116 1708 8168 1717
rect 8208 1708 8260 1760
rect 9404 1708 9456 1760
rect 9588 1751 9640 1760
rect 9588 1717 9597 1751
rect 9597 1717 9631 1751
rect 9631 1717 9640 1751
rect 9588 1708 9640 1717
rect 10140 1751 10192 1760
rect 10140 1717 10149 1751
rect 10149 1717 10183 1751
rect 10183 1717 10192 1751
rect 10140 1708 10192 1717
rect 10508 1751 10560 1760
rect 10508 1717 10517 1751
rect 10517 1717 10551 1751
rect 10551 1717 10560 1751
rect 10508 1708 10560 1717
rect 10692 1708 10744 1760
rect 11888 1751 11940 1760
rect 11888 1717 11897 1751
rect 11897 1717 11931 1751
rect 11931 1717 11940 1751
rect 11888 1708 11940 1717
rect 12164 1776 12216 1828
rect 12808 1776 12860 1828
rect 12532 1708 12584 1760
rect 13636 1776 13688 1828
rect 14096 1844 14148 1896
rect 14280 1844 14332 1896
rect 14464 1776 14516 1828
rect 14740 1819 14792 1828
rect 14740 1785 14749 1819
rect 14749 1785 14783 1819
rect 14783 1785 14792 1819
rect 14740 1776 14792 1785
rect 14924 1844 14976 1896
rect 15292 1844 15344 1896
rect 16028 1887 16080 1896
rect 16028 1853 16037 1887
rect 16037 1853 16071 1887
rect 16071 1853 16080 1887
rect 16028 1844 16080 1853
rect 16304 1912 16356 1964
rect 17040 1912 17092 1964
rect 20536 1955 20588 1964
rect 20536 1921 20545 1955
rect 20545 1921 20579 1955
rect 20579 1921 20588 1955
rect 20536 1912 20588 1921
rect 17500 1844 17552 1896
rect 12992 1751 13044 1760
rect 12992 1717 13001 1751
rect 13001 1717 13035 1751
rect 13035 1717 13044 1751
rect 12992 1708 13044 1717
rect 13084 1708 13136 1760
rect 13728 1708 13780 1760
rect 14188 1708 14240 1760
rect 16396 1708 16448 1760
rect 16488 1708 16540 1760
rect 3422 1606 3474 1658
rect 3486 1606 3538 1658
rect 3550 1606 3602 1658
rect 3614 1606 3666 1658
rect 3678 1606 3730 1658
rect 8367 1606 8419 1658
rect 8431 1606 8483 1658
rect 8495 1606 8547 1658
rect 8559 1606 8611 1658
rect 8623 1606 8675 1658
rect 13312 1606 13364 1658
rect 13376 1606 13428 1658
rect 13440 1606 13492 1658
rect 13504 1606 13556 1658
rect 13568 1606 13620 1658
rect 18257 1606 18309 1658
rect 18321 1606 18373 1658
rect 18385 1606 18437 1658
rect 18449 1606 18501 1658
rect 18513 1606 18565 1658
rect 1860 1547 1912 1556
rect 1860 1513 1869 1547
rect 1869 1513 1903 1547
rect 1903 1513 1912 1547
rect 1860 1504 1912 1513
rect 2504 1504 2556 1556
rect 4160 1504 4212 1556
rect 4344 1504 4396 1556
rect 4988 1547 5040 1556
rect 4988 1513 4997 1547
rect 4997 1513 5031 1547
rect 5031 1513 5040 1547
rect 4988 1504 5040 1513
rect 5080 1504 5132 1556
rect 480 1436 532 1488
rect 1032 1368 1084 1420
rect 20 1300 72 1352
rect 1768 1275 1820 1284
rect 1768 1241 1777 1275
rect 1777 1241 1811 1275
rect 1811 1241 1820 1275
rect 1768 1232 1820 1241
rect 2412 1232 2464 1284
rect 2596 1164 2648 1216
rect 3700 1300 3752 1352
rect 4896 1436 4948 1488
rect 5264 1436 5316 1488
rect 6092 1547 6144 1556
rect 6092 1513 6101 1547
rect 6101 1513 6135 1547
rect 6135 1513 6144 1547
rect 6092 1504 6144 1513
rect 6644 1547 6696 1556
rect 6644 1513 6653 1547
rect 6653 1513 6687 1547
rect 6687 1513 6696 1547
rect 6644 1504 6696 1513
rect 6828 1504 6880 1556
rect 9312 1504 9364 1556
rect 9772 1504 9824 1556
rect 10600 1504 10652 1556
rect 6000 1436 6052 1488
rect 5172 1368 5224 1420
rect 5356 1300 5408 1352
rect 4436 1232 4488 1284
rect 4528 1275 4580 1284
rect 4528 1241 4537 1275
rect 4537 1241 4571 1275
rect 4571 1241 4580 1275
rect 4528 1232 4580 1241
rect 4896 1275 4948 1284
rect 4896 1241 4905 1275
rect 4905 1241 4939 1275
rect 4939 1241 4948 1275
rect 4896 1232 4948 1241
rect 5264 1275 5316 1284
rect 5264 1241 5273 1275
rect 5273 1241 5307 1275
rect 5307 1241 5316 1275
rect 5264 1232 5316 1241
rect 5080 1164 5132 1216
rect 6368 1300 6420 1352
rect 6552 1300 6604 1352
rect 6736 1300 6788 1352
rect 7840 1343 7892 1352
rect 7840 1309 7849 1343
rect 7849 1309 7883 1343
rect 7883 1309 7892 1343
rect 7840 1300 7892 1309
rect 9864 1436 9916 1488
rect 10324 1436 10376 1488
rect 11980 1436 12032 1488
rect 10048 1354 10100 1406
rect 11612 1354 11664 1406
rect 11796 1368 11848 1420
rect 12256 1368 12308 1420
rect 12440 1504 12492 1556
rect 12624 1436 12676 1488
rect 13360 1436 13412 1488
rect 13636 1436 13688 1488
rect 13268 1368 13320 1420
rect 14096 1479 14148 1488
rect 14096 1445 14105 1479
rect 14105 1445 14139 1479
rect 14139 1445 14148 1479
rect 14096 1436 14148 1445
rect 9772 1300 9824 1352
rect 7564 1207 7616 1216
rect 7564 1173 7573 1207
rect 7573 1173 7607 1207
rect 7607 1173 7616 1207
rect 7564 1164 7616 1173
rect 9496 1232 9548 1284
rect 11060 1343 11112 1352
rect 11060 1309 11069 1343
rect 11069 1309 11103 1343
rect 11103 1309 11112 1343
rect 11060 1300 11112 1309
rect 11244 1300 11296 1352
rect 11520 1343 11572 1352
rect 11520 1309 11529 1343
rect 11529 1309 11563 1343
rect 11563 1309 11572 1343
rect 11520 1300 11572 1309
rect 11428 1232 11480 1284
rect 11704 1300 11756 1352
rect 12716 1300 12768 1352
rect 11888 1232 11940 1284
rect 12256 1232 12308 1284
rect 12440 1232 12492 1284
rect 12900 1232 12952 1284
rect 13544 1343 13596 1352
rect 13544 1309 13553 1343
rect 13553 1309 13587 1343
rect 13587 1309 13596 1343
rect 13544 1300 13596 1309
rect 14188 1368 14240 1420
rect 14648 1504 14700 1556
rect 15016 1504 15068 1556
rect 15384 1504 15436 1556
rect 15476 1504 15528 1556
rect 16580 1504 16632 1556
rect 16488 1436 16540 1488
rect 15016 1368 15068 1420
rect 17408 1504 17460 1556
rect 18052 1504 18104 1556
rect 16856 1436 16908 1488
rect 17132 1436 17184 1488
rect 16948 1368 17000 1420
rect 17316 1368 17368 1420
rect 13820 1232 13872 1284
rect 9036 1164 9088 1216
rect 9128 1207 9180 1216
rect 9128 1173 9137 1207
rect 9137 1173 9171 1207
rect 9171 1173 9180 1207
rect 9128 1164 9180 1173
rect 9680 1207 9732 1216
rect 9680 1173 9689 1207
rect 9689 1173 9723 1207
rect 9723 1173 9732 1207
rect 9680 1164 9732 1173
rect 9772 1164 9824 1216
rect 10600 1164 10652 1216
rect 11520 1164 11572 1216
rect 11704 1164 11756 1216
rect 12164 1164 12216 1216
rect 12716 1164 12768 1216
rect 16120 1300 16172 1352
rect 16304 1343 16356 1352
rect 16304 1309 16313 1343
rect 16313 1309 16347 1343
rect 16347 1309 16356 1343
rect 16304 1300 16356 1309
rect 16580 1300 16632 1352
rect 17132 1300 17184 1352
rect 17960 1343 18012 1352
rect 17960 1309 17969 1343
rect 17969 1309 18003 1343
rect 18003 1309 18012 1343
rect 17960 1300 18012 1309
rect 18880 1343 18932 1352
rect 18880 1309 18889 1343
rect 18889 1309 18923 1343
rect 18923 1309 18932 1343
rect 18880 1300 18932 1309
rect 19616 1411 19668 1420
rect 19616 1377 19625 1411
rect 19625 1377 19659 1411
rect 19659 1377 19668 1411
rect 19616 1368 19668 1377
rect 19800 1300 19852 1352
rect 15016 1164 15068 1216
rect 16304 1164 16356 1216
rect 16488 1164 16540 1216
rect 17776 1207 17828 1216
rect 17776 1173 17785 1207
rect 17785 1173 17819 1207
rect 17819 1173 17828 1207
rect 17776 1164 17828 1173
rect 5894 1062 5946 1114
rect 5958 1062 6010 1114
rect 6022 1062 6074 1114
rect 6086 1062 6138 1114
rect 6150 1062 6202 1114
rect 10839 1062 10891 1114
rect 10903 1062 10955 1114
rect 10967 1062 11019 1114
rect 11031 1062 11083 1114
rect 11095 1062 11147 1114
rect 15784 1062 15836 1114
rect 15848 1062 15900 1114
rect 15912 1062 15964 1114
rect 15976 1062 16028 1114
rect 16040 1062 16092 1114
rect 20729 1062 20781 1114
rect 20793 1062 20845 1114
rect 20857 1062 20909 1114
rect 20921 1062 20973 1114
rect 20985 1062 21037 1114
rect 5356 960 5408 1012
rect 7656 960 7708 1012
rect 9312 960 9364 1012
rect 10600 960 10652 1012
rect 11244 960 11296 1012
rect 11520 960 11572 1012
rect 11796 960 11848 1012
rect 14004 960 14056 1012
rect 14464 960 14516 1012
rect 14556 960 14608 1012
rect 14832 960 14884 1012
rect 15016 960 15068 1012
rect 17224 960 17276 1012
rect 18052 960 18104 1012
rect 17776 892 17828 944
rect 10232 824 10284 876
rect 10968 824 11020 876
rect 13268 824 13320 876
rect 10048 756 10100 808
rect 13544 756 13596 808
rect 13912 824 13964 876
rect 14740 756 14792 808
rect 15752 824 15804 876
rect 15844 824 15896 876
rect 4528 688 4580 740
rect 6092 688 6144 740
rect 10232 688 10284 740
rect 1768 620 1820 672
rect 3332 620 3384 672
rect 5264 620 5316 672
rect 6644 620 6696 672
rect 9680 620 9732 672
rect 11060 620 11112 672
rect 12532 688 12584 740
rect 13268 620 13320 672
rect 9128 552 9180 604
rect 10600 552 10652 604
rect 12256 552 12308 604
rect 13728 552 13780 604
rect 13912 688 13964 740
rect 20352 756 20404 808
rect 15384 688 15436 740
rect 15844 688 15896 740
rect 16028 688 16080 740
rect 16580 688 16632 740
rect 16764 688 16816 740
rect 19984 688 20036 740
rect 14280 620 14332 672
rect 20168 620 20220 672
rect 17868 552 17920 604
rect 18696 552 18748 604
rect 11152 484 11204 536
rect 2320 416 2372 468
rect 14280 416 14332 468
rect 14372 416 14424 468
rect 14832 416 14884 468
rect 14924 416 14976 468
rect 15108 416 15160 468
rect 15292 416 15344 468
rect 18236 416 18288 468
rect 11520 348 11572 400
rect 12440 280 12492 332
rect 13728 280 13780 332
rect 14188 348 14240 400
rect 19248 348 19300 400
rect 19432 280 19484 332
rect 13360 212 13412 264
rect 19156 212 19208 264
rect 10416 144 10468 196
rect 21180 144 21232 196
rect 10968 76 11020 128
rect 20444 76 20496 128
rect 5080 8 5132 60
rect 20628 8 20680 60
<< metal2 >>
rect 2410 44540 2466 45000
rect 2594 44540 2650 45000
rect 2778 44540 2834 45000
rect 2962 44540 3018 45000
rect 3146 44540 3202 45000
rect 3330 44540 3386 45000
rect 3514 44540 3570 45000
rect 3698 44540 3754 45000
rect 3882 44540 3938 45000
rect 4066 44540 4122 45000
rect 4250 44540 4306 45000
rect 4434 44540 4490 45000
rect 4618 44540 4674 45000
rect 4802 44540 4858 45000
rect 4986 44540 5042 45000
rect 5170 44540 5226 45000
rect 5354 44540 5410 45000
rect 5538 44540 5594 45000
rect 5722 44540 5778 45000
rect 5906 44540 5962 45000
rect 6090 44540 6146 45000
rect 6274 44540 6330 45000
rect 6458 44540 6514 45000
rect 6642 44540 6698 45000
rect 6826 44540 6882 45000
rect 7010 44540 7066 45000
rect 7194 44540 7250 45000
rect 7378 44540 7434 45000
rect 7562 44540 7618 45000
rect 7746 44540 7802 45000
rect 7930 44540 7986 45000
rect 8114 44540 8170 45000
rect 8298 44540 8354 45000
rect 8482 44540 8538 45000
rect 8666 44540 8722 45000
rect 8850 44540 8906 45000
rect 9034 44540 9090 45000
rect 9218 44540 9274 45000
rect 9402 44540 9458 45000
rect 9586 44540 9642 45000
rect 9770 44540 9826 45000
rect 9954 44540 10010 45000
rect 10138 44540 10194 45000
rect 10322 44540 10378 45000
rect 10506 44540 10562 45000
rect 10690 44540 10746 45000
rect 10874 44540 10930 45000
rect 11058 44540 11114 45000
rect 11242 44540 11298 45000
rect 11426 44540 11482 45000
rect 11610 44540 11666 45000
rect 11794 44540 11850 45000
rect 11978 44540 12034 45000
rect 12162 44540 12218 45000
rect 12346 44540 12402 45000
rect 12530 44540 12586 45000
rect 12714 44540 12770 45000
rect 12898 44540 12954 45000
rect 13082 44540 13138 45000
rect 13266 44540 13322 45000
rect 13450 44540 13506 45000
rect 13634 44540 13690 45000
rect 13818 44540 13874 45000
rect 14002 44540 14058 45000
rect 14186 44540 14242 45000
rect 14370 44540 14426 45000
rect 14554 44540 14610 45000
rect 14738 44540 14794 45000
rect 14922 44540 14978 45000
rect 15106 44540 15162 45000
rect 15290 44540 15346 45000
rect 15382 44568 15438 44577
rect 1308 43852 1360 43858
rect 1308 43794 1360 43800
rect 940 42220 992 42226
rect 940 42162 992 42168
rect 848 42084 900 42090
rect 848 42026 900 42032
rect 20 41676 72 41682
rect 20 41618 72 41624
rect 32 27418 60 41618
rect 202 41576 258 41585
rect 202 41511 258 41520
rect 216 27962 244 41511
rect 480 41472 532 41478
rect 480 41414 532 41420
rect 294 39808 350 39817
rect 294 39743 350 39752
rect 308 28150 336 39743
rect 388 36372 440 36378
rect 388 36314 440 36320
rect 296 28144 348 28150
rect 296 28086 348 28092
rect 294 27976 350 27985
rect 216 27934 294 27962
rect 294 27911 350 27920
rect 294 27432 350 27441
rect 32 27390 294 27418
rect 294 27367 350 27376
rect 400 26840 428 36314
rect 492 32881 520 41414
rect 756 40588 808 40594
rect 756 40530 808 40536
rect 664 36848 716 36854
rect 664 36790 716 36796
rect 478 32872 534 32881
rect 478 32807 534 32816
rect 572 31204 624 31210
rect 572 31146 624 31152
rect 584 29481 612 31146
rect 676 30938 704 36790
rect 768 36174 796 40530
rect 756 36168 808 36174
rect 756 36110 808 36116
rect 756 32904 808 32910
rect 756 32846 808 32852
rect 768 31929 796 32846
rect 754 31920 810 31929
rect 754 31855 810 31864
rect 664 30932 716 30938
rect 664 30874 716 30880
rect 756 30252 808 30258
rect 756 30194 808 30200
rect 570 29472 626 29481
rect 570 29407 626 29416
rect 768 29050 796 30194
rect 676 29022 796 29050
rect 572 28960 624 28966
rect 572 28902 624 28908
rect 216 26812 428 26840
rect 112 22704 164 22710
rect 112 22646 164 22652
rect 20 21412 72 21418
rect 20 21354 72 21360
rect 32 12170 60 21354
rect 124 19334 152 22646
rect 216 20126 244 26812
rect 584 26738 612 28902
rect 308 26710 612 26738
rect 308 20874 336 26710
rect 388 26172 440 26178
rect 388 26114 440 26120
rect 400 21350 428 26114
rect 676 25786 704 29022
rect 754 28928 810 28937
rect 754 28863 810 28872
rect 768 28558 796 28863
rect 756 28552 808 28558
rect 756 28494 808 28500
rect 756 28008 808 28014
rect 756 27950 808 27956
rect 768 26994 796 27950
rect 756 26988 808 26994
rect 756 26930 808 26936
rect 768 26024 796 26930
rect 860 26178 888 42026
rect 952 28422 980 42162
rect 1320 41414 1348 43794
rect 2320 43784 2372 43790
rect 2320 43726 2372 43732
rect 1492 43648 1544 43654
rect 1492 43590 1544 43596
rect 1504 43314 1532 43590
rect 1492 43308 1544 43314
rect 1492 43250 1544 43256
rect 2136 43308 2188 43314
rect 2136 43250 2188 43256
rect 1676 42696 1728 42702
rect 1676 42638 1728 42644
rect 1952 42696 2004 42702
rect 1952 42638 2004 42644
rect 1492 42560 1544 42566
rect 1492 42502 1544 42508
rect 1504 42362 1532 42502
rect 1492 42356 1544 42362
rect 1492 42298 1544 42304
rect 1688 42158 1716 42638
rect 1676 42152 1728 42158
rect 1676 42094 1728 42100
rect 1964 41449 1992 42638
rect 2148 41818 2176 43250
rect 2136 41812 2188 41818
rect 2136 41754 2188 41760
rect 2044 41540 2096 41546
rect 2044 41482 2096 41488
rect 1044 41386 1348 41414
rect 1950 41440 2006 41449
rect 1044 37466 1072 41386
rect 1950 41375 2006 41384
rect 1952 41200 2004 41206
rect 1780 41148 1952 41154
rect 1780 41142 2004 41148
rect 1780 41126 1992 41142
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1308 40112 1360 40118
rect 1228 40060 1308 40066
rect 1228 40054 1360 40060
rect 1228 40038 1348 40054
rect 1124 38344 1176 38350
rect 1228 38321 1256 40038
rect 1308 39976 1360 39982
rect 1308 39918 1360 39924
rect 1320 39273 1348 39918
rect 1412 39681 1440 40462
rect 1398 39672 1454 39681
rect 1398 39607 1454 39616
rect 1400 39432 1452 39438
rect 1400 39374 1452 39380
rect 1306 39264 1362 39273
rect 1306 39199 1362 39208
rect 1124 38286 1176 38292
rect 1214 38312 1270 38321
rect 1032 37460 1084 37466
rect 1032 37402 1084 37408
rect 1136 36689 1164 38286
rect 1214 38247 1270 38256
rect 1412 37913 1440 39374
rect 1492 38956 1544 38962
rect 1492 38898 1544 38904
rect 1398 37904 1454 37913
rect 1398 37839 1454 37848
rect 1400 37732 1452 37738
rect 1400 37674 1452 37680
rect 1216 37188 1268 37194
rect 1216 37130 1268 37136
rect 1228 36825 1256 37130
rect 1308 37120 1360 37126
rect 1306 37088 1308 37097
rect 1360 37088 1362 37097
rect 1306 37023 1362 37032
rect 1214 36816 1270 36825
rect 1214 36751 1270 36760
rect 1216 36712 1268 36718
rect 1122 36680 1178 36689
rect 1216 36654 1268 36660
rect 1122 36615 1178 36624
rect 1032 36168 1084 36174
rect 1032 36110 1084 36116
rect 1044 30161 1072 36110
rect 1228 36009 1256 36654
rect 1308 36644 1360 36650
rect 1308 36586 1360 36592
rect 1320 36281 1348 36586
rect 1306 36272 1362 36281
rect 1306 36207 1362 36216
rect 1214 36000 1270 36009
rect 1214 35935 1270 35944
rect 1412 35873 1440 37674
rect 1504 37369 1532 38898
rect 1584 38412 1636 38418
rect 1584 38354 1636 38360
rect 1490 37360 1546 37369
rect 1596 37330 1624 38354
rect 1676 38276 1728 38282
rect 1676 38218 1728 38224
rect 1490 37295 1546 37304
rect 1584 37324 1636 37330
rect 1584 37266 1636 37272
rect 1492 36780 1544 36786
rect 1492 36722 1544 36728
rect 1398 35864 1454 35873
rect 1398 35799 1454 35808
rect 1400 35760 1452 35766
rect 1214 35728 1270 35737
rect 1270 35708 1400 35714
rect 1270 35702 1452 35708
rect 1270 35686 1440 35702
rect 1214 35663 1270 35672
rect 1400 35624 1452 35630
rect 1400 35566 1452 35572
rect 1412 35154 1440 35566
rect 1124 35148 1176 35154
rect 1124 35090 1176 35096
rect 1400 35148 1452 35154
rect 1400 35090 1452 35096
rect 1136 31890 1164 35090
rect 1504 34785 1532 36722
rect 1596 36258 1624 37266
rect 1688 36825 1716 38218
rect 1780 36854 1808 41126
rect 2056 41120 2084 41482
rect 2332 41414 2360 43726
rect 2424 43450 2452 44540
rect 2412 43444 2464 43450
rect 2412 43386 2464 43392
rect 2504 43308 2556 43314
rect 2504 43250 2556 43256
rect 2516 42362 2544 43250
rect 2608 42362 2636 44540
rect 2792 43450 2820 44540
rect 2780 43444 2832 43450
rect 2780 43386 2832 43392
rect 2976 42702 3004 44540
rect 3056 43308 3108 43314
rect 3056 43250 3108 43256
rect 2964 42696 3016 42702
rect 2964 42638 3016 42644
rect 2688 42628 2740 42634
rect 2688 42570 2740 42576
rect 2504 42356 2556 42362
rect 2504 42298 2556 42304
rect 2596 42356 2648 42362
rect 2596 42298 2648 42304
rect 2700 41818 2728 42570
rect 2964 42560 3016 42566
rect 2964 42502 3016 42508
rect 2872 42152 2924 42158
rect 2872 42094 2924 42100
rect 2688 41812 2740 41818
rect 2688 41754 2740 41760
rect 2504 41608 2556 41614
rect 2504 41550 2556 41556
rect 2516 41414 2544 41550
rect 2332 41386 2452 41414
rect 2516 41386 2728 41414
rect 2424 41290 2452 41386
rect 2424 41262 2636 41290
rect 2056 41092 2544 41120
rect 2136 40928 2188 40934
rect 2136 40870 2188 40876
rect 1952 40452 2004 40458
rect 1952 40394 2004 40400
rect 1964 39409 1992 40394
rect 2044 39976 2096 39982
rect 2044 39918 2096 39924
rect 1950 39400 2006 39409
rect 1950 39335 2006 39344
rect 1952 38956 2004 38962
rect 1952 38898 2004 38904
rect 1860 37868 1912 37874
rect 1860 37810 1912 37816
rect 1768 36848 1820 36854
rect 1674 36816 1730 36825
rect 1768 36790 1820 36796
rect 1674 36751 1730 36760
rect 1596 36230 1716 36258
rect 1584 36168 1636 36174
rect 1584 36110 1636 36116
rect 1490 34776 1546 34785
rect 1490 34711 1546 34720
rect 1216 34604 1268 34610
rect 1216 34546 1268 34552
rect 1228 33153 1256 34546
rect 1492 34400 1544 34406
rect 1492 34342 1544 34348
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1308 33856 1360 33862
rect 1308 33798 1360 33804
rect 1320 33561 1348 33798
rect 1306 33552 1362 33561
rect 1306 33487 1362 33496
rect 1308 33448 1360 33454
rect 1308 33390 1360 33396
rect 1214 33144 1270 33153
rect 1214 33079 1270 33088
rect 1320 32978 1348 33390
rect 1308 32972 1360 32978
rect 1308 32914 1360 32920
rect 1216 32768 1268 32774
rect 1216 32710 1268 32716
rect 1124 31884 1176 31890
rect 1124 31826 1176 31832
rect 1228 31634 1256 32710
rect 1412 32609 1440 33934
rect 1504 32842 1532 34342
rect 1492 32836 1544 32842
rect 1492 32778 1544 32784
rect 1398 32600 1454 32609
rect 1308 32564 1360 32570
rect 1398 32535 1454 32544
rect 1308 32506 1360 32512
rect 1320 32201 1348 32506
rect 1400 32428 1452 32434
rect 1400 32370 1452 32376
rect 1306 32192 1362 32201
rect 1306 32127 1362 32136
rect 1412 31657 1440 32370
rect 1136 31606 1256 31634
rect 1398 31648 1454 31657
rect 1030 30152 1086 30161
rect 1030 30087 1086 30096
rect 1032 29776 1084 29782
rect 1032 29718 1084 29724
rect 1044 29510 1072 29718
rect 1032 29504 1084 29510
rect 1032 29446 1084 29452
rect 1044 29170 1072 29446
rect 1032 29164 1084 29170
rect 1032 29106 1084 29112
rect 1030 28792 1086 28801
rect 1030 28727 1086 28736
rect 940 28416 992 28422
rect 940 28358 992 28364
rect 1044 27878 1072 28727
rect 1032 27872 1084 27878
rect 1032 27814 1084 27820
rect 1136 27690 1164 31606
rect 1398 31583 1454 31592
rect 1398 31104 1454 31113
rect 1398 31039 1454 31048
rect 1308 30660 1360 30666
rect 1308 30602 1360 30608
rect 1214 29744 1270 29753
rect 1214 29679 1270 29688
rect 1228 28626 1256 29679
rect 1320 29306 1348 30602
rect 1412 30326 1440 31039
rect 1400 30320 1452 30326
rect 1400 30262 1452 30268
rect 1400 30048 1452 30054
rect 1400 29990 1452 29996
rect 1308 29300 1360 29306
rect 1308 29242 1360 29248
rect 1306 29064 1362 29073
rect 1306 28999 1362 29008
rect 1216 28620 1268 28626
rect 1216 28562 1268 28568
rect 1320 28506 1348 28999
rect 952 27662 1164 27690
rect 1228 28478 1348 28506
rect 1412 28506 1440 29990
rect 1504 29714 1532 32778
rect 1596 31482 1624 36110
rect 1688 35170 1716 36230
rect 1768 36168 1820 36174
rect 1768 36110 1820 36116
rect 1780 35578 1808 36110
rect 1872 35766 1900 37810
rect 1964 37641 1992 38898
rect 1950 37632 2006 37641
rect 1950 37567 2006 37576
rect 2056 37262 2084 39918
rect 2148 39817 2176 40870
rect 2134 39808 2190 39817
rect 2134 39743 2190 39752
rect 2136 39432 2188 39438
rect 2188 39380 2360 39386
rect 2136 39374 2360 39380
rect 2148 39358 2360 39374
rect 2332 38894 2360 39358
rect 2320 38888 2372 38894
rect 2320 38830 2372 38836
rect 2332 38418 2360 38830
rect 2320 38412 2372 38418
rect 2320 38354 2372 38360
rect 2320 37800 2372 37806
rect 2320 37742 2372 37748
rect 2044 37256 2096 37262
rect 2044 37198 2096 37204
rect 1952 36780 2004 36786
rect 1952 36722 2004 36728
rect 1860 35760 1912 35766
rect 1860 35702 1912 35708
rect 1780 35550 1900 35578
rect 1688 35142 1808 35170
rect 1676 35080 1728 35086
rect 1676 35022 1728 35028
rect 1688 33658 1716 35022
rect 1780 34746 1808 35142
rect 1768 34740 1820 34746
rect 1768 34682 1820 34688
rect 1768 34536 1820 34542
rect 1768 34478 1820 34484
rect 1676 33652 1728 33658
rect 1676 33594 1728 33600
rect 1780 31929 1808 34478
rect 1872 33590 1900 35550
rect 1964 34921 1992 36722
rect 2136 36576 2188 36582
rect 2136 36518 2188 36524
rect 1950 34912 2006 34921
rect 1950 34847 2006 34856
rect 1952 34604 2004 34610
rect 1952 34546 2004 34552
rect 1860 33584 1912 33590
rect 1860 33526 1912 33532
rect 1964 33289 1992 34546
rect 2044 33924 2096 33930
rect 2044 33866 2096 33872
rect 1950 33280 2006 33289
rect 1950 33215 2006 33224
rect 1952 33108 2004 33114
rect 1952 33050 2004 33056
rect 1860 32496 1912 32502
rect 1860 32438 1912 32444
rect 1872 32026 1900 32438
rect 1860 32020 1912 32026
rect 1860 31962 1912 31968
rect 1766 31920 1822 31929
rect 1766 31855 1822 31864
rect 1860 31816 1912 31822
rect 1780 31776 1860 31804
rect 1676 31680 1728 31686
rect 1676 31622 1728 31628
rect 1584 31476 1636 31482
rect 1584 31418 1636 31424
rect 1584 31272 1636 31278
rect 1584 31214 1636 31220
rect 1492 29708 1544 29714
rect 1492 29650 1544 29656
rect 1492 29572 1544 29578
rect 1492 29514 1544 29520
rect 1504 28665 1532 29514
rect 1596 29209 1624 31214
rect 1688 29714 1716 31622
rect 1780 30161 1808 31776
rect 1860 31758 1912 31764
rect 1964 31634 1992 33050
rect 2056 31736 2084 33866
rect 2148 32416 2176 36518
rect 2332 36281 2360 37742
rect 2410 37224 2466 37233
rect 2410 37159 2466 37168
rect 2318 36272 2374 36281
rect 2228 36236 2280 36242
rect 2318 36207 2374 36216
rect 2228 36178 2280 36184
rect 2240 35290 2268 36178
rect 2320 35692 2372 35698
rect 2320 35634 2372 35640
rect 2228 35284 2280 35290
rect 2228 35226 2280 35232
rect 2332 34950 2360 35634
rect 2424 35329 2452 37159
rect 2410 35320 2466 35329
rect 2410 35255 2466 35264
rect 2516 35222 2544 41092
rect 2608 36378 2636 41262
rect 2700 41206 2728 41386
rect 2688 41200 2740 41206
rect 2688 41142 2740 41148
rect 2780 41132 2832 41138
rect 2780 41074 2832 41080
rect 2686 40488 2742 40497
rect 2686 40423 2688 40432
rect 2740 40423 2742 40432
rect 2688 40394 2740 40400
rect 2688 40112 2740 40118
rect 2688 40054 2740 40060
rect 2700 38350 2728 40054
rect 2792 38729 2820 41074
rect 2778 38720 2834 38729
rect 2778 38655 2834 38664
rect 2688 38344 2740 38350
rect 2688 38286 2740 38292
rect 2780 37800 2832 37806
rect 2780 37742 2832 37748
rect 2792 37466 2820 37742
rect 2780 37460 2832 37466
rect 2780 37402 2832 37408
rect 2688 37256 2740 37262
rect 2688 37198 2740 37204
rect 2700 36802 2728 37198
rect 2700 36774 2820 36802
rect 2596 36372 2648 36378
rect 2596 36314 2648 36320
rect 2792 36258 2820 36774
rect 2884 36378 2912 42094
rect 2976 41750 3004 42502
rect 3068 41818 3096 43250
rect 3160 43246 3188 44540
rect 3148 43240 3200 43246
rect 3148 43182 3200 43188
rect 3344 42702 3372 44540
rect 3528 43450 3556 44540
rect 3516 43444 3568 43450
rect 3516 43386 3568 43392
rect 3712 43194 3740 44540
rect 3712 43166 3832 43194
rect 3422 43004 3730 43013
rect 3422 43002 3428 43004
rect 3484 43002 3508 43004
rect 3564 43002 3588 43004
rect 3644 43002 3668 43004
rect 3724 43002 3730 43004
rect 3484 42950 3486 43002
rect 3666 42950 3668 43002
rect 3422 42948 3428 42950
rect 3484 42948 3508 42950
rect 3564 42948 3588 42950
rect 3644 42948 3668 42950
rect 3724 42948 3730 42950
rect 3422 42939 3730 42948
rect 3700 42900 3752 42906
rect 3700 42842 3752 42848
rect 3608 42832 3660 42838
rect 3608 42774 3660 42780
rect 3332 42696 3384 42702
rect 3332 42638 3384 42644
rect 3148 42560 3200 42566
rect 3148 42502 3200 42508
rect 3160 41818 3188 42502
rect 3620 42294 3648 42774
rect 3608 42288 3660 42294
rect 3608 42230 3660 42236
rect 3240 42220 3292 42226
rect 3240 42162 3292 42168
rect 3332 42220 3384 42226
rect 3332 42162 3384 42168
rect 3252 41818 3280 42162
rect 3056 41812 3108 41818
rect 3056 41754 3108 41760
rect 3148 41812 3200 41818
rect 3148 41754 3200 41760
rect 3240 41812 3292 41818
rect 3240 41754 3292 41760
rect 2964 41744 3016 41750
rect 2964 41686 3016 41692
rect 3056 41608 3108 41614
rect 3054 41576 3056 41585
rect 3108 41576 3110 41585
rect 3054 41511 3110 41520
rect 3344 41274 3372 42162
rect 3712 42090 3740 42842
rect 3804 42770 3832 43166
rect 3896 42770 3924 44540
rect 3792 42764 3844 42770
rect 3792 42706 3844 42712
rect 3884 42764 3936 42770
rect 3884 42706 3936 42712
rect 3792 42628 3844 42634
rect 3792 42570 3844 42576
rect 3700 42084 3752 42090
rect 3700 42026 3752 42032
rect 3422 41916 3730 41925
rect 3422 41914 3428 41916
rect 3484 41914 3508 41916
rect 3564 41914 3588 41916
rect 3644 41914 3668 41916
rect 3724 41914 3730 41916
rect 3484 41862 3486 41914
rect 3666 41862 3668 41914
rect 3422 41860 3428 41862
rect 3484 41860 3508 41862
rect 3564 41860 3588 41862
rect 3644 41860 3668 41862
rect 3724 41860 3730 41862
rect 3422 41851 3730 41860
rect 3804 41274 3832 42570
rect 4080 42362 4108 44540
rect 4158 43888 4214 43897
rect 4158 43823 4214 43832
rect 4172 43450 4200 43823
rect 4160 43444 4212 43450
rect 4160 43386 4212 43392
rect 4160 43308 4212 43314
rect 4160 43250 4212 43256
rect 4068 42356 4120 42362
rect 4068 42298 4120 42304
rect 4068 42152 4120 42158
rect 4068 42094 4120 42100
rect 3976 42084 4028 42090
rect 3976 42026 4028 42032
rect 3988 41818 4016 42026
rect 3976 41812 4028 41818
rect 3976 41754 4028 41760
rect 3884 41608 3936 41614
rect 3884 41550 3936 41556
rect 3332 41268 3384 41274
rect 3332 41210 3384 41216
rect 3792 41268 3844 41274
rect 3792 41210 3844 41216
rect 3608 41132 3660 41138
rect 3608 41074 3660 41080
rect 3620 41041 3648 41074
rect 3606 41032 3662 41041
rect 3606 40967 3662 40976
rect 3422 40828 3730 40837
rect 3422 40826 3428 40828
rect 3484 40826 3508 40828
rect 3564 40826 3588 40828
rect 3644 40826 3668 40828
rect 3724 40826 3730 40828
rect 3484 40774 3486 40826
rect 3666 40774 3668 40826
rect 3422 40772 3428 40774
rect 3484 40772 3508 40774
rect 3564 40772 3588 40774
rect 3644 40772 3668 40774
rect 3724 40772 3730 40774
rect 3422 40763 3730 40772
rect 3056 40044 3108 40050
rect 3056 39986 3108 39992
rect 3068 38457 3096 39986
rect 3792 39840 3844 39846
rect 3792 39782 3844 39788
rect 3422 39740 3730 39749
rect 3422 39738 3428 39740
rect 3484 39738 3508 39740
rect 3564 39738 3588 39740
rect 3644 39738 3668 39740
rect 3724 39738 3730 39740
rect 3484 39686 3486 39738
rect 3666 39686 3668 39738
rect 3422 39684 3428 39686
rect 3484 39684 3508 39686
rect 3564 39684 3588 39686
rect 3644 39684 3668 39686
rect 3724 39684 3730 39686
rect 3422 39675 3730 39684
rect 3804 39574 3832 39782
rect 3792 39568 3844 39574
rect 3792 39510 3844 39516
rect 3792 39296 3844 39302
rect 3792 39238 3844 39244
rect 3422 38652 3730 38661
rect 3422 38650 3428 38652
rect 3484 38650 3508 38652
rect 3564 38650 3588 38652
rect 3644 38650 3668 38652
rect 3724 38650 3730 38652
rect 3484 38598 3486 38650
rect 3666 38598 3668 38650
rect 3422 38596 3428 38598
rect 3484 38596 3508 38598
rect 3564 38596 3588 38598
rect 3644 38596 3668 38598
rect 3724 38596 3730 38598
rect 3422 38587 3730 38596
rect 3054 38448 3110 38457
rect 3804 38418 3832 39238
rect 3896 38978 3924 41550
rect 4080 41414 4108 42094
rect 4172 41818 4200 43250
rect 4264 42770 4292 44540
rect 4344 43308 4396 43314
rect 4344 43250 4396 43256
rect 4356 42770 4384 43250
rect 4252 42764 4304 42770
rect 4252 42706 4304 42712
rect 4344 42764 4396 42770
rect 4344 42706 4396 42712
rect 4252 42628 4304 42634
rect 4448 42616 4476 44540
rect 4528 43444 4580 43450
rect 4632 43432 4660 44540
rect 4580 43404 4660 43432
rect 4528 43386 4580 43392
rect 4448 42588 4568 42616
rect 4252 42570 4304 42576
rect 4264 41818 4292 42570
rect 4344 42288 4396 42294
rect 4344 42230 4396 42236
rect 4160 41812 4212 41818
rect 4160 41754 4212 41760
rect 4252 41812 4304 41818
rect 4252 41754 4304 41760
rect 3988 41386 4108 41414
rect 4356 41414 4384 42230
rect 4540 42158 4568 42588
rect 4816 42362 4844 44540
rect 5000 42770 5028 44540
rect 4988 42764 5040 42770
rect 4988 42706 5040 42712
rect 4988 42628 5040 42634
rect 4988 42570 5040 42576
rect 4804 42356 4856 42362
rect 4804 42298 4856 42304
rect 4618 42256 4674 42265
rect 4618 42191 4674 42200
rect 4896 42220 4948 42226
rect 4528 42152 4580 42158
rect 4528 42094 4580 42100
rect 4356 41386 4476 41414
rect 3988 41274 4016 41386
rect 4448 41290 4476 41386
rect 3976 41268 4028 41274
rect 4448 41262 4568 41290
rect 3976 41210 4028 41216
rect 4068 41132 4120 41138
rect 4068 41074 4120 41080
rect 4344 41132 4396 41138
rect 4344 41074 4396 41080
rect 4436 41132 4488 41138
rect 4436 41074 4488 41080
rect 4080 40594 4108 41074
rect 4068 40588 4120 40594
rect 4068 40530 4120 40536
rect 4068 39976 4120 39982
rect 4068 39918 4120 39924
rect 4080 39438 4108 39918
rect 4068 39432 4120 39438
rect 4066 39400 4068 39409
rect 4120 39400 4122 39409
rect 4066 39335 4122 39344
rect 4252 39024 4304 39030
rect 4250 38992 4252 39001
rect 4304 38992 4306 39001
rect 3896 38950 4016 38978
rect 3884 38888 3936 38894
rect 3884 38830 3936 38836
rect 3054 38383 3110 38392
rect 3792 38412 3844 38418
rect 3792 38354 3844 38360
rect 3332 38208 3384 38214
rect 3332 38150 3384 38156
rect 3344 37942 3372 38150
rect 3896 38026 3924 38830
rect 3804 37998 3924 38026
rect 3804 37942 3832 37998
rect 3332 37936 3384 37942
rect 2962 37904 3018 37913
rect 3332 37878 3384 37884
rect 3792 37936 3844 37942
rect 3792 37878 3844 37884
rect 2962 37839 2964 37848
rect 3016 37839 3018 37848
rect 2964 37810 3016 37816
rect 3422 37564 3730 37573
rect 3422 37562 3428 37564
rect 3484 37562 3508 37564
rect 3564 37562 3588 37564
rect 3644 37562 3668 37564
rect 3724 37562 3730 37564
rect 3484 37510 3486 37562
rect 3666 37510 3668 37562
rect 3422 37508 3428 37510
rect 3484 37508 3508 37510
rect 3564 37508 3588 37510
rect 3644 37508 3668 37510
rect 3724 37508 3730 37510
rect 3422 37499 3730 37508
rect 3988 37448 4016 38950
rect 4250 38927 4306 38936
rect 4068 38820 4120 38826
rect 4068 38762 4120 38768
rect 4080 38457 4108 38762
rect 4160 38752 4212 38758
rect 4160 38694 4212 38700
rect 4066 38448 4122 38457
rect 4066 38383 4122 38392
rect 4172 38350 4200 38694
rect 4160 38344 4212 38350
rect 4160 38286 4212 38292
rect 4160 38208 4212 38214
rect 4160 38150 4212 38156
rect 4172 37942 4200 38150
rect 4160 37936 4212 37942
rect 4160 37878 4212 37884
rect 4160 37664 4212 37670
rect 4160 37606 4212 37612
rect 4068 37460 4120 37466
rect 3988 37420 4068 37448
rect 4068 37402 4120 37408
rect 3792 37392 3844 37398
rect 3792 37334 3844 37340
rect 3056 36916 3108 36922
rect 3056 36858 3108 36864
rect 2872 36372 2924 36378
rect 2872 36314 2924 36320
rect 2792 36230 3004 36258
rect 2596 36168 2648 36174
rect 2596 36110 2648 36116
rect 2780 36168 2832 36174
rect 2780 36110 2832 36116
rect 2608 36038 2636 36110
rect 2596 36032 2648 36038
rect 2596 35974 2648 35980
rect 2792 35834 2820 36110
rect 2872 36032 2924 36038
rect 2872 35974 2924 35980
rect 2780 35828 2832 35834
rect 2780 35770 2832 35776
rect 2596 35692 2648 35698
rect 2596 35634 2648 35640
rect 2504 35216 2556 35222
rect 2504 35158 2556 35164
rect 2320 34944 2372 34950
rect 2320 34886 2372 34892
rect 2332 34762 2360 34886
rect 2240 34734 2360 34762
rect 2240 32910 2268 34734
rect 2608 34678 2636 35634
rect 2780 35080 2832 35086
rect 2780 35022 2832 35028
rect 2596 34672 2648 34678
rect 2320 34604 2372 34610
rect 2320 34546 2372 34552
rect 2424 34598 2544 34626
rect 2596 34614 2648 34620
rect 2332 34066 2360 34546
rect 2424 34542 2452 34598
rect 2412 34536 2464 34542
rect 2412 34478 2464 34484
rect 2320 34060 2372 34066
rect 2320 34002 2372 34008
rect 2412 33312 2464 33318
rect 2412 33254 2464 33260
rect 2228 32904 2280 32910
rect 2228 32846 2280 32852
rect 2148 32388 2268 32416
rect 2136 32292 2188 32298
rect 2136 32234 2188 32240
rect 2148 31906 2176 32234
rect 2240 32008 2268 32388
rect 2424 32366 2452 33254
rect 2412 32360 2464 32366
rect 2412 32302 2464 32308
rect 2240 31980 2452 32008
rect 2148 31878 2360 31906
rect 2226 31784 2282 31793
rect 2136 31748 2188 31754
rect 2056 31708 2136 31736
rect 2226 31719 2282 31728
rect 2136 31690 2188 31696
rect 1964 31606 2084 31634
rect 1950 31512 2006 31521
rect 1950 31447 2006 31456
rect 1964 31346 1992 31447
rect 1952 31340 2004 31346
rect 1952 31282 2004 31288
rect 1860 30864 1912 30870
rect 1860 30806 1912 30812
rect 1872 30705 1900 30806
rect 1858 30696 1914 30705
rect 1858 30631 1914 30640
rect 1766 30152 1822 30161
rect 1766 30087 1822 30096
rect 1768 30048 1820 30054
rect 1768 29990 1820 29996
rect 1676 29708 1728 29714
rect 1676 29650 1728 29656
rect 1674 29608 1730 29617
rect 1674 29543 1676 29552
rect 1728 29543 1730 29552
rect 1676 29514 1728 29520
rect 1582 29200 1638 29209
rect 1582 29135 1638 29144
rect 1490 28656 1546 28665
rect 1674 28656 1730 28665
rect 1490 28591 1546 28600
rect 1596 28614 1674 28642
rect 1412 28478 1532 28506
rect 848 26172 900 26178
rect 848 26114 900 26120
rect 768 25996 888 26024
rect 756 25900 808 25906
rect 756 25842 808 25848
rect 492 25758 704 25786
rect 388 21344 440 21350
rect 388 21286 440 21292
rect 296 20868 348 20874
rect 296 20810 348 20816
rect 204 20120 256 20126
rect 204 20062 256 20068
rect 124 19306 336 19334
rect 204 16516 256 16522
rect 204 16458 256 16464
rect 112 13864 164 13870
rect 112 13806 164 13812
rect 20 12164 72 12170
rect 20 12106 72 12112
rect 32 11422 60 12106
rect 20 11416 72 11422
rect 20 11358 72 11364
rect 20 10736 72 10742
rect 20 10678 72 10684
rect 32 1358 60 10678
rect 124 9586 152 13806
rect 216 13326 244 16458
rect 308 15201 336 19306
rect 386 19000 442 19009
rect 386 18935 442 18944
rect 294 15192 350 15201
rect 294 15127 350 15136
rect 294 13832 350 13841
rect 294 13767 350 13776
rect 204 13320 256 13326
rect 204 13262 256 13268
rect 112 9580 164 9586
rect 112 9522 164 9528
rect 124 6322 152 9522
rect 308 7614 336 13767
rect 296 7608 348 7614
rect 296 7550 348 7556
rect 112 6316 164 6322
rect 112 6258 164 6264
rect 20 1352 72 1358
rect 20 1294 72 1300
rect 400 785 428 18935
rect 492 14929 520 25758
rect 664 25288 716 25294
rect 664 25230 716 25236
rect 676 24041 704 25230
rect 768 24857 796 25842
rect 754 24848 810 24857
rect 754 24783 810 24792
rect 860 24274 888 25996
rect 848 24268 900 24274
rect 848 24210 900 24216
rect 662 24032 718 24041
rect 662 23967 718 23976
rect 952 23882 980 27662
rect 1032 27600 1084 27606
rect 1032 27542 1084 27548
rect 584 23854 980 23882
rect 478 14920 534 14929
rect 478 14855 534 14864
rect 480 14816 532 14822
rect 480 14758 532 14764
rect 492 11506 520 14758
rect 584 14521 612 23854
rect 756 23724 808 23730
rect 756 23666 808 23672
rect 768 23497 796 23666
rect 754 23488 810 23497
rect 754 23423 810 23432
rect 756 23112 808 23118
rect 756 23054 808 23060
rect 768 22953 796 23054
rect 940 23044 992 23050
rect 940 22986 992 22992
rect 754 22944 810 22953
rect 754 22879 810 22888
rect 756 22636 808 22642
rect 756 22578 808 22584
rect 768 22409 796 22578
rect 754 22400 810 22409
rect 754 22335 810 22344
rect 848 22024 900 22030
rect 848 21966 900 21972
rect 860 21865 888 21966
rect 846 21856 902 21865
rect 846 21791 902 21800
rect 952 21593 980 22986
rect 1044 22778 1072 27542
rect 1124 27396 1176 27402
rect 1124 27338 1176 27344
rect 1136 27033 1164 27338
rect 1122 27024 1178 27033
rect 1122 26959 1178 26968
rect 1228 26874 1256 28478
rect 1400 28212 1452 28218
rect 1400 28154 1452 28160
rect 1308 28144 1360 28150
rect 1308 28086 1360 28092
rect 1320 27849 1348 28086
rect 1412 28014 1440 28154
rect 1400 28008 1452 28014
rect 1400 27950 1452 27956
rect 1306 27840 1362 27849
rect 1306 27775 1362 27784
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 1320 27062 1348 27231
rect 1308 27056 1360 27062
rect 1308 26998 1360 27004
rect 1136 26846 1256 26874
rect 1136 25673 1164 26846
rect 1216 26784 1268 26790
rect 1216 26726 1268 26732
rect 1306 26752 1362 26761
rect 1228 26489 1256 26726
rect 1306 26687 1362 26696
rect 1320 26586 1348 26687
rect 1308 26580 1360 26586
rect 1308 26522 1360 26528
rect 1214 26480 1270 26489
rect 1214 26415 1270 26424
rect 1308 26376 1360 26382
rect 1214 26344 1270 26353
rect 1308 26318 1360 26324
rect 1214 26279 1270 26288
rect 1122 25664 1178 25673
rect 1122 25599 1178 25608
rect 1122 25528 1178 25537
rect 1122 25463 1178 25472
rect 1032 22772 1084 22778
rect 1032 22714 1084 22720
rect 1136 22094 1164 25463
rect 1228 25401 1256 26279
rect 1214 25392 1270 25401
rect 1320 25362 1348 26318
rect 1412 25809 1440 27406
rect 1398 25800 1454 25809
rect 1398 25735 1454 25744
rect 1504 25537 1532 28478
rect 1596 28370 1624 28614
rect 1674 28591 1730 28600
rect 1674 28520 1730 28529
rect 1674 28455 1676 28464
rect 1728 28455 1730 28464
rect 1676 28426 1728 28432
rect 1596 28342 1716 28370
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1596 26246 1624 27270
rect 1584 26240 1636 26246
rect 1584 26182 1636 26188
rect 1688 26042 1716 28342
rect 1780 26489 1808 29990
rect 1766 26480 1822 26489
rect 1766 26415 1822 26424
rect 1780 26382 1808 26415
rect 1768 26376 1820 26382
rect 1768 26318 1820 26324
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 1872 25820 1900 30631
rect 1964 27520 1992 31282
rect 2056 29238 2084 31606
rect 2044 29232 2096 29238
rect 2044 29174 2096 29180
rect 2044 29130 2096 29136
rect 2044 29072 2096 29078
rect 2056 28218 2084 29072
rect 2044 28212 2096 28218
rect 2044 28154 2096 28160
rect 2044 28076 2096 28082
rect 2044 28018 2096 28024
rect 2056 27713 2084 28018
rect 2042 27704 2098 27713
rect 2042 27639 2098 27648
rect 1964 27492 2084 27520
rect 1952 27396 2004 27402
rect 1952 27338 2004 27344
rect 1964 26081 1992 27338
rect 2056 26908 2084 27492
rect 2148 26976 2176 31690
rect 2240 31686 2268 31719
rect 2228 31680 2280 31686
rect 2228 31622 2280 31628
rect 2240 31346 2268 31622
rect 2228 31340 2280 31346
rect 2228 31282 2280 31288
rect 2228 30184 2280 30190
rect 2228 30126 2280 30132
rect 2240 29850 2268 30126
rect 2228 29844 2280 29850
rect 2228 29786 2280 29792
rect 2228 29572 2280 29578
rect 2228 29514 2280 29520
rect 2240 27985 2268 29514
rect 2226 27976 2282 27985
rect 2332 27962 2360 31878
rect 2424 31346 2452 31980
rect 2412 31340 2464 31346
rect 2412 31282 2464 31288
rect 2516 31249 2544 34598
rect 2792 33833 2820 35022
rect 2778 33824 2834 33833
rect 2778 33759 2834 33768
rect 2884 33674 2912 35974
rect 2608 33646 2912 33674
rect 2608 32609 2636 33646
rect 2780 33516 2832 33522
rect 2780 33458 2832 33464
rect 2688 32836 2740 32842
rect 2688 32778 2740 32784
rect 2594 32600 2650 32609
rect 2594 32535 2650 32544
rect 2596 31952 2648 31958
rect 2596 31894 2648 31900
rect 2502 31240 2558 31249
rect 2502 31175 2558 31184
rect 2412 31136 2464 31142
rect 2412 31078 2464 31084
rect 2424 29073 2452 31078
rect 2608 30802 2636 31894
rect 2700 31754 2728 32778
rect 2792 32745 2820 33458
rect 2976 32978 3004 36230
rect 3068 34678 3096 36858
rect 3332 36712 3384 36718
rect 3332 36654 3384 36660
rect 3240 36576 3292 36582
rect 3240 36518 3292 36524
rect 3148 35692 3200 35698
rect 3148 35634 3200 35640
rect 3160 35154 3188 35634
rect 3148 35148 3200 35154
rect 3148 35090 3200 35096
rect 3056 34672 3108 34678
rect 3056 34614 3108 34620
rect 3068 33114 3096 34614
rect 3252 33998 3280 36518
rect 3344 35494 3372 36654
rect 3422 36476 3730 36485
rect 3422 36474 3428 36476
rect 3484 36474 3508 36476
rect 3564 36474 3588 36476
rect 3644 36474 3668 36476
rect 3724 36474 3730 36476
rect 3484 36422 3486 36474
rect 3666 36422 3668 36474
rect 3422 36420 3428 36422
rect 3484 36420 3508 36422
rect 3564 36420 3588 36422
rect 3644 36420 3668 36422
rect 3724 36420 3730 36422
rect 3422 36411 3730 36420
rect 3804 36038 3832 37334
rect 4068 37324 4120 37330
rect 4068 37266 4120 37272
rect 3884 36236 3936 36242
rect 3884 36178 3936 36184
rect 3792 36032 3844 36038
rect 3792 35974 3844 35980
rect 3896 35834 3924 36178
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 3884 35828 3936 35834
rect 3884 35770 3936 35776
rect 3332 35488 3384 35494
rect 3332 35430 3384 35436
rect 3422 35388 3730 35397
rect 3422 35386 3428 35388
rect 3484 35386 3508 35388
rect 3564 35386 3588 35388
rect 3644 35386 3668 35388
rect 3724 35386 3730 35388
rect 3484 35334 3486 35386
rect 3666 35334 3668 35386
rect 3422 35332 3428 35334
rect 3484 35332 3508 35334
rect 3564 35332 3588 35334
rect 3644 35332 3668 35334
rect 3724 35332 3730 35334
rect 3422 35323 3730 35332
rect 3792 35080 3844 35086
rect 3792 35022 3844 35028
rect 3424 34740 3476 34746
rect 3424 34682 3476 34688
rect 3332 34604 3384 34610
rect 3332 34546 3384 34552
rect 3344 34105 3372 34546
rect 3436 34406 3464 34682
rect 3804 34513 3832 35022
rect 3790 34504 3846 34513
rect 3790 34439 3846 34448
rect 3424 34400 3476 34406
rect 3424 34342 3476 34348
rect 3884 34400 3936 34406
rect 3884 34342 3936 34348
rect 3422 34300 3730 34309
rect 3422 34298 3428 34300
rect 3484 34298 3508 34300
rect 3564 34298 3588 34300
rect 3644 34298 3668 34300
rect 3724 34298 3730 34300
rect 3484 34246 3486 34298
rect 3666 34246 3668 34298
rect 3422 34244 3428 34246
rect 3484 34244 3508 34246
rect 3564 34244 3588 34246
rect 3644 34244 3668 34246
rect 3724 34244 3730 34246
rect 3422 34235 3730 34244
rect 3330 34096 3386 34105
rect 3330 34031 3386 34040
rect 3240 33992 3292 33998
rect 3240 33934 3292 33940
rect 3332 33856 3384 33862
rect 3332 33798 3384 33804
rect 3344 33658 3372 33798
rect 3332 33652 3384 33658
rect 3332 33594 3384 33600
rect 3240 33584 3292 33590
rect 3700 33584 3752 33590
rect 3698 33552 3700 33561
rect 3752 33552 3754 33561
rect 3292 33532 3372 33538
rect 3240 33526 3372 33532
rect 3252 33510 3372 33526
rect 3056 33108 3108 33114
rect 3056 33050 3108 33056
rect 2964 32972 3016 32978
rect 2964 32914 3016 32920
rect 2872 32904 2924 32910
rect 2872 32846 2924 32852
rect 2778 32736 2834 32745
rect 2778 32671 2834 32680
rect 2778 32600 2834 32609
rect 2778 32535 2834 32544
rect 2792 32434 2820 32535
rect 2780 32428 2832 32434
rect 2780 32370 2832 32376
rect 2700 31726 2820 31754
rect 2688 31680 2740 31686
rect 2688 31622 2740 31628
rect 2596 30796 2648 30802
rect 2596 30738 2648 30744
rect 2504 30728 2556 30734
rect 2504 30670 2556 30676
rect 2516 30433 2544 30670
rect 2502 30424 2558 30433
rect 2502 30359 2558 30368
rect 2410 29064 2466 29073
rect 2410 28999 2466 29008
rect 2516 28966 2544 30359
rect 2608 30122 2636 30738
rect 2700 30716 2728 31622
rect 2792 30954 2820 31726
rect 2884 31113 2912 32846
rect 3344 32842 3372 33510
rect 3698 33487 3754 33496
rect 3896 33454 3924 34342
rect 3988 33590 4016 36110
rect 4080 35601 4108 37266
rect 4172 36650 4200 37606
rect 4264 37262 4292 38927
rect 4252 37256 4304 37262
rect 4252 37198 4304 37204
rect 4252 36780 4304 36786
rect 4252 36722 4304 36728
rect 4160 36644 4212 36650
rect 4160 36586 4212 36592
rect 4172 36310 4200 36586
rect 4160 36304 4212 36310
rect 4160 36246 4212 36252
rect 4160 36032 4212 36038
rect 4158 36000 4160 36009
rect 4212 36000 4214 36009
rect 4158 35935 4214 35944
rect 4160 35624 4212 35630
rect 4066 35592 4122 35601
rect 4160 35566 4212 35572
rect 4066 35527 4122 35536
rect 4068 35012 4120 35018
rect 4068 34954 4120 34960
rect 4080 34105 4108 34954
rect 4066 34096 4122 34105
rect 4066 34031 4122 34040
rect 4172 33980 4200 35566
rect 4264 35193 4292 36722
rect 4250 35184 4306 35193
rect 4250 35119 4306 35128
rect 4080 33952 4200 33980
rect 4252 33992 4304 33998
rect 3976 33584 4028 33590
rect 3976 33526 4028 33532
rect 3884 33448 3936 33454
rect 3884 33390 3936 33396
rect 3422 33212 3730 33221
rect 3422 33210 3428 33212
rect 3484 33210 3508 33212
rect 3564 33210 3588 33212
rect 3644 33210 3668 33212
rect 3724 33210 3730 33212
rect 3484 33158 3486 33210
rect 3666 33158 3668 33210
rect 3422 33156 3428 33158
rect 3484 33156 3508 33158
rect 3564 33156 3588 33158
rect 3644 33156 3668 33158
rect 3724 33156 3730 33158
rect 3422 33147 3730 33156
rect 3882 32872 3938 32881
rect 3332 32836 3384 32842
rect 3882 32807 3884 32816
rect 3332 32778 3384 32784
rect 3936 32807 3938 32816
rect 3884 32778 3936 32784
rect 3056 32768 3108 32774
rect 3056 32710 3108 32716
rect 3068 32502 3096 32710
rect 3344 32502 3372 32778
rect 3056 32496 3108 32502
rect 3056 32438 3108 32444
rect 3332 32496 3384 32502
rect 3332 32438 3384 32444
rect 2964 32428 3016 32434
rect 2964 32370 3016 32376
rect 3884 32428 3936 32434
rect 3884 32370 3936 32376
rect 2976 31385 3004 32370
rect 3514 32328 3570 32337
rect 3514 32263 3516 32272
rect 3568 32263 3570 32272
rect 3516 32234 3568 32240
rect 3422 32124 3730 32133
rect 3422 32122 3428 32124
rect 3484 32122 3508 32124
rect 3564 32122 3588 32124
rect 3644 32122 3668 32124
rect 3724 32122 3730 32124
rect 3484 32070 3486 32122
rect 3666 32070 3668 32122
rect 3422 32068 3428 32070
rect 3484 32068 3508 32070
rect 3564 32068 3588 32070
rect 3644 32068 3668 32070
rect 3724 32068 3730 32070
rect 3422 32059 3730 32068
rect 3056 31816 3108 31822
rect 3056 31758 3108 31764
rect 3068 31414 3096 31758
rect 3608 31748 3660 31754
rect 3608 31690 3660 31696
rect 3792 31748 3844 31754
rect 3792 31690 3844 31696
rect 3056 31408 3108 31414
rect 2962 31376 3018 31385
rect 3056 31350 3108 31356
rect 2962 31311 3018 31320
rect 3332 31340 3384 31346
rect 3332 31282 3384 31288
rect 3240 31136 3292 31142
rect 2870 31104 2926 31113
rect 3240 31078 3292 31084
rect 2870 31039 2926 31048
rect 2792 30926 2912 30954
rect 2780 30728 2832 30734
rect 2700 30688 2780 30716
rect 2780 30670 2832 30676
rect 2778 30560 2834 30569
rect 2778 30495 2834 30504
rect 2596 30116 2648 30122
rect 2596 30058 2648 30064
rect 2688 30116 2740 30122
rect 2688 30058 2740 30064
rect 2700 29850 2728 30058
rect 2792 29889 2820 30495
rect 2778 29880 2834 29889
rect 2688 29844 2740 29850
rect 2778 29815 2834 29824
rect 2688 29786 2740 29792
rect 2780 29640 2832 29646
rect 2780 29582 2832 29588
rect 2596 29504 2648 29510
rect 2596 29446 2648 29452
rect 2608 29170 2636 29446
rect 2792 29345 2820 29582
rect 2778 29336 2834 29345
rect 2778 29271 2834 29280
rect 2884 29322 2912 30926
rect 2978 30252 3030 30258
rect 2978 30194 3030 30200
rect 2990 30138 3018 30194
rect 3252 30190 3280 31078
rect 2976 30110 3018 30138
rect 3222 30184 3280 30190
rect 3274 30144 3280 30184
rect 3222 30126 3274 30132
rect 2976 29481 3004 30110
rect 3344 29832 3372 31282
rect 3620 31142 3648 31690
rect 3804 31657 3832 31690
rect 3790 31648 3846 31657
rect 3790 31583 3846 31592
rect 3608 31136 3660 31142
rect 3608 31078 3660 31084
rect 3422 31036 3730 31045
rect 3422 31034 3428 31036
rect 3484 31034 3508 31036
rect 3564 31034 3588 31036
rect 3644 31034 3668 31036
rect 3724 31034 3730 31036
rect 3484 30982 3486 31034
rect 3666 30982 3668 31034
rect 3422 30980 3428 30982
rect 3484 30980 3508 30982
rect 3564 30980 3588 30982
rect 3644 30980 3668 30982
rect 3724 30980 3730 30982
rect 3422 30971 3730 30980
rect 3606 30832 3662 30841
rect 3606 30767 3662 30776
rect 3424 30728 3476 30734
rect 3424 30670 3476 30676
rect 3436 30297 3464 30670
rect 3620 30598 3648 30767
rect 3608 30592 3660 30598
rect 3608 30534 3660 30540
rect 3792 30592 3844 30598
rect 3792 30534 3844 30540
rect 3422 30288 3478 30297
rect 3422 30223 3478 30232
rect 3422 29948 3730 29957
rect 3422 29946 3428 29948
rect 3484 29946 3508 29948
rect 3564 29946 3588 29948
rect 3644 29946 3668 29948
rect 3724 29946 3730 29948
rect 3484 29894 3486 29946
rect 3666 29894 3668 29946
rect 3422 29892 3428 29894
rect 3484 29892 3508 29894
rect 3564 29892 3588 29894
rect 3644 29892 3668 29894
rect 3724 29892 3730 29894
rect 3422 29883 3730 29892
rect 3344 29804 3464 29832
rect 3330 29744 3386 29753
rect 3330 29679 3386 29688
rect 3344 29646 3372 29679
rect 3148 29640 3200 29646
rect 3148 29582 3200 29588
rect 3332 29640 3384 29646
rect 3332 29582 3384 29588
rect 2962 29472 3018 29481
rect 2962 29407 3018 29416
rect 2884 29294 3096 29322
rect 2596 29164 2648 29170
rect 2596 29106 2648 29112
rect 2504 28960 2556 28966
rect 2504 28902 2556 28908
rect 2594 28656 2650 28665
rect 2594 28591 2596 28600
rect 2648 28591 2650 28600
rect 2596 28562 2648 28568
rect 2596 28416 2648 28422
rect 2596 28358 2648 28364
rect 2410 28248 2466 28257
rect 2410 28183 2412 28192
rect 2464 28183 2466 28192
rect 2412 28154 2464 28160
rect 2332 27934 2544 27962
rect 2226 27911 2282 27920
rect 2412 27872 2464 27878
rect 2412 27814 2464 27820
rect 2424 27538 2452 27814
rect 2412 27532 2464 27538
rect 2412 27474 2464 27480
rect 2228 27396 2280 27402
rect 2228 27338 2280 27344
rect 2320 27396 2372 27402
rect 2320 27338 2372 27344
rect 2240 27130 2268 27338
rect 2228 27124 2280 27130
rect 2228 27066 2280 27072
rect 2148 26948 2268 26976
rect 2056 26880 2176 26908
rect 2044 26240 2096 26246
rect 2044 26182 2096 26188
rect 1950 26072 2006 26081
rect 1950 26007 2006 26016
rect 1964 25974 1992 26007
rect 1952 25968 2004 25974
rect 1952 25910 2004 25916
rect 1872 25792 1992 25820
rect 1490 25528 1546 25537
rect 1490 25463 1546 25472
rect 1214 25327 1270 25336
rect 1308 25356 1360 25362
rect 1308 25298 1360 25304
rect 1768 25288 1820 25294
rect 1768 25230 1820 25236
rect 1858 25256 1914 25265
rect 1308 25220 1360 25226
rect 1308 25162 1360 25168
rect 1320 25129 1348 25162
rect 1306 25120 1362 25129
rect 1306 25055 1362 25064
rect 1780 24954 1808 25230
rect 1858 25191 1914 25200
rect 1768 24948 1820 24954
rect 1768 24890 1820 24896
rect 1216 24812 1268 24818
rect 1216 24754 1268 24760
rect 1228 24313 1256 24754
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1308 24676 1360 24682
rect 1308 24618 1360 24624
rect 1320 24585 1348 24618
rect 1306 24576 1362 24585
rect 1306 24511 1362 24520
rect 1214 24304 1270 24313
rect 1214 24239 1270 24248
rect 1308 24132 1360 24138
rect 1308 24074 1360 24080
rect 1320 23769 1348 24074
rect 1306 23760 1362 23769
rect 1306 23695 1362 23704
rect 1306 23624 1362 23633
rect 1306 23559 1362 23568
rect 1320 22710 1348 23559
rect 1308 22704 1360 22710
rect 1412 22681 1440 24686
rect 1492 24268 1544 24274
rect 1544 24228 1624 24256
rect 1492 24210 1544 24216
rect 1490 23488 1546 23497
rect 1490 23423 1546 23432
rect 1308 22646 1360 22652
rect 1398 22672 1454 22681
rect 1398 22607 1454 22616
rect 1398 22128 1454 22137
rect 1136 22066 1348 22094
rect 1214 21992 1270 22001
rect 1214 21927 1270 21936
rect 1032 21888 1084 21894
rect 1032 21830 1084 21836
rect 938 21584 994 21593
rect 938 21519 994 21528
rect 1044 21468 1072 21830
rect 1122 21584 1178 21593
rect 1122 21519 1178 21528
rect 860 21440 1072 21468
rect 754 20496 810 20505
rect 754 20431 810 20440
rect 768 19446 796 20431
rect 756 19440 808 19446
rect 756 19382 808 19388
rect 860 18952 888 21440
rect 1032 21344 1084 21350
rect 1032 21286 1084 21292
rect 938 21176 994 21185
rect 938 21111 994 21120
rect 676 18924 888 18952
rect 676 16522 704 18924
rect 754 18864 810 18873
rect 754 18799 810 18808
rect 768 18766 796 18799
rect 756 18760 808 18766
rect 756 18702 808 18708
rect 754 18592 810 18601
rect 754 18527 810 18536
rect 768 18358 796 18527
rect 756 18352 808 18358
rect 756 18294 808 18300
rect 754 18184 810 18193
rect 754 18119 810 18128
rect 768 16561 796 18119
rect 848 17740 900 17746
rect 848 17682 900 17688
rect 754 16552 810 16561
rect 664 16516 716 16522
rect 754 16487 810 16496
rect 664 16458 716 16464
rect 662 16416 718 16425
rect 662 16351 718 16360
rect 676 14618 704 16351
rect 860 16266 888 17682
rect 768 16238 888 16266
rect 664 14612 716 14618
rect 664 14554 716 14560
rect 570 14512 626 14521
rect 570 14447 626 14456
rect 664 14476 716 14482
rect 664 14418 716 14424
rect 676 11676 704 14418
rect 768 11778 796 16238
rect 846 16144 902 16153
rect 846 16079 902 16088
rect 860 15162 888 16079
rect 848 15156 900 15162
rect 848 15098 900 15104
rect 846 14784 902 14793
rect 846 14719 902 14728
rect 860 11898 888 14719
rect 952 14498 980 21111
rect 1044 17954 1072 21286
rect 1136 21049 1164 21519
rect 1228 21418 1256 21927
rect 1216 21412 1268 21418
rect 1216 21354 1268 21360
rect 1122 21040 1178 21049
rect 1122 20975 1178 20984
rect 1124 20868 1176 20874
rect 1124 20810 1176 20816
rect 1136 18193 1164 20810
rect 1214 19408 1270 19417
rect 1320 19394 1348 22066
rect 1398 22063 1454 22072
rect 1412 19922 1440 22063
rect 1400 19916 1452 19922
rect 1400 19858 1452 19864
rect 1320 19366 1440 19394
rect 1214 19343 1270 19352
rect 1228 18834 1256 19343
rect 1308 19168 1360 19174
rect 1308 19110 1360 19116
rect 1216 18828 1268 18834
rect 1216 18770 1268 18776
rect 1216 18692 1268 18698
rect 1216 18634 1268 18640
rect 1228 18329 1256 18634
rect 1320 18426 1348 19110
rect 1308 18420 1360 18426
rect 1308 18362 1360 18368
rect 1214 18320 1270 18329
rect 1214 18255 1270 18264
rect 1122 18184 1178 18193
rect 1122 18119 1178 18128
rect 1044 17926 1256 17954
rect 1124 16720 1176 16726
rect 1124 16662 1176 16668
rect 1136 14822 1164 16662
rect 1124 14816 1176 14822
rect 1124 14758 1176 14764
rect 952 14470 1164 14498
rect 938 14376 994 14385
rect 938 14311 994 14320
rect 952 12442 980 14311
rect 940 12436 992 12442
rect 940 12378 992 12384
rect 848 11892 900 11898
rect 848 11834 900 11840
rect 1032 11824 1084 11830
rect 768 11750 980 11778
rect 1032 11766 1084 11772
rect 676 11648 888 11676
rect 492 11478 704 11506
rect 572 11416 624 11422
rect 572 11358 624 11364
rect 480 11280 532 11286
rect 480 11222 532 11228
rect 492 6798 520 11222
rect 584 8362 612 11358
rect 572 8356 624 8362
rect 572 8298 624 8304
rect 676 7698 704 11478
rect 860 11054 888 11648
rect 768 11026 888 11054
rect 768 8106 796 11026
rect 846 10976 902 10985
rect 846 10911 902 10920
rect 860 8401 888 10911
rect 846 8392 902 8401
rect 846 8327 902 8336
rect 846 8120 902 8129
rect 768 8078 846 8106
rect 846 8055 902 8064
rect 584 7670 704 7698
rect 584 7313 612 7670
rect 664 7608 716 7614
rect 952 7562 980 11750
rect 1044 10810 1072 11766
rect 1032 10804 1084 10810
rect 1032 10746 1084 10752
rect 1030 10704 1086 10713
rect 1030 10639 1086 10648
rect 1044 8294 1072 10639
rect 1032 8288 1084 8294
rect 1032 8230 1084 8236
rect 664 7550 716 7556
rect 570 7304 626 7313
rect 570 7239 626 7248
rect 480 6792 532 6798
rect 480 6734 532 6740
rect 570 6624 626 6633
rect 570 6559 626 6568
rect 584 4622 612 6559
rect 572 4616 624 4622
rect 572 4558 624 4564
rect 676 2854 704 7550
rect 756 7540 808 7546
rect 756 7482 808 7488
rect 860 7534 980 7562
rect 1030 7576 1086 7585
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 478 2680 534 2689
rect 478 2615 534 2624
rect 492 1494 520 2615
rect 768 1902 796 7482
rect 860 2009 888 7534
rect 1136 7546 1164 14470
rect 1228 14362 1256 17926
rect 1308 17808 1360 17814
rect 1308 17750 1360 17756
rect 1320 14482 1348 17750
rect 1412 14521 1440 19366
rect 1504 18465 1532 23423
rect 1596 22982 1624 24228
rect 1766 24032 1822 24041
rect 1766 23967 1822 23976
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1688 23225 1716 23666
rect 1674 23216 1730 23225
rect 1674 23151 1730 23160
rect 1584 22976 1636 22982
rect 1584 22918 1636 22924
rect 1676 22772 1728 22778
rect 1676 22714 1728 22720
rect 1582 22672 1638 22681
rect 1582 22607 1638 22616
rect 1596 22438 1624 22607
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1584 21684 1636 21690
rect 1584 21626 1636 21632
rect 1596 20602 1624 21626
rect 1688 21554 1716 22714
rect 1676 21548 1728 21554
rect 1676 21490 1728 21496
rect 1674 21040 1730 21049
rect 1674 20975 1730 20984
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1596 18902 1624 20538
rect 1688 19922 1716 20975
rect 1676 19916 1728 19922
rect 1676 19858 1728 19864
rect 1674 19272 1730 19281
rect 1674 19207 1730 19216
rect 1584 18896 1636 18902
rect 1584 18838 1636 18844
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1582 18320 1638 18329
rect 1582 18255 1638 18264
rect 1490 18048 1546 18057
rect 1490 17983 1546 17992
rect 1504 17678 1532 17983
rect 1596 17746 1624 18255
rect 1688 17882 1716 19207
rect 1780 19009 1808 23967
rect 1872 23594 1900 25191
rect 1860 23588 1912 23594
rect 1860 23530 1912 23536
rect 1964 23254 1992 25792
rect 1952 23248 2004 23254
rect 1952 23190 2004 23196
rect 1952 22976 2004 22982
rect 1952 22918 2004 22924
rect 1964 22098 1992 22918
rect 1952 22092 2004 22098
rect 1952 22034 2004 22040
rect 1964 21622 1992 22034
rect 2056 21690 2084 26182
rect 2148 25378 2176 26880
rect 2240 26246 2268 26948
rect 2228 26240 2280 26246
rect 2228 26182 2280 26188
rect 2332 26042 2360 27338
rect 2410 27160 2466 27169
rect 2410 27095 2466 27104
rect 2424 26994 2452 27095
rect 2412 26988 2464 26994
rect 2412 26930 2464 26936
rect 2516 26330 2544 27934
rect 2424 26302 2544 26330
rect 2320 26036 2372 26042
rect 2320 25978 2372 25984
rect 2228 25968 2280 25974
rect 2228 25910 2280 25916
rect 2240 25498 2268 25910
rect 2228 25492 2280 25498
rect 2228 25434 2280 25440
rect 2148 25350 2268 25378
rect 2136 25288 2188 25294
rect 2136 25230 2188 25236
rect 2148 24993 2176 25230
rect 2134 24984 2190 24993
rect 2134 24919 2190 24928
rect 2240 24868 2268 25350
rect 2148 24840 2268 24868
rect 2148 23798 2176 24840
rect 2228 24200 2280 24206
rect 2228 24142 2280 24148
rect 2136 23792 2188 23798
rect 2134 23760 2136 23769
rect 2188 23760 2190 23769
rect 2134 23695 2190 23704
rect 2240 23644 2268 24142
rect 2148 23616 2268 23644
rect 2148 22420 2176 23616
rect 2332 23322 2360 25978
rect 2424 25294 2452 26302
rect 2608 26246 2636 28358
rect 2792 26432 2820 29271
rect 2884 29170 2912 29294
rect 2964 29232 3016 29238
rect 2964 29174 3016 29180
rect 2872 29164 2924 29170
rect 2872 29106 2924 29112
rect 2872 28960 2924 28966
rect 2872 28902 2924 28908
rect 2700 26404 2820 26432
rect 2504 26240 2556 26246
rect 2504 26182 2556 26188
rect 2596 26240 2648 26246
rect 2596 26182 2648 26188
rect 2516 25906 2544 26182
rect 2596 26036 2648 26042
rect 2596 25978 2648 25984
rect 2504 25900 2556 25906
rect 2504 25842 2556 25848
rect 2504 25424 2556 25430
rect 2504 25366 2556 25372
rect 2412 25288 2464 25294
rect 2412 25230 2464 25236
rect 2516 24970 2544 25366
rect 2608 25158 2636 25978
rect 2596 25152 2648 25158
rect 2596 25094 2648 25100
rect 2700 24993 2728 26404
rect 2884 26330 2912 28902
rect 2976 27538 3004 29174
rect 3068 28257 3096 29294
rect 3054 28248 3110 28257
rect 3054 28183 3110 28192
rect 3068 28082 3096 28183
rect 3056 28076 3108 28082
rect 3056 28018 3108 28024
rect 3054 27976 3110 27985
rect 3054 27911 3056 27920
rect 3108 27911 3110 27920
rect 3056 27882 3108 27888
rect 3054 27840 3110 27849
rect 3054 27775 3110 27784
rect 3068 27674 3096 27775
rect 3056 27668 3108 27674
rect 3056 27610 3108 27616
rect 2964 27532 3016 27538
rect 2964 27474 3016 27480
rect 2964 27328 3016 27334
rect 2964 27270 3016 27276
rect 3160 27282 3188 29582
rect 3240 29572 3292 29578
rect 3240 29514 3292 29520
rect 3252 28937 3280 29514
rect 3332 29504 3384 29510
rect 3332 29446 3384 29452
rect 3238 28928 3294 28937
rect 3238 28863 3294 28872
rect 3240 28552 3292 28558
rect 3240 28494 3292 28500
rect 3252 27577 3280 28494
rect 3238 27568 3294 27577
rect 3238 27503 3294 27512
rect 3344 27305 3372 29446
rect 3436 29345 3464 29804
rect 3804 29714 3832 30534
rect 3792 29708 3844 29714
rect 3792 29650 3844 29656
rect 3422 29336 3478 29345
rect 3896 29306 3924 32370
rect 3988 30258 4016 33526
rect 4080 33300 4108 33952
rect 4252 33934 4304 33940
rect 4160 33856 4212 33862
rect 4160 33798 4212 33804
rect 4172 33425 4200 33798
rect 4158 33416 4214 33425
rect 4158 33351 4214 33360
rect 4080 33272 4200 33300
rect 4068 32904 4120 32910
rect 4068 32846 4120 32852
rect 4080 32570 4108 32846
rect 4068 32564 4120 32570
rect 4068 32506 4120 32512
rect 4068 32020 4120 32026
rect 4068 31962 4120 31968
rect 3976 30252 4028 30258
rect 3976 30194 4028 30200
rect 3976 30116 4028 30122
rect 3976 30058 4028 30064
rect 3988 30025 4016 30058
rect 3974 30016 4030 30025
rect 3974 29951 4030 29960
rect 3974 29744 4030 29753
rect 3974 29679 4030 29688
rect 3988 29646 4016 29679
rect 3976 29640 4028 29646
rect 3976 29582 4028 29588
rect 3422 29271 3478 29280
rect 3884 29300 3936 29306
rect 3884 29242 3936 29248
rect 3976 29300 4028 29306
rect 3976 29242 4028 29248
rect 3792 29096 3844 29102
rect 3792 29038 3844 29044
rect 3422 28860 3730 28869
rect 3422 28858 3428 28860
rect 3484 28858 3508 28860
rect 3564 28858 3588 28860
rect 3644 28858 3668 28860
rect 3724 28858 3730 28860
rect 3484 28806 3486 28858
rect 3666 28806 3668 28858
rect 3422 28804 3428 28806
rect 3484 28804 3508 28806
rect 3564 28804 3588 28806
rect 3644 28804 3668 28806
rect 3724 28804 3730 28806
rect 3422 28795 3730 28804
rect 3804 28121 3832 29038
rect 3884 29028 3936 29034
rect 3884 28970 3936 28976
rect 3790 28112 3846 28121
rect 3790 28047 3846 28056
rect 3422 27772 3730 27781
rect 3422 27770 3428 27772
rect 3484 27770 3508 27772
rect 3564 27770 3588 27772
rect 3644 27770 3668 27772
rect 3724 27770 3730 27772
rect 3484 27718 3486 27770
rect 3666 27718 3668 27770
rect 3422 27716 3428 27718
rect 3484 27716 3508 27718
rect 3564 27716 3588 27718
rect 3644 27716 3668 27718
rect 3724 27716 3730 27718
rect 3422 27707 3730 27716
rect 3700 27532 3752 27538
rect 3752 27492 3832 27520
rect 3700 27474 3752 27480
rect 3698 27432 3754 27441
rect 3698 27367 3754 27376
rect 3330 27296 3386 27305
rect 2792 26302 2912 26330
rect 2686 24984 2742 24993
rect 2516 24942 2636 24970
rect 2502 24712 2558 24721
rect 2502 24647 2504 24656
rect 2556 24647 2558 24656
rect 2504 24618 2556 24624
rect 2502 24304 2558 24313
rect 2502 24239 2558 24248
rect 2412 24064 2464 24070
rect 2412 24006 2464 24012
rect 2424 23662 2452 24006
rect 2412 23656 2464 23662
rect 2412 23598 2464 23604
rect 2320 23316 2372 23322
rect 2320 23258 2372 23264
rect 2332 23066 2360 23258
rect 2240 23038 2360 23066
rect 2516 23050 2544 24239
rect 2504 23044 2556 23050
rect 2240 22522 2268 23038
rect 2504 22986 2556 22992
rect 2320 22976 2372 22982
rect 2320 22918 2372 22924
rect 2332 22710 2360 22918
rect 2320 22704 2372 22710
rect 2320 22646 2372 22652
rect 2412 22636 2464 22642
rect 2412 22578 2464 22584
rect 2240 22494 2360 22522
rect 2148 22392 2268 22420
rect 2134 22128 2190 22137
rect 2134 22063 2190 22072
rect 2044 21684 2096 21690
rect 2044 21626 2096 21632
rect 1952 21616 2004 21622
rect 1952 21558 2004 21564
rect 1952 21344 2004 21350
rect 1950 21312 1952 21321
rect 2004 21312 2006 21321
rect 1950 21247 2006 21256
rect 2148 21162 2176 22063
rect 2056 21134 2176 21162
rect 1950 20632 2006 20641
rect 1860 20596 1912 20602
rect 1950 20567 2006 20576
rect 1860 20538 1912 20544
rect 1872 20466 1900 20538
rect 1860 20460 1912 20466
rect 1860 20402 1912 20408
rect 1858 19952 1914 19961
rect 1858 19887 1914 19896
rect 1766 19000 1822 19009
rect 1766 18935 1822 18944
rect 1768 18896 1820 18902
rect 1768 18838 1820 18844
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1582 17504 1638 17513
rect 1504 15706 1532 17478
rect 1582 17439 1638 17448
rect 1596 17338 1624 17439
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1780 16969 1808 18838
rect 1872 18698 1900 19887
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1964 18358 1992 20567
rect 2056 19938 2084 21134
rect 2240 20992 2268 22392
rect 2332 21486 2360 22494
rect 2424 21894 2452 22578
rect 2504 22568 2556 22574
rect 2504 22510 2556 22516
rect 2412 21888 2464 21894
rect 2412 21830 2464 21836
rect 2516 21690 2544 22510
rect 2504 21684 2556 21690
rect 2504 21626 2556 21632
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2320 21480 2372 21486
rect 2320 21422 2372 21428
rect 2424 21298 2452 21490
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2148 20964 2268 20992
rect 2332 21270 2452 21298
rect 2148 20074 2176 20964
rect 2228 20868 2280 20874
rect 2228 20810 2280 20816
rect 2240 20602 2268 20810
rect 2332 20754 2360 21270
rect 2516 20874 2544 21422
rect 2504 20868 2556 20874
rect 2504 20810 2556 20816
rect 2608 20754 2636 24942
rect 2686 24919 2742 24928
rect 2700 24886 2728 24919
rect 2688 24880 2740 24886
rect 2688 24822 2740 24828
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2700 24324 2728 24550
rect 2792 24392 2820 26302
rect 2872 25968 2924 25974
rect 2976 25956 3004 27270
rect 3160 27254 3280 27282
rect 3146 27160 3202 27169
rect 3252 27146 3280 27254
rect 3330 27231 3386 27240
rect 3252 27118 3372 27146
rect 3146 27095 3202 27104
rect 3056 26920 3108 26926
rect 3056 26862 3108 26868
rect 3068 26518 3096 26862
rect 3160 26858 3188 27095
rect 3240 26988 3292 26994
rect 3240 26930 3292 26936
rect 3148 26852 3200 26858
rect 3148 26794 3200 26800
rect 3252 26586 3280 26930
rect 3240 26580 3292 26586
rect 3240 26522 3292 26528
rect 3056 26512 3108 26518
rect 3056 26454 3108 26460
rect 3056 26376 3108 26382
rect 3054 26344 3056 26353
rect 3148 26376 3200 26382
rect 3108 26344 3110 26353
rect 3148 26318 3200 26324
rect 3054 26279 3110 26288
rect 2924 25928 3096 25956
rect 3160 25945 3188 26318
rect 2872 25910 2924 25916
rect 2870 25392 2926 25401
rect 2870 25327 2926 25336
rect 2884 24750 2912 25327
rect 2872 24744 2924 24750
rect 2924 24704 3004 24732
rect 2872 24686 2924 24692
rect 2792 24364 2912 24392
rect 2700 24296 2820 24324
rect 2792 23730 2820 24296
rect 2688 23724 2740 23730
rect 2688 23666 2740 23672
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2700 23322 2728 23666
rect 2688 23316 2740 23322
rect 2688 23258 2740 23264
rect 2688 23112 2740 23118
rect 2688 23054 2740 23060
rect 2332 20726 2452 20754
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2320 20256 2372 20262
rect 2320 20198 2372 20204
rect 2226 20088 2282 20097
rect 2148 20046 2226 20074
rect 2226 20023 2282 20032
rect 2056 19910 2268 19938
rect 2332 19922 2360 20198
rect 2134 19816 2190 19825
rect 2134 19751 2190 19760
rect 2148 19446 2176 19751
rect 2136 19440 2188 19446
rect 2136 19382 2188 19388
rect 2044 19168 2096 19174
rect 2096 19128 2176 19156
rect 2044 19110 2096 19116
rect 2042 18728 2098 18737
rect 2042 18663 2044 18672
rect 2096 18663 2098 18672
rect 2044 18634 2096 18640
rect 1952 18352 2004 18358
rect 1952 18294 2004 18300
rect 1952 18080 2004 18086
rect 1952 18022 2004 18028
rect 1860 17808 1912 17814
rect 1860 17750 1912 17756
rect 1582 16960 1638 16969
rect 1582 16895 1638 16904
rect 1766 16960 1822 16969
rect 1766 16895 1822 16904
rect 1596 16250 1624 16895
rect 1674 16824 1730 16833
rect 1674 16759 1730 16768
rect 1768 16788 1820 16794
rect 1584 16244 1636 16250
rect 1584 16186 1636 16192
rect 1688 16182 1716 16759
rect 1768 16730 1820 16736
rect 1780 16697 1808 16730
rect 1766 16688 1822 16697
rect 1766 16623 1822 16632
rect 1676 16176 1728 16182
rect 1676 16118 1728 16124
rect 1766 16008 1822 16017
rect 1766 15943 1822 15952
rect 1674 15872 1730 15881
rect 1674 15807 1730 15816
rect 1688 15706 1716 15807
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 1398 14512 1454 14521
rect 1308 14476 1360 14482
rect 1398 14447 1454 14456
rect 1308 14418 1360 14424
rect 1228 14334 1440 14362
rect 1306 13016 1362 13025
rect 1306 12951 1362 12960
rect 1320 10062 1348 12951
rect 1412 10985 1440 14334
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1504 11054 1532 13631
rect 1596 13530 1624 15263
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1584 13524 1636 13530
rect 1584 13466 1636 13472
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1596 12238 1624 13262
rect 1688 12986 1716 14962
rect 1780 14006 1808 15943
rect 1768 14000 1820 14006
rect 1768 13942 1820 13948
rect 1872 13258 1900 17750
rect 1964 17338 1992 18022
rect 2148 17954 2176 19128
rect 2056 17926 2176 17954
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2056 17202 2084 17926
rect 2240 17882 2268 19910
rect 2320 19916 2372 19922
rect 2320 19858 2372 19864
rect 2332 19174 2360 19858
rect 2320 19168 2372 19174
rect 2320 19110 2372 19116
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2228 17740 2280 17746
rect 2228 17682 2280 17688
rect 2136 17536 2188 17542
rect 2136 17478 2188 17484
rect 2148 17241 2176 17478
rect 2134 17232 2190 17241
rect 1952 17196 2004 17202
rect 1952 17138 2004 17144
rect 2044 17196 2096 17202
rect 2134 17167 2190 17176
rect 2044 17138 2096 17144
rect 1964 16250 1992 17138
rect 2056 16658 2084 17138
rect 2044 16652 2096 16658
rect 2044 16594 2096 16600
rect 2240 16538 2268 17682
rect 2332 17490 2360 18022
rect 2424 17746 2452 20726
rect 2516 20726 2636 20754
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2332 17462 2452 17490
rect 2318 17368 2374 17377
rect 2318 17303 2374 17312
rect 2332 17270 2360 17303
rect 2320 17264 2372 17270
rect 2320 17206 2372 17212
rect 2056 16510 2268 16538
rect 1952 16244 2004 16250
rect 1952 16186 2004 16192
rect 1952 16108 2004 16114
rect 1952 16050 2004 16056
rect 1964 15162 1992 16050
rect 2056 16017 2084 16510
rect 2320 16448 2372 16454
rect 2226 16416 2282 16425
rect 2320 16390 2372 16396
rect 2226 16351 2282 16360
rect 2240 16182 2268 16351
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2042 16008 2098 16017
rect 2042 15943 2098 15952
rect 2056 15502 2084 15943
rect 2136 15904 2188 15910
rect 2136 15846 2188 15852
rect 2148 15609 2176 15846
rect 2134 15600 2190 15609
rect 2134 15535 2190 15544
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2136 15496 2188 15502
rect 2136 15438 2188 15444
rect 1952 15156 2004 15162
rect 1952 15098 2004 15104
rect 1950 15056 2006 15065
rect 1950 14991 2006 15000
rect 2044 15020 2096 15026
rect 1964 14074 1992 14991
rect 2044 14962 2096 14968
rect 2056 14482 2084 14962
rect 2044 14476 2096 14482
rect 2044 14418 2096 14424
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2042 13968 2098 13977
rect 2042 13903 2098 13912
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1766 13152 1822 13161
rect 1766 13087 1822 13096
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1674 12336 1730 12345
rect 1674 12271 1730 12280
rect 1584 12232 1636 12238
rect 1584 12174 1636 12180
rect 1582 12064 1638 12073
rect 1582 11999 1638 12008
rect 1596 11234 1624 11999
rect 1688 11354 1716 12271
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1596 11206 1716 11234
rect 1504 11026 1624 11054
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1596 10810 1624 11026
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1308 10056 1360 10062
rect 1308 9998 1360 10004
rect 1306 9616 1362 9625
rect 1306 9551 1362 9560
rect 1214 8528 1270 8537
rect 1214 8463 1270 8472
rect 1030 7511 1086 7520
rect 1124 7540 1176 7546
rect 846 2000 902 2009
rect 846 1935 902 1944
rect 756 1896 808 1902
rect 756 1838 808 1844
rect 480 1488 532 1494
rect 480 1430 532 1436
rect 1044 1426 1072 7511
rect 1124 7482 1176 7488
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 1136 6866 1164 7278
rect 1124 6860 1176 6866
rect 1124 6802 1176 6808
rect 1136 5778 1164 6802
rect 1124 5772 1176 5778
rect 1124 5714 1176 5720
rect 1228 4826 1256 8463
rect 1320 5370 1348 9551
rect 1412 7954 1440 10746
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 10266 1532 10610
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1492 10124 1544 10130
rect 1492 10066 1544 10072
rect 1504 8634 1532 10066
rect 1582 9344 1638 9353
rect 1582 9279 1638 9288
rect 1492 8628 1544 8634
rect 1492 8570 1544 8576
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1400 7948 1452 7954
rect 1400 7890 1452 7896
rect 1398 7848 1454 7857
rect 1398 7783 1400 7792
rect 1452 7783 1454 7792
rect 1400 7754 1452 7760
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1412 6882 1440 7647
rect 1504 7002 1532 8434
rect 1596 7002 1624 9279
rect 1688 9160 1716 11206
rect 1780 9722 1808 13087
rect 1858 11792 1914 11801
rect 1964 11762 1992 13670
rect 2056 12646 2084 13903
rect 2148 13240 2176 15438
rect 2228 15156 2280 15162
rect 2228 15098 2280 15104
rect 2240 14414 2268 15098
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2228 14272 2280 14278
rect 2228 14214 2280 14220
rect 2240 13870 2268 14214
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2332 13734 2360 16390
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 2228 13252 2280 13258
rect 2148 13212 2228 13240
rect 2228 13194 2280 13200
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 1858 11727 1914 11736
rect 1952 11756 2004 11762
rect 1768 9716 1820 9722
rect 1768 9658 1820 9664
rect 1768 9172 1820 9178
rect 1688 9132 1768 9160
rect 1768 9114 1820 9120
rect 1766 9072 1822 9081
rect 1766 9007 1822 9016
rect 1674 8392 1730 8401
rect 1674 8327 1730 8336
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1412 6854 1532 6882
rect 1398 5808 1454 5817
rect 1398 5743 1454 5752
rect 1308 5364 1360 5370
rect 1308 5306 1360 5312
rect 1306 5264 1362 5273
rect 1306 5199 1362 5208
rect 1216 4820 1268 4826
rect 1216 4762 1268 4768
rect 1320 2038 1348 5199
rect 1412 2106 1440 5743
rect 1504 4154 1532 6854
rect 1584 6452 1636 6458
rect 1688 6440 1716 8327
rect 1780 7206 1808 9007
rect 1872 8634 1900 11727
rect 1952 11698 2004 11704
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1950 11520 2006 11529
rect 1950 11455 2006 11464
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 1872 7970 1900 8366
rect 1964 8090 1992 11455
rect 2056 11218 2084 11630
rect 2136 11552 2188 11558
rect 2136 11494 2188 11500
rect 2148 11286 2176 11494
rect 2136 11280 2188 11286
rect 2136 11222 2188 11228
rect 2044 11212 2096 11218
rect 2044 11154 2096 11160
rect 2042 11112 2098 11121
rect 2098 11070 2176 11098
rect 2042 11047 2098 11056
rect 2148 11014 2176 11070
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2056 8974 2084 10950
rect 2240 10849 2268 13194
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2332 12306 2360 12718
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2424 12170 2452 17462
rect 2516 16561 2544 20726
rect 2700 19854 2728 23054
rect 2792 22953 2820 23666
rect 2778 22944 2834 22953
rect 2778 22879 2834 22888
rect 2780 22636 2832 22642
rect 2780 22578 2832 22584
rect 2792 22234 2820 22578
rect 2780 22228 2832 22234
rect 2780 22170 2832 22176
rect 2780 22092 2832 22098
rect 2780 22034 2832 22040
rect 2792 20913 2820 22034
rect 2778 20904 2834 20913
rect 2778 20839 2834 20848
rect 2884 20806 2912 24364
rect 2976 24274 3004 24704
rect 2964 24268 3016 24274
rect 2964 24210 3016 24216
rect 2964 24064 3016 24070
rect 2964 24006 3016 24012
rect 2976 23866 3004 24006
rect 2964 23860 3016 23866
rect 2964 23802 3016 23808
rect 2962 23216 3018 23225
rect 2962 23151 3018 23160
rect 2976 22273 3004 23151
rect 2962 22264 3018 22273
rect 2962 22199 3018 22208
rect 3068 20874 3096 25928
rect 3146 25936 3202 25945
rect 3146 25871 3202 25880
rect 3240 25900 3292 25906
rect 3240 25842 3292 25848
rect 3148 25696 3200 25702
rect 3148 25638 3200 25644
rect 3160 23225 3188 25638
rect 3252 25430 3280 25842
rect 3240 25424 3292 25430
rect 3240 25366 3292 25372
rect 3240 24812 3292 24818
rect 3240 24754 3292 24760
rect 3252 24138 3280 24754
rect 3240 24132 3292 24138
rect 3240 24074 3292 24080
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3146 23216 3202 23225
rect 3146 23151 3202 23160
rect 3148 22704 3200 22710
rect 3148 22646 3200 22652
rect 3056 20868 3108 20874
rect 3056 20810 3108 20816
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 2688 19848 2740 19854
rect 2688 19790 2740 19796
rect 2700 19553 2728 19790
rect 2686 19544 2742 19553
rect 2686 19479 2742 19488
rect 2686 19408 2742 19417
rect 2686 19343 2742 19352
rect 2594 18864 2650 18873
rect 2594 18799 2650 18808
rect 2608 17082 2636 18799
rect 2700 18766 2728 19343
rect 2780 19168 2832 19174
rect 2780 19110 2832 19116
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2792 18630 2820 19110
rect 2780 18624 2832 18630
rect 2780 18566 2832 18572
rect 2884 18465 2912 20742
rect 2962 20496 3018 20505
rect 2962 20431 3018 20440
rect 2870 18456 2926 18465
rect 2870 18391 2926 18400
rect 2976 18306 3004 20431
rect 3068 18970 3096 20810
rect 3160 19689 3188 22646
rect 3252 21729 3280 23802
rect 3344 23304 3372 27118
rect 3608 27056 3660 27062
rect 3606 27024 3608 27033
rect 3660 27024 3662 27033
rect 3606 26959 3662 26968
rect 3712 26926 3740 27367
rect 3700 26920 3752 26926
rect 3700 26862 3752 26868
rect 3422 26684 3730 26693
rect 3422 26682 3428 26684
rect 3484 26682 3508 26684
rect 3564 26682 3588 26684
rect 3644 26682 3668 26684
rect 3724 26682 3730 26684
rect 3484 26630 3486 26682
rect 3666 26630 3668 26682
rect 3422 26628 3428 26630
rect 3484 26628 3508 26630
rect 3564 26628 3588 26630
rect 3644 26628 3668 26630
rect 3724 26628 3730 26630
rect 3422 26619 3730 26628
rect 3516 26240 3568 26246
rect 3608 26240 3660 26246
rect 3516 26182 3568 26188
rect 3606 26208 3608 26217
rect 3660 26208 3662 26217
rect 3528 25684 3556 26182
rect 3606 26143 3662 26152
rect 3700 25900 3752 25906
rect 3700 25842 3752 25848
rect 3712 25809 3740 25842
rect 3698 25800 3754 25809
rect 3698 25735 3754 25744
rect 3804 25752 3832 27492
rect 3896 26926 3924 28970
rect 3988 28150 4016 29242
rect 3976 28144 4028 28150
rect 3976 28086 4028 28092
rect 3988 27713 4016 28086
rect 3974 27704 4030 27713
rect 3974 27639 4030 27648
rect 3974 27568 4030 27577
rect 3974 27503 4030 27512
rect 3884 26920 3936 26926
rect 3884 26862 3936 26868
rect 3988 26518 4016 27503
rect 4080 27334 4108 31962
rect 4172 30938 4200 33272
rect 4264 33153 4292 33934
rect 4250 33144 4306 33153
rect 4356 33114 4384 41074
rect 4448 34202 4476 41074
rect 4540 38010 4568 41262
rect 4632 39030 4660 42191
rect 4896 42162 4948 42168
rect 4710 41848 4766 41857
rect 4710 41783 4766 41792
rect 4724 41614 4752 41783
rect 4712 41608 4764 41614
rect 4712 41550 4764 41556
rect 4908 41274 4936 42162
rect 5000 41274 5028 42570
rect 5184 42362 5212 44540
rect 5264 43308 5316 43314
rect 5264 43250 5316 43256
rect 5276 42906 5304 43250
rect 5264 42900 5316 42906
rect 5264 42842 5316 42848
rect 5368 42770 5396 44540
rect 5552 43450 5580 44540
rect 5632 43716 5684 43722
rect 5632 43658 5684 43664
rect 5540 43444 5592 43450
rect 5540 43386 5592 43392
rect 5448 43308 5500 43314
rect 5448 43250 5500 43256
rect 5356 42764 5408 42770
rect 5356 42706 5408 42712
rect 5172 42356 5224 42362
rect 5460 42344 5488 43250
rect 5172 42298 5224 42304
rect 5368 42316 5488 42344
rect 5172 42016 5224 42022
rect 5172 41958 5224 41964
rect 5184 41614 5212 41958
rect 5080 41608 5132 41614
rect 5080 41550 5132 41556
rect 5172 41608 5224 41614
rect 5172 41550 5224 41556
rect 5092 41290 5120 41550
rect 5172 41472 5224 41478
rect 5172 41414 5224 41420
rect 5184 41386 5304 41414
rect 4896 41268 4948 41274
rect 4896 41210 4948 41216
rect 4988 41268 5040 41274
rect 5092 41262 5212 41290
rect 5276 41274 5304 41386
rect 4988 41210 5040 41216
rect 5184 41154 5212 41262
rect 5264 41268 5316 41274
rect 5264 41210 5316 41216
rect 4988 41132 5040 41138
rect 4988 41074 5040 41080
rect 5080 41132 5132 41138
rect 5184 41126 5304 41154
rect 5080 41074 5132 41080
rect 4894 40624 4950 40633
rect 4894 40559 4950 40568
rect 4908 40050 4936 40559
rect 4896 40044 4948 40050
rect 4896 39986 4948 39992
rect 4712 39296 4764 39302
rect 4712 39238 4764 39244
rect 4620 39024 4672 39030
rect 4620 38966 4672 38972
rect 4632 38214 4660 38966
rect 4724 38894 4752 39238
rect 4802 39128 4858 39137
rect 4802 39063 4858 39072
rect 4816 39030 4844 39063
rect 4804 39024 4856 39030
rect 4804 38966 4856 38972
rect 4712 38888 4764 38894
rect 4712 38830 4764 38836
rect 4816 38350 4844 38966
rect 5000 38865 5028 41074
rect 4986 38856 5042 38865
rect 4986 38791 5042 38800
rect 4804 38344 4856 38350
rect 4804 38286 4856 38292
rect 4896 38344 4948 38350
rect 4896 38286 4948 38292
rect 4620 38208 4672 38214
rect 4620 38150 4672 38156
rect 4528 38004 4580 38010
rect 4528 37946 4580 37952
rect 4632 37890 4660 38150
rect 4540 37862 4660 37890
rect 4540 36145 4568 37862
rect 4618 36816 4674 36825
rect 4674 36774 4752 36802
rect 4618 36751 4674 36760
rect 4526 36136 4582 36145
rect 4526 36071 4582 36080
rect 4620 36100 4672 36106
rect 4620 36042 4672 36048
rect 4528 36032 4580 36038
rect 4528 35974 4580 35980
rect 4436 34196 4488 34202
rect 4436 34138 4488 34144
rect 4540 33590 4568 35974
rect 4632 35834 4660 36042
rect 4620 35828 4672 35834
rect 4620 35770 4672 35776
rect 4620 35692 4672 35698
rect 4620 35634 4672 35640
rect 4632 34950 4660 35634
rect 4724 35136 4752 36774
rect 4816 36174 4844 38286
rect 4908 38214 4936 38286
rect 4988 38276 5040 38282
rect 4988 38218 5040 38224
rect 4896 38208 4948 38214
rect 4896 38150 4948 38156
rect 4908 37874 4936 38150
rect 4896 37868 4948 37874
rect 4896 37810 4948 37816
rect 4804 36168 4856 36174
rect 4804 36110 4856 36116
rect 4908 36038 4936 37810
rect 5000 36106 5028 38218
rect 4988 36100 5040 36106
rect 4988 36042 5040 36048
rect 4896 36032 4948 36038
rect 4896 35974 4948 35980
rect 4724 35108 4844 35136
rect 4712 35012 4764 35018
rect 4712 34954 4764 34960
rect 4620 34944 4672 34950
rect 4620 34886 4672 34892
rect 4632 34678 4660 34886
rect 4620 34672 4672 34678
rect 4620 34614 4672 34620
rect 4724 34610 4752 34954
rect 4712 34604 4764 34610
rect 4712 34546 4764 34552
rect 4620 33992 4672 33998
rect 4620 33934 4672 33940
rect 4632 33862 4660 33934
rect 4620 33856 4672 33862
rect 4620 33798 4672 33804
rect 4528 33584 4580 33590
rect 4528 33526 4580 33532
rect 4436 33516 4488 33522
rect 4436 33458 4488 33464
rect 4448 33425 4476 33458
rect 4434 33416 4490 33425
rect 4434 33351 4490 33360
rect 4540 33300 4568 33526
rect 4448 33272 4568 33300
rect 4250 33079 4306 33088
rect 4344 33108 4396 33114
rect 4160 30932 4212 30938
rect 4160 30874 4212 30880
rect 4160 30184 4212 30190
rect 4160 30126 4212 30132
rect 4172 29889 4200 30126
rect 4158 29880 4214 29889
rect 4158 29815 4214 29824
rect 4160 29572 4212 29578
rect 4160 29514 4212 29520
rect 4172 28064 4200 29514
rect 4264 29306 4292 33079
rect 4344 33050 4396 33056
rect 4342 32464 4398 32473
rect 4342 32399 4344 32408
rect 4396 32399 4398 32408
rect 4344 32370 4396 32376
rect 4448 30274 4476 33272
rect 4816 33134 4844 35108
rect 4894 34640 4950 34649
rect 4894 34575 4950 34584
rect 4908 34406 4936 34575
rect 4896 34400 4948 34406
rect 4896 34342 4948 34348
rect 4908 34066 4936 34342
rect 4896 34060 4948 34066
rect 4896 34002 4948 34008
rect 5000 33522 5028 36042
rect 5092 35290 5120 41074
rect 5276 40662 5304 41126
rect 5368 41070 5396 42316
rect 5540 42220 5592 42226
rect 5540 42162 5592 42168
rect 5446 41848 5502 41857
rect 5552 41818 5580 42162
rect 5446 41783 5502 41792
rect 5540 41812 5592 41818
rect 5460 41750 5488 41783
rect 5540 41754 5592 41760
rect 5448 41744 5500 41750
rect 5448 41686 5500 41692
rect 5538 41712 5594 41721
rect 5538 41647 5594 41656
rect 5552 41614 5580 41647
rect 5448 41608 5500 41614
rect 5446 41576 5448 41585
rect 5540 41608 5592 41614
rect 5500 41576 5502 41585
rect 5540 41550 5592 41556
rect 5644 41562 5672 43658
rect 5736 42362 5764 44540
rect 5920 43738 5948 44540
rect 5828 43710 5948 43738
rect 6104 43738 6132 44540
rect 6288 43897 6316 44540
rect 6274 43888 6330 43897
rect 6274 43823 6330 43832
rect 6104 43710 6316 43738
rect 5828 43178 5856 43710
rect 5894 43548 6202 43557
rect 5894 43546 5900 43548
rect 5956 43546 5980 43548
rect 6036 43546 6060 43548
rect 6116 43546 6140 43548
rect 6196 43546 6202 43548
rect 5956 43494 5958 43546
rect 6138 43494 6140 43546
rect 5894 43492 5900 43494
rect 5956 43492 5980 43494
rect 6036 43492 6060 43494
rect 6116 43492 6140 43494
rect 6196 43492 6202 43494
rect 5894 43483 6202 43492
rect 5816 43172 5868 43178
rect 5816 43114 5868 43120
rect 5908 43104 5960 43110
rect 6000 43104 6052 43110
rect 5908 43046 5960 43052
rect 5998 43072 6000 43081
rect 6052 43072 6054 43081
rect 5920 42702 5948 43046
rect 5998 43007 6054 43016
rect 6288 42770 6316 43710
rect 6368 42900 6420 42906
rect 6368 42842 6420 42848
rect 6276 42764 6328 42770
rect 6276 42706 6328 42712
rect 5908 42696 5960 42702
rect 5908 42638 5960 42644
rect 5816 42628 5868 42634
rect 5816 42570 5868 42576
rect 5724 42356 5776 42362
rect 5724 42298 5776 42304
rect 5644 41534 5764 41562
rect 5446 41511 5502 41520
rect 5540 41472 5592 41478
rect 5540 41414 5592 41420
rect 5632 41472 5684 41478
rect 5632 41414 5684 41420
rect 5356 41064 5408 41070
rect 5356 41006 5408 41012
rect 5264 40656 5316 40662
rect 5264 40598 5316 40604
rect 5552 40610 5580 41414
rect 5644 40730 5672 41414
rect 5736 41018 5764 41534
rect 5828 41274 5856 42570
rect 5894 42460 6202 42469
rect 5894 42458 5900 42460
rect 5956 42458 5980 42460
rect 6036 42458 6060 42460
rect 6116 42458 6140 42460
rect 6196 42458 6202 42460
rect 5956 42406 5958 42458
rect 6138 42406 6140 42458
rect 5894 42404 5900 42406
rect 5956 42404 5980 42406
rect 6036 42404 6060 42406
rect 6116 42404 6140 42406
rect 6196 42404 6202 42406
rect 5894 42395 6202 42404
rect 6276 42220 6328 42226
rect 6276 42162 6328 42168
rect 5894 41372 6202 41381
rect 5894 41370 5900 41372
rect 5956 41370 5980 41372
rect 6036 41370 6060 41372
rect 6116 41370 6140 41372
rect 6196 41370 6202 41372
rect 5956 41318 5958 41370
rect 6138 41318 6140 41370
rect 5894 41316 5900 41318
rect 5956 41316 5980 41318
rect 6036 41316 6060 41318
rect 6116 41316 6140 41318
rect 6196 41316 6202 41318
rect 5894 41307 6202 41316
rect 5816 41268 5868 41274
rect 5816 41210 5868 41216
rect 6288 41070 6316 42162
rect 6380 41698 6408 42842
rect 6472 42770 6500 44540
rect 6460 42764 6512 42770
rect 6460 42706 6512 42712
rect 6552 42628 6604 42634
rect 6552 42570 6604 42576
rect 6380 41670 6500 41698
rect 6366 41576 6422 41585
rect 6366 41511 6422 41520
rect 6276 41064 6328 41070
rect 5736 40990 5856 41018
rect 6276 41006 6328 41012
rect 5724 40928 5776 40934
rect 5724 40870 5776 40876
rect 5632 40724 5684 40730
rect 5632 40666 5684 40672
rect 5736 40610 5764 40870
rect 5552 40582 5764 40610
rect 5828 40032 5856 40990
rect 5894 40284 6202 40293
rect 5894 40282 5900 40284
rect 5956 40282 5980 40284
rect 6036 40282 6060 40284
rect 6116 40282 6140 40284
rect 6196 40282 6202 40284
rect 5956 40230 5958 40282
rect 6138 40230 6140 40282
rect 5894 40228 5900 40230
rect 5956 40228 5980 40230
rect 6036 40228 6060 40230
rect 6116 40228 6140 40230
rect 6196 40228 6202 40230
rect 5894 40219 6202 40228
rect 5736 40004 5856 40032
rect 5448 39840 5500 39846
rect 5448 39782 5500 39788
rect 5540 39840 5592 39846
rect 5540 39782 5592 39788
rect 5460 39302 5488 39782
rect 5448 39296 5500 39302
rect 5448 39238 5500 39244
rect 5172 38956 5224 38962
rect 5172 38898 5224 38904
rect 5184 38282 5212 38898
rect 5262 38448 5318 38457
rect 5262 38383 5264 38392
rect 5316 38383 5318 38392
rect 5264 38354 5316 38360
rect 5172 38276 5224 38282
rect 5172 38218 5224 38224
rect 5264 38208 5316 38214
rect 5264 38150 5316 38156
rect 5276 37398 5304 38150
rect 5460 37992 5488 39238
rect 5552 39030 5580 39782
rect 5540 39024 5592 39030
rect 5540 38966 5592 38972
rect 5632 38956 5684 38962
rect 5632 38898 5684 38904
rect 5644 38350 5672 38898
rect 5632 38344 5684 38350
rect 5632 38286 5684 38292
rect 5460 37964 5672 37992
rect 5540 37868 5592 37874
rect 5540 37810 5592 37816
rect 5356 37800 5408 37806
rect 5356 37742 5408 37748
rect 5264 37392 5316 37398
rect 5264 37334 5316 37340
rect 5264 37256 5316 37262
rect 5262 37224 5264 37233
rect 5316 37224 5318 37233
rect 5262 37159 5318 37168
rect 5172 36712 5224 36718
rect 5172 36654 5224 36660
rect 5080 35284 5132 35290
rect 5080 35226 5132 35232
rect 4988 33516 5040 33522
rect 4988 33458 5040 33464
rect 4724 33106 4844 33134
rect 5184 33114 5212 36654
rect 5276 35086 5304 37159
rect 5368 36786 5396 37742
rect 5552 37369 5580 37810
rect 5538 37360 5594 37369
rect 5538 37295 5594 37304
rect 5448 37188 5500 37194
rect 5448 37130 5500 37136
rect 5540 37188 5592 37194
rect 5540 37130 5592 37136
rect 5460 36786 5488 37130
rect 5356 36780 5408 36786
rect 5356 36722 5408 36728
rect 5448 36780 5500 36786
rect 5448 36722 5500 36728
rect 5552 36666 5580 37130
rect 5368 36638 5580 36666
rect 5264 35080 5316 35086
rect 5264 35022 5316 35028
rect 5276 34746 5304 35022
rect 5264 34740 5316 34746
rect 5264 34682 5316 34688
rect 5264 34604 5316 34610
rect 5264 34546 5316 34552
rect 5276 33998 5304 34546
rect 5264 33992 5316 33998
rect 5262 33960 5264 33969
rect 5316 33960 5318 33969
rect 5262 33895 5318 33904
rect 5264 33448 5316 33454
rect 5264 33390 5316 33396
rect 4988 33108 5040 33114
rect 4618 32056 4674 32065
rect 4618 31991 4674 32000
rect 4632 31822 4660 31991
rect 4620 31816 4672 31822
rect 4620 31758 4672 31764
rect 4356 30258 4476 30274
rect 4344 30252 4476 30258
rect 4396 30246 4476 30252
rect 4344 30194 4396 30200
rect 4434 30152 4490 30161
rect 4434 30087 4490 30096
rect 4620 30116 4672 30122
rect 4342 29472 4398 29481
rect 4342 29407 4398 29416
rect 4252 29300 4304 29306
rect 4252 29242 4304 29248
rect 4252 29164 4304 29170
rect 4252 29106 4304 29112
rect 4264 28218 4292 29106
rect 4252 28212 4304 28218
rect 4252 28154 4304 28160
rect 4172 28036 4292 28064
rect 4160 27872 4212 27878
rect 4160 27814 4212 27820
rect 4068 27328 4120 27334
rect 4068 27270 4120 27276
rect 4080 26908 4108 27270
rect 4172 27062 4200 27814
rect 4160 27056 4212 27062
rect 4264 27033 4292 28036
rect 4160 26998 4212 27004
rect 4250 27024 4306 27033
rect 4250 26959 4306 26968
rect 4080 26880 4200 26908
rect 4068 26784 4120 26790
rect 4068 26726 4120 26732
rect 3976 26512 4028 26518
rect 3976 26454 4028 26460
rect 3804 25724 3924 25752
rect 3528 25656 3832 25684
rect 3422 25596 3730 25605
rect 3422 25594 3428 25596
rect 3484 25594 3508 25596
rect 3564 25594 3588 25596
rect 3644 25594 3668 25596
rect 3724 25594 3730 25596
rect 3484 25542 3486 25594
rect 3666 25542 3668 25594
rect 3422 25540 3428 25542
rect 3484 25540 3508 25542
rect 3564 25540 3588 25542
rect 3644 25540 3668 25542
rect 3724 25540 3730 25542
rect 3422 25531 3730 25540
rect 3422 24508 3730 24517
rect 3422 24506 3428 24508
rect 3484 24506 3508 24508
rect 3564 24506 3588 24508
rect 3644 24506 3668 24508
rect 3724 24506 3730 24508
rect 3484 24454 3486 24506
rect 3666 24454 3668 24506
rect 3422 24452 3428 24454
rect 3484 24452 3508 24454
rect 3564 24452 3588 24454
rect 3644 24452 3668 24454
rect 3724 24452 3730 24454
rect 3422 24443 3730 24452
rect 3700 24200 3752 24206
rect 3700 24142 3752 24148
rect 3712 23866 3740 24142
rect 3700 23860 3752 23866
rect 3700 23802 3752 23808
rect 3804 23662 3832 25656
rect 3792 23656 3844 23662
rect 3792 23598 3844 23604
rect 3896 23526 3924 25724
rect 3976 25356 4028 25362
rect 3976 25298 4028 25304
rect 3988 24954 4016 25298
rect 4080 25158 4108 26726
rect 4172 25974 4200 26880
rect 4160 25968 4212 25974
rect 4160 25910 4212 25916
rect 4264 25809 4292 26959
rect 4250 25800 4306 25809
rect 4250 25735 4306 25744
rect 4250 25528 4306 25537
rect 4250 25463 4306 25472
rect 4158 25392 4214 25401
rect 4158 25327 4214 25336
rect 4068 25152 4120 25158
rect 4068 25094 4120 25100
rect 3976 24948 4028 24954
rect 3976 24890 4028 24896
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 3422 23420 3730 23429
rect 3422 23418 3428 23420
rect 3484 23418 3508 23420
rect 3564 23418 3588 23420
rect 3644 23418 3668 23420
rect 3724 23418 3730 23420
rect 3484 23366 3486 23418
rect 3666 23366 3668 23418
rect 3422 23364 3428 23366
rect 3484 23364 3508 23366
rect 3564 23364 3588 23366
rect 3644 23364 3668 23366
rect 3724 23364 3730 23366
rect 3422 23355 3730 23364
rect 3344 23276 3464 23304
rect 3330 23080 3386 23089
rect 3330 23015 3386 23024
rect 3344 22778 3372 23015
rect 3332 22772 3384 22778
rect 3332 22714 3384 22720
rect 3436 22658 3464 23276
rect 3988 23225 4016 24550
rect 4080 24410 4108 25094
rect 4172 24954 4200 25327
rect 4264 25226 4292 25463
rect 4252 25220 4304 25226
rect 4252 25162 4304 25168
rect 4160 24948 4212 24954
rect 4160 24890 4212 24896
rect 4172 24818 4200 24890
rect 4160 24812 4212 24818
rect 4160 24754 4212 24760
rect 4158 24440 4214 24449
rect 4068 24404 4120 24410
rect 4158 24375 4214 24384
rect 4068 24346 4120 24352
rect 4172 24290 4200 24375
rect 4080 24262 4200 24290
rect 4080 24070 4108 24262
rect 4160 24132 4212 24138
rect 4160 24074 4212 24080
rect 4068 24064 4120 24070
rect 4068 24006 4120 24012
rect 4066 23352 4122 23361
rect 4066 23287 4122 23296
rect 3974 23216 4030 23225
rect 3700 23180 3752 23186
rect 3974 23151 4030 23160
rect 3700 23122 3752 23128
rect 3344 22630 3464 22658
rect 3608 22636 3660 22642
rect 3344 22216 3372 22630
rect 3608 22578 3660 22584
rect 3620 22545 3648 22578
rect 3606 22536 3662 22545
rect 3606 22471 3662 22480
rect 3712 22420 3740 23122
rect 4080 23118 4108 23287
rect 4068 23112 4120 23118
rect 4068 23054 4120 23060
rect 4068 22976 4120 22982
rect 4068 22918 4120 22924
rect 3974 22808 4030 22817
rect 3974 22743 3976 22752
rect 4028 22743 4030 22752
rect 3976 22714 4028 22720
rect 4080 22642 4108 22918
rect 3976 22636 4028 22642
rect 3976 22578 4028 22584
rect 4068 22636 4120 22642
rect 4068 22578 4120 22584
rect 3884 22568 3936 22574
rect 3884 22510 3936 22516
rect 3712 22392 3832 22420
rect 3422 22332 3730 22341
rect 3422 22330 3428 22332
rect 3484 22330 3508 22332
rect 3564 22330 3588 22332
rect 3644 22330 3668 22332
rect 3724 22330 3730 22332
rect 3484 22278 3486 22330
rect 3666 22278 3668 22330
rect 3422 22276 3428 22278
rect 3484 22276 3508 22278
rect 3564 22276 3588 22278
rect 3644 22276 3668 22278
rect 3724 22276 3730 22278
rect 3422 22267 3730 22276
rect 3344 22188 3556 22216
rect 3424 22024 3476 22030
rect 3424 21966 3476 21972
rect 3238 21720 3294 21729
rect 3238 21655 3294 21664
rect 3436 21593 3464 21966
rect 3422 21584 3478 21593
rect 3240 21548 3292 21554
rect 3422 21519 3478 21528
rect 3240 21490 3292 21496
rect 3252 20233 3280 21490
rect 3332 21344 3384 21350
rect 3528 21332 3556 22188
rect 3606 21992 3662 22001
rect 3606 21927 3662 21936
rect 3620 21894 3648 21927
rect 3608 21888 3660 21894
rect 3608 21830 3660 21836
rect 3804 21554 3832 22392
rect 3896 21622 3924 22510
rect 3988 22234 4016 22578
rect 4172 22488 4200 24074
rect 4080 22460 4200 22488
rect 3976 22228 4028 22234
rect 3976 22170 4028 22176
rect 3974 22128 4030 22137
rect 3974 22063 4030 22072
rect 3988 22030 4016 22063
rect 3976 22024 4028 22030
rect 3976 21966 4028 21972
rect 4080 21672 4108 22460
rect 4158 22400 4214 22409
rect 4158 22335 4214 22344
rect 4172 22166 4200 22335
rect 4160 22160 4212 22166
rect 4160 22102 4212 22108
rect 3988 21644 4108 21672
rect 3884 21616 3936 21622
rect 3884 21558 3936 21564
rect 3792 21548 3844 21554
rect 3792 21490 3844 21496
rect 3528 21304 3832 21332
rect 3332 21286 3384 21292
rect 3344 21128 3372 21286
rect 3422 21244 3730 21253
rect 3422 21242 3428 21244
rect 3484 21242 3508 21244
rect 3564 21242 3588 21244
rect 3644 21242 3668 21244
rect 3724 21242 3730 21244
rect 3484 21190 3486 21242
rect 3666 21190 3668 21242
rect 3422 21188 3428 21190
rect 3484 21188 3508 21190
rect 3564 21188 3588 21190
rect 3644 21188 3668 21190
rect 3724 21188 3730 21190
rect 3422 21179 3730 21188
rect 3344 21100 3464 21128
rect 3436 20942 3464 21100
rect 3700 21072 3752 21078
rect 3700 21014 3752 21020
rect 3424 20936 3476 20942
rect 3330 20904 3386 20913
rect 3424 20878 3476 20884
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3330 20839 3386 20848
rect 3238 20224 3294 20233
rect 3238 20159 3294 20168
rect 3238 20088 3294 20097
rect 3238 20023 3294 20032
rect 3344 20040 3372 20839
rect 3620 20602 3648 20878
rect 3608 20596 3660 20602
rect 3608 20538 3660 20544
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3528 20369 3556 20402
rect 3712 20369 3740 21014
rect 3514 20360 3570 20369
rect 3514 20295 3570 20304
rect 3698 20360 3754 20369
rect 3698 20295 3754 20304
rect 3422 20156 3730 20165
rect 3422 20154 3428 20156
rect 3484 20154 3508 20156
rect 3564 20154 3588 20156
rect 3644 20154 3668 20156
rect 3724 20154 3730 20156
rect 3484 20102 3486 20154
rect 3666 20102 3668 20154
rect 3422 20100 3428 20102
rect 3484 20100 3508 20102
rect 3564 20100 3588 20102
rect 3644 20100 3668 20102
rect 3724 20100 3730 20102
rect 3422 20091 3730 20100
rect 3700 20052 3752 20058
rect 3252 19786 3280 20023
rect 3344 20012 3464 20040
rect 3240 19780 3292 19786
rect 3240 19722 3292 19728
rect 3146 19680 3202 19689
rect 3146 19615 3202 19624
rect 3056 18964 3108 18970
rect 3056 18906 3108 18912
rect 3056 18760 3108 18766
rect 3056 18702 3108 18708
rect 3068 18601 3096 18702
rect 3160 18630 3188 19615
rect 3252 19514 3280 19722
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3344 19514 3372 19654
rect 3240 19508 3292 19514
rect 3240 19450 3292 19456
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3148 18624 3200 18630
rect 3054 18592 3110 18601
rect 3148 18566 3200 18572
rect 3054 18527 3110 18536
rect 3054 18456 3110 18465
rect 3054 18391 3110 18400
rect 3148 18420 3200 18426
rect 3068 18358 3096 18391
rect 3148 18362 3200 18368
rect 2884 18278 3004 18306
rect 3056 18352 3108 18358
rect 3056 18294 3108 18300
rect 2688 18080 2740 18086
rect 2884 18034 2912 18278
rect 2740 18028 2912 18034
rect 2688 18022 2912 18028
rect 2700 18006 2912 18022
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2700 17785 2728 17818
rect 2686 17776 2742 17785
rect 2686 17711 2742 17720
rect 3068 17134 3096 18294
rect 3160 17762 3188 18362
rect 3252 18358 3280 19450
rect 3330 19408 3386 19417
rect 3330 19343 3386 19352
rect 3344 18766 3372 19343
rect 3436 19174 3464 20012
rect 3700 19994 3752 20000
rect 3712 19718 3740 19994
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 3712 19446 3740 19654
rect 3700 19440 3752 19446
rect 3700 19382 3752 19388
rect 3424 19168 3476 19174
rect 3424 19110 3476 19116
rect 3422 19068 3730 19077
rect 3422 19066 3428 19068
rect 3484 19066 3508 19068
rect 3564 19066 3588 19068
rect 3644 19066 3668 19068
rect 3724 19066 3730 19068
rect 3484 19014 3486 19066
rect 3666 19014 3668 19066
rect 3422 19012 3428 19014
rect 3484 19012 3508 19014
rect 3564 19012 3588 19014
rect 3644 19012 3668 19014
rect 3724 19012 3730 19014
rect 3422 19003 3730 19012
rect 3700 18828 3752 18834
rect 3804 18816 3832 21304
rect 3988 21298 4016 21644
rect 4066 21584 4122 21593
rect 4066 21519 4122 21528
rect 4160 21548 4212 21554
rect 3896 21270 4016 21298
rect 3896 20534 3924 21270
rect 3974 21176 4030 21185
rect 3974 21111 4030 21120
rect 3884 20528 3936 20534
rect 3884 20470 3936 20476
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3752 18788 3832 18816
rect 3700 18770 3752 18776
rect 3332 18760 3384 18766
rect 3332 18702 3384 18708
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 3344 17762 3372 18702
rect 3606 18456 3662 18465
rect 3606 18391 3662 18400
rect 3620 18290 3648 18391
rect 3608 18284 3660 18290
rect 3608 18226 3660 18232
rect 3712 18068 3740 18770
rect 3896 18714 3924 19654
rect 3804 18686 3924 18714
rect 3804 18290 3832 18686
rect 3988 18442 4016 21111
rect 4080 20806 4108 21519
rect 4160 21490 4212 21496
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 4080 19922 4108 20198
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 4172 19825 4200 21490
rect 4264 20874 4292 25162
rect 4356 22778 4384 29407
rect 4448 29306 4476 30087
rect 4620 30058 4672 30064
rect 4632 29850 4660 30058
rect 4528 29844 4580 29850
rect 4528 29786 4580 29792
rect 4620 29844 4672 29850
rect 4620 29786 4672 29792
rect 4540 29578 4568 29786
rect 4724 29730 4752 33106
rect 4988 33050 5040 33056
rect 5172 33108 5224 33114
rect 5172 33050 5224 33056
rect 4804 32972 4856 32978
rect 4804 32914 4856 32920
rect 4816 32434 4844 32914
rect 4804 32428 4856 32434
rect 4804 32370 4856 32376
rect 4816 32201 4844 32370
rect 4896 32224 4948 32230
rect 4802 32192 4858 32201
rect 4896 32166 4948 32172
rect 4802 32127 4858 32136
rect 4804 31340 4856 31346
rect 4804 31282 4856 31288
rect 4816 30394 4844 31282
rect 4908 31278 4936 32166
rect 4896 31272 4948 31278
rect 4896 31214 4948 31220
rect 4804 30388 4856 30394
rect 4804 30330 4856 30336
rect 4802 30288 4858 30297
rect 4802 30223 4858 30232
rect 4632 29702 4752 29730
rect 4528 29572 4580 29578
rect 4528 29514 4580 29520
rect 4436 29300 4488 29306
rect 4436 29242 4488 29248
rect 4436 28756 4488 28762
rect 4488 28716 4568 28744
rect 4436 28698 4488 28704
rect 4540 28014 4568 28716
rect 4632 28558 4660 29702
rect 4816 29510 4844 30223
rect 4804 29504 4856 29510
rect 4804 29446 4856 29452
rect 4712 29300 4764 29306
rect 4712 29242 4764 29248
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 4618 28384 4674 28393
rect 4618 28319 4674 28328
rect 4528 28008 4580 28014
rect 4528 27950 4580 27956
rect 4436 27328 4488 27334
rect 4436 27270 4488 27276
rect 4344 22772 4396 22778
rect 4344 22714 4396 22720
rect 4448 22710 4476 27270
rect 4540 26382 4568 27950
rect 4632 27470 4660 28319
rect 4620 27464 4672 27470
rect 4620 27406 4672 27412
rect 4724 27334 4752 29242
rect 4804 29096 4856 29102
rect 4802 29064 4804 29073
rect 4856 29064 4858 29073
rect 4802 28999 4858 29008
rect 4804 28960 4856 28966
rect 4804 28902 4856 28908
rect 4816 28082 4844 28902
rect 4908 28762 4936 31214
rect 5000 29306 5028 33050
rect 5170 33008 5226 33017
rect 5170 32943 5226 32952
rect 5184 32774 5212 32943
rect 5172 32768 5224 32774
rect 5172 32710 5224 32716
rect 5172 31748 5224 31754
rect 5172 31690 5224 31696
rect 5184 31521 5212 31690
rect 5170 31512 5226 31521
rect 5170 31447 5226 31456
rect 5080 31340 5132 31346
rect 5080 31282 5132 31288
rect 5092 30734 5120 31282
rect 5276 31226 5304 33390
rect 5368 32230 5396 36638
rect 5644 35766 5672 37964
rect 5736 36553 5764 40004
rect 5894 39196 6202 39205
rect 5894 39194 5900 39196
rect 5956 39194 5980 39196
rect 6036 39194 6060 39196
rect 6116 39194 6140 39196
rect 6196 39194 6202 39196
rect 5956 39142 5958 39194
rect 6138 39142 6140 39194
rect 5894 39140 5900 39142
rect 5956 39140 5980 39142
rect 6036 39140 6060 39142
rect 6116 39140 6140 39142
rect 6196 39140 6202 39142
rect 5894 39131 6202 39140
rect 5816 38752 5868 38758
rect 5816 38694 5868 38700
rect 5722 36544 5778 36553
rect 5722 36479 5778 36488
rect 5632 35760 5684 35766
rect 5632 35702 5684 35708
rect 5724 35624 5776 35630
rect 5724 35566 5776 35572
rect 5448 34740 5500 34746
rect 5448 34682 5500 34688
rect 5460 32978 5488 34682
rect 5630 34504 5686 34513
rect 5630 34439 5686 34448
rect 5540 33856 5592 33862
rect 5540 33798 5592 33804
rect 5448 32972 5500 32978
rect 5448 32914 5500 32920
rect 5552 32910 5580 33798
rect 5540 32904 5592 32910
rect 5540 32846 5592 32852
rect 5644 32842 5672 34439
rect 5632 32836 5684 32842
rect 5632 32778 5684 32784
rect 5446 32600 5502 32609
rect 5446 32535 5502 32544
rect 5460 32502 5488 32535
rect 5448 32496 5500 32502
rect 5448 32438 5500 32444
rect 5540 32428 5592 32434
rect 5540 32370 5592 32376
rect 5356 32224 5408 32230
rect 5356 32166 5408 32172
rect 5448 32224 5500 32230
rect 5448 32166 5500 32172
rect 5460 31890 5488 32166
rect 5448 31884 5500 31890
rect 5448 31826 5500 31832
rect 5356 31816 5408 31822
rect 5356 31758 5408 31764
rect 5368 31482 5396 31758
rect 5448 31748 5500 31754
rect 5448 31690 5500 31696
rect 5356 31476 5408 31482
rect 5356 31418 5408 31424
rect 5460 31226 5488 31690
rect 5552 31414 5580 32370
rect 5540 31408 5592 31414
rect 5540 31350 5592 31356
rect 5276 31198 5488 31226
rect 5080 30728 5132 30734
rect 5080 30670 5132 30676
rect 5092 30297 5120 30670
rect 5172 30592 5224 30598
rect 5172 30534 5224 30540
rect 5078 30288 5134 30297
rect 5184 30258 5212 30534
rect 5078 30223 5134 30232
rect 5172 30252 5224 30258
rect 5172 30194 5224 30200
rect 5276 30054 5304 31198
rect 5356 31136 5408 31142
rect 5408 31096 5488 31124
rect 5356 31078 5408 31084
rect 5356 30728 5408 30734
rect 5356 30670 5408 30676
rect 5368 30433 5396 30670
rect 5354 30424 5410 30433
rect 5354 30359 5410 30368
rect 5356 30184 5408 30190
rect 5460 30161 5488 31096
rect 5632 30932 5684 30938
rect 5632 30874 5684 30880
rect 5538 30288 5594 30297
rect 5538 30223 5594 30232
rect 5356 30126 5408 30132
rect 5446 30152 5502 30161
rect 5080 30048 5132 30054
rect 5080 29990 5132 29996
rect 5264 30048 5316 30054
rect 5264 29990 5316 29996
rect 4988 29300 5040 29306
rect 4988 29242 5040 29248
rect 4896 28756 4948 28762
rect 4896 28698 4948 28704
rect 4988 28416 5040 28422
rect 4988 28358 5040 28364
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4816 27418 4844 28018
rect 5000 27538 5028 28358
rect 5092 28257 5120 29990
rect 5264 29640 5316 29646
rect 5264 29582 5316 29588
rect 5172 29572 5224 29578
rect 5172 29514 5224 29520
rect 5078 28248 5134 28257
rect 5078 28183 5134 28192
rect 5080 28144 5132 28150
rect 5080 28086 5132 28092
rect 4988 27532 5040 27538
rect 4988 27474 5040 27480
rect 5092 27470 5120 28086
rect 5080 27464 5132 27470
rect 4816 27390 5028 27418
rect 5080 27406 5132 27412
rect 4712 27328 4764 27334
rect 4896 27328 4948 27334
rect 4712 27270 4764 27276
rect 4816 27276 4896 27282
rect 4816 27270 4948 27276
rect 4816 27254 4936 27270
rect 4816 26994 4844 27254
rect 4804 26988 4856 26994
rect 4804 26930 4856 26936
rect 4710 26888 4766 26897
rect 4710 26823 4766 26832
rect 4724 26382 4752 26823
rect 4816 26586 4844 26930
rect 4804 26580 4856 26586
rect 4804 26522 4856 26528
rect 4896 26580 4948 26586
rect 4896 26522 4948 26528
rect 4528 26376 4580 26382
rect 4528 26318 4580 26324
rect 4712 26376 4764 26382
rect 4712 26318 4764 26324
rect 4540 25906 4568 26318
rect 4528 25900 4580 25906
rect 4528 25842 4580 25848
rect 4804 25832 4856 25838
rect 4804 25774 4856 25780
rect 4528 25696 4580 25702
rect 4528 25638 4580 25644
rect 4540 24750 4568 25638
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4620 25220 4672 25226
rect 4620 25162 4672 25168
rect 4528 24744 4580 24750
rect 4528 24686 4580 24692
rect 4632 24410 4660 25162
rect 4724 24954 4752 25230
rect 4816 25226 4844 25774
rect 4804 25220 4856 25226
rect 4804 25162 4856 25168
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 4908 24818 4936 26522
rect 5000 26353 5028 27390
rect 5184 27112 5212 29514
rect 5276 27316 5304 29582
rect 5368 29050 5396 30126
rect 5446 30087 5502 30096
rect 5446 29336 5502 29345
rect 5446 29271 5502 29280
rect 5460 29238 5488 29271
rect 5448 29232 5500 29238
rect 5552 29209 5580 30223
rect 5448 29174 5500 29180
rect 5538 29200 5594 29209
rect 5538 29135 5594 29144
rect 5368 29022 5488 29050
rect 5460 28558 5488 29022
rect 5540 28688 5592 28694
rect 5540 28630 5592 28636
rect 5356 28552 5408 28558
rect 5356 28494 5408 28500
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5368 28150 5396 28494
rect 5356 28144 5408 28150
rect 5356 28086 5408 28092
rect 5356 27328 5408 27334
rect 5276 27288 5356 27316
rect 5356 27270 5408 27276
rect 5092 27084 5212 27112
rect 4986 26344 5042 26353
rect 4986 26279 5042 26288
rect 4988 26240 5040 26246
rect 4988 26182 5040 26188
rect 4712 24812 4764 24818
rect 4712 24754 4764 24760
rect 4804 24812 4856 24818
rect 4804 24754 4856 24760
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 4620 24404 4672 24410
rect 4620 24346 4672 24352
rect 4724 24342 4752 24754
rect 4816 24698 4844 24754
rect 4816 24670 4936 24698
rect 4908 24410 4936 24670
rect 4896 24404 4948 24410
rect 4896 24346 4948 24352
rect 4712 24336 4764 24342
rect 4618 24304 4674 24313
rect 4712 24278 4764 24284
rect 4618 24239 4674 24248
rect 4632 24206 4660 24239
rect 4620 24200 4672 24206
rect 4620 24142 4672 24148
rect 4526 22944 4582 22953
rect 4526 22879 4582 22888
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4448 22030 4476 22646
rect 4436 22024 4488 22030
rect 4436 21966 4488 21972
rect 4540 21729 4568 22879
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 4632 22250 4660 22714
rect 4804 22568 4856 22574
rect 4724 22528 4804 22556
rect 4724 22409 4752 22528
rect 4804 22510 4856 22516
rect 4710 22400 4766 22409
rect 4908 22386 4936 24346
rect 5000 22642 5028 26182
rect 5092 25684 5120 27084
rect 5368 26994 5396 27270
rect 5460 27062 5488 28494
rect 5448 27056 5500 27062
rect 5448 26998 5500 27004
rect 5172 26988 5224 26994
rect 5172 26930 5224 26936
rect 5356 26988 5408 26994
rect 5356 26930 5408 26936
rect 5184 26042 5212 26930
rect 5354 26888 5410 26897
rect 5354 26823 5356 26832
rect 5408 26823 5410 26832
rect 5356 26794 5408 26800
rect 5448 26512 5500 26518
rect 5448 26454 5500 26460
rect 5172 26036 5224 26042
rect 5172 25978 5224 25984
rect 5264 26036 5316 26042
rect 5264 25978 5316 25984
rect 5170 25936 5226 25945
rect 5170 25871 5172 25880
rect 5224 25871 5226 25880
rect 5172 25842 5224 25848
rect 5172 25696 5224 25702
rect 5092 25656 5172 25684
rect 5092 25158 5120 25656
rect 5172 25638 5224 25644
rect 5276 25344 5304 25978
rect 5184 25316 5304 25344
rect 5080 25152 5132 25158
rect 5080 25094 5132 25100
rect 5092 24206 5120 25094
rect 5080 24200 5132 24206
rect 5080 24142 5132 24148
rect 5080 24064 5132 24070
rect 5184 24041 5212 25316
rect 5262 25256 5318 25265
rect 5460 25242 5488 26454
rect 5552 26042 5580 28630
rect 5644 26246 5672 30874
rect 5736 28694 5764 35566
rect 5828 34626 5856 38694
rect 6276 38412 6328 38418
rect 6276 38354 6328 38360
rect 5894 38108 6202 38117
rect 5894 38106 5900 38108
rect 5956 38106 5980 38108
rect 6036 38106 6060 38108
rect 6116 38106 6140 38108
rect 6196 38106 6202 38108
rect 5956 38054 5958 38106
rect 6138 38054 6140 38106
rect 5894 38052 5900 38054
rect 5956 38052 5980 38054
rect 6036 38052 6060 38054
rect 6116 38052 6140 38054
rect 6196 38052 6202 38054
rect 5894 38043 6202 38052
rect 6288 37942 6316 38354
rect 6276 37936 6328 37942
rect 6276 37878 6328 37884
rect 5908 37800 5960 37806
rect 6380 37777 6408 41511
rect 6472 38010 6500 41670
rect 6564 41274 6592 42570
rect 6656 41818 6684 44540
rect 6736 43308 6788 43314
rect 6736 43250 6788 43256
rect 6644 41812 6696 41818
rect 6644 41754 6696 41760
rect 6748 41274 6776 43250
rect 6840 42362 6868 44540
rect 6920 43172 6972 43178
rect 6920 43114 6972 43120
rect 6932 42702 6960 43114
rect 6920 42696 6972 42702
rect 6920 42638 6972 42644
rect 7024 42634 7052 44540
rect 7208 43602 7236 44540
rect 7208 43574 7328 43602
rect 7196 43376 7248 43382
rect 7196 43318 7248 43324
rect 7012 42628 7064 42634
rect 7012 42570 7064 42576
rect 6828 42356 6880 42362
rect 6828 42298 6880 42304
rect 7104 42220 7156 42226
rect 7104 42162 7156 42168
rect 6920 42152 6972 42158
rect 6920 42094 6972 42100
rect 6932 41596 6960 42094
rect 7012 42084 7064 42090
rect 7012 42026 7064 42032
rect 7024 41818 7052 42026
rect 7116 41818 7144 42162
rect 7012 41812 7064 41818
rect 7012 41754 7064 41760
rect 7104 41812 7156 41818
rect 7104 41754 7156 41760
rect 7208 41750 7236 43318
rect 7300 42906 7328 43574
rect 7392 43450 7420 44540
rect 7380 43444 7432 43450
rect 7380 43386 7432 43392
rect 7380 43240 7432 43246
rect 7380 43182 7432 43188
rect 7288 42900 7340 42906
rect 7288 42842 7340 42848
rect 7196 41744 7248 41750
rect 7196 41686 7248 41692
rect 7196 41608 7248 41614
rect 6932 41568 7144 41596
rect 7012 41472 7064 41478
rect 7012 41414 7064 41420
rect 7116 41414 7144 41568
rect 7248 41568 7328 41596
rect 7196 41550 7248 41556
rect 6932 41386 7052 41414
rect 7116 41386 7236 41414
rect 6552 41268 6604 41274
rect 6552 41210 6604 41216
rect 6736 41268 6788 41274
rect 6736 41210 6788 41216
rect 6932 41206 6960 41386
rect 6920 41200 6972 41206
rect 6920 41142 6972 41148
rect 7208 41002 7236 41386
rect 7196 40996 7248 41002
rect 7196 40938 7248 40944
rect 7194 40624 7250 40633
rect 7116 40582 7194 40610
rect 6644 39432 6696 39438
rect 6644 39374 6696 39380
rect 6552 38888 6604 38894
rect 6552 38830 6604 38836
rect 6460 38004 6512 38010
rect 6460 37946 6512 37952
rect 6458 37904 6514 37913
rect 6458 37839 6514 37848
rect 5908 37742 5960 37748
rect 6366 37768 6422 37777
rect 5920 37330 5948 37742
rect 6366 37703 6422 37712
rect 6368 37664 6420 37670
rect 6368 37606 6420 37612
rect 5908 37324 5960 37330
rect 5908 37266 5960 37272
rect 6380 37194 6408 37606
rect 6276 37188 6328 37194
rect 6276 37130 6328 37136
rect 6368 37188 6420 37194
rect 6368 37130 6420 37136
rect 5894 37020 6202 37029
rect 5894 37018 5900 37020
rect 5956 37018 5980 37020
rect 6036 37018 6060 37020
rect 6116 37018 6140 37020
rect 6196 37018 6202 37020
rect 5956 36966 5958 37018
rect 6138 36966 6140 37018
rect 5894 36964 5900 36966
rect 5956 36964 5980 36966
rect 6036 36964 6060 36966
rect 6116 36964 6140 36966
rect 6196 36964 6202 36966
rect 5894 36955 6202 36964
rect 6288 36922 6316 37130
rect 6276 36916 6328 36922
rect 6276 36858 6328 36864
rect 6380 36802 6408 37130
rect 6288 36774 6408 36802
rect 5894 35932 6202 35941
rect 5894 35930 5900 35932
rect 5956 35930 5980 35932
rect 6036 35930 6060 35932
rect 6116 35930 6140 35932
rect 6196 35930 6202 35932
rect 5956 35878 5958 35930
rect 6138 35878 6140 35930
rect 5894 35876 5900 35878
rect 5956 35876 5980 35878
rect 6036 35876 6060 35878
rect 6116 35876 6140 35878
rect 6196 35876 6202 35878
rect 5894 35867 6202 35876
rect 5906 35184 5962 35193
rect 5906 35119 5962 35128
rect 5920 34950 5948 35119
rect 5908 34944 5960 34950
rect 5908 34886 5960 34892
rect 5894 34844 6202 34853
rect 5894 34842 5900 34844
rect 5956 34842 5980 34844
rect 6036 34842 6060 34844
rect 6116 34842 6140 34844
rect 6196 34842 6202 34844
rect 5956 34790 5958 34842
rect 6138 34790 6140 34842
rect 5894 34788 5900 34790
rect 5956 34788 5980 34790
rect 6036 34788 6060 34790
rect 6116 34788 6140 34790
rect 6196 34788 6202 34790
rect 5894 34779 6202 34788
rect 5828 34598 6040 34626
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5920 33844 5948 34478
rect 6012 34116 6040 34598
rect 6288 34218 6316 36774
rect 6472 36666 6500 37839
rect 6380 36638 6500 36666
rect 6380 35630 6408 36638
rect 6564 36174 6592 38830
rect 6656 38654 6684 39374
rect 6920 38888 6972 38894
rect 6920 38830 6972 38836
rect 6932 38654 6960 38830
rect 6656 38626 6776 38654
rect 6644 37868 6696 37874
rect 6644 37810 6696 37816
rect 6656 36854 6684 37810
rect 6748 37670 6776 38626
rect 6840 38626 6960 38654
rect 6736 37664 6788 37670
rect 6736 37606 6788 37612
rect 6734 37360 6790 37369
rect 6734 37295 6790 37304
rect 6748 37194 6776 37295
rect 6736 37188 6788 37194
rect 6736 37130 6788 37136
rect 6644 36848 6696 36854
rect 6696 36808 6776 36836
rect 6644 36790 6696 36796
rect 6552 36168 6604 36174
rect 6552 36110 6604 36116
rect 6644 36168 6696 36174
rect 6644 36110 6696 36116
rect 6368 35624 6420 35630
rect 6368 35566 6420 35572
rect 6460 35284 6512 35290
rect 6460 35226 6512 35232
rect 6288 34190 6408 34218
rect 6012 34088 6316 34116
rect 5828 33816 5948 33844
rect 5828 31686 5856 33816
rect 5894 33756 6202 33765
rect 5894 33754 5900 33756
rect 5956 33754 5980 33756
rect 6036 33754 6060 33756
rect 6116 33754 6140 33756
rect 6196 33754 6202 33756
rect 5956 33702 5958 33754
rect 6138 33702 6140 33754
rect 5894 33700 5900 33702
rect 5956 33700 5980 33702
rect 6036 33700 6060 33702
rect 6116 33700 6140 33702
rect 6196 33700 6202 33702
rect 5894 33691 6202 33700
rect 6288 33590 6316 34088
rect 6276 33584 6328 33590
rect 6276 33526 6328 33532
rect 6380 33402 6408 34190
rect 6288 33374 6408 33402
rect 5894 32668 6202 32677
rect 5894 32666 5900 32668
rect 5956 32666 5980 32668
rect 6036 32666 6060 32668
rect 6116 32666 6140 32668
rect 6196 32666 6202 32668
rect 5956 32614 5958 32666
rect 6138 32614 6140 32666
rect 5894 32612 5900 32614
rect 5956 32612 5980 32614
rect 6036 32612 6060 32614
rect 6116 32612 6140 32614
rect 6196 32612 6202 32614
rect 5894 32603 6202 32612
rect 6288 32065 6316 33374
rect 6472 32910 6500 35226
rect 6564 34241 6592 36110
rect 6550 34232 6606 34241
rect 6550 34167 6606 34176
rect 6552 34128 6604 34134
rect 6552 34070 6604 34076
rect 6460 32904 6512 32910
rect 6460 32846 6512 32852
rect 6368 32836 6420 32842
rect 6368 32778 6420 32784
rect 6274 32056 6330 32065
rect 6274 31991 6330 32000
rect 6288 31890 6316 31991
rect 6276 31884 6328 31890
rect 6276 31826 6328 31832
rect 6276 31748 6328 31754
rect 6276 31690 6328 31696
rect 5816 31680 5868 31686
rect 5816 31622 5868 31628
rect 5828 31113 5856 31622
rect 5894 31580 6202 31589
rect 5894 31578 5900 31580
rect 5956 31578 5980 31580
rect 6036 31578 6060 31580
rect 6116 31578 6140 31580
rect 6196 31578 6202 31580
rect 5956 31526 5958 31578
rect 6138 31526 6140 31578
rect 5894 31524 5900 31526
rect 5956 31524 5980 31526
rect 6036 31524 6060 31526
rect 6116 31524 6140 31526
rect 6196 31524 6202 31526
rect 5894 31515 6202 31524
rect 6288 31385 6316 31690
rect 6274 31376 6330 31385
rect 6274 31311 6330 31320
rect 5814 31104 5870 31113
rect 5814 31039 5870 31048
rect 5894 30492 6202 30501
rect 5894 30490 5900 30492
rect 5956 30490 5980 30492
rect 6036 30490 6060 30492
rect 6116 30490 6140 30492
rect 6196 30490 6202 30492
rect 5956 30438 5958 30490
rect 6138 30438 6140 30490
rect 5894 30436 5900 30438
rect 5956 30436 5980 30438
rect 6036 30436 6060 30438
rect 6116 30436 6140 30438
rect 6196 30436 6202 30438
rect 5894 30427 6202 30436
rect 6380 29764 6408 32778
rect 6564 32348 6592 34070
rect 6656 33998 6684 36110
rect 6748 36038 6776 36808
rect 6840 36156 6868 38626
rect 6920 37120 6972 37126
rect 6920 37062 6972 37068
rect 6932 36378 6960 37062
rect 7012 36576 7064 36582
rect 7012 36518 7064 36524
rect 6920 36372 6972 36378
rect 6920 36314 6972 36320
rect 6920 36168 6972 36174
rect 6840 36128 6920 36156
rect 6920 36110 6972 36116
rect 6736 36032 6788 36038
rect 6736 35974 6788 35980
rect 6736 35488 6788 35494
rect 6736 35430 6788 35436
rect 6748 35086 6776 35430
rect 6736 35080 6788 35086
rect 6736 35022 6788 35028
rect 7024 35018 7052 36518
rect 6920 35012 6972 35018
rect 6920 34954 6972 34960
rect 7012 35012 7064 35018
rect 7012 34954 7064 34960
rect 6828 34944 6880 34950
rect 6828 34886 6880 34892
rect 6736 34740 6788 34746
rect 6736 34682 6788 34688
rect 6748 33998 6776 34682
rect 6840 34134 6868 34886
rect 6828 34128 6880 34134
rect 6828 34070 6880 34076
rect 6644 33992 6696 33998
rect 6644 33934 6696 33940
rect 6736 33992 6788 33998
rect 6736 33934 6788 33940
rect 6656 33046 6684 33934
rect 6748 33833 6776 33934
rect 6734 33824 6790 33833
rect 6734 33759 6790 33768
rect 6828 33584 6880 33590
rect 6828 33526 6880 33532
rect 6736 33312 6788 33318
rect 6736 33254 6788 33260
rect 6644 33040 6696 33046
rect 6644 32982 6696 32988
rect 6644 32904 6696 32910
rect 6644 32846 6696 32852
rect 6472 32320 6592 32348
rect 6380 29736 6433 29764
rect 6276 29640 6328 29646
rect 6196 29600 6276 29628
rect 6196 29492 6224 29600
rect 6405 29594 6433 29736
rect 6276 29582 6328 29588
rect 5828 29464 6224 29492
rect 6380 29566 6433 29594
rect 6274 29472 6330 29481
rect 5724 28688 5776 28694
rect 5724 28630 5776 28636
rect 5724 28552 5776 28558
rect 5724 28494 5776 28500
rect 5632 26240 5684 26246
rect 5632 26182 5684 26188
rect 5540 26036 5592 26042
rect 5540 25978 5592 25984
rect 5632 26036 5684 26042
rect 5632 25978 5684 25984
rect 5644 25294 5672 25978
rect 5736 25294 5764 28494
rect 5828 27470 5856 29464
rect 5894 29404 6202 29413
rect 6274 29407 6330 29416
rect 5894 29402 5900 29404
rect 5956 29402 5980 29404
rect 6036 29402 6060 29404
rect 6116 29402 6140 29404
rect 6196 29402 6202 29404
rect 5956 29350 5958 29402
rect 6138 29350 6140 29402
rect 5894 29348 5900 29350
rect 5956 29348 5980 29350
rect 6036 29348 6060 29350
rect 6116 29348 6140 29350
rect 6196 29348 6202 29350
rect 5894 29339 6202 29348
rect 5894 28316 6202 28325
rect 5894 28314 5900 28316
rect 5956 28314 5980 28316
rect 6036 28314 6060 28316
rect 6116 28314 6140 28316
rect 6196 28314 6202 28316
rect 5956 28262 5958 28314
rect 6138 28262 6140 28314
rect 5894 28260 5900 28262
rect 5956 28260 5980 28262
rect 6036 28260 6060 28262
rect 6116 28260 6140 28262
rect 6196 28260 6202 28262
rect 5894 28251 6202 28260
rect 5908 28212 5960 28218
rect 5908 28154 5960 28160
rect 5920 28121 5948 28154
rect 5906 28112 5962 28121
rect 5906 28047 5962 28056
rect 5816 27464 5868 27470
rect 5816 27406 5868 27412
rect 5894 27228 6202 27237
rect 5894 27226 5900 27228
rect 5956 27226 5980 27228
rect 6036 27226 6060 27228
rect 6116 27226 6140 27228
rect 6196 27226 6202 27228
rect 5956 27174 5958 27226
rect 6138 27174 6140 27226
rect 5894 27172 5900 27174
rect 5956 27172 5980 27174
rect 6036 27172 6060 27174
rect 6116 27172 6140 27174
rect 6196 27172 6202 27174
rect 5894 27163 6202 27172
rect 5816 26988 5868 26994
rect 5816 26930 5868 26936
rect 5828 26042 5856 26930
rect 6288 26217 6316 29407
rect 6380 27713 6408 29566
rect 6472 28801 6500 32320
rect 6552 32224 6604 32230
rect 6552 32166 6604 32172
rect 6564 30297 6592 32166
rect 6550 30288 6606 30297
rect 6550 30223 6606 30232
rect 6656 30122 6684 32846
rect 6748 32774 6776 33254
rect 6736 32768 6788 32774
rect 6736 32710 6788 32716
rect 6748 30734 6776 32710
rect 6736 30728 6788 30734
rect 6736 30670 6788 30676
rect 6644 30116 6696 30122
rect 6644 30058 6696 30064
rect 6552 30048 6604 30054
rect 6840 30002 6868 33526
rect 6932 32978 6960 34954
rect 6920 32972 6972 32978
rect 6920 32914 6972 32920
rect 7024 32910 7052 34954
rect 7116 34241 7144 40582
rect 7194 40559 7250 40568
rect 7300 38554 7328 41568
rect 7392 41274 7420 43182
rect 7472 42900 7524 42906
rect 7472 42842 7524 42848
rect 7484 41585 7512 42842
rect 7576 42362 7604 44540
rect 7564 42356 7616 42362
rect 7564 42298 7616 42304
rect 7760 42158 7788 44540
rect 7944 42752 7972 44540
rect 8024 42764 8076 42770
rect 7944 42724 8024 42752
rect 8024 42706 8076 42712
rect 8024 42628 8076 42634
rect 8024 42570 8076 42576
rect 8036 42362 8064 42570
rect 8128 42362 8156 44540
rect 8312 43058 8340 44540
rect 8496 43466 8524 44540
rect 8404 43438 8524 43466
rect 8680 43450 8708 44540
rect 8668 43444 8720 43450
rect 8404 43382 8432 43438
rect 8668 43386 8720 43392
rect 8392 43376 8444 43382
rect 8392 43318 8444 43324
rect 8576 43376 8628 43382
rect 8576 43318 8628 43324
rect 8588 43110 8616 43318
rect 8760 43240 8812 43246
rect 8760 43182 8812 43188
rect 8220 43030 8340 43058
rect 8576 43104 8628 43110
rect 8576 43046 8628 43052
rect 8220 42752 8248 43030
rect 8367 43004 8675 43013
rect 8367 43002 8373 43004
rect 8429 43002 8453 43004
rect 8509 43002 8533 43004
rect 8589 43002 8613 43004
rect 8669 43002 8675 43004
rect 8429 42950 8431 43002
rect 8611 42950 8613 43002
rect 8367 42948 8373 42950
rect 8429 42948 8453 42950
rect 8509 42948 8533 42950
rect 8589 42948 8613 42950
rect 8669 42948 8675 42950
rect 8367 42939 8675 42948
rect 8300 42764 8352 42770
rect 8220 42724 8300 42752
rect 8300 42706 8352 42712
rect 8024 42356 8076 42362
rect 8024 42298 8076 42304
rect 8116 42356 8168 42362
rect 8116 42298 8168 42304
rect 8208 42220 8260 42226
rect 8208 42162 8260 42168
rect 7748 42152 7800 42158
rect 7748 42094 7800 42100
rect 8220 41818 8248 42162
rect 8367 41916 8675 41925
rect 8367 41914 8373 41916
rect 8429 41914 8453 41916
rect 8509 41914 8533 41916
rect 8589 41914 8613 41916
rect 8669 41914 8675 41916
rect 8429 41862 8431 41914
rect 8611 41862 8613 41914
rect 8367 41860 8373 41862
rect 8429 41860 8453 41862
rect 8509 41860 8533 41862
rect 8589 41860 8613 41862
rect 8669 41860 8675 41862
rect 8367 41851 8675 41860
rect 8208 41812 8260 41818
rect 8208 41754 8260 41760
rect 8772 41750 8800 43182
rect 8864 42537 8892 44540
rect 9048 43314 9076 44540
rect 9036 43308 9088 43314
rect 9036 43250 9088 43256
rect 8944 43172 8996 43178
rect 8944 43114 8996 43120
rect 8850 42528 8906 42537
rect 8850 42463 8906 42472
rect 8956 42362 8984 43114
rect 9036 43104 9088 43110
rect 9036 43046 9088 43052
rect 8944 42356 8996 42362
rect 8944 42298 8996 42304
rect 8852 42220 8904 42226
rect 8852 42162 8904 42168
rect 8944 42220 8996 42226
rect 8944 42162 8996 42168
rect 8864 42129 8892 42162
rect 8850 42120 8906 42129
rect 8850 42055 8906 42064
rect 8760 41744 8812 41750
rect 8760 41686 8812 41692
rect 7748 41608 7800 41614
rect 7470 41576 7526 41585
rect 7748 41550 7800 41556
rect 8760 41608 8812 41614
rect 8760 41550 8812 41556
rect 7470 41511 7526 41520
rect 7380 41268 7432 41274
rect 7380 41210 7432 41216
rect 7564 40588 7616 40594
rect 7564 40530 7616 40536
rect 7576 39930 7604 40530
rect 7656 40384 7708 40390
rect 7656 40326 7708 40332
rect 7668 40186 7696 40326
rect 7656 40180 7708 40186
rect 7656 40122 7708 40128
rect 7576 39902 7696 39930
rect 7564 39840 7616 39846
rect 7564 39782 7616 39788
rect 7576 39642 7604 39782
rect 7564 39636 7616 39642
rect 7564 39578 7616 39584
rect 7380 39568 7432 39574
rect 7380 39510 7432 39516
rect 7392 38894 7420 39510
rect 7380 38888 7432 38894
rect 7380 38830 7432 38836
rect 7288 38548 7340 38554
rect 7288 38490 7340 38496
rect 7378 38040 7434 38049
rect 7378 37975 7434 37984
rect 7392 37874 7420 37975
rect 7380 37868 7432 37874
rect 7380 37810 7432 37816
rect 7472 37664 7524 37670
rect 7472 37606 7524 37612
rect 7484 37330 7512 37606
rect 7472 37324 7524 37330
rect 7472 37266 7524 37272
rect 7472 36780 7524 36786
rect 7472 36722 7524 36728
rect 7286 36680 7342 36689
rect 7286 36615 7342 36624
rect 7380 36644 7432 36650
rect 7300 35057 7328 36615
rect 7380 36586 7432 36592
rect 7286 35048 7342 35057
rect 7286 34983 7342 34992
rect 7392 34678 7420 36586
rect 7484 36378 7512 36722
rect 7564 36712 7616 36718
rect 7564 36654 7616 36660
rect 7472 36372 7524 36378
rect 7472 36314 7524 36320
rect 7576 36242 7604 36654
rect 7564 36236 7616 36242
rect 7564 36178 7616 36184
rect 7472 36168 7524 36174
rect 7472 36110 7524 36116
rect 7288 34672 7340 34678
rect 7288 34614 7340 34620
rect 7380 34672 7432 34678
rect 7380 34614 7432 34620
rect 7102 34232 7158 34241
rect 7102 34167 7158 34176
rect 7104 34128 7156 34134
rect 7104 34070 7156 34076
rect 7116 33386 7144 34070
rect 7196 33652 7248 33658
rect 7196 33594 7248 33600
rect 7104 33380 7156 33386
rect 7104 33322 7156 33328
rect 7104 32972 7156 32978
rect 7104 32914 7156 32920
rect 7012 32904 7064 32910
rect 7012 32846 7064 32852
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6932 32434 6960 32710
rect 7116 32434 7144 32914
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 7104 32428 7156 32434
rect 7104 32370 7156 32376
rect 6920 32020 6972 32026
rect 6972 31980 7052 32008
rect 6920 31962 6972 31968
rect 7024 31929 7052 31980
rect 7010 31920 7066 31929
rect 7010 31855 7066 31864
rect 7116 31822 7144 32370
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 7010 31648 7066 31657
rect 7010 31583 7066 31592
rect 6918 31240 6974 31249
rect 6918 31175 6974 31184
rect 6932 30326 6960 31175
rect 7024 30410 7052 31583
rect 7116 31346 7144 31758
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 7102 31240 7158 31249
rect 7102 31175 7104 31184
rect 7156 31175 7158 31184
rect 7104 31146 7156 31152
rect 7208 31142 7236 33594
rect 7300 33436 7328 34614
rect 7484 34066 7512 36110
rect 7564 34944 7616 34950
rect 7564 34886 7616 34892
rect 7576 34542 7604 34886
rect 7564 34536 7616 34542
rect 7564 34478 7616 34484
rect 7668 34388 7696 39902
rect 7760 35873 7788 41550
rect 8772 41414 8800 41550
rect 8772 41386 8892 41414
rect 7932 41132 7984 41138
rect 7932 41074 7984 41080
rect 7944 40089 7972 41074
rect 8760 41064 8812 41070
rect 8760 41006 8812 41012
rect 8367 40828 8675 40837
rect 8367 40826 8373 40828
rect 8429 40826 8453 40828
rect 8509 40826 8533 40828
rect 8589 40826 8613 40828
rect 8669 40826 8675 40828
rect 8429 40774 8431 40826
rect 8611 40774 8613 40826
rect 8367 40772 8373 40774
rect 8429 40772 8453 40774
rect 8509 40772 8533 40774
rect 8589 40772 8613 40774
rect 8669 40772 8675 40774
rect 8367 40763 8675 40772
rect 7930 40080 7986 40089
rect 7840 40054 7892 40060
rect 7930 40015 7986 40024
rect 7840 39996 7892 40002
rect 7852 39001 7880 39996
rect 7932 39840 7984 39846
rect 7932 39782 7984 39788
rect 7838 38992 7894 39001
rect 7944 38962 7972 39782
rect 8367 39740 8675 39749
rect 8367 39738 8373 39740
rect 8429 39738 8453 39740
rect 8509 39738 8533 39740
rect 8589 39738 8613 39740
rect 8669 39738 8675 39740
rect 8429 39686 8431 39738
rect 8611 39686 8613 39738
rect 8367 39684 8373 39686
rect 8429 39684 8453 39686
rect 8509 39684 8533 39686
rect 8589 39684 8613 39686
rect 8669 39684 8675 39686
rect 8367 39675 8675 39684
rect 7838 38927 7894 38936
rect 7932 38956 7984 38962
rect 7932 38898 7984 38904
rect 7840 38888 7892 38894
rect 7840 38830 7892 38836
rect 7746 35864 7802 35873
rect 7746 35799 7802 35808
rect 7748 35284 7800 35290
rect 7748 35226 7800 35232
rect 7760 34610 7788 35226
rect 7852 34610 7880 38830
rect 8367 38652 8675 38661
rect 8367 38650 8373 38652
rect 8429 38650 8453 38652
rect 8509 38650 8533 38652
rect 8589 38650 8613 38652
rect 8669 38650 8675 38652
rect 8429 38598 8431 38650
rect 8611 38598 8613 38650
rect 8367 38596 8373 38598
rect 8429 38596 8453 38598
rect 8509 38596 8533 38598
rect 8589 38596 8613 38598
rect 8669 38596 8675 38598
rect 8367 38587 8675 38596
rect 8772 37913 8800 41006
rect 8758 37904 8814 37913
rect 8758 37839 8814 37848
rect 7932 37664 7984 37670
rect 7932 37606 7984 37612
rect 8760 37664 8812 37670
rect 8760 37606 8812 37612
rect 7944 36242 7972 37606
rect 8367 37564 8675 37573
rect 8367 37562 8373 37564
rect 8429 37562 8453 37564
rect 8509 37562 8533 37564
rect 8589 37562 8613 37564
rect 8669 37562 8675 37564
rect 8429 37510 8431 37562
rect 8611 37510 8613 37562
rect 8367 37508 8373 37510
rect 8429 37508 8453 37510
rect 8509 37508 8533 37510
rect 8589 37508 8613 37510
rect 8669 37508 8675 37510
rect 8367 37499 8675 37508
rect 8484 37120 8536 37126
rect 8484 37062 8536 37068
rect 8496 36718 8524 37062
rect 8772 36786 8800 37606
rect 8760 36780 8812 36786
rect 8760 36722 8812 36728
rect 8024 36712 8076 36718
rect 8024 36654 8076 36660
rect 8484 36712 8536 36718
rect 8484 36654 8536 36660
rect 7932 36236 7984 36242
rect 7932 36178 7984 36184
rect 7932 35080 7984 35086
rect 7932 35022 7984 35028
rect 7748 34604 7800 34610
rect 7748 34546 7800 34552
rect 7840 34604 7892 34610
rect 7840 34546 7892 34552
rect 7852 34490 7880 34546
rect 7576 34360 7696 34388
rect 7760 34462 7880 34490
rect 7472 34060 7524 34066
rect 7472 34002 7524 34008
rect 7576 33640 7604 34360
rect 7656 34060 7708 34066
rect 7760 34048 7788 34462
rect 7944 34241 7972 35022
rect 8036 34746 8064 36654
rect 8206 36544 8262 36553
rect 8206 36479 8262 36488
rect 8024 34740 8076 34746
rect 8024 34682 8076 34688
rect 8220 34649 8248 36479
rect 8367 36476 8675 36485
rect 8367 36474 8373 36476
rect 8429 36474 8453 36476
rect 8509 36474 8533 36476
rect 8589 36474 8613 36476
rect 8669 36474 8675 36476
rect 8429 36422 8431 36474
rect 8611 36422 8613 36474
rect 8367 36420 8373 36422
rect 8429 36420 8453 36422
rect 8509 36420 8533 36422
rect 8589 36420 8613 36422
rect 8669 36420 8675 36422
rect 8367 36411 8675 36420
rect 8760 36100 8812 36106
rect 8760 36042 8812 36048
rect 8367 35388 8675 35397
rect 8367 35386 8373 35388
rect 8429 35386 8453 35388
rect 8509 35386 8533 35388
rect 8589 35386 8613 35388
rect 8669 35386 8675 35388
rect 8429 35334 8431 35386
rect 8611 35334 8613 35386
rect 8367 35332 8373 35334
rect 8429 35332 8453 35334
rect 8509 35332 8533 35334
rect 8589 35332 8613 35334
rect 8669 35332 8675 35334
rect 8367 35323 8675 35332
rect 8772 35222 8800 36042
rect 8760 35216 8812 35222
rect 8760 35158 8812 35164
rect 8760 35080 8812 35086
rect 8760 35022 8812 35028
rect 8300 34672 8352 34678
rect 8022 34640 8078 34649
rect 8206 34640 8262 34649
rect 8078 34598 8156 34626
rect 8022 34575 8078 34584
rect 7930 34232 7986 34241
rect 7930 34167 7986 34176
rect 8128 34066 8156 34598
rect 8300 34614 8352 34620
rect 8206 34575 8262 34584
rect 8312 34354 8340 34614
rect 8220 34326 8340 34354
rect 8220 34218 8248 34326
rect 8367 34300 8675 34309
rect 8367 34298 8373 34300
rect 8429 34298 8453 34300
rect 8509 34298 8533 34300
rect 8589 34298 8613 34300
rect 8669 34298 8675 34300
rect 8429 34246 8431 34298
rect 8611 34246 8613 34298
rect 8367 34244 8373 34246
rect 8429 34244 8453 34246
rect 8509 34244 8533 34246
rect 8589 34244 8613 34246
rect 8669 34244 8675 34246
rect 8367 34235 8675 34244
rect 8220 34190 8340 34218
rect 7708 34020 7788 34048
rect 7656 34002 7708 34008
rect 7656 33652 7708 33658
rect 7576 33612 7656 33640
rect 7656 33594 7708 33600
rect 7564 33516 7616 33522
rect 7564 33458 7616 33464
rect 7380 33448 7432 33454
rect 7300 33408 7380 33436
rect 7432 33408 7512 33436
rect 7380 33390 7432 33396
rect 7288 33040 7340 33046
rect 7288 32982 7340 32988
rect 7196 31136 7248 31142
rect 7196 31078 7248 31084
rect 7194 30696 7250 30705
rect 7194 30631 7196 30640
rect 7248 30631 7250 30640
rect 7196 30602 7248 30608
rect 7024 30382 7144 30410
rect 6920 30320 6972 30326
rect 6920 30262 6972 30268
rect 7012 30320 7064 30326
rect 7012 30262 7064 30268
rect 6552 29990 6604 29996
rect 6458 28792 6514 28801
rect 6458 28727 6514 28736
rect 6564 28676 6592 29990
rect 6656 29974 6868 30002
rect 6656 28778 6684 29974
rect 6920 29844 6972 29850
rect 6920 29786 6972 29792
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6748 28966 6776 29650
rect 6932 29458 6960 29786
rect 6840 29430 6960 29458
rect 6736 28960 6788 28966
rect 6736 28902 6788 28908
rect 6656 28750 6776 28778
rect 6840 28762 6868 29430
rect 7024 29034 7052 30262
rect 7116 29238 7144 30382
rect 7196 30388 7248 30394
rect 7196 30330 7248 30336
rect 7208 29714 7236 30330
rect 7196 29708 7248 29714
rect 7196 29650 7248 29656
rect 7196 29504 7248 29510
rect 7196 29446 7248 29452
rect 7208 29238 7236 29446
rect 7104 29232 7156 29238
rect 7104 29174 7156 29180
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 6920 29028 6972 29034
rect 6920 28970 6972 28976
rect 7012 29028 7064 29034
rect 7012 28970 7064 28976
rect 6932 28762 6960 28970
rect 6564 28648 6684 28676
rect 6460 28552 6512 28558
rect 6460 28494 6512 28500
rect 6552 28552 6604 28558
rect 6552 28494 6604 28500
rect 6366 27704 6422 27713
rect 6366 27639 6422 27648
rect 6368 27464 6420 27470
rect 6368 27406 6420 27412
rect 6274 26208 6330 26217
rect 5894 26140 6202 26149
rect 6274 26143 6330 26152
rect 5894 26138 5900 26140
rect 5956 26138 5980 26140
rect 6036 26138 6060 26140
rect 6116 26138 6140 26140
rect 6196 26138 6202 26140
rect 5956 26086 5958 26138
rect 6138 26086 6140 26138
rect 5894 26084 5900 26086
rect 5956 26084 5980 26086
rect 6036 26084 6060 26086
rect 6116 26084 6140 26086
rect 6196 26084 6202 26086
rect 5894 26075 6202 26084
rect 5816 26036 5868 26042
rect 5816 25978 5868 25984
rect 6276 26036 6328 26042
rect 6276 25978 6328 25984
rect 5816 25696 5868 25702
rect 5816 25638 5868 25644
rect 5828 25498 5856 25638
rect 5816 25492 5868 25498
rect 5816 25434 5868 25440
rect 5262 25191 5318 25200
rect 5368 25214 5488 25242
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5724 25288 5776 25294
rect 5724 25230 5776 25236
rect 5276 25158 5304 25191
rect 5264 25152 5316 25158
rect 5264 25094 5316 25100
rect 5264 24812 5316 24818
rect 5264 24754 5316 24760
rect 5276 24274 5304 24754
rect 5264 24268 5316 24274
rect 5264 24210 5316 24216
rect 5080 24006 5132 24012
rect 5170 24032 5226 24041
rect 5092 23730 5120 24006
rect 5170 23967 5226 23976
rect 5170 23896 5226 23905
rect 5170 23831 5226 23840
rect 5184 23730 5212 23831
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 5172 23724 5224 23730
rect 5172 23666 5224 23672
rect 5172 23520 5224 23526
rect 5172 23462 5224 23468
rect 5184 22982 5212 23462
rect 5368 23322 5396 25214
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 5460 24818 5488 25094
rect 5538 24848 5594 24857
rect 5448 24812 5500 24818
rect 5538 24783 5594 24792
rect 5448 24754 5500 24760
rect 5552 24313 5580 24783
rect 5538 24304 5594 24313
rect 5538 24239 5594 24248
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5356 23316 5408 23322
rect 5356 23258 5408 23264
rect 5264 23248 5316 23254
rect 5264 23190 5316 23196
rect 5172 22976 5224 22982
rect 5172 22918 5224 22924
rect 5172 22704 5224 22710
rect 5172 22646 5224 22652
rect 4988 22636 5040 22642
rect 4988 22578 5040 22584
rect 4710 22335 4766 22344
rect 4816 22358 4936 22386
rect 4632 22222 4752 22250
rect 4724 21894 4752 22222
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4526 21720 4582 21729
rect 4526 21655 4582 21664
rect 4436 21548 4488 21554
rect 4436 21490 4488 21496
rect 4252 20868 4304 20874
rect 4252 20810 4304 20816
rect 4264 19938 4292 20810
rect 4448 20330 4476 21490
rect 4620 21344 4672 21350
rect 4724 21321 4752 21830
rect 4620 21286 4672 21292
rect 4710 21312 4766 21321
rect 4632 20618 4660 21286
rect 4710 21247 4766 21256
rect 4632 20590 4752 20618
rect 4620 20528 4672 20534
rect 4540 20488 4620 20516
rect 4436 20324 4488 20330
rect 4436 20266 4488 20272
rect 4264 19910 4476 19938
rect 4158 19816 4214 19825
rect 4158 19751 4214 19760
rect 4252 19780 4304 19786
rect 3988 18414 4108 18442
rect 3976 18352 4028 18358
rect 3976 18294 4028 18300
rect 3792 18284 3844 18290
rect 3792 18226 3844 18232
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3804 18193 3832 18226
rect 3790 18184 3846 18193
rect 3790 18119 3846 18128
rect 3712 18040 3832 18068
rect 3422 17980 3730 17989
rect 3422 17978 3428 17980
rect 3484 17978 3508 17980
rect 3564 17978 3588 17980
rect 3644 17978 3668 17980
rect 3724 17978 3730 17980
rect 3484 17926 3486 17978
rect 3666 17926 3668 17978
rect 3422 17924 3428 17926
rect 3484 17924 3508 17926
rect 3564 17924 3588 17926
rect 3644 17924 3668 17926
rect 3724 17924 3730 17926
rect 3422 17915 3730 17924
rect 3514 17776 3570 17785
rect 3160 17734 3280 17762
rect 3344 17734 3464 17762
rect 3148 17672 3200 17678
rect 3148 17614 3200 17620
rect 2872 17128 2924 17134
rect 2608 17054 2728 17082
rect 2872 17070 2924 17076
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2594 16960 2650 16969
rect 2594 16895 2650 16904
rect 2502 16552 2558 16561
rect 2502 16487 2558 16496
rect 2516 16114 2544 16487
rect 2504 16108 2556 16114
rect 2504 16050 2556 16056
rect 2608 14414 2636 16895
rect 2700 16794 2728 17054
rect 2780 16992 2832 16998
rect 2780 16934 2832 16940
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 2686 16688 2742 16697
rect 2686 16623 2742 16632
rect 2700 15366 2728 16623
rect 2792 16114 2820 16934
rect 2884 16402 2912 17070
rect 2964 17060 3016 17066
rect 2964 17002 3016 17008
rect 2976 16590 3004 17002
rect 3054 16824 3110 16833
rect 3054 16759 3110 16768
rect 3068 16726 3096 16759
rect 3056 16720 3108 16726
rect 3056 16662 3108 16668
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2884 16374 3004 16402
rect 2870 16144 2926 16153
rect 2780 16108 2832 16114
rect 2870 16079 2926 16088
rect 2780 16050 2832 16056
rect 2884 15994 2912 16079
rect 2792 15966 2912 15994
rect 2792 15502 2820 15966
rect 2780 15496 2832 15502
rect 2780 15438 2832 15444
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2688 15088 2740 15094
rect 2688 15030 2740 15036
rect 2700 14657 2728 15030
rect 2686 14648 2742 14657
rect 2686 14583 2742 14592
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 13870 2544 14214
rect 2594 14104 2650 14113
rect 2594 14039 2650 14048
rect 2504 13864 2556 13870
rect 2504 13806 2556 13812
rect 2516 13297 2544 13806
rect 2502 13288 2558 13297
rect 2502 13223 2558 13232
rect 2608 12646 2636 14039
rect 2596 12640 2648 12646
rect 2596 12582 2648 12588
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2594 12200 2650 12209
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2412 12164 2464 12170
rect 2594 12135 2650 12144
rect 2412 12106 2464 12112
rect 2332 11762 2360 12106
rect 2608 11830 2636 12135
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2226 10840 2282 10849
rect 2226 10775 2282 10784
rect 2228 10736 2280 10742
rect 2332 10724 2360 11154
rect 2504 11144 2556 11150
rect 2502 11112 2504 11121
rect 2556 11112 2558 11121
rect 2502 11047 2558 11056
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2502 10976 2558 10985
rect 2280 10696 2360 10724
rect 2228 10678 2280 10684
rect 2226 10568 2282 10577
rect 2226 10503 2282 10512
rect 2240 9926 2268 10503
rect 2318 10432 2374 10441
rect 2318 10367 2374 10376
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2044 8968 2096 8974
rect 2044 8910 2096 8916
rect 2042 8664 2098 8673
rect 2042 8599 2098 8608
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1872 7942 1992 7970
rect 1858 7848 1914 7857
rect 1858 7783 1860 7792
rect 1912 7783 1914 7792
rect 1860 7754 1912 7760
rect 1872 7410 1900 7754
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1636 6412 1716 6440
rect 1584 6394 1636 6400
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1688 4434 1716 5578
rect 1780 4622 1808 6598
rect 1858 6352 1914 6361
rect 1858 6287 1914 6296
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1688 4406 1808 4434
rect 1504 4126 1624 4154
rect 1596 3194 1624 4126
rect 1780 3534 1808 4406
rect 1872 3942 1900 6287
rect 1964 5681 1992 7942
rect 2056 7886 2084 8599
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2042 7440 2098 7449
rect 2042 7375 2098 7384
rect 2056 7002 2084 7375
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2148 6390 2176 9318
rect 2240 8974 2268 9862
rect 2332 9178 2360 10367
rect 2424 9654 2452 10950
rect 2502 10911 2558 10920
rect 2516 10810 2544 10911
rect 2504 10804 2556 10810
rect 2504 10746 2556 10752
rect 2594 10296 2650 10305
rect 2516 10254 2594 10282
rect 2412 9648 2464 9654
rect 2412 9590 2464 9596
rect 2320 9172 2372 9178
rect 2320 9114 2372 9120
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2516 8838 2544 10254
rect 2594 10231 2650 10240
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2504 8832 2556 8838
rect 2318 8800 2374 8809
rect 2504 8774 2556 8780
rect 2318 8735 2374 8744
rect 2226 8528 2282 8537
rect 2226 8463 2282 8472
rect 2240 7478 2268 8463
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2226 7032 2282 7041
rect 2226 6967 2282 6976
rect 2240 6866 2268 6967
rect 2228 6860 2280 6866
rect 2228 6802 2280 6808
rect 2226 6760 2282 6769
rect 2226 6695 2282 6704
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 2044 6316 2096 6322
rect 2044 6258 2096 6264
rect 1950 5672 2006 5681
rect 1950 5607 2006 5616
rect 1952 5228 2004 5234
rect 1952 5170 2004 5176
rect 1964 4554 1992 5170
rect 2056 4826 2084 6258
rect 2136 5228 2188 5234
rect 2240 5216 2268 6695
rect 2332 6458 2360 8735
rect 2516 8566 2544 8774
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2410 8392 2466 8401
rect 2410 8327 2466 8336
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2318 6216 2374 6225
rect 2318 6151 2374 6160
rect 2332 5234 2360 6151
rect 2424 5710 2452 8327
rect 2504 8288 2556 8294
rect 2504 8230 2556 8236
rect 2516 6780 2544 8230
rect 2608 7546 2636 9930
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2700 7449 2728 12582
rect 2792 10674 2820 15438
rect 2872 15360 2924 15366
rect 2872 15302 2924 15308
rect 2884 13870 2912 15302
rect 2976 15094 3004 16374
rect 2964 15088 3016 15094
rect 2964 15030 3016 15036
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2884 12073 2912 12786
rect 2976 12782 3004 14894
rect 3068 14074 3096 16458
rect 3160 16250 3188 17614
rect 3148 16244 3200 16250
rect 3148 16186 3200 16192
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3160 15502 3188 16050
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3148 14816 3200 14822
rect 3148 14758 3200 14764
rect 3160 14550 3188 14758
rect 3148 14544 3200 14550
rect 3148 14486 3200 14492
rect 3148 14408 3200 14414
rect 3148 14350 3200 14356
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3160 13546 3188 14350
rect 3252 13920 3280 17734
rect 3332 17672 3384 17678
rect 3332 17614 3384 17620
rect 3344 16794 3372 17614
rect 3436 17066 3464 17734
rect 3514 17711 3570 17720
rect 3528 17678 3556 17711
rect 3516 17672 3568 17678
rect 3516 17614 3568 17620
rect 3608 17604 3660 17610
rect 3608 17546 3660 17552
rect 3620 17338 3648 17546
rect 3608 17332 3660 17338
rect 3608 17274 3660 17280
rect 3424 17060 3476 17066
rect 3424 17002 3476 17008
rect 3422 16892 3730 16901
rect 3422 16890 3428 16892
rect 3484 16890 3508 16892
rect 3564 16890 3588 16892
rect 3644 16890 3668 16892
rect 3724 16890 3730 16892
rect 3484 16838 3486 16890
rect 3666 16838 3668 16890
rect 3422 16836 3428 16838
rect 3484 16836 3508 16838
rect 3564 16836 3588 16838
rect 3644 16836 3668 16838
rect 3724 16836 3730 16838
rect 3422 16827 3730 16836
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3804 16590 3832 18040
rect 3896 17338 3924 18226
rect 3988 17542 4016 18294
rect 3976 17536 4028 17542
rect 3976 17478 4028 17484
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3988 16674 4016 17478
rect 3896 16646 4016 16674
rect 3792 16584 3844 16590
rect 3422 16552 3478 16561
rect 3332 16516 3384 16522
rect 3792 16526 3844 16532
rect 3422 16487 3478 16496
rect 3332 16458 3384 16464
rect 3344 14929 3372 16458
rect 3436 16182 3464 16487
rect 3804 16425 3832 16526
rect 3790 16416 3846 16425
rect 3896 16402 3924 16646
rect 3976 16584 4028 16590
rect 3974 16552 3976 16561
rect 4028 16552 4030 16561
rect 3974 16487 4030 16496
rect 3896 16374 4016 16402
rect 3790 16351 3846 16360
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3792 15904 3844 15910
rect 3884 15904 3936 15910
rect 3792 15846 3844 15852
rect 3882 15872 3884 15881
rect 3936 15872 3938 15881
rect 3422 15804 3730 15813
rect 3422 15802 3428 15804
rect 3484 15802 3508 15804
rect 3564 15802 3588 15804
rect 3644 15802 3668 15804
rect 3724 15802 3730 15804
rect 3484 15750 3486 15802
rect 3666 15750 3668 15802
rect 3422 15748 3428 15750
rect 3484 15748 3508 15750
rect 3564 15748 3588 15750
rect 3644 15748 3668 15750
rect 3724 15748 3730 15750
rect 3422 15739 3730 15748
rect 3804 15722 3832 15846
rect 3882 15807 3938 15816
rect 3804 15694 3924 15722
rect 3896 15366 3924 15694
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3884 15360 3936 15366
rect 3884 15302 3936 15308
rect 3330 14920 3386 14929
rect 3330 14855 3386 14864
rect 3422 14716 3730 14725
rect 3422 14714 3428 14716
rect 3484 14714 3508 14716
rect 3564 14714 3588 14716
rect 3644 14714 3668 14716
rect 3724 14714 3730 14716
rect 3484 14662 3486 14714
rect 3666 14662 3668 14714
rect 3422 14660 3428 14662
rect 3484 14660 3508 14662
rect 3564 14660 3588 14662
rect 3644 14660 3668 14662
rect 3724 14660 3730 14662
rect 3422 14651 3730 14660
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3332 13932 3384 13938
rect 3252 13892 3332 13920
rect 3332 13874 3384 13880
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3528 13716 3556 13874
rect 3712 13734 3740 14418
rect 3068 13518 3188 13546
rect 3344 13688 3556 13716
rect 3700 13728 3752 13734
rect 3344 13530 3372 13688
rect 3700 13670 3752 13676
rect 3422 13628 3730 13637
rect 3422 13626 3428 13628
rect 3484 13626 3508 13628
rect 3564 13626 3588 13628
rect 3644 13626 3668 13628
rect 3724 13626 3730 13628
rect 3484 13574 3486 13626
rect 3666 13574 3668 13626
rect 3422 13572 3428 13574
rect 3484 13572 3508 13574
rect 3564 13572 3588 13574
rect 3644 13572 3668 13574
rect 3724 13572 3730 13574
rect 3422 13563 3730 13572
rect 3332 13524 3384 13530
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2964 12096 3016 12102
rect 2870 12064 2926 12073
rect 2964 12038 3016 12044
rect 2870 11999 2926 12008
rect 2872 11824 2924 11830
rect 2872 11766 2924 11772
rect 2884 11054 2912 11766
rect 2976 11150 3004 12038
rect 2964 11144 3016 11150
rect 2964 11086 3016 11092
rect 2884 11026 3004 11054
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2780 10668 2832 10674
rect 2780 10610 2832 10616
rect 2884 10062 2912 10678
rect 2976 10130 3004 11026
rect 3068 10198 3096 13518
rect 3332 13466 3384 13472
rect 3700 13456 3752 13462
rect 3700 13398 3752 13404
rect 3148 13252 3200 13258
rect 3148 13194 3200 13200
rect 3160 11558 3188 13194
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3238 13016 3294 13025
rect 3238 12951 3294 12960
rect 3252 12850 3280 12951
rect 3620 12850 3648 13126
rect 3712 12850 3740 13398
rect 3804 12918 3832 15302
rect 3884 15088 3936 15094
rect 3884 15030 3936 15036
rect 3896 13841 3924 15030
rect 3988 14940 4016 16374
rect 4080 15094 4108 18414
rect 4172 17270 4200 19751
rect 4252 19722 4304 19728
rect 4264 19378 4292 19722
rect 4344 19508 4396 19514
rect 4344 19450 4396 19456
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4264 18290 4292 19314
rect 4356 18970 4384 19450
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4448 18850 4476 19910
rect 4356 18822 4476 18850
rect 4356 18426 4384 18822
rect 4436 18760 4488 18766
rect 4436 18702 4488 18708
rect 4344 18420 4396 18426
rect 4344 18362 4396 18368
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4250 18184 4306 18193
rect 4448 18170 4476 18702
rect 4306 18142 4476 18170
rect 4250 18119 4306 18128
rect 4250 17912 4306 17921
rect 4250 17847 4306 17856
rect 4160 17264 4212 17270
rect 4160 17206 4212 17212
rect 4264 17202 4292 17847
rect 4448 17678 4476 18142
rect 4436 17672 4488 17678
rect 4436 17614 4488 17620
rect 4540 17270 4568 20488
rect 4620 20470 4672 20476
rect 4724 20466 4752 20590
rect 4712 20460 4764 20466
rect 4712 20402 4764 20408
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4632 19446 4660 19654
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 4632 18358 4660 19382
rect 4712 19372 4764 19378
rect 4712 19314 4764 19320
rect 4620 18352 4672 18358
rect 4620 18294 4672 18300
rect 4528 17264 4580 17270
rect 4528 17206 4580 17212
rect 4252 17196 4304 17202
rect 4252 17138 4304 17144
rect 4158 16824 4214 16833
rect 4158 16759 4214 16768
rect 4068 15088 4120 15094
rect 4068 15030 4120 15036
rect 3988 14912 4108 14940
rect 4080 14482 4108 14912
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4066 14104 4122 14113
rect 4066 14039 4122 14048
rect 4080 14006 4108 14039
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4172 13938 4200 16759
rect 4264 15094 4292 17138
rect 4528 17128 4580 17134
rect 4342 17096 4398 17105
rect 4528 17070 4580 17076
rect 4342 17031 4398 17040
rect 4356 16289 4384 17031
rect 4342 16280 4398 16289
rect 4342 16215 4398 16224
rect 4344 16040 4396 16046
rect 4344 15982 4396 15988
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3882 13832 3938 13841
rect 3882 13767 3938 13776
rect 4068 13796 4120 13802
rect 4068 13738 4120 13744
rect 3976 13728 4028 13734
rect 3896 13688 3976 13716
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3608 12844 3660 12850
rect 3608 12786 3660 12792
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3252 11762 3280 12786
rect 3896 12696 3924 13688
rect 3976 13670 4028 13676
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 3988 13433 4016 13466
rect 3974 13424 4030 13433
rect 3974 13359 4030 13368
rect 3974 13288 4030 13297
rect 4080 13274 4108 13738
rect 4030 13246 4108 13274
rect 3974 13223 4030 13232
rect 4066 12880 4122 12889
rect 4122 12838 4200 12866
rect 4066 12815 4122 12824
rect 4068 12776 4120 12782
rect 4068 12718 4120 12724
rect 3344 12668 3924 12696
rect 3344 11778 3372 12668
rect 3882 12608 3938 12617
rect 3938 12566 4016 12594
rect 3422 12540 3730 12549
rect 3882 12543 3938 12552
rect 3422 12538 3428 12540
rect 3484 12538 3508 12540
rect 3564 12538 3588 12540
rect 3644 12538 3668 12540
rect 3724 12538 3730 12540
rect 3484 12486 3486 12538
rect 3666 12486 3668 12538
rect 3422 12484 3428 12486
rect 3484 12484 3508 12486
rect 3564 12484 3588 12486
rect 3644 12484 3668 12486
rect 3724 12484 3730 12486
rect 3422 12475 3730 12484
rect 3790 12438 3846 12447
rect 3790 12373 3846 12382
rect 3608 12232 3660 12238
rect 3608 12174 3660 12180
rect 3240 11756 3292 11762
rect 3344 11750 3556 11778
rect 3620 11762 3648 12174
rect 3240 11698 3292 11704
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3148 11552 3200 11558
rect 3148 11494 3200 11500
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 3252 11354 3280 11494
rect 3240 11348 3292 11354
rect 3240 11290 3292 11296
rect 3344 11150 3372 11630
rect 3528 11626 3556 11750
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3422 11452 3730 11461
rect 3422 11450 3428 11452
rect 3484 11450 3508 11452
rect 3564 11450 3588 11452
rect 3644 11450 3668 11452
rect 3724 11450 3730 11452
rect 3484 11398 3486 11450
rect 3666 11398 3668 11450
rect 3422 11396 3428 11398
rect 3484 11396 3508 11398
rect 3564 11396 3588 11398
rect 3644 11396 3668 11398
rect 3724 11396 3730 11398
rect 3422 11387 3730 11396
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 3332 11144 3384 11150
rect 3332 11086 3384 11092
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 2964 10124 3016 10130
rect 2964 10066 3016 10072
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2780 9716 2832 9722
rect 2780 9658 2832 9664
rect 2792 9625 2820 9658
rect 2778 9616 2834 9625
rect 2778 9551 2834 9560
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 7596 2820 9454
rect 2884 8430 2912 9862
rect 2976 8634 3004 9862
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2962 8392 3018 8401
rect 2962 8327 3018 8336
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2884 7750 2912 8230
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2792 7568 2912 7596
rect 2686 7440 2742 7449
rect 2686 7375 2742 7384
rect 2884 7342 2912 7568
rect 2872 7336 2924 7342
rect 2686 7304 2742 7313
rect 2976 7313 3004 8327
rect 3068 7546 3096 9386
rect 3160 8974 3188 10610
rect 3252 9722 3280 10950
rect 3344 10266 3372 11086
rect 3528 10606 3556 11222
rect 3608 11076 3660 11082
rect 3608 11018 3660 11024
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3620 10470 3648 11018
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3422 10364 3730 10373
rect 3422 10362 3428 10364
rect 3484 10362 3508 10364
rect 3564 10362 3588 10364
rect 3644 10362 3668 10364
rect 3724 10362 3730 10364
rect 3484 10310 3486 10362
rect 3666 10310 3668 10362
rect 3422 10308 3428 10310
rect 3484 10308 3508 10310
rect 3564 10308 3588 10310
rect 3644 10308 3668 10310
rect 3724 10308 3730 10310
rect 3422 10299 3730 10308
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3424 10260 3476 10266
rect 3424 10202 3476 10208
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3344 9625 3372 9658
rect 3330 9616 3386 9625
rect 3330 9551 3386 9560
rect 3436 9466 3464 10202
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3528 9586 3556 10066
rect 3516 9580 3568 9586
rect 3516 9522 3568 9528
rect 3344 9438 3464 9466
rect 3238 9344 3294 9353
rect 3238 9279 3294 9288
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3160 8634 3188 8774
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3146 8256 3202 8265
rect 3146 8191 3202 8200
rect 3160 7546 3188 8191
rect 3252 7970 3280 9279
rect 3344 9160 3372 9438
rect 3422 9276 3730 9285
rect 3422 9274 3428 9276
rect 3484 9274 3508 9276
rect 3564 9274 3588 9276
rect 3644 9274 3668 9276
rect 3724 9274 3730 9276
rect 3484 9222 3486 9274
rect 3666 9222 3668 9274
rect 3422 9220 3428 9222
rect 3484 9220 3508 9222
rect 3564 9220 3588 9222
rect 3644 9220 3668 9222
rect 3724 9220 3730 9222
rect 3422 9211 3730 9220
rect 3344 9132 3464 9160
rect 3436 8537 3464 9132
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3422 8528 3478 8537
rect 3422 8463 3424 8472
rect 3476 8463 3478 8472
rect 3424 8434 3476 8440
rect 3528 8276 3556 8978
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3712 8498 3740 8774
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3344 8248 3556 8276
rect 3344 8072 3372 8248
rect 3422 8188 3730 8197
rect 3422 8186 3428 8188
rect 3484 8186 3508 8188
rect 3564 8186 3588 8188
rect 3644 8186 3668 8188
rect 3724 8186 3730 8188
rect 3484 8134 3486 8186
rect 3666 8134 3668 8186
rect 3422 8132 3428 8134
rect 3484 8132 3508 8134
rect 3564 8132 3588 8134
rect 3644 8132 3668 8134
rect 3724 8132 3730 8134
rect 3422 8123 3730 8132
rect 3344 8044 3464 8072
rect 3252 7942 3372 7970
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3148 7540 3200 7546
rect 3148 7482 3200 7488
rect 2872 7278 2924 7284
rect 2962 7304 3018 7313
rect 2686 7239 2742 7248
rect 2780 7268 2832 7274
rect 2596 6792 2648 6798
rect 2516 6752 2596 6780
rect 2596 6734 2648 6740
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2410 5400 2466 5409
rect 2410 5335 2466 5344
rect 2424 5234 2452 5335
rect 2188 5188 2268 5216
rect 2320 5228 2372 5234
rect 2136 5170 2188 5176
rect 2320 5170 2372 5176
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2228 5092 2280 5098
rect 2228 5034 2280 5040
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 1952 4548 2004 4554
rect 1952 4490 2004 4496
rect 2240 4010 2268 5034
rect 2332 4078 2360 5170
rect 2424 4154 2452 5170
rect 2516 4622 2544 5510
rect 2608 5234 2636 6054
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2424 4146 2544 4154
rect 2424 4140 2556 4146
rect 2424 4126 2504 4140
rect 2504 4082 2556 4088
rect 2320 4072 2372 4078
rect 2320 4014 2372 4020
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1768 3528 1820 3534
rect 1768 3470 1820 3476
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1688 2650 1716 3334
rect 1780 3058 1808 3470
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1676 2644 1728 2650
rect 1676 2586 1728 2592
rect 1780 2514 1808 2994
rect 1858 2680 1914 2689
rect 1858 2615 1914 2624
rect 1768 2508 1820 2514
rect 1768 2450 1820 2456
rect 1400 2100 1452 2106
rect 1400 2042 1452 2048
rect 1308 2032 1360 2038
rect 1308 1974 1360 1980
rect 1872 1562 1900 2615
rect 1860 1556 1912 1562
rect 1860 1498 1912 1504
rect 1032 1420 1084 1426
rect 1032 1362 1084 1368
rect 1768 1284 1820 1290
rect 1768 1226 1820 1232
rect 386 776 442 785
rect 386 711 442 720
rect 1780 678 1808 1226
rect 1768 672 1820 678
rect 1768 614 1820 620
rect 2332 474 2360 4014
rect 2608 3738 2636 5034
rect 2700 4826 2728 7239
rect 2780 7210 2832 7216
rect 2792 5914 2820 7210
rect 2884 6254 2912 7278
rect 2962 7239 3018 7248
rect 2962 7168 3018 7177
rect 2962 7103 3018 7112
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 2870 5944 2926 5953
rect 2780 5908 2832 5914
rect 2870 5879 2926 5888
rect 2780 5850 2832 5856
rect 2884 5273 2912 5879
rect 2870 5264 2926 5273
rect 2870 5199 2926 5208
rect 2780 5160 2832 5166
rect 2884 5148 2912 5199
rect 2832 5120 2912 5148
rect 2780 5102 2832 5108
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2792 4154 2820 4966
rect 2700 4126 2820 4154
rect 2700 4078 2728 4126
rect 2884 4078 2912 5120
rect 2976 4154 3004 7103
rect 3252 7041 3280 7822
rect 3344 7750 3372 7942
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3436 7290 3464 8044
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3528 7818 3556 7958
rect 3698 7848 3754 7857
rect 3516 7812 3568 7818
rect 3698 7783 3754 7792
rect 3516 7754 3568 7760
rect 3344 7262 3464 7290
rect 3238 7032 3294 7041
rect 3238 6967 3294 6976
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 3068 6662 3096 6802
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3240 6180 3292 6186
rect 3240 6122 3292 6128
rect 3068 5817 3096 6122
rect 3146 6080 3202 6089
rect 3146 6015 3202 6024
rect 3054 5808 3110 5817
rect 3054 5743 3110 5752
rect 3054 5536 3110 5545
rect 3054 5471 3110 5480
rect 3068 4758 3096 5471
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2976 4126 3096 4154
rect 2688 4072 2740 4078
rect 2688 4014 2740 4020
rect 2872 4072 2924 4078
rect 2872 4014 2924 4020
rect 2780 4004 2832 4010
rect 2780 3946 2832 3952
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2596 3732 2648 3738
rect 2596 3674 2648 3680
rect 2594 3632 2650 3641
rect 2594 3567 2650 3576
rect 2410 3496 2466 3505
rect 2410 3431 2466 3440
rect 2424 2038 2452 3431
rect 2502 2680 2558 2689
rect 2502 2615 2558 2624
rect 2412 2032 2464 2038
rect 2412 1974 2464 1980
rect 2516 1562 2544 2615
rect 2608 2038 2636 3567
rect 2792 3126 2820 3946
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2976 2650 3004 3946
rect 3068 3194 3096 4126
rect 3160 3738 3188 6015
rect 3252 5914 3280 6122
rect 3344 6118 3372 7262
rect 3712 7206 3740 7783
rect 3804 7721 3832 12373
rect 3988 12322 4016 12566
rect 3896 12294 4016 12322
rect 3896 11898 3924 12294
rect 3976 12232 4028 12238
rect 3976 12174 4028 12180
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3896 10130 3924 11562
rect 3988 11218 4016 12174
rect 4080 11801 4108 12718
rect 4172 12442 4200 12838
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4066 11792 4122 11801
rect 4066 11727 4122 11736
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 4080 11354 4108 11562
rect 4172 11529 4200 11630
rect 4158 11520 4214 11529
rect 4158 11455 4214 11464
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 4066 11248 4122 11257
rect 3976 11212 4028 11218
rect 4122 11206 4200 11234
rect 4066 11183 4122 11192
rect 3976 11154 4028 11160
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 3988 10305 4016 10639
rect 3974 10296 4030 10305
rect 4172 10266 4200 11206
rect 4264 10742 4292 14894
rect 4356 14278 4384 15982
rect 4540 15910 4568 17070
rect 4620 16108 4672 16114
rect 4724 16096 4752 19314
rect 4816 19242 4844 22358
rect 5000 22216 5028 22578
rect 5080 22432 5132 22438
rect 5080 22374 5132 22380
rect 4908 22188 5028 22216
rect 4908 21690 4936 22188
rect 5092 22094 5120 22374
rect 5000 22066 5120 22094
rect 5000 22030 5028 22066
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 4896 21684 4948 21690
rect 4896 21626 4948 21632
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4908 19718 4936 20878
rect 5000 20874 5028 21830
rect 5080 21616 5132 21622
rect 5080 21558 5132 21564
rect 4988 20868 5040 20874
rect 4988 20810 5040 20816
rect 5000 20641 5028 20810
rect 4986 20632 5042 20641
rect 4986 20567 5042 20576
rect 5092 20312 5120 21558
rect 5184 20942 5212 22646
rect 5172 20936 5224 20942
rect 5172 20878 5224 20884
rect 5092 20284 5212 20312
rect 5078 20224 5134 20233
rect 5078 20159 5134 20168
rect 4986 19952 5042 19961
rect 4986 19887 5042 19896
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4896 19236 4948 19242
rect 4896 19178 4948 19184
rect 4908 18986 4936 19178
rect 4816 18958 4936 18986
rect 4816 16164 4844 18958
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4908 18290 4936 18770
rect 4896 18284 4948 18290
rect 4896 18226 4948 18232
rect 4908 17678 4936 18226
rect 4896 17672 4948 17678
rect 4896 17614 4948 17620
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4908 17134 4936 17206
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4896 16516 4948 16522
rect 5000 16504 5028 19887
rect 5092 18426 5120 20159
rect 5184 19922 5212 20284
rect 5276 20097 5304 23190
rect 5356 23180 5408 23186
rect 5356 23122 5408 23128
rect 5262 20088 5318 20097
rect 5262 20023 5318 20032
rect 5172 19916 5224 19922
rect 5172 19858 5224 19864
rect 5262 19680 5318 19689
rect 5262 19615 5318 19624
rect 5276 19446 5304 19615
rect 5264 19440 5316 19446
rect 5264 19382 5316 19388
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5172 18964 5224 18970
rect 5172 18906 5224 18912
rect 5184 18698 5212 18906
rect 5172 18692 5224 18698
rect 5172 18634 5224 18640
rect 5080 18420 5132 18426
rect 5080 18362 5132 18368
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 5092 17610 5120 18226
rect 5080 17604 5132 17610
rect 5080 17546 5132 17552
rect 5172 17536 5224 17542
rect 5078 17504 5134 17513
rect 5172 17478 5224 17484
rect 5078 17439 5134 17448
rect 5092 16590 5120 17439
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 4948 16476 5028 16504
rect 4896 16458 4948 16464
rect 4908 16425 4936 16458
rect 4894 16416 4950 16425
rect 4894 16351 4950 16360
rect 4816 16136 4936 16164
rect 4672 16068 4844 16096
rect 4620 16050 4672 16056
rect 4712 15972 4764 15978
rect 4712 15914 4764 15920
rect 4528 15904 4580 15910
rect 4528 15846 4580 15852
rect 4540 15638 4568 15846
rect 4528 15632 4580 15638
rect 4528 15574 4580 15580
rect 4540 15026 4568 15574
rect 4528 15020 4580 15026
rect 4528 14962 4580 14968
rect 4724 14958 4752 15914
rect 4712 14952 4764 14958
rect 4618 14920 4674 14929
rect 4712 14894 4764 14900
rect 4618 14855 4674 14864
rect 4632 14362 4660 14855
rect 4710 14512 4766 14521
rect 4816 14482 4844 16068
rect 4710 14447 4712 14456
rect 4764 14447 4766 14456
rect 4804 14476 4856 14482
rect 4712 14418 4764 14424
rect 4804 14418 4856 14424
rect 4802 14376 4858 14385
rect 4632 14334 4802 14362
rect 4344 14272 4396 14278
rect 4344 14214 4396 14220
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4434 13968 4490 13977
rect 4434 13903 4436 13912
rect 4488 13903 4490 13912
rect 4436 13874 4488 13880
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 13258 4476 13670
rect 4540 13326 4568 14214
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4436 13252 4488 13258
rect 4436 13194 4488 13200
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4356 12986 4384 13126
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4632 12696 4660 14334
rect 4802 14311 4858 14320
rect 4712 13796 4764 13802
rect 4712 13738 4764 13744
rect 4356 12668 4660 12696
rect 4356 10742 4384 12668
rect 4448 12566 4660 12594
rect 4448 12306 4476 12566
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4436 12300 4488 12306
rect 4436 12242 4488 12248
rect 4436 12096 4488 12102
rect 4434 12064 4436 12073
rect 4488 12064 4490 12073
rect 4434 11999 4490 12008
rect 4540 11762 4568 12378
rect 4528 11756 4580 11762
rect 4528 11698 4580 11704
rect 4632 11540 4660 12566
rect 4724 11608 4752 13738
rect 4804 13728 4856 13734
rect 4804 13670 4856 13676
rect 4816 13326 4844 13670
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4816 12782 4844 13262
rect 4804 12776 4856 12782
rect 4804 12718 4856 12724
rect 4816 11676 4844 12718
rect 4908 12345 4936 16136
rect 5080 15020 5132 15026
rect 5080 14962 5132 14968
rect 5092 13938 5120 14962
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 4988 13320 5040 13326
rect 4986 13288 4988 13297
rect 5040 13288 5042 13297
rect 4986 13223 5042 13232
rect 5080 13184 5132 13190
rect 5080 13126 5132 13132
rect 4986 13016 5042 13025
rect 4986 12951 5042 12960
rect 5000 12918 5028 12951
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4986 12608 5042 12617
rect 4986 12543 5042 12552
rect 4894 12336 4950 12345
rect 4894 12271 4950 12280
rect 4896 11892 4948 11898
rect 5000 11880 5028 12543
rect 4948 11852 5028 11880
rect 4896 11834 4948 11840
rect 4816 11648 4936 11676
rect 4724 11580 4844 11608
rect 4526 11520 4582 11529
rect 4632 11512 4752 11540
rect 4526 11455 4582 11464
rect 4540 11354 4568 11455
rect 4724 11354 4752 11512
rect 4528 11348 4580 11354
rect 4712 11348 4764 11354
rect 4580 11308 4660 11336
rect 4528 11290 4580 11296
rect 4526 11248 4582 11257
rect 4436 11212 4488 11218
rect 4526 11183 4582 11192
rect 4436 11154 4488 11160
rect 4448 10810 4476 11154
rect 4540 10985 4568 11183
rect 4632 11014 4660 11308
rect 4712 11290 4764 11296
rect 4712 11212 4764 11218
rect 4816 11200 4844 11580
rect 4908 11529 4936 11648
rect 4894 11520 4950 11529
rect 4894 11455 4950 11464
rect 4894 11384 4950 11393
rect 4894 11319 4950 11328
rect 4764 11172 4844 11200
rect 4712 11154 4764 11160
rect 4620 11008 4672 11014
rect 4526 10976 4582 10985
rect 4620 10950 4672 10956
rect 4526 10911 4582 10920
rect 4436 10804 4488 10810
rect 4436 10746 4488 10752
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4724 10266 4752 11154
rect 4802 11112 4858 11121
rect 4802 11047 4858 11056
rect 4816 10606 4844 11047
rect 4908 10985 4936 11319
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 4894 10976 4950 10985
rect 4894 10911 4950 10920
rect 5000 10810 5028 11086
rect 4988 10804 5040 10810
rect 4988 10746 5040 10752
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 5092 10690 5120 13126
rect 5184 12442 5212 17478
rect 5276 16114 5304 19110
rect 5368 17542 5396 23122
rect 5460 23066 5488 24142
rect 5644 23186 5672 25230
rect 5736 24410 5764 25230
rect 5828 24410 5856 25434
rect 5894 25052 6202 25061
rect 5894 25050 5900 25052
rect 5956 25050 5980 25052
rect 6036 25050 6060 25052
rect 6116 25050 6140 25052
rect 6196 25050 6202 25052
rect 5956 24998 5958 25050
rect 6138 24998 6140 25050
rect 5894 24996 5900 24998
rect 5956 24996 5980 24998
rect 6036 24996 6060 24998
rect 6116 24996 6140 24998
rect 6196 24996 6202 24998
rect 5894 24987 6202 24996
rect 6184 24948 6236 24954
rect 6184 24890 6236 24896
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5724 24404 5776 24410
rect 5724 24346 5776 24352
rect 5816 24404 5868 24410
rect 5816 24346 5868 24352
rect 5920 24290 5948 24754
rect 6000 24744 6052 24750
rect 6000 24686 6052 24692
rect 6012 24410 6040 24686
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 5736 24262 5948 24290
rect 5632 23180 5684 23186
rect 5632 23122 5684 23128
rect 5460 23038 5672 23066
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5460 21554 5488 22918
rect 5540 22092 5592 22098
rect 5540 22034 5592 22040
rect 5552 21978 5580 22034
rect 5552 21950 5598 21978
rect 5570 21876 5598 21950
rect 5644 21894 5672 23038
rect 5552 21848 5598 21876
rect 5632 21888 5684 21894
rect 5552 21690 5580 21848
rect 5632 21830 5684 21836
rect 5540 21684 5592 21690
rect 5736 21672 5764 24262
rect 6196 24206 6224 24890
rect 6184 24200 6236 24206
rect 5540 21626 5592 21632
rect 5644 21644 5764 21672
rect 5828 24160 6184 24188
rect 5448 21548 5500 21554
rect 5448 21490 5500 21496
rect 5460 20505 5488 21490
rect 5644 21298 5672 21644
rect 5828 21570 5856 24160
rect 6184 24142 6236 24148
rect 5894 23964 6202 23973
rect 5894 23962 5900 23964
rect 5956 23962 5980 23964
rect 6036 23962 6060 23964
rect 6116 23962 6140 23964
rect 6196 23962 6202 23964
rect 5956 23910 5958 23962
rect 6138 23910 6140 23962
rect 5894 23908 5900 23910
rect 5956 23908 5980 23910
rect 6036 23908 6060 23910
rect 6116 23908 6140 23910
rect 6196 23908 6202 23910
rect 5894 23899 6202 23908
rect 6288 23730 6316 25978
rect 6380 24954 6408 27406
rect 6368 24948 6420 24954
rect 6368 24890 6420 24896
rect 6472 24834 6500 28494
rect 6564 28218 6592 28494
rect 6552 28212 6604 28218
rect 6552 28154 6604 28160
rect 6656 28098 6684 28648
rect 6748 28642 6776 28750
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 6920 28756 6972 28762
rect 6920 28698 6972 28704
rect 6748 28614 6868 28642
rect 6380 24806 6500 24834
rect 6564 28070 6684 28098
rect 6276 23724 6328 23730
rect 6276 23666 6328 23672
rect 6380 23526 6408 24806
rect 6458 24576 6514 24585
rect 6458 24511 6514 24520
rect 6472 23662 6500 24511
rect 6460 23656 6512 23662
rect 6460 23598 6512 23604
rect 6368 23520 6420 23526
rect 5998 23488 6054 23497
rect 6368 23462 6420 23468
rect 5998 23423 6054 23432
rect 6012 23254 6040 23423
rect 6000 23248 6052 23254
rect 6000 23190 6052 23196
rect 6274 22944 6330 22953
rect 5894 22876 6202 22885
rect 6274 22879 6330 22888
rect 5894 22874 5900 22876
rect 5956 22874 5980 22876
rect 6036 22874 6060 22876
rect 6116 22874 6140 22876
rect 6196 22874 6202 22876
rect 5956 22822 5958 22874
rect 6138 22822 6140 22874
rect 5894 22820 5900 22822
rect 5956 22820 5980 22822
rect 6036 22820 6060 22822
rect 6116 22820 6140 22822
rect 6196 22820 6202 22822
rect 5894 22811 6202 22820
rect 5908 22636 5960 22642
rect 5908 22578 5960 22584
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 5920 22098 5948 22578
rect 6012 22166 6040 22578
rect 6000 22160 6052 22166
rect 6000 22102 6052 22108
rect 5908 22092 5960 22098
rect 5908 22034 5960 22040
rect 6184 22024 6236 22030
rect 6184 21966 6236 21972
rect 6196 21894 6224 21966
rect 6184 21888 6236 21894
rect 6184 21830 6236 21836
rect 5894 21788 6202 21797
rect 5894 21786 5900 21788
rect 5956 21786 5980 21788
rect 6036 21786 6060 21788
rect 6116 21786 6140 21788
rect 6196 21786 6202 21788
rect 5956 21734 5958 21786
rect 6138 21734 6140 21786
rect 5894 21732 5900 21734
rect 5956 21732 5980 21734
rect 6036 21732 6060 21734
rect 6116 21732 6140 21734
rect 6196 21732 6202 21734
rect 5894 21723 6202 21732
rect 5552 21270 5672 21298
rect 5736 21542 5856 21570
rect 5446 20496 5502 20505
rect 5446 20431 5502 20440
rect 5552 19553 5580 21270
rect 5736 21128 5764 21542
rect 5906 21312 5962 21321
rect 5906 21247 5962 21256
rect 5644 21100 5764 21128
rect 5644 19718 5672 21100
rect 5920 20942 5948 21247
rect 5816 20936 5868 20942
rect 5816 20878 5868 20884
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5722 20768 5778 20777
rect 5722 20703 5778 20712
rect 5736 19854 5764 20703
rect 5828 20330 5856 20878
rect 5894 20700 6202 20709
rect 5894 20698 5900 20700
rect 5956 20698 5980 20700
rect 6036 20698 6060 20700
rect 6116 20698 6140 20700
rect 6196 20698 6202 20700
rect 5956 20646 5958 20698
rect 6138 20646 6140 20698
rect 5894 20644 5900 20646
rect 5956 20644 5980 20646
rect 6036 20644 6060 20646
rect 6116 20644 6140 20646
rect 6196 20644 6202 20646
rect 5894 20635 6202 20644
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5724 19848 5776 19854
rect 5776 19808 5856 19836
rect 5724 19790 5776 19796
rect 5632 19712 5684 19718
rect 5632 19654 5684 19660
rect 5538 19544 5594 19553
rect 5538 19479 5594 19488
rect 5644 19378 5672 19654
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5460 17785 5488 18566
rect 5446 17776 5502 17785
rect 5446 17711 5502 17720
rect 5724 17604 5776 17610
rect 5724 17546 5776 17552
rect 5356 17536 5408 17542
rect 5356 17478 5408 17484
rect 5448 17536 5500 17542
rect 5448 17478 5500 17484
rect 5356 16720 5408 16726
rect 5356 16662 5408 16668
rect 5368 16522 5396 16662
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 5460 16153 5488 17478
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5446 16144 5502 16153
rect 5264 16108 5316 16114
rect 5446 16079 5502 16088
rect 5264 16050 5316 16056
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5172 12300 5224 12306
rect 5276 12288 5304 16050
rect 5446 15600 5502 15609
rect 5446 15535 5502 15544
rect 5460 15502 5488 15535
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5448 15360 5500 15366
rect 5552 15337 5580 16526
rect 5448 15302 5500 15308
rect 5538 15328 5594 15337
rect 5460 14618 5488 15302
rect 5538 15263 5594 15272
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5644 13818 5672 17138
rect 5460 13790 5672 13818
rect 5356 13320 5408 13326
rect 5356 13262 5408 13268
rect 5368 12434 5396 13262
rect 5368 12406 5421 12434
rect 5393 12356 5421 12406
rect 5224 12260 5304 12288
rect 5368 12328 5421 12356
rect 5172 12242 5224 12248
rect 5184 11218 5212 12242
rect 5368 12152 5396 12328
rect 5276 12124 5396 12152
rect 5172 11212 5224 11218
rect 5172 11154 5224 11160
rect 5170 11112 5226 11121
rect 5170 11047 5226 11056
rect 5184 10810 5212 11047
rect 5276 10810 5304 12124
rect 5354 12064 5410 12073
rect 5354 11999 5410 12008
rect 5368 11898 5396 11999
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5264 10804 5316 10810
rect 5264 10746 5316 10752
rect 4804 10600 4856 10606
rect 4804 10542 4856 10548
rect 3974 10231 4030 10240
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4804 10260 4856 10266
rect 4804 10202 4856 10208
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 4436 10056 4488 10062
rect 4620 10056 4672 10062
rect 4436 9998 4488 10004
rect 4526 10024 4582 10033
rect 4068 9920 4120 9926
rect 3988 9880 4068 9908
rect 3988 9194 4016 9880
rect 4068 9862 4120 9868
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4066 9752 4122 9761
rect 4122 9710 4292 9738
rect 4066 9687 4122 9696
rect 4160 9648 4212 9654
rect 4158 9616 4160 9625
rect 4212 9616 4214 9625
rect 4158 9551 4214 9560
rect 4160 9512 4212 9518
rect 4160 9454 4212 9460
rect 3896 9166 4016 9194
rect 4066 9208 4122 9217
rect 3896 8022 3924 9166
rect 4066 9143 4122 9152
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 3884 8016 3936 8022
rect 3884 7958 3936 7964
rect 3790 7712 3846 7721
rect 3790 7647 3846 7656
rect 3988 7562 4016 9007
rect 4080 8430 4108 9143
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 4080 8129 4108 8366
rect 4066 8120 4122 8129
rect 4172 8090 4200 9454
rect 4264 9178 4292 9710
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4356 8974 4384 9862
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4252 8900 4304 8906
rect 4252 8842 4304 8848
rect 4066 8055 4122 8064
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4066 7984 4122 7993
rect 4264 7954 4292 8842
rect 4448 8537 4476 9998
rect 4620 9998 4672 10004
rect 4526 9959 4582 9968
rect 4434 8528 4490 8537
rect 4434 8463 4436 8472
rect 4488 8463 4490 8472
rect 4436 8434 4488 8440
rect 4540 8378 4568 9959
rect 4632 9926 4660 9998
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4710 9888 4766 9897
rect 4710 9823 4766 9832
rect 4724 9518 4752 9823
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4448 8350 4568 8378
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4066 7919 4122 7928
rect 4252 7948 4304 7954
rect 4080 7750 4108 7919
rect 4252 7890 4304 7896
rect 4158 7848 4214 7857
rect 4158 7783 4214 7792
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 3988 7534 4108 7562
rect 3882 7440 3938 7449
rect 3882 7375 3884 7384
rect 3936 7375 3938 7384
rect 3884 7346 3936 7352
rect 3976 7336 4028 7342
rect 3974 7304 3976 7313
rect 4028 7304 4030 7313
rect 3974 7239 4030 7248
rect 3700 7200 3752 7206
rect 3700 7142 3752 7148
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 3422 7100 3730 7109
rect 3422 7098 3428 7100
rect 3484 7098 3508 7100
rect 3564 7098 3588 7100
rect 3644 7098 3668 7100
rect 3724 7098 3730 7100
rect 3484 7046 3486 7098
rect 3666 7046 3668 7098
rect 3422 7044 3428 7046
rect 3484 7044 3508 7046
rect 3564 7044 3588 7046
rect 3644 7044 3668 7046
rect 3724 7044 3730 7046
rect 3422 7035 3730 7044
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6322 3832 6598
rect 3896 6458 3924 7142
rect 3974 6896 4030 6905
rect 3974 6831 4030 6840
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3332 6112 3384 6118
rect 3882 6080 3938 6089
rect 3332 6054 3384 6060
rect 3804 6038 3882 6066
rect 3422 6012 3730 6021
rect 3422 6010 3428 6012
rect 3484 6010 3508 6012
rect 3564 6010 3588 6012
rect 3644 6010 3668 6012
rect 3724 6010 3730 6012
rect 3484 5958 3486 6010
rect 3666 5958 3668 6010
rect 3422 5956 3428 5958
rect 3484 5956 3508 5958
rect 3564 5956 3588 5958
rect 3644 5956 3668 5958
rect 3724 5956 3730 5958
rect 3422 5947 3730 5956
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3436 5386 3464 5510
rect 3252 5358 3464 5386
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3056 3188 3108 3194
rect 3056 3130 3108 3136
rect 3252 3126 3280 5358
rect 3378 5228 3430 5234
rect 3378 5170 3430 5176
rect 3390 5114 3418 5170
rect 3344 5086 3418 5114
rect 3344 4826 3372 5086
rect 3422 4924 3730 4933
rect 3422 4922 3428 4924
rect 3484 4922 3508 4924
rect 3564 4922 3588 4924
rect 3644 4922 3668 4924
rect 3724 4922 3730 4924
rect 3484 4870 3486 4922
rect 3666 4870 3668 4922
rect 3422 4868 3428 4870
rect 3484 4868 3508 4870
rect 3564 4868 3588 4870
rect 3644 4868 3668 4870
rect 3724 4868 3730 4870
rect 3422 4859 3730 4868
rect 3332 4820 3384 4826
rect 3332 4762 3384 4768
rect 3516 4820 3568 4826
rect 3516 4762 3568 4768
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3344 3466 3372 4626
rect 3528 4154 3556 4762
rect 3804 4729 3832 6038
rect 3882 6015 3938 6024
rect 3988 5914 4016 6831
rect 4080 6633 4108 7534
rect 4172 7410 4200 7783
rect 4356 7546 4384 8230
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4158 7168 4214 7177
rect 4158 7103 4214 7112
rect 4066 6624 4122 6633
rect 4066 6559 4122 6568
rect 4066 6488 4122 6497
rect 4066 6423 4122 6432
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 4080 5658 4108 6423
rect 4172 5778 4200 7103
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3988 5630 4108 5658
rect 4158 5672 4214 5681
rect 3896 5370 3924 5578
rect 3988 5370 4016 5630
rect 4158 5607 4214 5616
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 3884 5364 3936 5370
rect 3884 5306 3936 5312
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3988 5098 4016 5306
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3988 4826 4016 5034
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3606 4720 3662 4729
rect 3606 4655 3662 4664
rect 3790 4720 3846 4729
rect 3790 4655 3846 4664
rect 3620 4622 3648 4655
rect 4080 4622 4108 5510
rect 4172 5166 4200 5607
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 3608 4616 3660 4622
rect 4068 4616 4120 4622
rect 3608 4558 3660 4564
rect 3974 4584 4030 4593
rect 4068 4558 4120 4564
rect 3974 4519 4030 4528
rect 3790 4448 3846 4457
rect 3790 4383 3846 4392
rect 3436 4146 3556 4154
rect 3424 4140 3556 4146
rect 3476 4126 3556 4140
rect 3424 4082 3476 4088
rect 3422 3836 3730 3845
rect 3422 3834 3428 3836
rect 3484 3834 3508 3836
rect 3564 3834 3588 3836
rect 3644 3834 3668 3836
rect 3724 3834 3730 3836
rect 3484 3782 3486 3834
rect 3666 3782 3668 3834
rect 3422 3780 3428 3782
rect 3484 3780 3508 3782
rect 3564 3780 3588 3782
rect 3644 3780 3668 3782
rect 3724 3780 3730 3782
rect 3422 3771 3730 3780
rect 3332 3460 3384 3466
rect 3332 3402 3384 3408
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 3068 2854 3096 2994
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3422 2748 3730 2757
rect 3422 2746 3428 2748
rect 3484 2746 3508 2748
rect 3564 2746 3588 2748
rect 3644 2746 3668 2748
rect 3724 2746 3730 2748
rect 3484 2694 3486 2746
rect 3666 2694 3668 2746
rect 3422 2692 3428 2694
rect 3484 2692 3508 2694
rect 3564 2692 3588 2694
rect 3644 2692 3668 2694
rect 3724 2692 3730 2694
rect 3422 2683 3730 2692
rect 3804 2650 3832 4383
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3896 3194 3924 4014
rect 3988 3738 4016 4519
rect 4172 4321 4200 5102
rect 4158 4312 4214 4321
rect 4158 4247 4214 4256
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4080 3618 4108 3975
rect 4158 3904 4214 3913
rect 4158 3839 4214 3848
rect 3988 3590 4108 3618
rect 3988 3466 4016 3590
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 4172 3194 4200 3839
rect 4264 3777 4292 7278
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 6390 4384 6802
rect 4344 6384 4396 6390
rect 4344 6326 4396 6332
rect 4448 5710 4476 8350
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4540 7478 4568 8230
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6458 4568 6734
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4526 6352 4582 6361
rect 4526 6287 4582 6296
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4434 5264 4490 5273
rect 4540 5234 4568 6287
rect 4434 5199 4436 5208
rect 4488 5199 4490 5208
rect 4528 5228 4580 5234
rect 4436 5170 4488 5176
rect 4528 5170 4580 5176
rect 4526 4992 4582 5001
rect 4526 4927 4582 4936
rect 4540 4622 4568 4927
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4250 3768 4306 3777
rect 4356 3738 4384 4490
rect 4448 3738 4476 4490
rect 4250 3703 4306 3712
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4436 3732 4488 3738
rect 4436 3674 4488 3680
rect 4540 3618 4568 4558
rect 4448 3590 4568 3618
rect 3884 3188 3936 3194
rect 4160 3188 4212 3194
rect 3884 3130 3936 3136
rect 4080 3148 4160 3176
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3790 2544 3846 2553
rect 4080 2514 4108 3148
rect 4160 3130 4212 3136
rect 4342 2680 4398 2689
rect 4448 2650 4476 3590
rect 4528 3528 4580 3534
rect 4632 3516 4660 9318
rect 4724 9081 4752 9454
rect 4710 9072 4766 9081
rect 4710 9007 4766 9016
rect 4710 8936 4766 8945
rect 4710 8871 4766 8880
rect 4724 8634 4752 8871
rect 4816 8673 4844 10202
rect 4908 9518 4936 10678
rect 5092 10662 5304 10690
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5092 9926 5120 9998
rect 5080 9920 5132 9926
rect 5080 9862 5132 9868
rect 4896 9512 4948 9518
rect 4896 9454 4948 9460
rect 5078 9480 5134 9489
rect 4988 9444 5040 9450
rect 5078 9415 5134 9424
rect 4988 9386 5040 9392
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4802 8664 4858 8673
rect 4712 8628 4764 8634
rect 4802 8599 4858 8608
rect 4712 8570 4764 8576
rect 4908 8344 4936 9318
rect 5000 8634 5028 9386
rect 5092 8974 5120 9415
rect 5184 9178 5212 10406
rect 5276 9552 5304 10662
rect 5368 9722 5396 11698
rect 5460 11626 5488 13790
rect 5632 13728 5684 13734
rect 5538 13696 5594 13705
rect 5632 13670 5684 13676
rect 5538 13631 5594 13640
rect 5552 12424 5580 13631
rect 5644 12714 5672 13670
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5630 12608 5686 12617
rect 5736 12594 5764 17546
rect 5828 17218 5856 19808
rect 5894 19612 6202 19621
rect 5894 19610 5900 19612
rect 5956 19610 5980 19612
rect 6036 19610 6060 19612
rect 6116 19610 6140 19612
rect 6196 19610 6202 19612
rect 5956 19558 5958 19610
rect 6138 19558 6140 19610
rect 5894 19556 5900 19558
rect 5956 19556 5980 19558
rect 6036 19556 6060 19558
rect 6116 19556 6140 19558
rect 6196 19556 6202 19558
rect 5894 19547 6202 19556
rect 5894 18524 6202 18533
rect 5894 18522 5900 18524
rect 5956 18522 5980 18524
rect 6036 18522 6060 18524
rect 6116 18522 6140 18524
rect 6196 18522 6202 18524
rect 5956 18470 5958 18522
rect 6138 18470 6140 18522
rect 5894 18468 5900 18470
rect 5956 18468 5980 18470
rect 6036 18468 6060 18470
rect 6116 18468 6140 18470
rect 6196 18468 6202 18470
rect 5894 18459 6202 18468
rect 5906 18320 5962 18329
rect 5906 18255 5962 18264
rect 5920 17542 5948 18255
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5894 17436 6202 17445
rect 5894 17434 5900 17436
rect 5956 17434 5980 17436
rect 6036 17434 6060 17436
rect 6116 17434 6140 17436
rect 6196 17434 6202 17436
rect 5956 17382 5958 17434
rect 6138 17382 6140 17434
rect 5894 17380 5900 17382
rect 5956 17380 5980 17382
rect 6036 17380 6060 17382
rect 6116 17380 6140 17382
rect 6196 17380 6202 17382
rect 5894 17371 6202 17380
rect 6288 17320 6316 22879
rect 6380 22234 6408 23462
rect 6460 23180 6512 23186
rect 6460 23122 6512 23128
rect 6368 22228 6420 22234
rect 6368 22170 6420 22176
rect 6366 22128 6422 22137
rect 6366 22063 6422 22072
rect 6380 22030 6408 22063
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 6368 20868 6420 20874
rect 6368 20810 6420 20816
rect 6380 20777 6408 20810
rect 6366 20768 6422 20777
rect 6366 20703 6422 20712
rect 6368 19848 6420 19854
rect 6368 19790 6420 19796
rect 6380 19417 6408 19790
rect 6366 19408 6422 19417
rect 6366 19343 6422 19352
rect 6196 17292 6316 17320
rect 6000 17264 6052 17270
rect 5828 17202 5948 17218
rect 6000 17206 6052 17212
rect 5828 17196 5960 17202
rect 5828 17190 5908 17196
rect 5908 17138 5960 17144
rect 5920 16969 5948 17138
rect 6012 16998 6040 17206
rect 6000 16992 6052 16998
rect 5906 16960 5962 16969
rect 6000 16934 6052 16940
rect 5906 16895 5962 16904
rect 6196 16454 6224 17292
rect 6380 16538 6408 19343
rect 6472 18766 6500 23122
rect 6564 23118 6592 28070
rect 6840 27962 6868 28614
rect 6656 27934 6868 27962
rect 6656 23746 6684 27934
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6840 27470 6868 27814
rect 6828 27464 6880 27470
rect 6828 27406 6880 27412
rect 6734 27160 6790 27169
rect 6734 27095 6736 27104
rect 6788 27095 6790 27104
rect 6736 27066 6788 27072
rect 6840 26450 6868 27406
rect 6920 27056 6972 27062
rect 6920 26998 6972 27004
rect 6828 26444 6880 26450
rect 6828 26386 6880 26392
rect 6932 26081 6960 26998
rect 7024 26518 7052 28970
rect 7104 28960 7156 28966
rect 7104 28902 7156 28908
rect 7116 28626 7144 28902
rect 7104 28620 7156 28626
rect 7104 28562 7156 28568
rect 7300 28014 7328 32982
rect 7484 32502 7512 33408
rect 7576 33318 7604 33458
rect 7564 33312 7616 33318
rect 7564 33254 7616 33260
rect 7656 33312 7708 33318
rect 7656 33254 7708 33260
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7472 32496 7524 32502
rect 7378 32464 7434 32473
rect 7472 32438 7524 32444
rect 7378 32399 7380 32408
rect 7432 32399 7434 32408
rect 7380 32370 7432 32376
rect 7380 31748 7432 31754
rect 7380 31690 7432 31696
rect 7392 31657 7420 31690
rect 7378 31648 7434 31657
rect 7378 31583 7434 31592
rect 7380 31136 7432 31142
rect 7380 31078 7432 31084
rect 7392 29753 7420 31078
rect 7378 29744 7434 29753
rect 7378 29679 7434 29688
rect 7392 29578 7420 29679
rect 7380 29572 7432 29578
rect 7380 29514 7432 29520
rect 7380 29232 7432 29238
rect 7380 29174 7432 29180
rect 7288 28008 7340 28014
rect 7288 27950 7340 27956
rect 7288 27872 7340 27878
rect 7288 27814 7340 27820
rect 7194 27704 7250 27713
rect 7194 27639 7250 27648
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 7116 26586 7144 27406
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7012 26512 7064 26518
rect 7012 26454 7064 26460
rect 7012 26240 7064 26246
rect 7012 26182 7064 26188
rect 6918 26072 6974 26081
rect 6918 26007 6974 26016
rect 6734 25528 6790 25537
rect 6932 25498 6960 26007
rect 7024 25838 7052 26182
rect 7104 25968 7156 25974
rect 7104 25910 7156 25916
rect 7012 25832 7064 25838
rect 7012 25774 7064 25780
rect 7012 25696 7064 25702
rect 7012 25638 7064 25644
rect 7024 25498 7052 25638
rect 6734 25463 6790 25472
rect 6920 25492 6972 25498
rect 6748 25294 6776 25463
rect 6920 25434 6972 25440
rect 7012 25492 7064 25498
rect 7012 25434 7064 25440
rect 6736 25288 6788 25294
rect 6736 25230 6788 25236
rect 6828 25288 6880 25294
rect 6828 25230 6880 25236
rect 6840 24886 6868 25230
rect 6828 24880 6880 24886
rect 6734 24848 6790 24857
rect 6828 24822 6880 24828
rect 6734 24783 6736 24792
rect 6788 24783 6790 24792
rect 6736 24754 6788 24760
rect 6840 24274 6868 24822
rect 6828 24268 6880 24274
rect 6828 24210 6880 24216
rect 6656 23718 6776 23746
rect 6644 23656 6696 23662
rect 6644 23598 6696 23604
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 6656 21536 6684 23598
rect 6748 23186 6776 23718
rect 6828 23588 6880 23594
rect 6828 23530 6880 23536
rect 6840 23254 6868 23530
rect 6828 23248 6880 23254
rect 6828 23190 6880 23196
rect 6736 23180 6788 23186
rect 6736 23122 6788 23128
rect 6828 23112 6880 23118
rect 6748 23060 6828 23066
rect 6748 23054 6880 23060
rect 6748 23038 6868 23054
rect 6748 22148 6776 23038
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 6840 22250 6868 22578
rect 6932 22438 6960 25434
rect 7012 25356 7064 25362
rect 7012 25298 7064 25304
rect 7024 24342 7052 25298
rect 7116 24410 7144 25910
rect 7208 24834 7236 27639
rect 7300 27033 7328 27814
rect 7286 27024 7342 27033
rect 7286 26959 7342 26968
rect 7288 26580 7340 26586
rect 7288 26522 7340 26528
rect 7300 25945 7328 26522
rect 7286 25936 7342 25945
rect 7286 25871 7342 25880
rect 7288 25832 7340 25838
rect 7288 25774 7340 25780
rect 7300 25430 7328 25774
rect 7392 25430 7420 29174
rect 7288 25424 7340 25430
rect 7288 25366 7340 25372
rect 7380 25424 7432 25430
rect 7380 25366 7432 25372
rect 7484 25242 7512 32438
rect 7576 30598 7604 33050
rect 7668 31482 7696 33254
rect 7760 33114 7788 34020
rect 7932 34060 7984 34066
rect 8116 34060 8168 34066
rect 7984 34020 8064 34048
rect 7932 34002 7984 34008
rect 7840 33652 7892 33658
rect 7840 33594 7892 33600
rect 7748 33108 7800 33114
rect 7748 33050 7800 33056
rect 7852 31940 7880 33594
rect 8036 33454 8064 34020
rect 8116 34002 8168 34008
rect 8024 33448 8076 33454
rect 8024 33390 8076 33396
rect 8036 32570 8064 33390
rect 8312 33266 8340 34190
rect 8576 34196 8628 34202
rect 8576 34138 8628 34144
rect 8588 33969 8616 34138
rect 8772 34134 8800 35022
rect 8864 34626 8892 41386
rect 8956 34746 8984 42162
rect 9048 41290 9076 43046
rect 9232 42684 9260 44540
rect 9416 43314 9444 44540
rect 9404 43308 9456 43314
rect 9404 43250 9456 43256
rect 9496 43308 9548 43314
rect 9600 43296 9628 44540
rect 9680 43716 9732 43722
rect 9680 43658 9732 43664
rect 9548 43268 9628 43296
rect 9496 43250 9548 43256
rect 9692 43246 9720 43658
rect 9680 43240 9732 43246
rect 9680 43182 9732 43188
rect 9680 43104 9732 43110
rect 9680 43046 9732 43052
rect 9692 42838 9720 43046
rect 9680 42832 9732 42838
rect 9680 42774 9732 42780
rect 9496 42696 9548 42702
rect 9232 42656 9496 42684
rect 9496 42638 9548 42644
rect 9632 42566 9688 42571
rect 9128 42560 9180 42566
rect 9126 42528 9128 42537
rect 9632 42562 9732 42566
rect 9688 42560 9732 42562
rect 9180 42528 9182 42537
rect 9688 42506 9732 42508
rect 9632 42502 9732 42506
rect 9632 42497 9688 42502
rect 9126 42463 9182 42472
rect 9588 42356 9640 42362
rect 9588 42298 9640 42304
rect 9496 42220 9548 42226
rect 9496 42162 9548 42168
rect 9508 42106 9536 42162
rect 9416 42078 9536 42106
rect 9128 41608 9180 41614
rect 9126 41576 9128 41585
rect 9180 41576 9182 41585
rect 9126 41511 9182 41520
rect 9048 41262 9260 41290
rect 9232 38654 9260 41262
rect 9416 38865 9444 42078
rect 9496 42016 9548 42022
rect 9496 41958 9548 41964
rect 9508 41818 9536 41958
rect 9496 41812 9548 41818
rect 9496 41754 9548 41760
rect 9600 41414 9628 42298
rect 9784 42294 9812 44540
rect 9864 43852 9916 43858
rect 9864 43794 9916 43800
rect 9876 43314 9904 43794
rect 9968 43432 9996 44540
rect 10152 43858 10180 44540
rect 10140 43852 10192 43858
rect 10140 43794 10192 43800
rect 10140 43648 10192 43654
rect 10336 43602 10364 44540
rect 10140 43590 10192 43596
rect 9968 43404 10088 43432
rect 9864 43308 9916 43314
rect 9864 43250 9916 43256
rect 9864 43104 9916 43110
rect 9864 43046 9916 43052
rect 9772 42288 9824 42294
rect 9772 42230 9824 42236
rect 9772 42016 9824 42022
rect 9772 41958 9824 41964
rect 9784 41721 9812 41958
rect 9770 41712 9826 41721
rect 9770 41647 9826 41656
rect 9508 41386 9628 41414
rect 9402 38856 9458 38865
rect 9402 38791 9458 38800
rect 9232 38626 9352 38654
rect 9128 38208 9180 38214
rect 9128 38150 9180 38156
rect 9036 37732 9088 37738
rect 9036 37674 9088 37680
rect 9048 37252 9076 37674
rect 9036 37246 9088 37252
rect 9036 37188 9088 37194
rect 9036 37120 9088 37126
rect 9036 37062 9088 37068
rect 9048 36786 9076 37062
rect 9036 36780 9088 36786
rect 9036 36722 9088 36728
rect 9036 36576 9088 36582
rect 9036 36518 9088 36524
rect 9048 36174 9076 36518
rect 9036 36168 9088 36174
rect 9036 36110 9088 36116
rect 9048 35086 9076 36110
rect 9036 35080 9088 35086
rect 9036 35022 9088 35028
rect 9048 34785 9076 35022
rect 9034 34776 9090 34785
rect 8944 34740 8996 34746
rect 9140 34746 9168 38150
rect 9220 37664 9272 37670
rect 9220 37606 9272 37612
rect 9034 34711 9090 34720
rect 9128 34740 9180 34746
rect 8944 34682 8996 34688
rect 9128 34682 9180 34688
rect 8864 34598 9168 34626
rect 8852 34536 8904 34542
rect 8852 34478 8904 34484
rect 8944 34536 8996 34542
rect 8944 34478 8996 34484
rect 8864 34202 8892 34478
rect 8852 34196 8904 34202
rect 8852 34138 8904 34144
rect 8760 34128 8812 34134
rect 8760 34070 8812 34076
rect 8668 34060 8720 34066
rect 8668 34002 8720 34008
rect 8574 33960 8630 33969
rect 8574 33895 8630 33904
rect 8484 33856 8536 33862
rect 8484 33798 8536 33804
rect 8496 33318 8524 33798
rect 8220 33238 8340 33266
rect 8484 33312 8536 33318
rect 8680 33300 8708 34002
rect 8760 33992 8812 33998
rect 8760 33934 8812 33940
rect 8772 33658 8800 33934
rect 8956 33862 8984 34478
rect 9036 34468 9088 34474
rect 9036 34410 9088 34416
rect 8944 33856 8996 33862
rect 9048 33833 9076 34410
rect 8944 33798 8996 33804
rect 9034 33824 9090 33833
rect 8760 33652 8812 33658
rect 8760 33594 8812 33600
rect 8850 33552 8906 33561
rect 8956 33522 8984 33798
rect 9034 33759 9090 33768
rect 8850 33487 8852 33496
rect 8904 33487 8906 33496
rect 8944 33516 8996 33522
rect 8852 33458 8904 33464
rect 8944 33458 8996 33464
rect 8680 33272 8800 33300
rect 8484 33254 8536 33260
rect 8220 33114 8248 33238
rect 8367 33212 8675 33221
rect 8367 33210 8373 33212
rect 8429 33210 8453 33212
rect 8509 33210 8533 33212
rect 8589 33210 8613 33212
rect 8669 33210 8675 33212
rect 8429 33158 8431 33210
rect 8611 33158 8613 33210
rect 8367 33156 8373 33158
rect 8429 33156 8453 33158
rect 8509 33156 8533 33158
rect 8589 33156 8613 33158
rect 8669 33156 8675 33158
rect 8367 33147 8675 33156
rect 8208 33108 8260 33114
rect 8208 33050 8260 33056
rect 8576 33040 8628 33046
rect 8574 33008 8576 33017
rect 8628 33008 8630 33017
rect 8574 32943 8630 32952
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 8024 32564 8076 32570
rect 8024 32506 8076 32512
rect 7852 31912 7972 31940
rect 7840 31680 7892 31686
rect 7840 31622 7892 31628
rect 7656 31476 7708 31482
rect 7656 31418 7708 31424
rect 7564 30592 7616 30598
rect 7564 30534 7616 30540
rect 7562 30424 7618 30433
rect 7668 30394 7696 31418
rect 7852 30802 7880 31622
rect 7944 31498 7972 31912
rect 8022 31784 8078 31793
rect 8128 31770 8156 32846
rect 8367 32124 8675 32133
rect 8367 32122 8373 32124
rect 8429 32122 8453 32124
rect 8509 32122 8533 32124
rect 8589 32122 8613 32124
rect 8669 32122 8675 32124
rect 8429 32070 8431 32122
rect 8611 32070 8613 32122
rect 8367 32068 8373 32070
rect 8429 32068 8453 32070
rect 8509 32068 8533 32070
rect 8589 32068 8613 32070
rect 8669 32068 8675 32070
rect 8367 32059 8675 32068
rect 8078 31742 8156 31770
rect 8022 31719 8078 31728
rect 8114 31512 8170 31521
rect 7944 31470 8114 31498
rect 8114 31447 8170 31456
rect 8206 31376 8262 31385
rect 8206 31311 8208 31320
rect 8260 31311 8262 31320
rect 8208 31282 8260 31288
rect 8208 31136 8260 31142
rect 8208 31078 8260 31084
rect 8114 30968 8170 30977
rect 8220 30938 8248 31078
rect 8367 31036 8675 31045
rect 8367 31034 8373 31036
rect 8429 31034 8453 31036
rect 8509 31034 8533 31036
rect 8589 31034 8613 31036
rect 8669 31034 8675 31036
rect 8429 30982 8431 31034
rect 8611 30982 8613 31034
rect 8367 30980 8373 30982
rect 8429 30980 8453 30982
rect 8509 30980 8533 30982
rect 8589 30980 8613 30982
rect 8669 30980 8675 30982
rect 8367 30971 8675 30980
rect 8114 30903 8170 30912
rect 8208 30932 8260 30938
rect 7840 30796 7892 30802
rect 7840 30738 7892 30744
rect 7840 30660 7892 30666
rect 7840 30602 7892 30608
rect 7932 30660 7984 30666
rect 7932 30602 7984 30608
rect 7562 30359 7618 30368
rect 7656 30388 7708 30394
rect 7576 30258 7604 30359
rect 7656 30330 7708 30336
rect 7564 30252 7616 30258
rect 7564 30194 7616 30200
rect 7576 29238 7604 30194
rect 7656 29504 7708 29510
rect 7656 29446 7708 29452
rect 7668 29306 7696 29446
rect 7656 29300 7708 29306
rect 7656 29242 7708 29248
rect 7564 29232 7616 29238
rect 7564 29174 7616 29180
rect 7746 29200 7802 29209
rect 7746 29135 7802 29144
rect 7656 28008 7708 28014
rect 7656 27950 7708 27956
rect 7564 26988 7616 26994
rect 7564 26930 7616 26936
rect 7576 26586 7604 26930
rect 7564 26580 7616 26586
rect 7564 26522 7616 26528
rect 7564 26308 7616 26314
rect 7564 26250 7616 26256
rect 7576 25809 7604 26250
rect 7562 25800 7618 25809
rect 7562 25735 7618 25744
rect 7392 25214 7512 25242
rect 7208 24806 7328 24834
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 7196 24404 7248 24410
rect 7196 24346 7248 24352
rect 7012 24336 7064 24342
rect 7012 24278 7064 24284
rect 7102 23896 7158 23905
rect 7102 23831 7158 23840
rect 7116 23662 7144 23831
rect 7104 23656 7156 23662
rect 7104 23598 7156 23604
rect 6920 22432 6972 22438
rect 6920 22374 6972 22380
rect 6840 22222 6960 22250
rect 6748 22120 6868 22148
rect 6736 21548 6788 21554
rect 6656 21508 6736 21536
rect 6656 20913 6684 21508
rect 6736 21490 6788 21496
rect 6642 20904 6698 20913
rect 6642 20839 6698 20848
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6748 20398 6776 20538
rect 6736 20392 6788 20398
rect 6736 20334 6788 20340
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6550 19544 6606 19553
rect 6550 19479 6606 19488
rect 6564 18970 6592 19479
rect 6748 18970 6776 19926
rect 6840 19428 6868 22120
rect 6932 19530 6960 22222
rect 6932 19502 7052 19530
rect 6840 19400 6960 19428
rect 6828 19236 6880 19242
rect 6828 19178 6880 19184
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6288 16510 6408 16538
rect 5816 16448 5868 16454
rect 5816 16390 5868 16396
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 5828 15502 5856 16390
rect 5894 16348 6202 16357
rect 5894 16346 5900 16348
rect 5956 16346 5980 16348
rect 6036 16346 6060 16348
rect 6116 16346 6140 16348
rect 6196 16346 6202 16348
rect 5956 16294 5958 16346
rect 6138 16294 6140 16346
rect 5894 16292 5900 16294
rect 5956 16292 5980 16294
rect 6036 16292 6060 16294
rect 6116 16292 6140 16294
rect 6196 16292 6202 16294
rect 5894 16283 6202 16292
rect 6000 16040 6052 16046
rect 5920 16000 6000 16028
rect 5920 15881 5948 16000
rect 6000 15982 6052 15988
rect 6184 15904 6236 15910
rect 5906 15872 5962 15881
rect 6184 15846 6236 15852
rect 5906 15807 5962 15816
rect 6196 15706 6224 15846
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6288 15502 6316 16510
rect 6368 16448 6420 16454
rect 6368 16390 6420 16396
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 5828 14414 5856 15438
rect 5894 15260 6202 15269
rect 5894 15258 5900 15260
rect 5956 15258 5980 15260
rect 6036 15258 6060 15260
rect 6116 15258 6140 15260
rect 6196 15258 6202 15260
rect 5956 15206 5958 15258
rect 6138 15206 6140 15258
rect 5894 15204 5900 15206
rect 5956 15204 5980 15206
rect 6036 15204 6060 15206
rect 6116 15204 6140 15206
rect 6196 15204 6202 15206
rect 5894 15195 6202 15204
rect 6182 14784 6238 14793
rect 6182 14719 6238 14728
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5828 13802 5856 14350
rect 6196 14346 6224 14719
rect 6288 14657 6316 15438
rect 6274 14648 6330 14657
rect 6274 14583 6330 14592
rect 6184 14340 6236 14346
rect 6184 14282 6236 14288
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 5894 14172 6202 14181
rect 5894 14170 5900 14172
rect 5956 14170 5980 14172
rect 6036 14170 6060 14172
rect 6116 14170 6140 14172
rect 6196 14170 6202 14172
rect 5956 14118 5958 14170
rect 6138 14118 6140 14170
rect 5894 14116 5900 14118
rect 5956 14116 5980 14118
rect 6036 14116 6060 14118
rect 6116 14116 6140 14118
rect 6196 14116 6202 14118
rect 5894 14107 6202 14116
rect 6092 13864 6144 13870
rect 6092 13806 6144 13812
rect 5816 13796 5868 13802
rect 5816 13738 5868 13744
rect 5828 13546 5856 13738
rect 5998 13560 6054 13569
rect 5828 13518 5998 13546
rect 5998 13495 6054 13504
rect 5814 13424 5870 13433
rect 6104 13394 6132 13806
rect 5814 13359 5870 13368
rect 6092 13388 6144 13394
rect 5828 12730 5856 13359
rect 6092 13330 6144 13336
rect 5894 13084 6202 13093
rect 5894 13082 5900 13084
rect 5956 13082 5980 13084
rect 6036 13082 6060 13084
rect 6116 13082 6140 13084
rect 6196 13082 6202 13084
rect 5956 13030 5958 13082
rect 6138 13030 6140 13082
rect 5894 13028 5900 13030
rect 5956 13028 5980 13030
rect 6036 13028 6060 13030
rect 6116 13028 6140 13030
rect 6196 13028 6202 13030
rect 5894 13019 6202 13028
rect 5828 12702 5948 12730
rect 5686 12566 5764 12594
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5630 12543 5686 12552
rect 5724 12436 5776 12442
rect 5552 12396 5638 12424
rect 5610 12356 5638 12396
rect 5724 12378 5776 12384
rect 5610 12328 5672 12356
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5552 12073 5580 12174
rect 5538 12064 5594 12073
rect 5538 11999 5594 12008
rect 5538 11928 5594 11937
rect 5644 11898 5672 12328
rect 5736 12238 5764 12378
rect 5828 12306 5856 12582
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5920 12084 5948 12702
rect 5722 12064 5778 12073
rect 5722 11999 5778 12008
rect 5828 12056 5948 12084
rect 5538 11863 5540 11872
rect 5592 11863 5594 11872
rect 5632 11892 5684 11898
rect 5540 11834 5592 11840
rect 5632 11834 5684 11840
rect 5736 11812 5764 11999
rect 5828 11880 5856 12056
rect 5894 11996 6202 12005
rect 5894 11994 5900 11996
rect 5956 11994 5980 11996
rect 6036 11994 6060 11996
rect 6116 11994 6140 11996
rect 6196 11994 6202 11996
rect 5956 11942 5958 11994
rect 6138 11942 6140 11994
rect 5894 11940 5900 11942
rect 5956 11940 5980 11942
rect 6036 11940 6060 11942
rect 6116 11940 6140 11942
rect 6196 11940 6202 11942
rect 5894 11931 6202 11940
rect 5828 11852 6224 11880
rect 5736 11784 5948 11812
rect 6196 11801 6224 11852
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5446 11384 5502 11393
rect 5552 11370 5580 11698
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5502 11342 5580 11370
rect 5446 11319 5502 11328
rect 5644 11268 5672 11494
rect 5460 11240 5672 11268
rect 5460 11121 5488 11240
rect 5736 11200 5764 11630
rect 5920 11626 5948 11784
rect 6182 11792 6238 11801
rect 6092 11756 6144 11762
rect 6182 11727 6184 11736
rect 6092 11698 6144 11704
rect 6236 11727 6238 11736
rect 6184 11698 6236 11704
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5908 11620 5960 11626
rect 5908 11562 5960 11568
rect 5828 11506 5856 11562
rect 5828 11478 6040 11506
rect 6012 11234 6040 11478
rect 6104 11393 6132 11698
rect 6288 11626 6316 14214
rect 6380 14113 6408 16390
rect 6472 16250 6500 18702
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6564 16454 6592 17614
rect 6656 16794 6684 18702
rect 6840 17954 6868 19178
rect 6748 17926 6868 17954
rect 6644 16788 6696 16794
rect 6644 16730 6696 16736
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6460 16244 6512 16250
rect 6460 16186 6512 16192
rect 6564 16046 6592 16390
rect 6748 16046 6776 17926
rect 6932 17746 6960 19400
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6920 17740 6972 17746
rect 6920 17682 6972 17688
rect 6840 17338 6868 17682
rect 6828 17332 6880 17338
rect 6828 17274 6880 17280
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6472 15042 6500 15982
rect 6564 15201 6592 15982
rect 6748 15745 6776 15982
rect 6734 15736 6790 15745
rect 6734 15671 6790 15680
rect 6642 15600 6698 15609
rect 6698 15558 6776 15586
rect 6642 15535 6698 15544
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6550 15192 6606 15201
rect 6550 15127 6606 15136
rect 6550 15056 6606 15065
rect 6472 15014 6550 15042
rect 6550 14991 6606 15000
rect 6656 14958 6684 15302
rect 6552 14952 6604 14958
rect 6552 14894 6604 14900
rect 6644 14952 6696 14958
rect 6644 14894 6696 14900
rect 6460 14884 6512 14890
rect 6460 14826 6512 14832
rect 6366 14104 6422 14113
rect 6366 14039 6422 14048
rect 6472 13546 6500 14826
rect 6564 13938 6592 14894
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6380 13518 6500 13546
rect 6380 13394 6408 13518
rect 6460 13456 6512 13462
rect 6460 13398 6512 13404
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6472 13274 6500 13398
rect 6380 13246 6500 13274
rect 6380 13025 6408 13246
rect 6564 13190 6592 13874
rect 6644 13456 6696 13462
rect 6644 13398 6696 13404
rect 6552 13184 6604 13190
rect 6458 13152 6514 13161
rect 6552 13126 6604 13132
rect 6458 13087 6514 13096
rect 6366 13016 6422 13025
rect 6366 12951 6422 12960
rect 6366 12744 6422 12753
rect 6366 12679 6368 12688
rect 6420 12679 6422 12688
rect 6368 12650 6420 12656
rect 6368 12368 6420 12374
rect 6368 12310 6420 12316
rect 6380 11694 6408 12310
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6090 11384 6146 11393
rect 6090 11319 6146 11328
rect 5644 11172 5764 11200
rect 6010 11206 6040 11234
rect 5558 11144 5610 11150
rect 5446 11112 5502 11121
rect 5446 11047 5502 11056
rect 5552 11092 5558 11132
rect 5552 11086 5610 11092
rect 5552 10520 5580 11086
rect 5460 10492 5580 10520
rect 5460 10198 5488 10492
rect 5538 10432 5594 10441
rect 5538 10367 5594 10376
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5448 9920 5500 9926
rect 5552 9908 5580 10367
rect 5644 10062 5672 11172
rect 6010 11132 6038 11206
rect 6010 11104 6040 11132
rect 5736 11070 5948 11098
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5552 9880 5672 9908
rect 5448 9862 5500 9868
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5460 9636 5488 9862
rect 5354 9616 5410 9625
rect 5460 9608 5580 9636
rect 5448 9570 5500 9576
rect 5410 9560 5448 9568
rect 5264 9546 5316 9552
rect 5354 9551 5448 9560
rect 5368 9540 5448 9551
rect 5552 9518 5580 9608
rect 5448 9512 5500 9518
rect 5540 9512 5592 9518
rect 5316 9494 5396 9500
rect 5264 9488 5396 9494
rect 5276 9472 5396 9488
rect 5368 9353 5396 9472
rect 5540 9454 5592 9460
rect 5354 9344 5410 9353
rect 5354 9279 5410 9288
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5080 8968 5132 8974
rect 5080 8910 5132 8916
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 4724 8316 4936 8344
rect 4724 7274 4752 8316
rect 5172 8288 5224 8294
rect 4908 8248 5172 8276
rect 4908 7886 4936 8248
rect 4896 7880 4948 7886
rect 4802 7848 4858 7857
rect 4896 7822 4948 7828
rect 4802 7783 4858 7792
rect 4712 7268 4764 7274
rect 4712 7210 4764 7216
rect 4816 6848 4844 7783
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4908 7342 4936 7686
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4724 6820 4844 6848
rect 4724 6712 4752 6820
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4724 6684 4844 6712
rect 4710 6624 4766 6633
rect 4710 6559 4766 6568
rect 4724 6322 4752 6559
rect 4712 6316 4764 6322
rect 4712 6258 4764 6264
rect 4724 4729 4752 6258
rect 4710 4720 4766 4729
rect 4710 4655 4766 4664
rect 4580 3488 4660 3516
rect 4528 3470 4580 3476
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4342 2615 4398 2624
rect 4436 2644 4488 2650
rect 3790 2479 3846 2488
rect 4068 2508 4120 2514
rect 3804 2446 3832 2479
rect 4068 2450 4120 2456
rect 3424 2440 3476 2446
rect 3344 2400 3424 2428
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 2596 2032 2648 2038
rect 2596 1974 2648 1980
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 2504 1556 2556 1562
rect 2504 1498 2556 1504
rect 2412 1284 2464 1290
rect 2412 1226 2464 1232
rect 2320 468 2372 474
rect 2320 410 2372 416
rect 2424 160 2452 1226
rect 2596 1216 2648 1222
rect 2596 1158 2648 1164
rect 2608 160 2636 1158
rect 2792 160 2820 1838
rect 2976 160 3004 2314
rect 3240 1964 3292 1970
rect 3240 1906 3292 1912
rect 2410 -300 2466 160
rect 2594 -300 2650 160
rect 2778 -300 2834 160
rect 2962 -300 3018 160
rect 3146 82 3202 160
rect 3252 82 3280 1906
rect 3344 1272 3372 2400
rect 3424 2382 3476 2388
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 4158 2408 4214 2417
rect 4068 2372 4120 2378
rect 4158 2343 4214 2352
rect 4068 2314 4120 2320
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3988 2088 4016 2246
rect 3896 2060 4016 2088
rect 3422 1660 3730 1669
rect 3422 1658 3428 1660
rect 3484 1658 3508 1660
rect 3564 1658 3588 1660
rect 3644 1658 3668 1660
rect 3724 1658 3730 1660
rect 3484 1606 3486 1658
rect 3666 1606 3668 1658
rect 3422 1604 3428 1606
rect 3484 1604 3508 1606
rect 3564 1604 3588 1606
rect 3644 1604 3668 1606
rect 3724 1604 3730 1606
rect 3422 1595 3730 1604
rect 3700 1352 3752 1358
rect 3700 1294 3752 1300
rect 3344 1244 3556 1272
rect 3332 672 3384 678
rect 3332 614 3384 620
rect 3344 160 3372 614
rect 3528 160 3556 1244
rect 3712 160 3740 1294
rect 3896 649 3924 2060
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 3882 640 3938 649
rect 3882 575 3938 584
rect 3146 54 3280 82
rect 3146 -300 3202 54
rect 3330 -300 3386 160
rect 3514 -300 3570 160
rect 3698 -300 3754 160
rect 3882 82 3938 160
rect 3988 82 4016 1906
rect 4080 160 4108 2314
rect 4172 2106 4200 2343
rect 4160 2100 4212 2106
rect 4160 2042 4212 2048
rect 4160 1964 4212 1970
rect 4160 1906 4212 1912
rect 4172 1562 4200 1906
rect 4356 1562 4384 2615
rect 4436 2586 4488 2592
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4540 2020 4568 2382
rect 4448 1992 4568 2020
rect 4160 1556 4212 1562
rect 4160 1498 4212 1504
rect 4344 1556 4396 1562
rect 4344 1498 4396 1504
rect 4448 1442 4476 1992
rect 4632 1952 4660 2926
rect 4540 1924 4660 1952
rect 4540 1766 4568 1924
rect 4712 1896 4764 1902
rect 4632 1856 4712 1884
rect 4528 1760 4580 1766
rect 4528 1702 4580 1708
rect 4356 1414 4476 1442
rect 3882 54 4016 82
rect 3882 -300 3938 54
rect 4066 -300 4122 160
rect 4250 82 4306 160
rect 4356 82 4384 1414
rect 4436 1284 4488 1290
rect 4436 1226 4488 1232
rect 4528 1284 4580 1290
rect 4528 1226 4580 1232
rect 4448 160 4476 1226
rect 4540 746 4568 1226
rect 4528 740 4580 746
rect 4528 682 4580 688
rect 4632 160 4660 1856
rect 4712 1838 4764 1844
rect 4816 1850 4844 6684
rect 4908 6089 4936 6734
rect 5000 6458 5028 7210
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4986 6352 5042 6361
rect 4986 6287 5042 6296
rect 4894 6080 4950 6089
rect 4894 6015 4950 6024
rect 5000 5930 5028 6287
rect 4908 5902 5028 5930
rect 4908 3176 4936 5902
rect 5092 5702 5120 8248
rect 5172 8230 5224 8236
rect 5172 8084 5224 8090
rect 5276 8072 5304 8774
rect 5224 8044 5304 8072
rect 5172 8026 5224 8032
rect 5262 7984 5318 7993
rect 5262 7919 5318 7928
rect 5170 7712 5226 7721
rect 5170 7647 5226 7656
rect 5184 6322 5212 7647
rect 5276 7410 5304 7919
rect 5264 7404 5316 7410
rect 5264 7346 5316 7352
rect 5276 7206 5304 7346
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5262 6896 5318 6905
rect 5262 6831 5318 6840
rect 5276 6798 5304 6831
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5092 5674 5212 5702
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4986 4856 5042 4865
rect 4986 4791 4988 4800
rect 5040 4791 5042 4800
rect 4988 4762 5040 4768
rect 5092 3942 5120 5578
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4908 3148 5120 3176
rect 4986 3088 5042 3097
rect 4986 3023 5042 3032
rect 4896 2848 4948 2854
rect 4896 2790 4948 2796
rect 4908 2106 4936 2790
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 5000 1970 5028 3023
rect 4988 1964 5040 1970
rect 4988 1906 5040 1912
rect 4816 1822 5028 1850
rect 5000 1562 5028 1822
rect 5092 1562 5120 3148
rect 5184 2650 5212 5674
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5170 2408 5226 2417
rect 5170 2343 5226 2352
rect 5184 1902 5212 2343
rect 5172 1896 5224 1902
rect 5172 1838 5224 1844
rect 4988 1556 5040 1562
rect 4988 1498 5040 1504
rect 5080 1556 5132 1562
rect 5080 1498 5132 1504
rect 5276 1494 5304 6598
rect 5368 5409 5396 9279
rect 5558 9172 5610 9178
rect 5552 9120 5558 9160
rect 5552 9114 5610 9120
rect 5552 7886 5580 9114
rect 5644 7970 5672 9880
rect 5736 8498 5764 11070
rect 5920 11014 5948 11070
rect 6012 11014 6040 11104
rect 5816 11008 5868 11014
rect 5816 10950 5868 10956
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 5828 10606 5856 10950
rect 5894 10908 6202 10917
rect 5894 10906 5900 10908
rect 5956 10906 5980 10908
rect 6036 10906 6060 10908
rect 6116 10906 6140 10908
rect 6196 10906 6202 10908
rect 5956 10854 5958 10906
rect 6138 10854 6140 10906
rect 5894 10852 5900 10854
rect 5956 10852 5980 10854
rect 6036 10852 6060 10854
rect 6116 10852 6140 10854
rect 6196 10852 6202 10854
rect 5894 10843 6202 10852
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5920 10452 5948 10610
rect 6012 10470 6040 10678
rect 6184 10600 6236 10606
rect 6184 10542 6236 10548
rect 5828 10424 5948 10452
rect 6000 10464 6052 10470
rect 5828 8974 5856 10424
rect 6000 10406 6052 10412
rect 6012 10130 6040 10406
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6196 9926 6224 10542
rect 6184 9920 6236 9926
rect 6184 9862 6236 9868
rect 5894 9820 6202 9829
rect 5894 9818 5900 9820
rect 5956 9818 5980 9820
rect 6036 9818 6060 9820
rect 6116 9818 6140 9820
rect 6196 9818 6202 9820
rect 5956 9766 5958 9818
rect 6138 9766 6140 9818
rect 5894 9764 5900 9766
rect 5956 9764 5980 9766
rect 6036 9764 6060 9766
rect 6116 9764 6140 9766
rect 6196 9764 6202 9766
rect 5894 9755 6202 9764
rect 6182 9616 6238 9625
rect 6104 9574 6182 9602
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5998 9480 6054 9489
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5920 8820 5948 9454
rect 5998 9415 6054 9424
rect 6012 8906 6040 9415
rect 6104 9042 6132 9574
rect 6182 9551 6238 9560
rect 6288 9466 6316 11562
rect 6380 11121 6408 11630
rect 6366 11112 6422 11121
rect 6366 11047 6422 11056
rect 6368 11008 6420 11014
rect 6368 10950 6420 10956
rect 6380 10674 6408 10950
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6380 9586 6408 10610
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6196 9438 6316 9466
rect 6196 9217 6224 9438
rect 6276 9376 6328 9382
rect 6276 9318 6328 9324
rect 6182 9208 6238 9217
rect 6182 9143 6238 9152
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 5828 8792 5948 8820
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 5722 8256 5778 8265
rect 5722 8191 5778 8200
rect 5736 8090 5764 8191
rect 5828 8129 5856 8792
rect 5894 8732 6202 8741
rect 5894 8730 5900 8732
rect 5956 8730 5980 8732
rect 6036 8730 6060 8732
rect 6116 8730 6140 8732
rect 6196 8730 6202 8732
rect 5956 8678 5958 8730
rect 6138 8678 6140 8730
rect 5894 8676 5900 8678
rect 5956 8676 5980 8678
rect 6036 8676 6060 8678
rect 6116 8676 6140 8678
rect 6196 8676 6202 8678
rect 5894 8667 6202 8676
rect 6092 8560 6144 8566
rect 6090 8528 6092 8537
rect 6144 8528 6146 8537
rect 5908 8492 5960 8498
rect 6090 8463 6146 8472
rect 5908 8434 5960 8440
rect 5814 8120 5870 8129
rect 5724 8084 5776 8090
rect 5814 8055 5870 8064
rect 5724 8026 5776 8032
rect 5644 7942 5764 7970
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5552 7002 5580 7346
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5644 6866 5672 7822
rect 5736 7460 5764 7942
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 5828 7528 5856 7890
rect 5920 7750 5948 8434
rect 5998 8256 6054 8265
rect 5998 8191 6054 8200
rect 6012 7818 6040 8191
rect 6104 7954 6132 8463
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 8129 6224 8366
rect 6182 8120 6238 8129
rect 6182 8055 6184 8064
rect 6236 8055 6238 8064
rect 6184 8026 6236 8032
rect 6092 7948 6144 7954
rect 6092 7890 6144 7896
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5894 7644 6202 7653
rect 5894 7642 5900 7644
rect 5956 7642 5980 7644
rect 6036 7642 6060 7644
rect 6116 7642 6140 7644
rect 6196 7642 6202 7644
rect 5956 7590 5958 7642
rect 6138 7590 6140 7642
rect 5894 7588 5900 7590
rect 5956 7588 5980 7590
rect 6036 7588 6060 7590
rect 6116 7588 6140 7590
rect 6196 7588 6202 7590
rect 5894 7579 6202 7588
rect 5828 7500 6040 7528
rect 5736 7432 5948 7460
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5630 6488 5686 6497
rect 5630 6423 5632 6432
rect 5684 6423 5686 6432
rect 5632 6394 5684 6400
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5540 5704 5592 5710
rect 5538 5672 5540 5681
rect 5592 5672 5594 5681
rect 5538 5607 5594 5616
rect 5540 5568 5592 5574
rect 5540 5510 5592 5516
rect 5354 5400 5410 5409
rect 5354 5335 5410 5344
rect 5448 5364 5500 5370
rect 5448 5306 5500 5312
rect 5356 5228 5408 5234
rect 5460 5216 5488 5306
rect 5552 5234 5580 5510
rect 5408 5188 5488 5216
rect 5540 5228 5592 5234
rect 5356 5170 5408 5176
rect 5540 5170 5592 5176
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 4282 5396 4966
rect 5446 4720 5502 4729
rect 5446 4655 5502 4664
rect 5460 4554 5488 4655
rect 5448 4548 5500 4554
rect 5448 4490 5500 4496
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5460 3670 5488 4490
rect 5644 4298 5672 6258
rect 5552 4270 5672 4298
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5356 3392 5408 3398
rect 5356 3334 5408 3340
rect 5368 2650 5396 3334
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5460 2428 5488 3402
rect 5552 3126 5580 4270
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5540 3120 5592 3126
rect 5540 3062 5592 3068
rect 5644 2854 5672 3878
rect 5736 3534 5764 7142
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5828 6322 5856 6734
rect 5920 6662 5948 7432
rect 6012 6798 6040 7500
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 6104 6905 6132 7278
rect 6090 6896 6146 6905
rect 6090 6831 6146 6840
rect 6196 6798 6224 7346
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 6184 6792 6236 6798
rect 6184 6734 6236 6740
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5894 6556 6202 6565
rect 5894 6554 5900 6556
rect 5956 6554 5980 6556
rect 6036 6554 6060 6556
rect 6116 6554 6140 6556
rect 6196 6554 6202 6556
rect 5956 6502 5958 6554
rect 6138 6502 6140 6554
rect 5894 6500 5900 6502
rect 5956 6500 5980 6502
rect 6036 6500 6060 6502
rect 6116 6500 6140 6502
rect 6196 6500 6202 6502
rect 5894 6491 6202 6500
rect 6288 6458 6316 9318
rect 6380 9178 6408 9522
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6380 7290 6408 8910
rect 6472 7857 6500 13087
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11286 6592 12038
rect 6656 11354 6684 13398
rect 6748 13161 6776 15558
rect 6840 15473 6868 16730
rect 6826 15464 6882 15473
rect 6826 15399 6882 15408
rect 6826 15056 6882 15065
rect 6826 14991 6882 15000
rect 6734 13152 6790 13161
rect 6734 13087 6790 13096
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6644 11348 6696 11354
rect 6644 11290 6696 11296
rect 6552 11280 6604 11286
rect 6552 11222 6604 11228
rect 6644 11144 6696 11150
rect 6550 11112 6606 11121
rect 6644 11086 6696 11092
rect 6550 11047 6606 11056
rect 6564 9722 6592 11047
rect 6656 10674 6684 11086
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6748 10418 6776 12922
rect 6840 12374 6868 14991
rect 6932 14890 6960 17682
rect 7024 16794 7052 19502
rect 7116 17882 7144 23598
rect 7208 22574 7236 24346
rect 7300 23100 7328 24806
rect 7392 23168 7420 25214
rect 7472 25152 7524 25158
rect 7472 25094 7524 25100
rect 7484 24954 7512 25094
rect 7472 24948 7524 24954
rect 7472 24890 7524 24896
rect 7668 24449 7696 27950
rect 7760 26330 7788 29135
rect 7852 28506 7880 30602
rect 7944 28694 7972 30602
rect 8128 30598 8156 30903
rect 8772 30920 8800 33272
rect 8850 33144 8906 33153
rect 8850 33079 8906 33088
rect 8864 32978 8892 33079
rect 9034 33008 9090 33017
rect 8852 32972 8904 32978
rect 8852 32914 8904 32920
rect 8956 32966 9034 32994
rect 8956 32842 8984 32966
rect 9034 32943 9090 32952
rect 9034 32872 9090 32881
rect 8944 32836 8996 32842
rect 8864 32796 8944 32824
rect 8864 31754 8892 32796
rect 9034 32807 9090 32816
rect 8944 32778 8996 32784
rect 8944 32360 8996 32366
rect 8944 32302 8996 32308
rect 8956 31793 8984 32302
rect 8942 31784 8998 31793
rect 8852 31748 8904 31754
rect 8942 31719 8998 31728
rect 8852 31690 8904 31696
rect 8208 30874 8260 30880
rect 8680 30892 8800 30920
rect 8300 30728 8352 30734
rect 8206 30696 8262 30705
rect 8300 30670 8352 30676
rect 8484 30728 8536 30734
rect 8484 30670 8536 30676
rect 8206 30631 8262 30640
rect 8116 30592 8168 30598
rect 8036 30552 8116 30580
rect 7932 28688 7984 28694
rect 7932 28630 7984 28636
rect 7852 28478 7972 28506
rect 7840 27668 7892 27674
rect 7840 27610 7892 27616
rect 7852 26926 7880 27610
rect 7944 26994 7972 28478
rect 8036 27146 8064 30552
rect 8116 30534 8168 30540
rect 8116 30048 8168 30054
rect 8116 29990 8168 29996
rect 8128 28529 8156 29990
rect 8220 29646 8248 30631
rect 8312 30394 8340 30670
rect 8300 30388 8352 30394
rect 8300 30330 8352 30336
rect 8496 30190 8524 30670
rect 8576 30592 8628 30598
rect 8576 30534 8628 30540
rect 8588 30190 8616 30534
rect 8680 30258 8708 30892
rect 8852 30864 8904 30870
rect 8852 30806 8904 30812
rect 8668 30252 8720 30258
rect 8668 30194 8720 30200
rect 8484 30184 8536 30190
rect 8484 30126 8536 30132
rect 8576 30184 8628 30190
rect 8576 30126 8628 30132
rect 8760 30048 8812 30054
rect 8760 29990 8812 29996
rect 8367 29948 8675 29957
rect 8367 29946 8373 29948
rect 8429 29946 8453 29948
rect 8509 29946 8533 29948
rect 8589 29946 8613 29948
rect 8669 29946 8675 29948
rect 8429 29894 8431 29946
rect 8611 29894 8613 29946
rect 8367 29892 8373 29894
rect 8429 29892 8453 29894
rect 8509 29892 8533 29894
rect 8589 29892 8613 29894
rect 8669 29892 8675 29894
rect 8367 29883 8675 29892
rect 8208 29640 8260 29646
rect 8208 29582 8260 29588
rect 8300 29572 8352 29578
rect 8300 29514 8352 29520
rect 8208 29300 8260 29306
rect 8208 29242 8260 29248
rect 8114 28520 8170 28529
rect 8114 28455 8170 28464
rect 8220 28404 8248 29242
rect 8312 29073 8340 29514
rect 8298 29064 8354 29073
rect 8298 28999 8354 29008
rect 8367 28860 8675 28869
rect 8367 28858 8373 28860
rect 8429 28858 8453 28860
rect 8509 28858 8533 28860
rect 8589 28858 8613 28860
rect 8669 28858 8675 28860
rect 8429 28806 8431 28858
rect 8611 28806 8613 28858
rect 8367 28804 8373 28806
rect 8429 28804 8453 28806
rect 8509 28804 8533 28806
rect 8589 28804 8613 28806
rect 8669 28804 8675 28806
rect 8367 28795 8675 28804
rect 8772 28762 8800 29990
rect 8760 28756 8812 28762
rect 8760 28698 8812 28704
rect 8298 28656 8354 28665
rect 8298 28591 8354 28600
rect 8312 28422 8340 28591
rect 8668 28552 8720 28558
rect 8668 28494 8720 28500
rect 8128 28376 8248 28404
rect 8300 28416 8352 28422
rect 8128 27538 8156 28376
rect 8300 28358 8352 28364
rect 8680 28218 8708 28494
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 8208 28144 8260 28150
rect 8208 28086 8260 28092
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 8036 27118 8156 27146
rect 8128 27062 8156 27118
rect 8116 27056 8168 27062
rect 8220 27033 8248 28086
rect 8367 27772 8675 27781
rect 8367 27770 8373 27772
rect 8429 27770 8453 27772
rect 8509 27770 8533 27772
rect 8589 27770 8613 27772
rect 8669 27770 8675 27772
rect 8429 27718 8431 27770
rect 8611 27718 8613 27770
rect 8367 27716 8373 27718
rect 8429 27716 8453 27718
rect 8509 27716 8533 27718
rect 8589 27716 8613 27718
rect 8669 27716 8675 27718
rect 8367 27707 8675 27716
rect 8392 27464 8444 27470
rect 8392 27406 8444 27412
rect 8668 27464 8720 27470
rect 8668 27406 8720 27412
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 8116 26998 8168 27004
rect 8206 27024 8262 27033
rect 7932 26988 7984 26994
rect 8206 26959 8262 26968
rect 7932 26930 7984 26936
rect 7840 26920 7892 26926
rect 7840 26862 7892 26868
rect 8312 26738 8340 27270
rect 8404 27130 8432 27406
rect 8392 27124 8444 27130
rect 8392 27066 8444 27072
rect 8680 26772 8708 27406
rect 8760 27056 8812 27062
rect 8760 26998 8812 27004
rect 8680 26744 8733 26772
rect 8310 26710 8340 26738
rect 8310 26602 8338 26710
rect 8367 26684 8675 26693
rect 8367 26682 8373 26684
rect 8429 26682 8453 26684
rect 8509 26682 8533 26684
rect 8589 26682 8613 26684
rect 8669 26682 8675 26684
rect 8429 26630 8431 26682
rect 8611 26630 8613 26682
rect 8367 26628 8373 26630
rect 8429 26628 8453 26630
rect 8509 26628 8533 26630
rect 8589 26628 8613 26630
rect 8669 26628 8675 26630
rect 8367 26619 8675 26628
rect 8310 26574 8340 26602
rect 8114 26344 8170 26353
rect 7760 26302 7880 26330
rect 7852 26217 7880 26302
rect 8024 26308 8076 26314
rect 8114 26279 8116 26288
rect 8024 26250 8076 26256
rect 8168 26279 8170 26288
rect 8116 26250 8168 26256
rect 7838 26208 7894 26217
rect 7838 26143 7894 26152
rect 7840 26036 7892 26042
rect 7840 25978 7892 25984
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7760 24993 7788 25842
rect 7852 25430 7880 25978
rect 7932 25968 7984 25974
rect 7932 25910 7984 25916
rect 7840 25424 7892 25430
rect 7840 25366 7892 25372
rect 7838 25120 7894 25129
rect 7838 25055 7894 25064
rect 7746 24984 7802 24993
rect 7746 24919 7802 24928
rect 7654 24440 7710 24449
rect 7654 24375 7710 24384
rect 7852 24256 7880 25055
rect 7944 24954 7972 25910
rect 7932 24948 7984 24954
rect 7932 24890 7984 24896
rect 8036 24834 8064 26250
rect 8312 25974 8340 26574
rect 8705 26568 8733 26744
rect 8680 26540 8733 26568
rect 8680 26382 8708 26540
rect 8668 26376 8720 26382
rect 8574 26344 8630 26353
rect 8668 26318 8720 26324
rect 8574 26279 8630 26288
rect 8300 25968 8352 25974
rect 8300 25910 8352 25916
rect 8588 25786 8616 26279
rect 7760 24228 7880 24256
rect 7944 24806 8064 24834
rect 8128 25758 8616 25786
rect 7564 24064 7616 24070
rect 7564 24006 7616 24012
rect 7470 23760 7526 23769
rect 7576 23730 7604 24006
rect 7470 23695 7526 23704
rect 7564 23724 7616 23730
rect 7484 23662 7512 23695
rect 7564 23666 7616 23672
rect 7472 23656 7524 23662
rect 7472 23598 7524 23604
rect 7472 23180 7524 23186
rect 7392 23140 7472 23168
rect 7576 23168 7604 23666
rect 7656 23180 7708 23186
rect 7576 23140 7656 23168
rect 7472 23122 7524 23128
rect 7656 23122 7708 23128
rect 7300 23072 7420 23100
rect 7196 22568 7248 22574
rect 7196 22510 7248 22516
rect 7196 22432 7248 22438
rect 7196 22374 7248 22380
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 7208 17762 7236 22374
rect 7392 22094 7420 23072
rect 7484 22273 7512 23122
rect 7564 22772 7616 22778
rect 7564 22714 7616 22720
rect 7470 22264 7526 22273
rect 7470 22199 7526 22208
rect 7392 22066 7512 22094
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7380 21344 7432 21350
rect 7380 21286 7432 21292
rect 7300 20874 7328 21286
rect 7392 21146 7420 21286
rect 7380 21140 7432 21146
rect 7380 21082 7432 21088
rect 7288 20868 7340 20874
rect 7288 20810 7340 20816
rect 7484 20777 7512 22066
rect 7470 20768 7526 20777
rect 7470 20703 7526 20712
rect 7286 20632 7342 20641
rect 7286 20567 7342 20576
rect 7300 19514 7328 20567
rect 7380 20460 7432 20466
rect 7380 20402 7432 20408
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7392 20369 7420 20402
rect 7378 20360 7434 20369
rect 7378 20295 7434 20304
rect 7392 19961 7420 20295
rect 7484 20058 7512 20402
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7378 19952 7434 19961
rect 7378 19887 7434 19896
rect 7378 19816 7434 19825
rect 7378 19751 7434 19760
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7286 18864 7342 18873
rect 7286 18799 7342 18808
rect 7300 18766 7328 18799
rect 7392 18766 7420 19751
rect 7576 19174 7604 22714
rect 7654 22536 7710 22545
rect 7654 22471 7710 22480
rect 7668 21690 7696 22471
rect 7656 21684 7708 21690
rect 7656 21626 7708 21632
rect 7668 19378 7696 21626
rect 7760 21622 7788 24228
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7852 22574 7880 24074
rect 7944 23633 7972 24806
rect 8128 23712 8156 25758
rect 8208 25696 8260 25702
rect 8680 25684 8708 26318
rect 8680 25656 8733 25684
rect 8208 25638 8260 25644
rect 8220 25498 8248 25638
rect 8367 25596 8675 25605
rect 8367 25594 8373 25596
rect 8429 25594 8453 25596
rect 8509 25594 8533 25596
rect 8589 25594 8613 25596
rect 8669 25594 8675 25596
rect 8429 25542 8431 25594
rect 8611 25542 8613 25594
rect 8367 25540 8373 25542
rect 8429 25540 8453 25542
rect 8509 25540 8533 25542
rect 8589 25540 8613 25542
rect 8669 25540 8675 25542
rect 8367 25531 8675 25540
rect 8208 25492 8260 25498
rect 8705 25480 8733 25656
rect 8208 25434 8260 25440
rect 8588 25452 8733 25480
rect 8588 25294 8616 25452
rect 8772 25378 8800 26998
rect 8680 25350 8800 25378
rect 8576 25288 8628 25294
rect 8576 25230 8628 25236
rect 8208 25220 8260 25226
rect 8208 25162 8260 25168
rect 8220 24834 8248 25162
rect 8220 24818 8524 24834
rect 8220 24812 8536 24818
rect 8220 24806 8484 24812
rect 8220 24206 8248 24806
rect 8484 24754 8536 24760
rect 8680 24596 8708 25350
rect 8760 25220 8812 25226
rect 8760 25162 8812 25168
rect 8772 24993 8800 25162
rect 8758 24984 8814 24993
rect 8758 24919 8814 24928
rect 8680 24568 8800 24596
rect 8367 24508 8675 24517
rect 8367 24506 8373 24508
rect 8429 24506 8453 24508
rect 8509 24506 8533 24508
rect 8589 24506 8613 24508
rect 8669 24506 8675 24508
rect 8429 24454 8431 24506
rect 8611 24454 8613 24506
rect 8367 24452 8373 24454
rect 8429 24452 8453 24454
rect 8509 24452 8533 24454
rect 8589 24452 8613 24454
rect 8669 24452 8675 24454
rect 8367 24443 8675 24452
rect 8772 24410 8800 24568
rect 8760 24404 8812 24410
rect 8760 24346 8812 24352
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 8220 24041 8248 24142
rect 8206 24032 8262 24041
rect 8206 23967 8262 23976
rect 8312 23882 8340 24142
rect 8036 23684 8156 23712
rect 8220 23854 8340 23882
rect 7930 23624 7986 23633
rect 7930 23559 7986 23568
rect 7840 22568 7892 22574
rect 8036 22556 8064 23684
rect 8220 23610 8248 23854
rect 7840 22510 7892 22516
rect 7944 22528 8064 22556
rect 8128 23582 8248 23610
rect 7840 22228 7892 22234
rect 7840 22170 7892 22176
rect 7748 21616 7800 21622
rect 7748 21558 7800 21564
rect 7656 19372 7708 19378
rect 7656 19314 7708 19320
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7564 18964 7616 18970
rect 7564 18906 7616 18912
rect 7288 18760 7340 18766
rect 7288 18702 7340 18708
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7116 17734 7236 17762
rect 7116 17678 7144 17734
rect 7104 17672 7156 17678
rect 7104 17614 7156 17620
rect 7116 16833 7144 17614
rect 7196 17536 7248 17542
rect 7196 17478 7248 17484
rect 7102 16824 7158 16833
rect 7012 16788 7064 16794
rect 7102 16759 7158 16768
rect 7012 16730 7064 16736
rect 7104 16652 7156 16658
rect 7104 16594 7156 16600
rect 7012 16516 7064 16522
rect 7012 16458 7064 16464
rect 7024 15978 7052 16458
rect 7012 15972 7064 15978
rect 7012 15914 7064 15920
rect 7010 15736 7066 15745
rect 7010 15671 7066 15680
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6920 14408 6972 14414
rect 6920 14350 6972 14356
rect 6932 13433 6960 14350
rect 6918 13424 6974 13433
rect 6918 13359 6974 13368
rect 6920 13320 6972 13326
rect 7024 13308 7052 15671
rect 6972 13280 7052 13308
rect 6920 13262 6972 13268
rect 6828 12368 6880 12374
rect 6828 12310 6880 12316
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6840 11898 6868 12038
rect 6828 11892 6880 11898
rect 6828 11834 6880 11840
rect 6826 11792 6882 11801
rect 6826 11727 6882 11736
rect 6840 11626 6868 11727
rect 6932 11626 6960 13262
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 7024 13025 7052 13126
rect 7010 13016 7066 13025
rect 7010 12951 7066 12960
rect 7116 12102 7144 16594
rect 7208 16046 7236 17478
rect 7300 17218 7328 18702
rect 7470 18320 7526 18329
rect 7470 18255 7472 18264
rect 7524 18255 7526 18264
rect 7472 18226 7524 18232
rect 7472 17876 7524 17882
rect 7472 17818 7524 17824
rect 7390 17672 7442 17678
rect 7390 17614 7442 17620
rect 7392 17338 7420 17614
rect 7380 17332 7432 17338
rect 7380 17274 7432 17280
rect 7300 17190 7420 17218
rect 7288 16992 7340 16998
rect 7288 16934 7340 16940
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7208 14414 7236 15982
rect 7300 15026 7328 16934
rect 7392 16658 7420 17190
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7300 14521 7328 14962
rect 7392 14958 7420 16186
rect 7484 16114 7512 17818
rect 7576 17134 7604 18906
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7668 18086 7696 18566
rect 7656 18080 7708 18086
rect 7656 18022 7708 18028
rect 7564 17128 7616 17134
rect 7564 17070 7616 17076
rect 7576 16522 7604 17070
rect 7564 16516 7616 16522
rect 7564 16458 7616 16464
rect 7668 16250 7696 18022
rect 7760 16590 7788 21558
rect 7852 20466 7880 22170
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7944 19334 7972 22528
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 8036 22137 8064 22374
rect 8022 22128 8078 22137
rect 8022 22063 8078 22072
rect 8128 22001 8156 23582
rect 8208 23520 8260 23526
rect 8208 23462 8260 23468
rect 8220 23322 8248 23462
rect 8367 23420 8675 23429
rect 8367 23418 8373 23420
rect 8429 23418 8453 23420
rect 8509 23418 8533 23420
rect 8589 23418 8613 23420
rect 8669 23418 8675 23420
rect 8429 23366 8431 23418
rect 8611 23366 8613 23418
rect 8367 23364 8373 23366
rect 8429 23364 8453 23366
rect 8509 23364 8533 23366
rect 8589 23364 8613 23366
rect 8669 23364 8675 23366
rect 8367 23355 8675 23364
rect 8208 23316 8260 23322
rect 8208 23258 8260 23264
rect 8668 23248 8720 23254
rect 8668 23190 8720 23196
rect 8208 23180 8260 23186
rect 8208 23122 8260 23128
rect 8114 21992 8170 22001
rect 8114 21927 8170 21936
rect 8220 21622 8248 23122
rect 8680 22420 8708 23190
rect 8760 22976 8812 22982
rect 8760 22918 8812 22924
rect 8680 22392 8733 22420
rect 8367 22332 8675 22341
rect 8367 22330 8373 22332
rect 8429 22330 8453 22332
rect 8509 22330 8533 22332
rect 8589 22330 8613 22332
rect 8669 22330 8675 22332
rect 8429 22278 8431 22330
rect 8611 22278 8613 22330
rect 8367 22276 8373 22278
rect 8429 22276 8453 22278
rect 8509 22276 8533 22278
rect 8589 22276 8613 22278
rect 8669 22276 8675 22278
rect 8367 22267 8675 22276
rect 8705 22216 8733 22392
rect 8496 22188 8733 22216
rect 8208 21616 8260 21622
rect 8128 21576 8208 21604
rect 8024 20800 8076 20806
rect 8024 20742 8076 20748
rect 7852 19306 7972 19334
rect 7852 18873 7880 19306
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 7838 18864 7894 18873
rect 7838 18799 7894 18808
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7852 17513 7880 18362
rect 7838 17504 7894 17513
rect 7838 17439 7894 17448
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7656 16244 7708 16250
rect 7656 16186 7708 16192
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7656 16108 7708 16114
rect 7656 16050 7708 16056
rect 7668 15722 7696 16050
rect 7576 15706 7696 15722
rect 7564 15700 7696 15706
rect 7616 15694 7696 15700
rect 7564 15642 7616 15648
rect 7470 15600 7526 15609
rect 7470 15535 7526 15544
rect 7484 15502 7512 15535
rect 7760 15502 7788 16526
rect 7838 16416 7894 16425
rect 7838 16351 7894 16360
rect 7472 15496 7524 15502
rect 7472 15438 7524 15444
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7380 14952 7432 14958
rect 7380 14894 7432 14900
rect 7286 14512 7342 14521
rect 7286 14447 7342 14456
rect 7196 14408 7248 14414
rect 7196 14350 7248 14356
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7208 13920 7236 14350
rect 7300 14113 7328 14350
rect 7286 14104 7342 14113
rect 7286 14039 7342 14048
rect 7392 13938 7420 14894
rect 7484 14414 7512 15438
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7288 13932 7340 13938
rect 7208 13892 7288 13920
rect 7288 13874 7340 13880
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7194 13832 7250 13841
rect 7194 13767 7250 13776
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11892 7064 11898
rect 7012 11834 7064 11840
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6840 10690 6868 11562
rect 6932 11286 6960 11562
rect 7024 11393 7052 11834
rect 7104 11620 7156 11626
rect 7104 11562 7156 11568
rect 7010 11384 7066 11393
rect 7010 11319 7066 11328
rect 6920 11280 6972 11286
rect 6920 11222 6972 11228
rect 7116 11064 7144 11562
rect 6932 11036 7144 11064
rect 6932 10810 6960 11036
rect 7102 10976 7158 10985
rect 7024 10934 7102 10962
rect 7024 10810 7052 10934
rect 7102 10911 7158 10920
rect 7208 10860 7236 13767
rect 7286 13696 7342 13705
rect 7286 13631 7342 13640
rect 7116 10832 7236 10860
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6840 10662 6960 10690
rect 6656 10390 6776 10418
rect 6826 10432 6882 10441
rect 6552 9716 6604 9722
rect 6552 9658 6604 9664
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6564 9178 6592 9522
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6552 9036 6604 9042
rect 6552 8978 6604 8984
rect 6564 8673 6592 8978
rect 6550 8664 6606 8673
rect 6550 8599 6606 8608
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6458 7848 6514 7857
rect 6458 7783 6514 7792
rect 6458 7576 6514 7585
rect 6458 7511 6514 7520
rect 6472 7410 6500 7511
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6380 7262 6500 7290
rect 6368 7200 6420 7206
rect 6368 7142 6420 7148
rect 6380 6934 6408 7142
rect 6368 6928 6420 6934
rect 6368 6870 6420 6876
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 6092 6316 6144 6322
rect 6092 6258 6144 6264
rect 5828 5778 5856 6258
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5920 5534 5948 6054
rect 5828 5506 5948 5534
rect 6104 5534 6132 6258
rect 6380 6225 6408 6734
rect 6472 6730 6500 7262
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6472 6497 6500 6666
rect 6458 6488 6514 6497
rect 6458 6423 6514 6432
rect 6564 6225 6592 8026
rect 6366 6216 6422 6225
rect 6366 6151 6422 6160
rect 6550 6216 6606 6225
rect 6550 6151 6606 6160
rect 6368 6112 6420 6118
rect 6420 6072 6592 6100
rect 6368 6054 6420 6060
rect 6458 5944 6514 5953
rect 6458 5879 6514 5888
rect 6368 5636 6420 5642
rect 6368 5578 6420 5584
rect 6104 5506 6316 5534
rect 5828 4214 5856 5506
rect 5894 5468 6202 5477
rect 5894 5466 5900 5468
rect 5956 5466 5980 5468
rect 6036 5466 6060 5468
rect 6116 5466 6140 5468
rect 6196 5466 6202 5468
rect 5956 5414 5958 5466
rect 6138 5414 6140 5466
rect 5894 5412 5900 5414
rect 5956 5412 5980 5414
rect 6036 5412 6060 5414
rect 6116 5412 6140 5414
rect 6196 5412 6202 5414
rect 5894 5403 6202 5412
rect 6288 5370 6316 5506
rect 6276 5364 6328 5370
rect 6276 5306 6328 5312
rect 6380 5250 6408 5578
rect 6288 5222 6408 5250
rect 5894 4380 6202 4389
rect 5894 4378 5900 4380
rect 5956 4378 5980 4380
rect 6036 4378 6060 4380
rect 6116 4378 6140 4380
rect 6196 4378 6202 4380
rect 5956 4326 5958 4378
rect 6138 4326 6140 4378
rect 5894 4324 5900 4326
rect 5956 4324 5980 4326
rect 6036 4324 6060 4326
rect 6116 4324 6140 4326
rect 6196 4324 6202 4326
rect 5894 4315 6202 4324
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5368 2400 5488 2428
rect 5632 2440 5684 2446
rect 4896 1488 4948 1494
rect 5264 1488 5316 1494
rect 4948 1436 5028 1442
rect 4896 1430 5028 1436
rect 5264 1430 5316 1436
rect 4908 1414 5028 1430
rect 4896 1284 4948 1290
rect 4896 1226 4948 1232
rect 4908 660 4936 1226
rect 4816 632 4936 660
rect 4816 160 4844 632
rect 5000 160 5028 1414
rect 5172 1420 5224 1426
rect 5172 1362 5224 1368
rect 5080 1216 5132 1222
rect 5080 1158 5132 1164
rect 4250 54 4384 82
rect 4250 -300 4306 54
rect 4434 -300 4490 160
rect 4618 -300 4674 160
rect 4802 -300 4858 160
rect 4986 -300 5042 160
rect 5092 66 5120 1158
rect 5184 160 5212 1362
rect 5368 1358 5396 2400
rect 5632 2382 5684 2388
rect 5540 2372 5592 2378
rect 5460 2332 5540 2360
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 5264 1284 5316 1290
rect 5264 1226 5316 1232
rect 5276 678 5304 1226
rect 5354 1184 5410 1193
rect 5354 1119 5410 1128
rect 5368 1018 5396 1119
rect 5356 1012 5408 1018
rect 5356 954 5408 960
rect 5264 672 5316 678
rect 5264 614 5316 620
rect 5080 60 5132 66
rect 5080 2 5132 8
rect 5170 -300 5226 160
rect 5354 82 5410 160
rect 5460 82 5488 2332
rect 5540 2314 5592 2320
rect 5540 1964 5592 1970
rect 5540 1906 5592 1912
rect 5552 1329 5580 1906
rect 5538 1320 5594 1329
rect 5538 1255 5594 1264
rect 5644 1204 5672 2382
rect 5552 1176 5672 1204
rect 5552 160 5580 1176
rect 5736 160 5764 2994
rect 5828 2990 5856 4014
rect 6288 3398 6316 5222
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4826 6408 5102
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6276 3392 6328 3398
rect 6276 3334 6328 3340
rect 5894 3292 6202 3301
rect 5894 3290 5900 3292
rect 5956 3290 5980 3292
rect 6036 3290 6060 3292
rect 6116 3290 6140 3292
rect 6196 3290 6202 3292
rect 5956 3238 5958 3290
rect 6138 3238 6140 3290
rect 5894 3236 5900 3238
rect 5956 3236 5980 3238
rect 6036 3236 6060 3238
rect 6116 3236 6140 3238
rect 6196 3236 6202 3238
rect 5894 3227 6202 3236
rect 6274 3224 6330 3233
rect 6274 3159 6330 3168
rect 6182 3088 6238 3097
rect 6182 3023 6238 3032
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 6196 2310 6224 3023
rect 6288 2582 6316 3159
rect 6276 2576 6328 2582
rect 6276 2518 6328 2524
rect 6380 2530 6408 3674
rect 6472 2650 6500 5879
rect 6564 3641 6592 6072
rect 6550 3632 6606 3641
rect 6550 3567 6606 3576
rect 6656 3058 6684 10390
rect 6826 10367 6882 10376
rect 6840 10266 6868 10367
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6748 9586 6776 9862
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 5545 6776 9318
rect 6840 6866 6868 9658
rect 6932 9625 6960 10662
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6918 9616 6974 9625
rect 6918 9551 6974 9560
rect 6920 9104 6972 9110
rect 6918 9072 6920 9081
rect 6972 9072 6974 9081
rect 6918 9007 6974 9016
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 7313 6960 8774
rect 7024 7886 7052 9998
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 7024 7546 7052 7686
rect 7012 7540 7064 7546
rect 7012 7482 7064 7488
rect 7116 7410 7144 10832
rect 7194 10432 7250 10441
rect 7194 10367 7250 10376
rect 7208 10266 7236 10367
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7300 10198 7328 13631
rect 7378 13560 7434 13569
rect 7378 13495 7434 13504
rect 7392 12646 7420 13495
rect 7484 12850 7512 14214
rect 7576 12986 7604 15302
rect 7746 15056 7802 15065
rect 7746 14991 7802 15000
rect 7654 14920 7710 14929
rect 7654 14855 7710 14864
rect 7564 12980 7616 12986
rect 7564 12922 7616 12928
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7380 12640 7432 12646
rect 7380 12582 7432 12588
rect 7392 12306 7420 12582
rect 7562 12336 7618 12345
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7484 12294 7562 12322
rect 7380 12096 7432 12102
rect 7380 12038 7432 12044
rect 7392 11762 7420 12038
rect 7380 11756 7432 11762
rect 7380 11698 7432 11704
rect 7484 11286 7512 12294
rect 7562 12271 7618 12280
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7380 11280 7432 11286
rect 7380 11222 7432 11228
rect 7472 11280 7524 11286
rect 7472 11222 7524 11228
rect 7288 10192 7340 10198
rect 7288 10134 7340 10140
rect 7196 9988 7248 9994
rect 7196 9930 7248 9936
rect 7208 9761 7236 9930
rect 7194 9752 7250 9761
rect 7194 9687 7250 9696
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7300 9489 7328 9590
rect 7286 9480 7342 9489
rect 7286 9415 7342 9424
rect 7214 8968 7266 8974
rect 7392 8956 7420 11222
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7484 10674 7512 11086
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 9558 7512 10406
rect 7576 9926 7604 11630
rect 7668 10985 7696 14855
rect 7760 14414 7788 14991
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 7746 14240 7802 14249
rect 7746 14175 7802 14184
rect 7760 11778 7788 14175
rect 7852 13326 7880 16351
rect 7944 15366 7972 19110
rect 8036 18442 8064 20742
rect 8128 19242 8156 21576
rect 8208 21558 8260 21564
rect 8208 21480 8260 21486
rect 8208 21422 8260 21428
rect 8220 21146 8248 21422
rect 8496 21332 8524 22188
rect 8772 22030 8800 22918
rect 8864 22778 8892 30806
rect 8956 29714 8984 31719
rect 8944 29708 8996 29714
rect 8944 29650 8996 29656
rect 8956 28014 8984 29650
rect 9048 28064 9076 32807
rect 9140 30326 9168 34598
rect 9128 30320 9180 30326
rect 9128 30262 9180 30268
rect 9126 30152 9182 30161
rect 9126 30087 9182 30096
rect 9140 28234 9168 30087
rect 9232 29306 9260 37606
rect 9324 35476 9352 38626
rect 9508 37670 9536 41386
rect 9876 39681 9904 43046
rect 9956 42764 10008 42770
rect 9956 42706 10008 42712
rect 9968 42129 9996 42706
rect 10060 42226 10088 43404
rect 10152 42906 10180 43590
rect 10244 43574 10364 43602
rect 10244 43489 10272 43574
rect 10230 43480 10286 43489
rect 10230 43415 10286 43424
rect 10416 43376 10468 43382
rect 10244 43336 10416 43364
rect 10140 42900 10192 42906
rect 10140 42842 10192 42848
rect 10140 42696 10192 42702
rect 10138 42664 10140 42673
rect 10192 42664 10194 42673
rect 10138 42599 10194 42608
rect 10140 42560 10192 42566
rect 10140 42502 10192 42508
rect 10048 42220 10100 42226
rect 10048 42162 10100 42168
rect 9954 42120 10010 42129
rect 9954 42055 10010 42064
rect 9956 41540 10008 41546
rect 9956 41482 10008 41488
rect 9862 39672 9918 39681
rect 9862 39607 9918 39616
rect 9588 39364 9640 39370
rect 9588 39306 9640 39312
rect 9600 37738 9628 39306
rect 9680 38480 9732 38486
rect 9968 38434 9996 41482
rect 9680 38422 9732 38428
rect 9692 38185 9720 38422
rect 9876 38406 9996 38434
rect 9772 38344 9824 38350
rect 9772 38286 9824 38292
rect 9678 38176 9734 38185
rect 9678 38111 9734 38120
rect 9680 38004 9732 38010
rect 9680 37946 9732 37952
rect 9588 37732 9640 37738
rect 9588 37674 9640 37680
rect 9496 37664 9548 37670
rect 9496 37606 9548 37612
rect 9692 37398 9720 37946
rect 9680 37392 9732 37398
rect 9680 37334 9732 37340
rect 9402 37224 9458 37233
rect 9402 37159 9404 37168
rect 9456 37159 9458 37168
rect 9404 37130 9456 37136
rect 9680 36780 9732 36786
rect 9680 36722 9732 36728
rect 9692 36666 9720 36722
rect 9784 36718 9812 38286
rect 9508 36638 9720 36666
rect 9772 36712 9824 36718
rect 9772 36654 9824 36660
rect 9402 36272 9458 36281
rect 9402 36207 9458 36216
rect 9416 36174 9444 36207
rect 9404 36168 9456 36174
rect 9404 36110 9456 36116
rect 9508 35737 9536 36638
rect 9588 36576 9640 36582
rect 9588 36518 9640 36524
rect 9494 35728 9550 35737
rect 9494 35663 9550 35672
rect 9600 35630 9628 36518
rect 9770 35864 9826 35873
rect 9770 35799 9826 35808
rect 9784 35766 9812 35799
rect 9876 35766 9904 38406
rect 9956 38276 10008 38282
rect 9956 38218 10008 38224
rect 9968 38010 9996 38218
rect 9956 38004 10008 38010
rect 9956 37946 10008 37952
rect 10046 37904 10102 37913
rect 10046 37839 10048 37848
rect 10100 37839 10102 37848
rect 10048 37810 10100 37816
rect 9956 37256 10008 37262
rect 9956 37198 10008 37204
rect 9968 36122 9996 37198
rect 10060 36786 10088 37810
rect 10048 36780 10100 36786
rect 10048 36722 10100 36728
rect 9968 36094 10088 36122
rect 9956 36032 10008 36038
rect 9956 35974 10008 35980
rect 9772 35760 9824 35766
rect 9772 35702 9824 35708
rect 9864 35760 9916 35766
rect 9864 35702 9916 35708
rect 9588 35624 9640 35630
rect 9588 35566 9640 35572
rect 9324 35448 9720 35476
rect 9324 35278 9628 35306
rect 9324 35222 9352 35278
rect 9312 35216 9364 35222
rect 9312 35158 9364 35164
rect 9496 35216 9548 35222
rect 9496 35158 9548 35164
rect 9312 34400 9364 34406
rect 9312 34342 9364 34348
rect 9324 34202 9352 34342
rect 9312 34196 9364 34202
rect 9312 34138 9364 34144
rect 9404 33992 9456 33998
rect 9310 33960 9366 33969
rect 9366 33940 9404 33946
rect 9366 33934 9456 33940
rect 9366 33918 9444 33934
rect 9310 33895 9366 33904
rect 9508 33862 9536 35158
rect 9496 33856 9548 33862
rect 9496 33798 9548 33804
rect 9496 33312 9548 33318
rect 9496 33254 9548 33260
rect 9312 33108 9364 33114
rect 9312 33050 9364 33056
rect 9324 32570 9352 33050
rect 9312 32564 9364 32570
rect 9312 32506 9364 32512
rect 9404 32496 9456 32502
rect 9404 32438 9456 32444
rect 9416 31929 9444 32438
rect 9508 32314 9536 33254
rect 9600 33017 9628 35278
rect 9692 33946 9720 35448
rect 9968 35329 9996 35974
rect 9954 35320 10010 35329
rect 9954 35255 10010 35264
rect 9954 35048 10010 35057
rect 9876 35006 9954 35034
rect 9772 34944 9824 34950
rect 9772 34886 9824 34892
rect 9784 34066 9812 34886
rect 9876 34610 9904 35006
rect 9954 34983 10010 34992
rect 9956 34944 10008 34950
rect 9956 34886 10008 34892
rect 9968 34746 9996 34886
rect 9956 34740 10008 34746
rect 9956 34682 10008 34688
rect 9864 34604 9916 34610
rect 9864 34546 9916 34552
rect 9956 34536 10008 34542
rect 9956 34478 10008 34484
rect 9968 34202 9996 34478
rect 9956 34196 10008 34202
rect 9956 34138 10008 34144
rect 9772 34060 9824 34066
rect 9772 34002 9824 34008
rect 9692 33918 9812 33946
rect 9586 33008 9642 33017
rect 9586 32943 9642 32952
rect 9680 32428 9732 32434
rect 9680 32370 9732 32376
rect 9508 32286 9628 32314
rect 9496 32224 9548 32230
rect 9496 32166 9548 32172
rect 9402 31920 9458 31929
rect 9312 31884 9364 31890
rect 9402 31855 9458 31864
rect 9312 31826 9364 31832
rect 9324 30802 9352 31826
rect 9404 31748 9456 31754
rect 9404 31690 9456 31696
rect 9416 31657 9444 31690
rect 9402 31648 9458 31657
rect 9402 31583 9458 31592
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9416 30938 9444 31214
rect 9404 30932 9456 30938
rect 9404 30874 9456 30880
rect 9312 30796 9364 30802
rect 9312 30738 9364 30744
rect 9312 29640 9364 29646
rect 9312 29582 9364 29588
rect 9220 29300 9272 29306
rect 9220 29242 9272 29248
rect 9140 28206 9260 28234
rect 9128 28076 9180 28082
rect 9048 28036 9128 28064
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 8956 24886 8984 27950
rect 9048 25537 9076 28036
rect 9128 28018 9180 28024
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9140 27033 9168 27406
rect 9126 27024 9182 27033
rect 9126 26959 9182 26968
rect 9128 26580 9180 26586
rect 9128 26522 9180 26528
rect 9034 25528 9090 25537
rect 9034 25463 9036 25472
rect 9088 25463 9090 25472
rect 9036 25434 9088 25440
rect 9036 25152 9088 25158
rect 9036 25094 9088 25100
rect 8944 24880 8996 24886
rect 8944 24822 8996 24828
rect 8956 24410 8984 24822
rect 8944 24404 8996 24410
rect 8944 24346 8996 24352
rect 8852 22772 8904 22778
rect 8852 22714 8904 22720
rect 8852 22432 8904 22438
rect 8852 22374 8904 22380
rect 8760 22024 8812 22030
rect 8760 21966 8812 21972
rect 8864 21876 8892 22374
rect 8312 21304 8524 21332
rect 8772 21848 8892 21876
rect 8312 21298 8340 21304
rect 8310 21270 8340 21298
rect 8310 21162 8338 21270
rect 8367 21244 8675 21253
rect 8367 21242 8373 21244
rect 8429 21242 8453 21244
rect 8509 21242 8533 21244
rect 8589 21242 8613 21244
rect 8669 21242 8675 21244
rect 8429 21190 8431 21242
rect 8611 21190 8613 21242
rect 8367 21188 8373 21190
rect 8429 21188 8453 21190
rect 8509 21188 8533 21190
rect 8589 21188 8613 21190
rect 8669 21188 8675 21190
rect 8367 21179 8675 21188
rect 8208 21140 8260 21146
rect 8310 21134 8340 21162
rect 8208 21082 8260 21088
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8220 20398 8248 20742
rect 8312 20602 8340 21134
rect 8668 20936 8720 20942
rect 8666 20904 8668 20913
rect 8720 20904 8722 20913
rect 8772 20874 8800 21848
rect 8852 21548 8904 21554
rect 8852 21490 8904 21496
rect 8666 20839 8722 20848
rect 8760 20868 8812 20874
rect 8760 20810 8812 20816
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8760 20460 8812 20466
rect 8760 20402 8812 20408
rect 8208 20392 8260 20398
rect 8208 20334 8260 20340
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8668 20256 8720 20262
rect 8720 20204 8733 20244
rect 8668 20198 8733 20204
rect 8220 20074 8248 20198
rect 8367 20156 8675 20165
rect 8367 20154 8373 20156
rect 8429 20154 8453 20156
rect 8509 20154 8533 20156
rect 8589 20154 8613 20156
rect 8669 20154 8675 20156
rect 8429 20102 8431 20154
rect 8611 20102 8613 20154
rect 8367 20100 8373 20102
rect 8429 20100 8453 20102
rect 8509 20100 8533 20102
rect 8589 20100 8613 20102
rect 8669 20100 8675 20102
rect 8367 20091 8675 20100
rect 8220 20046 8340 20074
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8220 18630 8248 19790
rect 8312 19310 8340 20046
rect 8705 20040 8733 20198
rect 8680 20012 8733 20040
rect 8576 19984 8628 19990
rect 8576 19926 8628 19932
rect 8588 19378 8616 19926
rect 8680 19922 8708 20012
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8668 19372 8720 19378
rect 8772 19360 8800 20402
rect 8864 20380 8892 21490
rect 8956 20534 8984 24346
rect 9048 23322 9076 25094
rect 9036 23316 9088 23322
rect 9036 23258 9088 23264
rect 9034 23080 9090 23089
rect 9034 23015 9036 23024
rect 9088 23015 9090 23024
rect 9036 22986 9088 22992
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 9048 22681 9076 22714
rect 9034 22672 9090 22681
rect 9034 22607 9090 22616
rect 9034 22536 9090 22545
rect 9034 22471 9090 22480
rect 9048 21729 9076 22471
rect 9034 21720 9090 21729
rect 9034 21655 9090 21664
rect 9036 21616 9088 21622
rect 9036 21558 9088 21564
rect 9048 21146 9076 21558
rect 9036 21140 9088 21146
rect 9036 21082 9088 21088
rect 9036 20868 9088 20874
rect 9036 20810 9088 20816
rect 8944 20528 8996 20534
rect 8944 20470 8996 20476
rect 8864 20352 8984 20380
rect 8852 20256 8904 20262
rect 8852 20198 8904 20204
rect 8864 19990 8892 20198
rect 8852 19984 8904 19990
rect 8852 19926 8904 19932
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8864 19378 8892 19654
rect 8956 19514 8984 20352
rect 8944 19508 8996 19514
rect 8944 19450 8996 19456
rect 8942 19408 8998 19417
rect 8720 19332 8800 19360
rect 8668 19314 8720 19320
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8367 19068 8675 19077
rect 8367 19066 8373 19068
rect 8429 19066 8453 19068
rect 8509 19066 8533 19068
rect 8589 19066 8613 19068
rect 8669 19066 8675 19068
rect 8429 19014 8431 19066
rect 8611 19014 8613 19066
rect 8367 19012 8373 19014
rect 8429 19012 8453 19014
rect 8509 19012 8533 19014
rect 8589 19012 8613 19014
rect 8669 19012 8675 19014
rect 8367 19003 8675 19012
rect 8300 18964 8352 18970
rect 8300 18906 8352 18912
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8036 18414 8248 18442
rect 8024 17536 8076 17542
rect 8024 17478 8076 17484
rect 8036 17338 8064 17478
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 8116 16244 8168 16250
rect 8036 16204 8116 16232
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 8036 14929 8064 16204
rect 8116 16186 8168 16192
rect 8114 16144 8170 16153
rect 8114 16079 8170 16088
rect 8022 14920 8078 14929
rect 8022 14855 8078 14864
rect 7930 14512 7986 14521
rect 7986 14470 8064 14498
rect 7930 14447 7986 14456
rect 7930 13832 7986 13841
rect 7930 13767 7986 13776
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7852 12986 7880 13126
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7760 11750 7880 11778
rect 7748 11688 7800 11694
rect 7748 11630 7800 11636
rect 7654 10976 7710 10985
rect 7654 10911 7710 10920
rect 7654 10840 7710 10849
rect 7654 10775 7710 10784
rect 7668 10033 7696 10775
rect 7654 10024 7710 10033
rect 7654 9959 7710 9968
rect 7564 9920 7616 9926
rect 7564 9862 7616 9868
rect 7654 9752 7710 9761
rect 7760 9722 7788 11630
rect 7654 9687 7710 9696
rect 7748 9716 7800 9722
rect 7484 9530 7604 9558
rect 7470 9480 7526 9489
rect 7470 9415 7526 9424
rect 7266 8928 7420 8956
rect 7214 8910 7266 8916
rect 7392 8838 7420 8928
rect 7380 8832 7432 8838
rect 7194 8800 7250 8809
rect 7380 8774 7432 8780
rect 7194 8735 7250 8744
rect 7104 7404 7156 7410
rect 7104 7346 7156 7352
rect 6918 7304 6974 7313
rect 6918 7239 6974 7248
rect 7104 7268 7156 7274
rect 6932 7002 6960 7239
rect 7104 7210 7156 7216
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 5914 6868 6598
rect 6932 5914 6960 6802
rect 7116 6633 7144 7210
rect 7102 6624 7158 6633
rect 7102 6559 7158 6568
rect 7010 6216 7066 6225
rect 7116 6186 7144 6559
rect 7010 6151 7066 6160
rect 7104 6180 7156 6186
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6918 5808 6974 5817
rect 6840 5766 6918 5794
rect 6734 5536 6790 5545
rect 6734 5471 6790 5480
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6748 4690 6776 5306
rect 6840 5234 6868 5766
rect 6918 5743 6974 5752
rect 7024 5370 7052 6151
rect 7104 6122 7156 6128
rect 7208 5846 7236 8735
rect 7484 8242 7512 9415
rect 7576 8809 7604 9530
rect 7562 8800 7618 8809
rect 7562 8735 7618 8744
rect 7562 8528 7618 8537
rect 7562 8463 7618 8472
rect 7300 8214 7512 8242
rect 7300 6882 7328 8214
rect 7470 8120 7526 8129
rect 7470 8055 7526 8064
rect 7484 7857 7512 8055
rect 7470 7848 7526 7857
rect 7470 7783 7526 7792
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7484 6914 7512 7686
rect 7576 7177 7604 8463
rect 7668 7868 7696 9687
rect 7748 9658 7800 9664
rect 7748 9580 7800 9586
rect 7748 9522 7800 9528
rect 7760 8566 7788 9522
rect 7852 9382 7880 11750
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7838 9072 7894 9081
rect 7838 9007 7894 9016
rect 7852 8566 7880 9007
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7748 8288 7800 8294
rect 7748 8230 7800 8236
rect 7760 8129 7788 8230
rect 7746 8120 7802 8129
rect 7746 8055 7802 8064
rect 7748 7880 7800 7886
rect 7668 7840 7748 7868
rect 7748 7822 7800 7828
rect 7944 7818 7972 13767
rect 8036 11665 8064 14470
rect 8128 12850 8156 16079
rect 8220 13841 8248 18414
rect 8312 18290 8340 18906
rect 8300 18284 8352 18290
rect 8300 18226 8352 18232
rect 8367 17980 8675 17989
rect 8367 17978 8373 17980
rect 8429 17978 8453 17980
rect 8509 17978 8533 17980
rect 8589 17978 8613 17980
rect 8669 17978 8675 17980
rect 8429 17926 8431 17978
rect 8611 17926 8613 17978
rect 8367 17924 8373 17926
rect 8429 17924 8453 17926
rect 8509 17924 8533 17926
rect 8589 17924 8613 17926
rect 8669 17924 8675 17926
rect 8367 17915 8675 17924
rect 8772 16998 8800 19332
rect 8852 19372 8904 19378
rect 8942 19343 8998 19352
rect 8852 19314 8904 19320
rect 8852 17740 8904 17746
rect 8852 17682 8904 17688
rect 8864 17338 8892 17682
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8760 16992 8812 16998
rect 8760 16934 8812 16940
rect 8367 16892 8675 16901
rect 8367 16890 8373 16892
rect 8429 16890 8453 16892
rect 8509 16890 8533 16892
rect 8589 16890 8613 16892
rect 8669 16890 8675 16892
rect 8429 16838 8431 16890
rect 8611 16838 8613 16890
rect 8367 16836 8373 16838
rect 8429 16836 8453 16838
rect 8509 16836 8533 16838
rect 8589 16836 8613 16838
rect 8669 16836 8675 16838
rect 8367 16827 8675 16836
rect 8956 16640 8984 19343
rect 8864 16612 8984 16640
rect 8758 16144 8814 16153
rect 8758 16079 8814 16088
rect 8772 15910 8800 16079
rect 8760 15904 8812 15910
rect 8760 15846 8812 15852
rect 8367 15804 8675 15813
rect 8367 15802 8373 15804
rect 8429 15802 8453 15804
rect 8509 15802 8533 15804
rect 8589 15802 8613 15804
rect 8669 15802 8675 15804
rect 8429 15750 8431 15802
rect 8611 15750 8613 15802
rect 8367 15748 8373 15750
rect 8429 15748 8453 15750
rect 8509 15748 8533 15750
rect 8589 15748 8613 15750
rect 8669 15748 8675 15750
rect 8367 15739 8675 15748
rect 8668 15428 8720 15434
rect 8668 15370 8720 15376
rect 8680 15337 8708 15370
rect 8666 15328 8722 15337
rect 8666 15263 8722 15272
rect 8300 15020 8352 15026
rect 8300 14962 8352 14968
rect 8312 14770 8340 14962
rect 8574 14920 8630 14929
rect 8574 14855 8576 14864
rect 8628 14855 8630 14864
rect 8576 14826 8628 14832
rect 8310 14742 8340 14770
rect 8310 14634 8338 14742
rect 8367 14716 8675 14725
rect 8367 14714 8373 14716
rect 8429 14714 8453 14716
rect 8509 14714 8533 14716
rect 8589 14714 8613 14716
rect 8669 14714 8675 14716
rect 8429 14662 8431 14714
rect 8611 14662 8613 14714
rect 8367 14660 8373 14662
rect 8429 14660 8453 14662
rect 8509 14660 8533 14662
rect 8589 14660 8613 14662
rect 8669 14660 8675 14662
rect 8367 14651 8675 14660
rect 8310 14606 8340 14634
rect 8206 13832 8262 13841
rect 8206 13767 8262 13776
rect 8208 13728 8260 13734
rect 8312 13682 8340 14606
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8680 13802 8708 14350
rect 8772 14249 8800 15846
rect 8864 15194 8892 16612
rect 8944 16516 8996 16522
rect 8944 16458 8996 16464
rect 8956 15570 8984 16458
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 8864 15166 8984 15194
rect 8758 14240 8814 14249
rect 8758 14175 8814 14184
rect 8852 14068 8904 14074
rect 8772 14028 8852 14056
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8208 13670 8260 13676
rect 8220 13530 8248 13670
rect 8310 13654 8340 13682
rect 8310 13546 8338 13654
rect 8367 13628 8675 13637
rect 8367 13626 8373 13628
rect 8429 13626 8453 13628
rect 8509 13626 8533 13628
rect 8589 13626 8613 13628
rect 8669 13626 8675 13628
rect 8429 13574 8431 13626
rect 8611 13574 8613 13626
rect 8367 13572 8373 13574
rect 8429 13572 8453 13574
rect 8509 13572 8533 13574
rect 8589 13572 8613 13574
rect 8669 13572 8675 13574
rect 8367 13563 8675 13572
rect 8208 13524 8260 13530
rect 8310 13518 8340 13546
rect 8312 13512 8340 13518
rect 8312 13484 8432 13512
rect 8208 13466 8260 13472
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8298 13152 8354 13161
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8022 11656 8078 11665
rect 8022 11591 8078 11600
rect 8036 11014 8064 11591
rect 8128 11150 8156 12786
rect 8220 12442 8248 13126
rect 8298 13087 8354 13096
rect 8312 12986 8340 13087
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8404 12866 8432 13484
rect 8666 13424 8722 13433
rect 8666 13359 8722 13368
rect 8680 12986 8708 13359
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8312 12838 8432 12866
rect 8312 12594 8340 12838
rect 8668 12776 8720 12782
rect 8666 12744 8668 12753
rect 8720 12744 8722 12753
rect 8666 12679 8722 12688
rect 8310 12566 8340 12594
rect 8310 12458 8338 12566
rect 8367 12540 8675 12549
rect 8367 12538 8373 12540
rect 8429 12538 8453 12540
rect 8509 12538 8533 12540
rect 8589 12538 8613 12540
rect 8669 12538 8675 12540
rect 8429 12486 8431 12538
rect 8611 12486 8613 12538
rect 8367 12484 8373 12486
rect 8429 12484 8453 12486
rect 8509 12484 8533 12486
rect 8589 12484 8613 12486
rect 8669 12484 8675 12486
rect 8367 12475 8675 12484
rect 8208 12436 8260 12442
rect 8310 12430 8340 12458
rect 8208 12378 8260 12384
rect 8208 12300 8260 12306
rect 8208 12242 8260 12248
rect 8116 11144 8168 11150
rect 8116 11086 8168 11092
rect 8024 11008 8076 11014
rect 8024 10950 8076 10956
rect 8116 10736 8168 10742
rect 8022 10704 8078 10713
rect 8116 10678 8168 10684
rect 8022 10639 8078 10648
rect 8036 10606 8064 10639
rect 8024 10600 8076 10606
rect 8024 10542 8076 10548
rect 8022 10432 8078 10441
rect 8022 10367 8078 10376
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7562 7168 7618 7177
rect 7562 7103 7618 7112
rect 7482 6886 7512 6914
rect 7668 6914 7696 7686
rect 7852 7546 7880 7754
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7852 7002 7880 7346
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7840 6996 7892 7002
rect 7840 6938 7892 6944
rect 7944 6934 7972 7278
rect 7932 6928 7984 6934
rect 7668 6886 7788 6914
rect 7300 6854 7418 6882
rect 7390 6848 7418 6854
rect 7390 6820 7420 6848
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7300 6633 7328 6734
rect 7286 6624 7342 6633
rect 7286 6559 7342 6568
rect 7286 6488 7342 6497
rect 7286 6423 7342 6432
rect 7300 6390 7328 6423
rect 7288 6384 7340 6390
rect 7288 6326 7340 6332
rect 7392 6304 7420 6820
rect 7482 6798 7510 6886
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7760 6440 7788 6886
rect 7932 6870 7984 6876
rect 7930 6760 7986 6769
rect 7930 6695 7986 6704
rect 7668 6412 7788 6440
rect 7392 6276 7512 6304
rect 7286 6080 7342 6089
rect 7286 6015 7342 6024
rect 7196 5840 7248 5846
rect 7196 5782 7248 5788
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 7010 4856 7066 4865
rect 6932 4814 7010 4842
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6734 4584 6790 4593
rect 6734 4519 6736 4528
rect 6788 4519 6790 4528
rect 6736 4490 6788 4496
rect 6828 4480 6880 4486
rect 6734 4448 6790 4457
rect 6828 4422 6880 4428
rect 6734 4383 6790 4392
rect 6748 3942 6776 4383
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6736 3528 6788 3534
rect 6840 3505 6868 4422
rect 6736 3470 6788 3476
rect 6826 3496 6882 3505
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 6748 2961 6776 3470
rect 6826 3431 6882 3440
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6734 2952 6790 2961
rect 6552 2916 6604 2922
rect 6734 2887 6790 2896
rect 6552 2858 6604 2864
rect 6460 2644 6512 2650
rect 6460 2586 6512 2592
rect 6380 2502 6500 2530
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 6276 2372 6328 2378
rect 6276 2314 6328 2320
rect 5908 2304 5960 2310
rect 5828 2264 5908 2292
rect 5354 54 5488 82
rect 5354 -300 5410 54
rect 5538 -300 5594 160
rect 5722 -300 5778 160
rect 5828 82 5856 2264
rect 5908 2246 5960 2252
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 5894 2204 6202 2213
rect 5894 2202 5900 2204
rect 5956 2202 5980 2204
rect 6036 2202 6060 2204
rect 6116 2202 6140 2204
rect 6196 2202 6202 2204
rect 5956 2150 5958 2202
rect 6138 2150 6140 2202
rect 5894 2148 5900 2150
rect 5956 2148 5980 2150
rect 6036 2148 6060 2150
rect 6116 2148 6140 2150
rect 6196 2148 6202 2150
rect 5894 2139 6202 2148
rect 6090 2000 6146 2009
rect 6090 1935 6146 1944
rect 6000 1760 6052 1766
rect 6000 1702 6052 1708
rect 6012 1494 6040 1702
rect 6104 1562 6132 1935
rect 6288 1834 6316 2314
rect 6276 1828 6328 1834
rect 6276 1770 6328 1776
rect 6092 1556 6144 1562
rect 6092 1498 6144 1504
rect 6000 1488 6052 1494
rect 6380 1442 6408 2382
rect 6000 1430 6052 1436
rect 6288 1414 6408 1442
rect 6472 1442 6500 2502
rect 6564 2106 6592 2858
rect 6644 2848 6696 2854
rect 6644 2790 6696 2796
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6656 2446 6684 2790
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6552 2100 6604 2106
rect 6552 2042 6604 2048
rect 6642 2000 6698 2009
rect 6642 1935 6698 1944
rect 6656 1562 6684 1935
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 6472 1414 6592 1442
rect 5894 1116 6202 1125
rect 5894 1114 5900 1116
rect 5956 1114 5980 1116
rect 6036 1114 6060 1116
rect 6116 1114 6140 1116
rect 6196 1114 6202 1116
rect 5956 1062 5958 1114
rect 6138 1062 6140 1114
rect 5894 1060 5900 1062
rect 5956 1060 5980 1062
rect 6036 1060 6060 1062
rect 6116 1060 6140 1062
rect 6196 1060 6202 1062
rect 5894 1051 6202 1060
rect 6092 740 6144 746
rect 6092 682 6144 688
rect 6104 160 6132 682
rect 6288 160 6316 1414
rect 6564 1358 6592 1414
rect 6748 1358 6776 2790
rect 6840 2106 6868 3334
rect 6932 3210 6960 4814
rect 7116 4826 7144 5510
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7208 4826 7236 5170
rect 7010 4791 7066 4800
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7300 4457 7328 6015
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7286 4448 7342 4457
rect 7286 4383 7342 4392
rect 7288 4208 7340 4214
rect 7288 4150 7340 4156
rect 7300 4049 7328 4150
rect 7286 4040 7342 4049
rect 7286 3975 7342 3984
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7012 3528 7064 3534
rect 7012 3470 7064 3476
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7024 3369 7052 3470
rect 7010 3360 7066 3369
rect 7010 3295 7066 3304
rect 6932 3182 7052 3210
rect 6918 3088 6974 3097
rect 6918 3023 6974 3032
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 6932 1970 6960 3023
rect 7024 2650 7052 3182
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7010 2408 7066 2417
rect 7010 2343 7066 2352
rect 7024 2106 7052 2343
rect 7012 2100 7064 2106
rect 7012 2042 7064 2048
rect 6920 1964 6972 1970
rect 6920 1906 6972 1912
rect 6826 1864 6882 1873
rect 7116 1850 7144 3470
rect 7208 3233 7236 3606
rect 7194 3224 7250 3233
rect 7392 3194 7420 5170
rect 7484 4078 7512 6276
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7576 4758 7604 6054
rect 7668 5409 7696 6412
rect 7944 6304 7972 6695
rect 7760 6276 7972 6304
rect 7654 5400 7710 5409
rect 7654 5335 7710 5344
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7668 5001 7696 5238
rect 7654 4992 7710 5001
rect 7654 4927 7710 4936
rect 7564 4752 7616 4758
rect 7564 4694 7616 4700
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7760 3738 7788 6276
rect 7930 6216 7986 6225
rect 7930 6151 7986 6160
rect 7944 5370 7972 6151
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7852 5273 7880 5306
rect 7838 5264 7894 5273
rect 7838 5199 7894 5208
rect 7838 3904 7894 3913
rect 7838 3839 7894 3848
rect 7852 3738 7880 3839
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 8036 3618 8064 10367
rect 8128 10062 8156 10678
rect 8220 10130 8248 12242
rect 8312 12238 8340 12430
rect 8668 12368 8720 12374
rect 8668 12310 8720 12316
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8576 12232 8628 12238
rect 8576 12174 8628 12180
rect 8588 12073 8616 12174
rect 8574 12064 8630 12073
rect 8574 11999 8630 12008
rect 8680 11830 8708 12310
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8367 11452 8675 11461
rect 8367 11450 8373 11452
rect 8429 11450 8453 11452
rect 8509 11450 8533 11452
rect 8589 11450 8613 11452
rect 8669 11450 8675 11452
rect 8429 11398 8431 11450
rect 8611 11398 8613 11450
rect 8367 11396 8373 11398
rect 8429 11396 8453 11398
rect 8509 11396 8533 11398
rect 8589 11396 8613 11398
rect 8669 11396 8675 11398
rect 8367 11387 8675 11396
rect 8392 11076 8444 11082
rect 8392 11018 8444 11024
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10418 8340 10950
rect 8404 10742 8432 11018
rect 8392 10736 8444 10742
rect 8392 10678 8444 10684
rect 8310 10390 8340 10418
rect 8576 10464 8628 10470
rect 8628 10424 8733 10452
rect 8576 10406 8628 10412
rect 8310 10282 8338 10390
rect 8367 10364 8675 10373
rect 8367 10362 8373 10364
rect 8429 10362 8453 10364
rect 8509 10362 8533 10364
rect 8589 10362 8613 10364
rect 8669 10362 8675 10364
rect 8429 10310 8431 10362
rect 8611 10310 8613 10362
rect 8367 10308 8373 10310
rect 8429 10308 8453 10310
rect 8509 10308 8533 10310
rect 8589 10308 8613 10310
rect 8669 10308 8675 10310
rect 8367 10299 8675 10308
rect 8310 10254 8340 10282
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8220 9897 8248 10066
rect 8312 10062 8340 10254
rect 8705 10248 8733 10424
rect 8772 10418 8800 14028
rect 8852 14010 8904 14016
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 8864 12238 8892 13738
rect 8852 12232 8904 12238
rect 8852 12174 8904 12180
rect 8852 11824 8904 11830
rect 8852 11766 8904 11772
rect 8864 10810 8892 11766
rect 8852 10804 8904 10810
rect 8852 10746 8904 10752
rect 8772 10390 8892 10418
rect 8496 10220 8733 10248
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8392 9920 8444 9926
rect 8206 9888 8262 9897
rect 8392 9862 8444 9868
rect 8206 9823 8262 9832
rect 8114 9752 8170 9761
rect 8298 9752 8354 9761
rect 8114 9687 8170 9696
rect 8220 9710 8298 9738
rect 8128 7920 8156 9687
rect 8220 9217 8248 9710
rect 8404 9722 8432 9862
rect 8298 9687 8354 9696
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8496 9586 8524 10220
rect 8758 10160 8814 10169
rect 8758 10095 8760 10104
rect 8812 10095 8814 10104
rect 8760 10066 8812 10072
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8588 9466 8616 9998
rect 8666 9752 8722 9761
rect 8722 9710 8800 9738
rect 8666 9687 8722 9696
rect 8312 9438 8616 9466
rect 8312 9330 8340 9438
rect 8404 9382 8432 9438
rect 8310 9302 8340 9330
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8206 9208 8262 9217
rect 8310 9194 8338 9302
rect 8367 9276 8675 9285
rect 8367 9274 8373 9276
rect 8429 9274 8453 9276
rect 8509 9274 8533 9276
rect 8589 9274 8613 9276
rect 8669 9274 8675 9276
rect 8429 9222 8431 9274
rect 8611 9222 8613 9274
rect 8367 9220 8373 9222
rect 8429 9220 8453 9222
rect 8509 9220 8533 9222
rect 8589 9220 8613 9222
rect 8669 9220 8675 9222
rect 8367 9211 8675 9220
rect 8310 9166 8340 9194
rect 8206 9143 8262 9152
rect 8206 9072 8262 9081
rect 8206 9007 8208 9016
rect 8260 9007 8262 9016
rect 8208 8978 8260 8984
rect 8312 8922 8340 9166
rect 8574 9072 8630 9081
rect 8574 9007 8630 9016
rect 8220 8894 8340 8922
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8116 7914 8168 7920
rect 8116 7856 8168 7862
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 7576 3590 8064 3618
rect 7194 3159 7250 3168
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7472 3052 7524 3058
rect 6826 1799 6882 1808
rect 7024 1822 7144 1850
rect 7208 3012 7472 3040
rect 6840 1562 6868 1799
rect 6920 1760 6972 1766
rect 6920 1702 6972 1708
rect 6828 1556 6880 1562
rect 6828 1498 6880 1504
rect 6368 1352 6420 1358
rect 6552 1352 6604 1358
rect 6420 1312 6500 1340
rect 6368 1294 6420 1300
rect 6472 160 6500 1312
rect 6552 1294 6604 1300
rect 6736 1352 6788 1358
rect 6736 1294 6788 1300
rect 6932 1034 6960 1702
rect 6840 1006 6960 1034
rect 6644 672 6696 678
rect 6644 614 6696 620
rect 6656 160 6684 614
rect 6840 160 6868 1006
rect 7024 160 7052 1822
rect 7208 160 7236 3012
rect 7472 2994 7524 3000
rect 7576 2938 7604 3590
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7484 2910 7604 2938
rect 7286 2680 7342 2689
rect 7286 2615 7342 2624
rect 7300 2446 7328 2615
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7392 160 7420 2858
rect 7484 2650 7512 2910
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7472 2644 7524 2650
rect 7472 2586 7524 2592
rect 7470 2272 7526 2281
rect 7470 2207 7526 2216
rect 7484 1834 7512 2207
rect 7576 1970 7604 2790
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 7668 1850 7696 3470
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7760 1970 7788 3334
rect 7944 3233 7972 3470
rect 7930 3224 7986 3233
rect 7930 3159 7986 3168
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 8024 3052 8076 3058
rect 8128 3040 8156 7754
rect 8220 7478 8248 8894
rect 8392 8832 8444 8838
rect 8392 8774 8444 8780
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8312 8242 8340 8502
rect 8404 8401 8432 8774
rect 8496 8673 8524 8910
rect 8482 8664 8538 8673
rect 8482 8599 8538 8608
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8390 8392 8446 8401
rect 8390 8327 8446 8336
rect 8496 8276 8524 8502
rect 8588 8498 8616 9007
rect 8772 8634 8800 9710
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8668 8492 8720 8498
rect 8720 8452 8800 8480
rect 8668 8434 8720 8440
rect 8496 8248 8733 8276
rect 8310 8214 8340 8242
rect 8310 8106 8338 8214
rect 8367 8188 8675 8197
rect 8367 8186 8373 8188
rect 8429 8186 8453 8188
rect 8509 8186 8533 8188
rect 8589 8186 8613 8188
rect 8669 8186 8675 8188
rect 8429 8134 8431 8186
rect 8611 8134 8613 8186
rect 8367 8132 8373 8134
rect 8429 8132 8453 8134
rect 8509 8132 8533 8134
rect 8589 8132 8613 8134
rect 8669 8132 8675 8134
rect 8367 8123 8675 8132
rect 8310 8090 8340 8106
rect 8300 8084 8352 8090
rect 8705 8072 8733 8248
rect 8300 8026 8352 8032
rect 8680 8044 8733 8072
rect 8300 7880 8352 7886
rect 8680 7857 8708 8044
rect 8300 7822 8352 7828
rect 8666 7848 8722 7857
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8208 7200 8260 7206
rect 8312 7154 8340 7822
rect 8666 7783 8722 7792
rect 8666 7712 8722 7721
rect 8666 7647 8722 7656
rect 8680 7188 8708 7647
rect 8680 7160 8733 7188
rect 8208 7142 8260 7148
rect 8220 6458 8248 7142
rect 8310 7126 8340 7154
rect 8310 7018 8338 7126
rect 8367 7100 8675 7109
rect 8367 7098 8373 7100
rect 8429 7098 8453 7100
rect 8509 7098 8533 7100
rect 8589 7098 8613 7100
rect 8669 7098 8675 7100
rect 8429 7046 8431 7098
rect 8611 7046 8613 7098
rect 8367 7044 8373 7046
rect 8429 7044 8453 7046
rect 8509 7044 8533 7046
rect 8589 7044 8613 7046
rect 8669 7044 8675 7046
rect 8367 7035 8675 7044
rect 8310 6990 8340 7018
rect 8312 6984 8340 6990
rect 8705 6984 8733 7160
rect 8312 6956 8432 6984
rect 8404 6914 8432 6956
rect 8312 6886 8432 6914
rect 8588 6956 8733 6984
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8312 6202 8340 6886
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8390 6624 8446 6633
rect 8390 6559 8446 6568
rect 8220 6174 8340 6202
rect 8220 4865 8248 6174
rect 8404 6100 8432 6559
rect 8496 6458 8524 6802
rect 8484 6452 8536 6458
rect 8484 6394 8536 6400
rect 8588 6225 8616 6956
rect 8772 6914 8800 8452
rect 8680 6886 8800 6914
rect 8574 6216 8630 6225
rect 8574 6151 8630 6160
rect 8312 6072 8432 6100
rect 8680 6100 8708 6886
rect 8680 6072 8800 6100
rect 8312 6066 8340 6072
rect 8310 6038 8340 6066
rect 8310 5930 8338 6038
rect 8367 6012 8675 6021
rect 8367 6010 8373 6012
rect 8429 6010 8453 6012
rect 8509 6010 8533 6012
rect 8589 6010 8613 6012
rect 8669 6010 8675 6012
rect 8429 5958 8431 6010
rect 8611 5958 8613 6010
rect 8367 5956 8373 5958
rect 8429 5956 8453 5958
rect 8509 5956 8533 5958
rect 8589 5956 8613 5958
rect 8669 5956 8675 5958
rect 8367 5947 8675 5956
rect 8310 5902 8340 5930
rect 8312 4978 8340 5902
rect 8666 5808 8722 5817
rect 8392 5772 8444 5778
rect 8666 5743 8722 5752
rect 8392 5714 8444 5720
rect 8404 5234 8432 5714
rect 8680 5234 8708 5743
rect 8772 5642 8800 6072
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8668 5228 8720 5234
rect 8720 5188 8800 5216
rect 8668 5170 8720 5176
rect 8310 4950 8340 4978
rect 8206 4856 8262 4865
rect 8310 4842 8338 4950
rect 8367 4924 8675 4933
rect 8367 4922 8373 4924
rect 8429 4922 8453 4924
rect 8509 4922 8533 4924
rect 8589 4922 8613 4924
rect 8669 4922 8675 4924
rect 8429 4870 8431 4922
rect 8611 4870 8613 4922
rect 8367 4868 8373 4870
rect 8429 4868 8453 4870
rect 8509 4868 8533 4870
rect 8589 4868 8613 4870
rect 8669 4868 8675 4870
rect 8367 4859 8675 4868
rect 8310 4814 8340 4842
rect 8206 4791 8262 4800
rect 8312 4706 8340 4814
rect 8220 4678 8340 4706
rect 8220 3176 8248 4678
rect 8772 4146 8800 5188
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8367 3836 8675 3845
rect 8367 3834 8373 3836
rect 8429 3834 8453 3836
rect 8509 3834 8533 3836
rect 8589 3834 8613 3836
rect 8669 3834 8675 3836
rect 8429 3782 8431 3834
rect 8611 3782 8613 3834
rect 8367 3780 8373 3782
rect 8429 3780 8453 3782
rect 8509 3780 8533 3782
rect 8589 3780 8613 3782
rect 8669 3780 8675 3782
rect 8367 3771 8675 3780
rect 8390 3632 8446 3641
rect 8390 3567 8446 3576
rect 8300 3188 8352 3194
rect 8220 3148 8300 3176
rect 8300 3130 8352 3136
rect 8404 3126 8432 3567
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8864 3058 8892 10390
rect 8300 3052 8352 3058
rect 8076 3012 8156 3040
rect 8220 3012 8300 3040
rect 8024 2994 8076 3000
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7852 2106 7880 2790
rect 7840 2100 7892 2106
rect 7840 2042 7892 2048
rect 7748 1964 7800 1970
rect 7748 1906 7800 1912
rect 7472 1828 7524 1834
rect 7668 1822 7788 1850
rect 7472 1770 7524 1776
rect 7656 1760 7708 1766
rect 7656 1702 7708 1708
rect 7564 1216 7616 1222
rect 7564 1158 7616 1164
rect 7576 785 7604 1158
rect 7668 1018 7696 1702
rect 7656 1012 7708 1018
rect 7656 954 7708 960
rect 7562 776 7618 785
rect 7562 711 7618 720
rect 7484 190 7604 218
rect 5906 82 5962 160
rect 5828 54 5962 82
rect 5906 -300 5962 54
rect 6090 -300 6146 160
rect 6274 -300 6330 160
rect 6458 -300 6514 160
rect 6642 -300 6698 160
rect 6826 -300 6882 160
rect 7010 -300 7066 160
rect 7194 -300 7250 160
rect 7378 -300 7434 160
rect 7484 105 7512 190
rect 7576 160 7604 190
rect 7760 160 7788 1822
rect 7840 1828 7892 1834
rect 7840 1770 7892 1776
rect 7852 1358 7880 1770
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 7944 160 7972 2994
rect 8220 2938 8248 3012
rect 8300 2994 8352 3000
rect 8576 3052 8628 3058
rect 8852 3052 8904 3058
rect 8628 3012 8800 3040
rect 8576 2994 8628 3000
rect 8036 2910 8248 2938
rect 8036 1442 8064 2910
rect 8116 2848 8168 2854
rect 8392 2848 8444 2854
rect 8116 2790 8168 2796
rect 8220 2808 8392 2836
rect 8128 2038 8156 2790
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 8220 1970 8248 2808
rect 8392 2790 8444 2796
rect 8367 2748 8675 2757
rect 8367 2746 8373 2748
rect 8429 2746 8453 2748
rect 8509 2746 8533 2748
rect 8589 2746 8613 2748
rect 8669 2746 8675 2748
rect 8429 2694 8431 2746
rect 8611 2694 8613 2746
rect 8367 2692 8373 2694
rect 8429 2692 8453 2694
rect 8509 2692 8533 2694
rect 8589 2692 8613 2694
rect 8669 2692 8675 2694
rect 8367 2683 8675 2692
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 8404 2446 8432 2586
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8588 2038 8616 2246
rect 8484 2032 8536 2038
rect 8482 2000 8484 2009
rect 8576 2032 8628 2038
rect 8536 2000 8538 2009
rect 8208 1964 8260 1970
rect 8576 1974 8628 1980
rect 8482 1935 8538 1944
rect 8208 1906 8260 1912
rect 8116 1760 8168 1766
rect 8208 1760 8260 1766
rect 8116 1702 8168 1708
rect 8206 1728 8208 1737
rect 8260 1728 8262 1737
rect 8128 1601 8156 1702
rect 8206 1663 8262 1672
rect 8367 1660 8675 1669
rect 8367 1658 8373 1660
rect 8429 1658 8453 1660
rect 8509 1658 8533 1660
rect 8589 1658 8613 1660
rect 8669 1658 8675 1660
rect 8429 1606 8431 1658
rect 8611 1606 8613 1658
rect 8367 1604 8373 1606
rect 8429 1604 8453 1606
rect 8509 1604 8533 1606
rect 8589 1604 8613 1606
rect 8669 1604 8675 1606
rect 8114 1592 8170 1601
rect 8367 1595 8675 1604
rect 8772 1578 8800 3012
rect 8956 3040 8984 15166
rect 9048 14006 9076 20810
rect 9140 20584 9168 26522
rect 9232 26042 9260 28206
rect 9220 26036 9272 26042
rect 9220 25978 9272 25984
rect 9220 25696 9272 25702
rect 9220 25638 9272 25644
rect 9232 25294 9260 25638
rect 9220 25288 9272 25294
rect 9220 25230 9272 25236
rect 9220 25152 9272 25158
rect 9324 25129 9352 29582
rect 9404 29232 9456 29238
rect 9404 29174 9456 29180
rect 9416 29073 9444 29174
rect 9402 29064 9458 29073
rect 9402 28999 9458 29008
rect 9404 28416 9456 28422
rect 9404 28358 9456 28364
rect 9416 28150 9444 28358
rect 9404 28144 9456 28150
rect 9404 28086 9456 28092
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9416 26246 9444 26862
rect 9404 26240 9456 26246
rect 9404 26182 9456 26188
rect 9404 26036 9456 26042
rect 9404 25978 9456 25984
rect 9416 25158 9444 25978
rect 9404 25152 9456 25158
rect 9220 25094 9272 25100
rect 9310 25120 9366 25129
rect 9232 24596 9260 25094
rect 9508 25106 9536 32166
rect 9600 30394 9628 32286
rect 9692 32201 9720 32370
rect 9678 32192 9734 32201
rect 9678 32127 9734 32136
rect 9784 32042 9812 33918
rect 9954 33824 10010 33833
rect 9954 33759 10010 33768
rect 9864 32768 9916 32774
rect 9864 32710 9916 32716
rect 9692 32014 9812 32042
rect 9692 30580 9720 32014
rect 9876 31328 9904 32710
rect 9968 32065 9996 33759
rect 9954 32056 10010 32065
rect 9954 31991 10010 32000
rect 10060 31668 10088 36094
rect 10152 35834 10180 42502
rect 10244 41546 10272 43336
rect 10416 43318 10468 43324
rect 10324 42696 10376 42702
rect 10520 42684 10548 44540
rect 10704 43874 10732 44540
rect 10612 43846 10732 43874
rect 10612 43450 10640 43846
rect 10888 43738 10916 44540
rect 10704 43710 10916 43738
rect 11072 43738 11100 44540
rect 11256 43874 11284 44540
rect 11256 43846 11376 43874
rect 11072 43710 11284 43738
rect 10600 43444 10652 43450
rect 10600 43386 10652 43392
rect 10598 43344 10654 43353
rect 10598 43279 10654 43288
rect 10376 42656 10548 42684
rect 10324 42638 10376 42644
rect 10612 42226 10640 43279
rect 10704 42684 10732 43710
rect 10839 43548 11147 43557
rect 10839 43546 10845 43548
rect 10901 43546 10925 43548
rect 10981 43546 11005 43548
rect 11061 43546 11085 43548
rect 11141 43546 11147 43548
rect 10901 43494 10903 43546
rect 11083 43494 11085 43546
rect 10839 43492 10845 43494
rect 10901 43492 10925 43494
rect 10981 43492 11005 43494
rect 11061 43492 11085 43494
rect 11141 43492 11147 43494
rect 10839 43483 11147 43492
rect 10784 43308 10836 43314
rect 10784 43250 10836 43256
rect 10796 42945 10824 43250
rect 11152 43104 11204 43110
rect 11152 43046 11204 43052
rect 10782 42936 10838 42945
rect 10782 42871 10838 42880
rect 10876 42900 10928 42906
rect 10876 42842 10928 42848
rect 10888 42786 10916 42842
rect 10888 42758 11008 42786
rect 10876 42696 10928 42702
rect 10704 42656 10876 42684
rect 10876 42638 10928 42644
rect 10980 42548 11008 42758
rect 11164 42566 11192 43046
rect 10704 42520 11008 42548
rect 11152 42560 11204 42566
rect 10600 42220 10652 42226
rect 10600 42162 10652 42168
rect 10324 42084 10376 42090
rect 10324 42026 10376 42032
rect 10232 41540 10284 41546
rect 10232 41482 10284 41488
rect 10336 41414 10364 42026
rect 10416 42016 10468 42022
rect 10416 41958 10468 41964
rect 10244 41386 10364 41414
rect 10244 37942 10272 41386
rect 10324 38412 10376 38418
rect 10324 38354 10376 38360
rect 10336 38010 10364 38354
rect 10428 38214 10456 41958
rect 10508 38344 10560 38350
rect 10598 38312 10654 38321
rect 10560 38292 10598 38298
rect 10508 38286 10598 38292
rect 10520 38270 10598 38286
rect 10598 38247 10654 38256
rect 10416 38208 10468 38214
rect 10508 38208 10560 38214
rect 10416 38150 10468 38156
rect 10506 38176 10508 38185
rect 10560 38176 10562 38185
rect 10506 38111 10562 38120
rect 10324 38004 10376 38010
rect 10324 37946 10376 37952
rect 10232 37936 10284 37942
rect 10232 37878 10284 37884
rect 10416 36848 10468 36854
rect 10416 36790 10468 36796
rect 10428 36417 10456 36790
rect 10414 36408 10470 36417
rect 10414 36343 10470 36352
rect 10324 36032 10376 36038
rect 10324 35974 10376 35980
rect 10336 35873 10364 35974
rect 10322 35864 10378 35873
rect 10140 35828 10192 35834
rect 10140 35770 10192 35776
rect 10232 35828 10284 35834
rect 10322 35799 10378 35808
rect 10232 35770 10284 35776
rect 10140 35692 10192 35698
rect 10140 35634 10192 35640
rect 10152 34649 10180 35634
rect 10138 34640 10194 34649
rect 10138 34575 10194 34584
rect 10140 34196 10192 34202
rect 10140 34138 10192 34144
rect 10152 31822 10180 34138
rect 10244 32230 10272 35770
rect 10324 35284 10376 35290
rect 10324 35226 10376 35232
rect 10336 35018 10364 35226
rect 10324 35012 10376 35018
rect 10324 34954 10376 34960
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 10336 33998 10364 34682
rect 10428 34202 10456 36343
rect 10520 35873 10548 38111
rect 10600 38004 10652 38010
rect 10600 37946 10652 37952
rect 10612 37874 10640 37946
rect 10600 37868 10652 37874
rect 10600 37810 10652 37816
rect 10600 37460 10652 37466
rect 10600 37402 10652 37408
rect 10506 35864 10562 35873
rect 10506 35799 10562 35808
rect 10508 35760 10560 35766
rect 10508 35702 10560 35708
rect 10520 35193 10548 35702
rect 10612 35630 10640 37402
rect 10600 35624 10652 35630
rect 10600 35566 10652 35572
rect 10600 35284 10652 35290
rect 10600 35226 10652 35232
rect 10506 35184 10562 35193
rect 10506 35119 10562 35128
rect 10612 34490 10640 35226
rect 10520 34462 10640 34490
rect 10416 34196 10468 34202
rect 10416 34138 10468 34144
rect 10324 33992 10376 33998
rect 10324 33934 10376 33940
rect 10520 33114 10548 34462
rect 10600 34400 10652 34406
rect 10600 34342 10652 34348
rect 10508 33108 10560 33114
rect 10508 33050 10560 33056
rect 10232 32224 10284 32230
rect 10232 32166 10284 32172
rect 10508 32224 10560 32230
rect 10508 32166 10560 32172
rect 10230 32056 10286 32065
rect 10230 31991 10286 32000
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10060 31640 10180 31668
rect 9784 31300 9904 31328
rect 10048 31340 10100 31346
rect 9784 31210 9812 31300
rect 10048 31282 10100 31288
rect 9772 31204 9824 31210
rect 9772 31146 9824 31152
rect 9864 31204 9916 31210
rect 9916 31164 9996 31192
rect 9864 31146 9916 31152
rect 9770 30832 9826 30841
rect 9770 30767 9826 30776
rect 9784 30734 9812 30767
rect 9772 30728 9824 30734
rect 9772 30670 9824 30676
rect 9692 30552 9812 30580
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9600 28744 9628 30330
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9692 29306 9720 29990
rect 9680 29300 9732 29306
rect 9680 29242 9732 29248
rect 9600 28716 9720 28744
rect 9586 28656 9642 28665
rect 9586 28591 9642 28600
rect 9600 28558 9628 28591
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9404 25094 9456 25100
rect 9310 25055 9366 25064
rect 9506 25078 9536 25106
rect 9506 24970 9534 25078
rect 9404 24948 9456 24954
rect 9506 24942 9536 24970
rect 9692 24954 9720 28716
rect 9784 25129 9812 30552
rect 9864 29504 9916 29510
rect 9864 29446 9916 29452
rect 9876 29306 9904 29446
rect 9864 29300 9916 29306
rect 9864 29242 9916 29248
rect 9862 28928 9918 28937
rect 9862 28863 9918 28872
rect 9876 26194 9904 28863
rect 9968 28404 9996 31164
rect 10060 30734 10088 31282
rect 10048 30728 10100 30734
rect 10048 30670 10100 30676
rect 10060 30054 10088 30670
rect 10048 30048 10100 30054
rect 10048 29990 10100 29996
rect 10048 29504 10100 29510
rect 10048 29446 10100 29452
rect 10060 28558 10088 29446
rect 10048 28552 10100 28558
rect 10048 28494 10100 28500
rect 9968 28393 10054 28404
rect 9968 28384 10102 28393
rect 9968 28376 10046 28384
rect 10026 28342 10046 28376
rect 10046 28319 10102 28328
rect 9956 27124 10008 27130
rect 9956 27066 10008 27072
rect 9968 26353 9996 27066
rect 9954 26344 10010 26353
rect 10060 26330 10088 28319
rect 10152 26586 10180 31640
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 10060 26302 10180 26330
rect 9954 26279 10010 26288
rect 10048 26240 10100 26246
rect 9876 26166 9996 26194
rect 10048 26182 10100 26188
rect 9862 26072 9918 26081
rect 9862 26007 9918 26016
rect 9770 25120 9826 25129
rect 9770 25055 9826 25064
rect 9404 24890 9456 24896
rect 9416 24818 9444 24890
rect 9508 24834 9536 24942
rect 9680 24948 9732 24954
rect 9680 24890 9732 24896
rect 9770 24848 9826 24857
rect 9404 24812 9456 24818
rect 9508 24806 9628 24834
rect 9404 24754 9456 24760
rect 9232 24568 9352 24596
rect 9218 23624 9274 23633
rect 9218 23559 9274 23568
rect 9232 23254 9260 23559
rect 9324 23497 9352 24568
rect 9310 23488 9366 23497
rect 9310 23423 9366 23432
rect 9220 23248 9272 23254
rect 9220 23190 9272 23196
rect 9312 22976 9364 22982
rect 9312 22918 9364 22924
rect 9218 22808 9274 22817
rect 9218 22743 9220 22752
rect 9272 22743 9274 22752
rect 9220 22714 9272 22720
rect 9220 22500 9272 22506
rect 9220 22442 9272 22448
rect 9232 22030 9260 22442
rect 9324 22098 9352 22918
rect 9416 22778 9444 24754
rect 9496 24744 9548 24750
rect 9496 24686 9548 24692
rect 9508 24410 9536 24686
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9496 24064 9548 24070
rect 9496 24006 9548 24012
rect 9508 23866 9536 24006
rect 9496 23860 9548 23866
rect 9496 23802 9548 23808
rect 9496 23316 9548 23322
rect 9496 23258 9548 23264
rect 9508 23118 9536 23258
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9404 22772 9456 22778
rect 9404 22714 9456 22720
rect 9312 22092 9364 22098
rect 9312 22034 9364 22040
rect 9220 22024 9272 22030
rect 9220 21966 9272 21972
rect 9416 21672 9444 22714
rect 9508 22574 9536 23054
rect 9600 22778 9628 24806
rect 9770 24783 9826 24792
rect 9784 24290 9812 24783
rect 9692 24262 9812 24290
rect 9588 22772 9640 22778
rect 9588 22714 9640 22720
rect 9588 22636 9640 22642
rect 9588 22578 9640 22584
rect 9496 22568 9548 22574
rect 9496 22510 9548 22516
rect 9600 22234 9628 22578
rect 9588 22228 9640 22234
rect 9588 22170 9640 22176
rect 9416 21644 9628 21672
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9404 21480 9456 21486
rect 9310 21448 9366 21457
rect 9404 21422 9456 21428
rect 9310 21383 9312 21392
rect 9364 21383 9366 21392
rect 9312 21354 9364 21360
rect 9140 20556 9352 20584
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9140 19514 9168 19790
rect 9128 19508 9180 19514
rect 9128 19450 9180 19456
rect 9220 18624 9272 18630
rect 9220 18566 9272 18572
rect 9232 17134 9260 18566
rect 9324 18193 9352 20556
rect 9416 19174 9444 21422
rect 9508 19854 9536 21490
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9404 19168 9456 19174
rect 9404 19110 9456 19116
rect 9496 19168 9548 19174
rect 9496 19110 9548 19116
rect 9402 19000 9458 19009
rect 9402 18935 9458 18944
rect 9310 18184 9366 18193
rect 9310 18119 9366 18128
rect 9416 17728 9444 18935
rect 9508 18426 9536 19110
rect 9496 18420 9548 18426
rect 9496 18362 9548 18368
rect 9600 18290 9628 21644
rect 9692 19446 9720 24262
rect 9772 24200 9824 24206
rect 9772 24142 9824 24148
rect 9784 23798 9812 24142
rect 9876 24018 9904 26007
rect 9968 25242 9996 26166
rect 10060 26042 10088 26182
rect 10152 26081 10180 26302
rect 10138 26072 10194 26081
rect 10048 26036 10100 26042
rect 10138 26007 10194 26016
rect 10048 25978 10100 25984
rect 10140 25968 10192 25974
rect 10140 25910 10192 25916
rect 10046 25800 10102 25809
rect 10046 25735 10102 25744
rect 10060 25362 10088 25735
rect 10152 25401 10180 25910
rect 10138 25392 10194 25401
rect 10048 25356 10100 25362
rect 10138 25327 10194 25336
rect 10048 25298 10100 25304
rect 9968 25214 10088 25242
rect 9956 25152 10008 25158
rect 9956 25094 10008 25100
rect 9968 24585 9996 25094
rect 10060 24857 10088 25214
rect 10140 25152 10192 25158
rect 10140 25094 10192 25100
rect 10046 24848 10102 24857
rect 10046 24783 10102 24792
rect 9954 24576 10010 24585
rect 9954 24511 10010 24520
rect 10152 24426 10180 25094
rect 9968 24398 10180 24426
rect 9968 24138 9996 24398
rect 9956 24132 10008 24138
rect 9956 24074 10008 24080
rect 10140 24132 10192 24138
rect 10140 24074 10192 24080
rect 10152 24018 10180 24074
rect 9876 23990 10180 24018
rect 9954 23896 10010 23905
rect 10244 23882 10272 31991
rect 10520 31754 10548 32166
rect 10336 31726 10548 31754
rect 10336 31346 10364 31726
rect 10414 31512 10470 31521
rect 10414 31447 10416 31456
rect 10468 31447 10470 31456
rect 10416 31418 10468 31424
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10508 31136 10560 31142
rect 10508 31078 10560 31084
rect 10324 30932 10376 30938
rect 10324 30874 10376 30880
rect 10336 29073 10364 30874
rect 10416 30592 10468 30598
rect 10416 30534 10468 30540
rect 10428 29714 10456 30534
rect 10416 29708 10468 29714
rect 10416 29650 10468 29656
rect 10520 29306 10548 31078
rect 10612 30734 10640 34342
rect 10600 30728 10652 30734
rect 10600 30670 10652 30676
rect 10600 30592 10652 30598
rect 10600 30534 10652 30540
rect 10508 29300 10560 29306
rect 10508 29242 10560 29248
rect 10322 29064 10378 29073
rect 10322 28999 10378 29008
rect 10416 29028 10468 29034
rect 10416 28970 10468 28976
rect 10324 28960 10376 28966
rect 10324 28902 10376 28908
rect 10336 28665 10364 28902
rect 10322 28656 10378 28665
rect 10322 28591 10378 28600
rect 10324 28552 10376 28558
rect 10324 28494 10376 28500
rect 10336 28150 10364 28494
rect 10324 28144 10376 28150
rect 10324 28086 10376 28092
rect 10324 27668 10376 27674
rect 10324 27610 10376 27616
rect 10336 26314 10364 27610
rect 10324 26308 10376 26314
rect 10324 26250 10376 26256
rect 10322 26208 10378 26217
rect 10322 26143 10378 26152
rect 10336 24818 10364 26143
rect 10428 24954 10456 28970
rect 10508 28416 10560 28422
rect 10508 28358 10560 28364
rect 10520 27606 10548 28358
rect 10508 27600 10560 27606
rect 10508 27542 10560 27548
rect 10520 26874 10548 27542
rect 10612 27130 10640 30534
rect 10704 29238 10732 42520
rect 11256 42548 11284 43710
rect 11348 42838 11376 43846
rect 11336 42832 11388 42838
rect 11336 42774 11388 42780
rect 11336 42696 11388 42702
rect 11440 42684 11468 44540
rect 11520 43988 11572 43994
rect 11520 43930 11572 43936
rect 11532 43450 11560 43930
rect 11624 43874 11652 44540
rect 11808 44010 11836 44540
rect 11808 43982 11928 44010
rect 11624 43846 11836 43874
rect 11704 43648 11756 43654
rect 11704 43590 11756 43596
rect 11520 43444 11572 43450
rect 11520 43386 11572 43392
rect 11716 43382 11744 43590
rect 11808 43382 11836 43846
rect 11704 43376 11756 43382
rect 11704 43318 11756 43324
rect 11796 43376 11848 43382
rect 11796 43318 11848 43324
rect 11612 43172 11664 43178
rect 11612 43114 11664 43120
rect 11388 42656 11468 42684
rect 11336 42638 11388 42644
rect 11428 42560 11480 42566
rect 11256 42520 11376 42548
rect 11152 42502 11204 42508
rect 10839 42460 11147 42469
rect 10839 42458 10845 42460
rect 10901 42458 10925 42460
rect 10981 42458 11005 42460
rect 11061 42458 11085 42460
rect 11141 42458 11147 42460
rect 10901 42406 10903 42458
rect 11083 42406 11085 42458
rect 10839 42404 10845 42406
rect 10901 42404 10925 42406
rect 10981 42404 11005 42406
rect 11061 42404 11085 42406
rect 11141 42404 11147 42406
rect 10839 42395 11147 42404
rect 11348 42226 11376 42520
rect 11428 42502 11480 42508
rect 11520 42560 11572 42566
rect 11520 42502 11572 42508
rect 11336 42220 11388 42226
rect 11336 42162 11388 42168
rect 10839 41372 11147 41381
rect 10839 41370 10845 41372
rect 10901 41370 10925 41372
rect 10981 41370 11005 41372
rect 11061 41370 11085 41372
rect 11141 41370 11147 41372
rect 10901 41318 10903 41370
rect 11083 41318 11085 41370
rect 10839 41316 10845 41318
rect 10901 41316 10925 41318
rect 10981 41316 11005 41318
rect 11061 41316 11085 41318
rect 11141 41316 11147 41318
rect 10839 41307 11147 41316
rect 10839 40284 11147 40293
rect 10839 40282 10845 40284
rect 10901 40282 10925 40284
rect 10981 40282 11005 40284
rect 11061 40282 11085 40284
rect 11141 40282 11147 40284
rect 10901 40230 10903 40282
rect 11083 40230 11085 40282
rect 10839 40228 10845 40230
rect 10901 40228 10925 40230
rect 10981 40228 11005 40230
rect 11061 40228 11085 40230
rect 11141 40228 11147 40230
rect 10839 40219 11147 40228
rect 11336 40044 11388 40050
rect 11336 39986 11388 39992
rect 10839 39196 11147 39205
rect 10839 39194 10845 39196
rect 10901 39194 10925 39196
rect 10981 39194 11005 39196
rect 11061 39194 11085 39196
rect 11141 39194 11147 39196
rect 10901 39142 10903 39194
rect 11083 39142 11085 39194
rect 10839 39140 10845 39142
rect 10901 39140 10925 39142
rect 10981 39140 11005 39142
rect 11061 39140 11085 39142
rect 11141 39140 11147 39142
rect 10839 39131 11147 39140
rect 11244 39092 11296 39098
rect 11244 39034 11296 39040
rect 10784 38344 10836 38350
rect 10784 38286 10836 38292
rect 10796 38214 10824 38286
rect 10784 38208 10836 38214
rect 10784 38150 10836 38156
rect 10839 38108 11147 38117
rect 10839 38106 10845 38108
rect 10901 38106 10925 38108
rect 10981 38106 11005 38108
rect 11061 38106 11085 38108
rect 11141 38106 11147 38108
rect 10901 38054 10903 38106
rect 11083 38054 11085 38106
rect 10839 38052 10845 38054
rect 10901 38052 10925 38054
rect 10981 38052 11005 38054
rect 11061 38052 11085 38054
rect 11141 38052 11147 38054
rect 10839 38043 11147 38052
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 10796 37262 10824 37810
rect 11256 37262 11284 39034
rect 10784 37256 10836 37262
rect 10784 37198 10836 37204
rect 11244 37256 11296 37262
rect 11244 37198 11296 37204
rect 10839 37020 11147 37029
rect 10839 37018 10845 37020
rect 10901 37018 10925 37020
rect 10981 37018 11005 37020
rect 11061 37018 11085 37020
rect 11141 37018 11147 37020
rect 10901 36966 10903 37018
rect 11083 36966 11085 37018
rect 10839 36964 10845 36966
rect 10901 36964 10925 36966
rect 10981 36964 11005 36966
rect 11061 36964 11085 36966
rect 11141 36964 11147 36966
rect 10839 36955 11147 36964
rect 11348 36666 11376 39986
rect 11440 39982 11468 42502
rect 11532 41414 11560 42502
rect 11624 42294 11652 43114
rect 11900 42702 11928 43982
rect 11992 43314 12020 44540
rect 12072 43920 12124 43926
rect 12072 43862 12124 43868
rect 11980 43308 12032 43314
rect 11980 43250 12032 43256
rect 11980 43104 12032 43110
rect 11980 43046 12032 43052
rect 11888 42696 11940 42702
rect 11702 42664 11758 42673
rect 11888 42638 11940 42644
rect 11702 42599 11758 42608
rect 11612 42288 11664 42294
rect 11612 42230 11664 42236
rect 11716 41546 11744 42599
rect 11796 42560 11848 42566
rect 11796 42502 11848 42508
rect 11704 41540 11756 41546
rect 11704 41482 11756 41488
rect 11808 41414 11836 42502
rect 11532 41386 11652 41414
rect 11428 39976 11480 39982
rect 11428 39918 11480 39924
rect 11428 39432 11480 39438
rect 11428 39374 11480 39380
rect 11440 36786 11468 39374
rect 11520 38208 11572 38214
rect 11520 38150 11572 38156
rect 11532 38010 11560 38150
rect 11520 38004 11572 38010
rect 11520 37946 11572 37952
rect 11518 37904 11574 37913
rect 11518 37839 11574 37848
rect 11532 37806 11560 37839
rect 11520 37800 11572 37806
rect 11520 37742 11572 37748
rect 11520 37460 11572 37466
rect 11520 37402 11572 37408
rect 11428 36780 11480 36786
rect 11428 36722 11480 36728
rect 11256 36638 11376 36666
rect 11256 36242 11284 36638
rect 11336 36576 11388 36582
rect 11336 36518 11388 36524
rect 11244 36236 11296 36242
rect 11244 36178 11296 36184
rect 10839 35932 11147 35941
rect 10839 35930 10845 35932
rect 10901 35930 10925 35932
rect 10981 35930 11005 35932
rect 11061 35930 11085 35932
rect 11141 35930 11147 35932
rect 10901 35878 10903 35930
rect 11083 35878 11085 35930
rect 10839 35876 10845 35878
rect 10901 35876 10925 35878
rect 10981 35876 11005 35878
rect 11061 35876 11085 35878
rect 11141 35876 11147 35878
rect 10839 35867 11147 35876
rect 10784 35828 10836 35834
rect 10784 35770 10836 35776
rect 10796 35562 10824 35770
rect 10784 35556 10836 35562
rect 10784 35498 10836 35504
rect 10876 35556 10928 35562
rect 10876 35498 10928 35504
rect 10888 34950 10916 35498
rect 11256 35154 11284 36178
rect 11244 35148 11296 35154
rect 11244 35090 11296 35096
rect 11348 35034 11376 36518
rect 11428 36032 11480 36038
rect 11428 35974 11480 35980
rect 11440 35290 11468 35974
rect 11428 35284 11480 35290
rect 11428 35226 11480 35232
rect 11428 35148 11480 35154
rect 11428 35090 11480 35096
rect 11256 35006 11376 35034
rect 10876 34944 10928 34950
rect 10876 34886 10928 34892
rect 10839 34844 11147 34853
rect 10839 34842 10845 34844
rect 10901 34842 10925 34844
rect 10981 34842 11005 34844
rect 11061 34842 11085 34844
rect 11141 34842 11147 34844
rect 10901 34790 10903 34842
rect 11083 34790 11085 34842
rect 10839 34788 10845 34790
rect 10901 34788 10925 34790
rect 10981 34788 11005 34790
rect 11061 34788 11085 34790
rect 11141 34788 11147 34790
rect 10839 34779 11147 34788
rect 11060 34536 11112 34542
rect 11060 34478 11112 34484
rect 11072 33969 11100 34478
rect 11058 33960 11114 33969
rect 11256 33930 11284 35006
rect 11336 34944 11388 34950
rect 11336 34886 11388 34892
rect 11058 33895 11114 33904
rect 11244 33924 11296 33930
rect 11244 33866 11296 33872
rect 10839 33756 11147 33765
rect 10839 33754 10845 33756
rect 10901 33754 10925 33756
rect 10981 33754 11005 33756
rect 11061 33754 11085 33756
rect 11141 33754 11147 33756
rect 10901 33702 10903 33754
rect 11083 33702 11085 33754
rect 10839 33700 10845 33702
rect 10901 33700 10925 33702
rect 10981 33700 11005 33702
rect 11061 33700 11085 33702
rect 11141 33700 11147 33702
rect 10839 33691 11147 33700
rect 11256 33522 11284 33866
rect 11244 33516 11296 33522
rect 11244 33458 11296 33464
rect 11256 33153 11284 33458
rect 11242 33144 11298 33153
rect 11242 33079 11298 33088
rect 11152 32904 11204 32910
rect 11204 32864 11284 32892
rect 11152 32846 11204 32852
rect 10839 32668 11147 32677
rect 10839 32666 10845 32668
rect 10901 32666 10925 32668
rect 10981 32666 11005 32668
rect 11061 32666 11085 32668
rect 11141 32666 11147 32668
rect 10901 32614 10903 32666
rect 11083 32614 11085 32666
rect 10839 32612 10845 32614
rect 10901 32612 10925 32614
rect 10981 32612 11005 32614
rect 11061 32612 11085 32614
rect 11141 32612 11147 32614
rect 10839 32603 11147 32612
rect 10784 32428 10836 32434
rect 10784 32370 10836 32376
rect 10796 31668 10824 32370
rect 11060 32224 11112 32230
rect 11058 32192 11060 32201
rect 11112 32192 11114 32201
rect 11058 32127 11114 32136
rect 10778 31640 10824 31668
rect 10778 31464 10806 31640
rect 10839 31580 11147 31589
rect 10839 31578 10845 31580
rect 10901 31578 10925 31580
rect 10981 31578 11005 31580
rect 11061 31578 11085 31580
rect 11141 31578 11147 31580
rect 10901 31526 10903 31578
rect 11083 31526 11085 31578
rect 10839 31524 10845 31526
rect 10901 31524 10925 31526
rect 10981 31524 11005 31526
rect 11061 31524 11085 31526
rect 11141 31524 11147 31526
rect 10839 31515 11147 31524
rect 10778 31436 10824 31464
rect 10796 31385 10824 31436
rect 10782 31376 10838 31385
rect 10782 31311 10838 31320
rect 11152 31340 11204 31346
rect 10796 30705 10824 31311
rect 11152 31282 11204 31288
rect 11058 31240 11114 31249
rect 11058 31175 11114 31184
rect 11072 30734 11100 31175
rect 11164 30938 11192 31282
rect 11256 30938 11284 32864
rect 11152 30932 11204 30938
rect 11152 30874 11204 30880
rect 11244 30932 11296 30938
rect 11244 30874 11296 30880
rect 11060 30728 11112 30734
rect 10782 30696 10838 30705
rect 11060 30670 11112 30676
rect 10782 30631 10838 30640
rect 11348 30598 11376 34886
rect 11440 34678 11468 35090
rect 11428 34672 11480 34678
rect 11428 34614 11480 34620
rect 11532 34524 11560 37402
rect 11624 36038 11652 41386
rect 11716 41386 11836 41414
rect 11612 36032 11664 36038
rect 11612 35974 11664 35980
rect 11612 35624 11664 35630
rect 11612 35566 11664 35572
rect 11624 35086 11652 35566
rect 11612 35080 11664 35086
rect 11612 35022 11664 35028
rect 11624 34649 11652 35022
rect 11716 34746 11744 41386
rect 11888 37868 11940 37874
rect 11888 37810 11940 37816
rect 11796 37120 11848 37126
rect 11796 37062 11848 37068
rect 11808 36582 11836 37062
rect 11796 36576 11848 36582
rect 11796 36518 11848 36524
rect 11900 36174 11928 37810
rect 11888 36168 11940 36174
rect 11888 36110 11940 36116
rect 11888 36032 11940 36038
rect 11888 35974 11940 35980
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11808 35154 11836 35566
rect 11900 35290 11928 35974
rect 11888 35284 11940 35290
rect 11888 35226 11940 35232
rect 11796 35148 11848 35154
rect 11796 35090 11848 35096
rect 11704 34740 11756 34746
rect 11704 34682 11756 34688
rect 11808 34649 11836 35090
rect 11610 34640 11666 34649
rect 11610 34575 11666 34584
rect 11794 34640 11850 34649
rect 11794 34575 11850 34584
rect 11440 34496 11560 34524
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 10839 30492 11147 30501
rect 10839 30490 10845 30492
rect 10901 30490 10925 30492
rect 10981 30490 11005 30492
rect 11061 30490 11085 30492
rect 11141 30490 11147 30492
rect 10901 30438 10903 30490
rect 11083 30438 11085 30490
rect 10839 30436 10845 30438
rect 10901 30436 10925 30438
rect 10981 30436 11005 30438
rect 11061 30436 11085 30438
rect 11141 30436 11147 30438
rect 10839 30427 11147 30436
rect 10876 30048 10928 30054
rect 10876 29990 10928 29996
rect 10888 29646 10916 29990
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 11244 29572 11296 29578
rect 11244 29514 11296 29520
rect 10839 29404 11147 29413
rect 10839 29402 10845 29404
rect 10901 29402 10925 29404
rect 10981 29402 11005 29404
rect 11061 29402 11085 29404
rect 11141 29402 11147 29404
rect 10901 29350 10903 29402
rect 11083 29350 11085 29402
rect 10839 29348 10845 29350
rect 10901 29348 10925 29350
rect 10981 29348 11005 29350
rect 11061 29348 11085 29350
rect 11141 29348 11147 29350
rect 10839 29339 11147 29348
rect 10692 29232 10744 29238
rect 10692 29174 10744 29180
rect 11256 29073 11284 29514
rect 11336 29232 11388 29238
rect 11336 29174 11388 29180
rect 11242 29064 11298 29073
rect 11242 28999 11298 29008
rect 11244 28960 11296 28966
rect 11244 28902 11296 28908
rect 10690 28520 10746 28529
rect 10690 28455 10746 28464
rect 10704 28422 10732 28455
rect 10692 28416 10744 28422
rect 10692 28358 10744 28364
rect 10839 28316 11147 28325
rect 10839 28314 10845 28316
rect 10901 28314 10925 28316
rect 10981 28314 11005 28316
rect 11061 28314 11085 28316
rect 11141 28314 11147 28316
rect 10901 28262 10903 28314
rect 11083 28262 11085 28314
rect 10839 28260 10845 28262
rect 10901 28260 10925 28262
rect 10981 28260 11005 28262
rect 11061 28260 11085 28262
rect 11141 28260 11147 28262
rect 10839 28251 11147 28260
rect 10784 28144 10836 28150
rect 10784 28086 10836 28092
rect 10876 28144 10928 28150
rect 10876 28086 10928 28092
rect 10796 27470 10824 28086
rect 10784 27464 10836 27470
rect 10784 27406 10836 27412
rect 10888 27316 10916 28086
rect 10704 27288 10916 27316
rect 10600 27124 10652 27130
rect 10600 27066 10652 27072
rect 10704 27062 10732 27288
rect 10839 27228 11147 27237
rect 10839 27226 10845 27228
rect 10901 27226 10925 27228
rect 10981 27226 11005 27228
rect 11061 27226 11085 27228
rect 11141 27226 11147 27228
rect 10901 27174 10903 27226
rect 11083 27174 11085 27226
rect 10839 27172 10845 27174
rect 10901 27172 10925 27174
rect 10981 27172 11005 27174
rect 11061 27172 11085 27174
rect 11141 27172 11147 27174
rect 10839 27163 11147 27172
rect 10692 27056 10744 27062
rect 10692 26998 10744 27004
rect 10966 27024 11022 27033
rect 10966 26959 11022 26968
rect 10980 26926 11008 26959
rect 10968 26920 11020 26926
rect 10520 26846 10732 26874
rect 10968 26862 11020 26868
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10520 25401 10548 26726
rect 10600 26308 10652 26314
rect 10600 26250 10652 26256
rect 10612 25786 10640 26250
rect 10704 25906 10732 26846
rect 10968 26784 11020 26790
rect 10968 26726 11020 26732
rect 11060 26784 11112 26790
rect 11060 26726 11112 26732
rect 10980 26382 11008 26726
rect 11072 26450 11100 26726
rect 11060 26444 11112 26450
rect 11060 26386 11112 26392
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10839 26140 11147 26149
rect 10839 26138 10845 26140
rect 10901 26138 10925 26140
rect 10981 26138 11005 26140
rect 11061 26138 11085 26140
rect 11141 26138 11147 26140
rect 10901 26086 10903 26138
rect 11083 26086 11085 26138
rect 10839 26084 10845 26086
rect 10901 26084 10925 26086
rect 10981 26084 11005 26086
rect 11061 26084 11085 26086
rect 11141 26084 11147 26086
rect 10839 26075 11147 26084
rect 11256 25974 11284 28902
rect 11244 25968 11296 25974
rect 11244 25910 11296 25916
rect 11348 25922 11376 29174
rect 11440 26217 11468 34496
rect 11992 34082 12020 43046
rect 12084 42838 12112 43862
rect 12176 43296 12204 44540
rect 12360 43314 12388 44540
rect 12440 43784 12492 43790
rect 12440 43726 12492 43732
rect 12256 43308 12308 43314
rect 12176 43268 12256 43296
rect 12256 43250 12308 43256
rect 12348 43308 12400 43314
rect 12348 43250 12400 43256
rect 12072 42832 12124 42838
rect 12072 42774 12124 42780
rect 12072 42696 12124 42702
rect 12072 42638 12124 42644
rect 12084 37330 12112 42638
rect 12256 42628 12308 42634
rect 12256 42570 12308 42576
rect 12162 42256 12218 42265
rect 12162 42191 12218 42200
rect 12176 42022 12204 42191
rect 12164 42016 12216 42022
rect 12164 41958 12216 41964
rect 12268 38350 12296 42570
rect 12348 42560 12400 42566
rect 12348 42502 12400 42508
rect 12360 42362 12388 42502
rect 12348 42356 12400 42362
rect 12348 42298 12400 42304
rect 12348 42220 12400 42226
rect 12348 42162 12400 42168
rect 12360 41993 12388 42162
rect 12346 41984 12402 41993
rect 12346 41919 12402 41928
rect 12452 41750 12480 43726
rect 12544 43602 12572 44540
rect 12544 43574 12664 43602
rect 12636 42770 12664 43574
rect 12728 43314 12756 44540
rect 12912 43382 12940 44540
rect 12900 43376 12952 43382
rect 12900 43318 12952 43324
rect 12716 43308 12768 43314
rect 12716 43250 12768 43256
rect 12716 43172 12768 43178
rect 12716 43114 12768 43120
rect 12624 42764 12676 42770
rect 12624 42706 12676 42712
rect 12532 42696 12584 42702
rect 12532 42638 12584 42644
rect 12440 41744 12492 41750
rect 12440 41686 12492 41692
rect 12348 41540 12400 41546
rect 12348 41482 12400 41488
rect 12256 38344 12308 38350
rect 12256 38286 12308 38292
rect 12164 38276 12216 38282
rect 12164 38218 12216 38224
rect 12072 37324 12124 37330
rect 12072 37266 12124 37272
rect 12072 37120 12124 37126
rect 12072 37062 12124 37068
rect 12084 35630 12112 37062
rect 12176 35873 12204 38218
rect 12360 36310 12388 41482
rect 12438 41032 12494 41041
rect 12438 40967 12494 40976
rect 12452 40390 12480 40967
rect 12440 40384 12492 40390
rect 12440 40326 12492 40332
rect 12452 38962 12480 40326
rect 12440 38956 12492 38962
rect 12440 38898 12492 38904
rect 12438 38312 12494 38321
rect 12438 38247 12440 38256
rect 12492 38247 12494 38256
rect 12440 38218 12492 38224
rect 12452 37913 12480 38218
rect 12438 37904 12494 37913
rect 12438 37839 12494 37848
rect 12544 37274 12572 42638
rect 12624 42560 12676 42566
rect 12624 42502 12676 42508
rect 12636 41818 12664 42502
rect 12624 41812 12676 41818
rect 12624 41754 12676 41760
rect 12728 41414 12756 43114
rect 12992 43104 13044 43110
rect 12992 43046 13044 43052
rect 12900 42900 12952 42906
rect 12900 42842 12952 42848
rect 12808 42696 12860 42702
rect 12808 42638 12860 42644
rect 12820 42129 12848 42638
rect 12806 42120 12862 42129
rect 12806 42055 12862 42064
rect 12808 41540 12860 41546
rect 12808 41482 12860 41488
rect 12636 41386 12756 41414
rect 12636 39506 12664 41386
rect 12820 41120 12848 41482
rect 12728 41092 12848 41120
rect 12624 39500 12676 39506
rect 12624 39442 12676 39448
rect 12728 37913 12756 41092
rect 12808 40996 12860 41002
rect 12808 40938 12860 40944
rect 12820 40050 12848 40938
rect 12808 40044 12860 40050
rect 12808 39986 12860 39992
rect 12912 38654 12940 42842
rect 12820 38626 12940 38654
rect 12714 37904 12770 37913
rect 12714 37839 12770 37848
rect 12544 37246 12664 37274
rect 12438 36816 12494 36825
rect 12438 36751 12494 36760
rect 12348 36304 12400 36310
rect 12452 36281 12480 36751
rect 12348 36246 12400 36252
rect 12438 36272 12494 36281
rect 12438 36207 12494 36216
rect 12162 35864 12218 35873
rect 12162 35799 12218 35808
rect 12162 35728 12218 35737
rect 12162 35663 12218 35672
rect 12072 35624 12124 35630
rect 12072 35566 12124 35572
rect 12072 35216 12124 35222
rect 12072 35158 12124 35164
rect 11532 34054 12020 34082
rect 11532 27674 11560 34054
rect 11612 33924 11664 33930
rect 11612 33866 11664 33872
rect 11624 32434 11652 33866
rect 11796 33856 11848 33862
rect 11796 33798 11848 33804
rect 11808 33046 11836 33798
rect 12084 33590 12112 35158
rect 12176 34610 12204 35663
rect 12256 35284 12308 35290
rect 12256 35226 12308 35232
rect 12268 35068 12296 35226
rect 12440 35080 12492 35086
rect 12268 35040 12440 35068
rect 12440 35022 12492 35028
rect 12532 35080 12584 35086
rect 12532 35022 12584 35028
rect 12544 34921 12572 35022
rect 12254 34912 12310 34921
rect 12254 34847 12310 34856
rect 12530 34912 12586 34921
rect 12530 34847 12586 34856
rect 12164 34604 12216 34610
rect 12164 34546 12216 34552
rect 12176 33930 12204 34546
rect 12268 34406 12296 34847
rect 12532 34672 12584 34678
rect 12532 34614 12584 34620
rect 12256 34400 12308 34406
rect 12256 34342 12308 34348
rect 12544 34066 12572 34614
rect 12532 34060 12584 34066
rect 12532 34002 12584 34008
rect 12636 33946 12664 37246
rect 12716 36576 12768 36582
rect 12716 36518 12768 36524
rect 12728 35698 12756 36518
rect 12716 35692 12768 35698
rect 12716 35634 12768 35640
rect 12820 35494 12848 38626
rect 13004 38185 13032 43046
rect 13096 42684 13124 44540
rect 13280 43450 13308 44540
rect 13464 44010 13492 44540
rect 13464 43982 13584 44010
rect 13556 43926 13584 43982
rect 13544 43920 13596 43926
rect 13544 43862 13596 43868
rect 13648 43654 13676 44540
rect 13832 43897 13860 44540
rect 13818 43888 13874 43897
rect 13818 43823 13874 43832
rect 13820 43716 13872 43722
rect 13820 43658 13872 43664
rect 13636 43648 13688 43654
rect 13636 43590 13688 43596
rect 13268 43444 13320 43450
rect 13268 43386 13320 43392
rect 13542 43208 13598 43217
rect 13542 43143 13598 43152
rect 13636 43172 13688 43178
rect 13556 43110 13584 43143
rect 13636 43114 13688 43120
rect 13544 43104 13596 43110
rect 13544 43046 13596 43052
rect 13312 43004 13620 43013
rect 13312 43002 13318 43004
rect 13374 43002 13398 43004
rect 13454 43002 13478 43004
rect 13534 43002 13558 43004
rect 13614 43002 13620 43004
rect 13374 42950 13376 43002
rect 13556 42950 13558 43002
rect 13312 42948 13318 42950
rect 13374 42948 13398 42950
rect 13454 42948 13478 42950
rect 13534 42948 13558 42950
rect 13614 42948 13620 42950
rect 13312 42939 13620 42948
rect 13452 42832 13504 42838
rect 13452 42774 13504 42780
rect 13176 42696 13228 42702
rect 13096 42656 13176 42684
rect 13176 42638 13228 42644
rect 13464 42362 13492 42774
rect 13648 42702 13676 43114
rect 13728 43104 13780 43110
rect 13728 43046 13780 43052
rect 13636 42696 13688 42702
rect 13636 42638 13688 42644
rect 13544 42560 13596 42566
rect 13544 42502 13596 42508
rect 13556 42362 13584 42502
rect 13740 42362 13768 43046
rect 13452 42356 13504 42362
rect 13452 42298 13504 42304
rect 13544 42356 13596 42362
rect 13544 42298 13596 42304
rect 13728 42356 13780 42362
rect 13728 42298 13780 42304
rect 13832 42242 13860 43658
rect 13910 43344 13966 43353
rect 13910 43279 13966 43288
rect 13648 42214 13860 42242
rect 13648 42158 13676 42214
rect 13636 42152 13688 42158
rect 13096 42078 13308 42106
rect 13924 42106 13952 43279
rect 14016 42809 14044 44540
rect 14200 44033 14228 44540
rect 14186 44024 14242 44033
rect 14186 43959 14242 43968
rect 14188 43648 14240 43654
rect 14188 43590 14240 43596
rect 14200 43382 14228 43590
rect 14384 43466 14412 44540
rect 14384 43450 14504 43466
rect 14384 43444 14516 43450
rect 14384 43438 14464 43444
rect 14464 43386 14516 43392
rect 14188 43376 14240 43382
rect 14188 43318 14240 43324
rect 14280 43104 14332 43110
rect 14280 43046 14332 43052
rect 14464 43104 14516 43110
rect 14464 43046 14516 43052
rect 14186 42936 14242 42945
rect 14108 42894 14186 42922
rect 14002 42800 14058 42809
rect 14002 42735 14058 42744
rect 14004 42560 14056 42566
rect 14004 42502 14056 42508
rect 13636 42094 13688 42100
rect 13096 41562 13124 42078
rect 13280 42022 13308 42078
rect 13832 42078 13952 42106
rect 13176 42016 13228 42022
rect 13176 41958 13228 41964
rect 13268 42016 13320 42022
rect 13268 41958 13320 41964
rect 13188 41721 13216 41958
rect 13312 41916 13620 41925
rect 13312 41914 13318 41916
rect 13374 41914 13398 41916
rect 13454 41914 13478 41916
rect 13534 41914 13558 41916
rect 13614 41914 13620 41916
rect 13374 41862 13376 41914
rect 13556 41862 13558 41914
rect 13312 41860 13318 41862
rect 13374 41860 13398 41862
rect 13454 41860 13478 41862
rect 13534 41860 13558 41862
rect 13614 41860 13620 41862
rect 13312 41851 13620 41860
rect 13832 41750 13860 42078
rect 13912 42016 13964 42022
rect 13912 41958 13964 41964
rect 13820 41744 13872 41750
rect 13174 41712 13230 41721
rect 13174 41647 13230 41656
rect 13556 41670 13768 41698
rect 13820 41686 13872 41692
rect 13556 41614 13584 41670
rect 13544 41608 13596 41614
rect 13096 41534 13216 41562
rect 13544 41550 13596 41556
rect 13636 41608 13688 41614
rect 13636 41550 13688 41556
rect 13084 40724 13136 40730
rect 13084 40666 13136 40672
rect 13096 39137 13124 40666
rect 13082 39128 13138 39137
rect 13082 39063 13138 39072
rect 13084 38956 13136 38962
rect 13084 38898 13136 38904
rect 12990 38176 13046 38185
rect 12990 38111 13046 38120
rect 12992 37664 13044 37670
rect 12992 37606 13044 37612
rect 12900 36576 12952 36582
rect 12900 36518 12952 36524
rect 12808 35488 12860 35494
rect 12808 35430 12860 35436
rect 12716 35080 12768 35086
rect 12716 35022 12768 35028
rect 12726 35006 12756 35022
rect 12728 34746 12756 35006
rect 12806 34776 12862 34785
rect 12716 34740 12768 34746
rect 12806 34711 12862 34720
rect 12716 34682 12768 34688
rect 12716 34400 12768 34406
rect 12716 34342 12768 34348
rect 12164 33924 12216 33930
rect 12164 33866 12216 33872
rect 12544 33918 12664 33946
rect 12072 33584 12124 33590
rect 12072 33526 12124 33532
rect 12348 33312 12400 33318
rect 12348 33254 12400 33260
rect 11796 33040 11848 33046
rect 11978 33008 12034 33017
rect 11796 32982 11848 32988
rect 11704 32972 11756 32978
rect 11704 32914 11756 32920
rect 11900 32966 11978 32994
rect 11612 32428 11664 32434
rect 11612 32370 11664 32376
rect 11612 31816 11664 31822
rect 11716 31804 11744 32914
rect 11664 31776 11744 31804
rect 11612 31758 11664 31764
rect 11612 30388 11664 30394
rect 11612 30330 11664 30336
rect 11624 29510 11652 30330
rect 11716 30161 11744 31776
rect 11796 31680 11848 31686
rect 11796 31622 11848 31628
rect 11808 31482 11836 31622
rect 11796 31476 11848 31482
rect 11796 31418 11848 31424
rect 11796 31340 11848 31346
rect 11796 31282 11848 31288
rect 11808 31249 11836 31282
rect 11794 31240 11850 31249
rect 11794 31175 11850 31184
rect 11900 30802 11928 32966
rect 12360 32978 12388 33254
rect 12544 33114 12572 33918
rect 12624 33856 12676 33862
rect 12624 33798 12676 33804
rect 12440 33108 12492 33114
rect 12440 33050 12492 33056
rect 12532 33108 12584 33114
rect 12532 33050 12584 33056
rect 11978 32943 12034 32952
rect 12348 32972 12400 32978
rect 12452 32960 12480 33050
rect 12532 32972 12584 32978
rect 12452 32932 12532 32960
rect 12348 32914 12400 32920
rect 12532 32914 12584 32920
rect 12164 32904 12216 32910
rect 12084 32852 12164 32858
rect 12084 32846 12216 32852
rect 12084 32830 12204 32846
rect 11980 32224 12032 32230
rect 11980 32166 12032 32172
rect 11992 31754 12020 32166
rect 12084 31929 12112 32830
rect 12440 32768 12492 32774
rect 12440 32710 12492 32716
rect 12164 32224 12216 32230
rect 12164 32166 12216 32172
rect 12070 31920 12126 31929
rect 12070 31855 12126 31864
rect 11980 31748 12032 31754
rect 11980 31690 12032 31696
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 11888 30660 11940 30666
rect 11888 30602 11940 30608
rect 11796 30592 11848 30598
rect 11796 30534 11848 30540
rect 11702 30152 11758 30161
rect 11702 30087 11758 30096
rect 11702 29744 11758 29753
rect 11702 29679 11704 29688
rect 11756 29679 11758 29688
rect 11704 29650 11756 29656
rect 11808 29646 11836 30534
rect 11796 29640 11848 29646
rect 11796 29582 11848 29588
rect 11612 29504 11664 29510
rect 11612 29446 11664 29452
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11716 29306 11744 29446
rect 11704 29300 11756 29306
rect 11704 29242 11756 29248
rect 11900 28994 11928 30602
rect 11992 30394 12020 31690
rect 12084 31482 12112 31855
rect 12176 31482 12204 32166
rect 12452 31686 12480 32710
rect 12532 31816 12584 31822
rect 12532 31758 12584 31764
rect 12440 31680 12492 31686
rect 12440 31622 12492 31628
rect 12072 31476 12124 31482
rect 12072 31418 12124 31424
rect 12164 31476 12216 31482
rect 12164 31418 12216 31424
rect 11980 30388 12032 30394
rect 11980 30330 12032 30336
rect 11980 30252 12032 30258
rect 11980 30194 12032 30200
rect 11808 28966 11928 28994
rect 11612 28960 11664 28966
rect 11612 28902 11664 28908
rect 11624 28540 11652 28902
rect 11808 28665 11836 28966
rect 11794 28656 11850 28665
rect 11794 28591 11850 28600
rect 11704 28552 11756 28558
rect 11624 28512 11704 28540
rect 11704 28494 11756 28500
rect 11888 28552 11940 28558
rect 11888 28494 11940 28500
rect 11612 28416 11664 28422
rect 11612 28358 11664 28364
rect 11624 28150 11652 28358
rect 11716 28150 11744 28494
rect 11612 28144 11664 28150
rect 11612 28086 11664 28092
rect 11704 28144 11756 28150
rect 11704 28086 11756 28092
rect 11794 28112 11850 28121
rect 11794 28047 11850 28056
rect 11612 28008 11664 28014
rect 11612 27950 11664 27956
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11520 27668 11572 27674
rect 11520 27610 11572 27616
rect 11520 27464 11572 27470
rect 11520 27406 11572 27412
rect 11426 26208 11482 26217
rect 11426 26143 11482 26152
rect 11532 26042 11560 27406
rect 11624 26246 11652 27950
rect 11716 26314 11744 27950
rect 11806 27928 11834 28047
rect 11900 27928 11928 28494
rect 11992 28422 12020 30194
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11806 27900 11836 27928
rect 11900 27900 12020 27928
rect 11808 27826 11836 27900
rect 11808 27798 11928 27826
rect 11794 26752 11850 26761
rect 11794 26687 11850 26696
rect 11808 26382 11836 26687
rect 11796 26376 11848 26382
rect 11796 26318 11848 26324
rect 11704 26308 11756 26314
rect 11704 26250 11756 26256
rect 11900 26246 11928 27798
rect 11992 27334 12020 27900
rect 12084 27554 12112 31418
rect 12452 31414 12480 31622
rect 12544 31482 12572 31758
rect 12532 31476 12584 31482
rect 12532 31418 12584 31424
rect 12348 31408 12400 31414
rect 12348 31350 12400 31356
rect 12440 31408 12492 31414
rect 12440 31350 12492 31356
rect 12256 30796 12308 30802
rect 12256 30738 12308 30744
rect 12268 29306 12296 30738
rect 12360 30734 12388 31350
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 12348 30728 12400 30734
rect 12348 30670 12400 30676
rect 12438 30560 12494 30569
rect 12438 30495 12494 30504
rect 12452 29594 12480 30495
rect 12360 29566 12480 29594
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12162 29064 12218 29073
rect 12162 28999 12218 29008
rect 12256 29028 12308 29034
rect 12176 27860 12204 28999
rect 12256 28970 12308 28976
rect 12268 28014 12296 28970
rect 12256 28008 12308 28014
rect 12256 27950 12308 27956
rect 12176 27832 12296 27860
rect 12268 27674 12296 27832
rect 12360 27713 12388 29566
rect 12440 29504 12492 29510
rect 12440 29446 12492 29452
rect 12452 28393 12480 29446
rect 12438 28384 12494 28393
rect 12438 28319 12494 28328
rect 12440 28008 12492 28014
rect 12544 27996 12572 31282
rect 12492 27968 12572 27996
rect 12440 27950 12492 27956
rect 12346 27704 12402 27713
rect 12256 27668 12308 27674
rect 12346 27639 12402 27648
rect 12256 27610 12308 27616
rect 12084 27526 12388 27554
rect 12072 27464 12124 27470
rect 12072 27406 12124 27412
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 12084 27062 12112 27406
rect 12256 27396 12308 27402
rect 12256 27338 12308 27344
rect 12164 27328 12216 27334
rect 12164 27270 12216 27276
rect 12072 27056 12124 27062
rect 12072 26998 12124 27004
rect 12176 26738 12204 27270
rect 12268 26858 12296 27338
rect 12360 27033 12388 27526
rect 12346 27024 12402 27033
rect 12346 26959 12402 26968
rect 12452 26926 12480 27950
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12440 26920 12492 26926
rect 12440 26862 12492 26868
rect 12256 26852 12308 26858
rect 12256 26794 12308 26800
rect 12348 26784 12400 26790
rect 12346 26752 12348 26761
rect 12400 26752 12402 26761
rect 12176 26710 12296 26738
rect 12162 26616 12218 26625
rect 12162 26551 12218 26560
rect 11980 26512 12032 26518
rect 11980 26454 12032 26460
rect 11992 26353 12020 26454
rect 11978 26344 12034 26353
rect 11978 26279 12034 26288
rect 11612 26240 11664 26246
rect 11612 26182 11664 26188
rect 11888 26240 11940 26246
rect 11888 26182 11940 26188
rect 11980 26240 12032 26246
rect 11980 26182 12032 26188
rect 11520 26036 11572 26042
rect 11624 26024 11652 26182
rect 11624 25996 11744 26024
rect 11520 25978 11572 25984
rect 10692 25900 10744 25906
rect 11348 25894 11652 25922
rect 10692 25842 10744 25848
rect 11334 25800 11390 25809
rect 10612 25758 10824 25786
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 10692 25696 10744 25702
rect 10692 25638 10744 25644
rect 10506 25392 10562 25401
rect 10506 25327 10562 25336
rect 10612 25158 10640 25638
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10416 24948 10468 24954
rect 10416 24890 10468 24896
rect 10600 24948 10652 24954
rect 10600 24890 10652 24896
rect 10508 24880 10560 24886
rect 10414 24848 10470 24857
rect 10324 24812 10376 24818
rect 10508 24822 10560 24828
rect 10414 24783 10470 24792
rect 10324 24754 10376 24760
rect 10324 24676 10376 24682
rect 10324 24618 10376 24624
rect 10336 24206 10364 24618
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10010 23854 10086 23882
rect 9954 23831 10010 23840
rect 9772 23792 9824 23798
rect 9772 23734 9824 23740
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 9784 23497 9812 23734
rect 9770 23488 9826 23497
rect 9770 23423 9826 23432
rect 9968 23322 9996 23734
rect 10058 23662 10086 23854
rect 10152 23854 10272 23882
rect 10048 23656 10100 23662
rect 10048 23598 10100 23604
rect 9956 23316 10008 23322
rect 9956 23258 10008 23264
rect 10152 23168 10180 23854
rect 10322 23352 10378 23361
rect 10322 23287 10378 23296
rect 9968 23140 10180 23168
rect 9772 22772 9824 22778
rect 9772 22714 9824 22720
rect 9784 22030 9812 22714
rect 9862 22672 9918 22681
rect 9862 22607 9918 22616
rect 9772 22024 9824 22030
rect 9772 21966 9824 21972
rect 9770 21856 9826 21865
rect 9770 21791 9826 21800
rect 9680 19440 9732 19446
rect 9680 19382 9732 19388
rect 9692 18952 9720 19382
rect 9784 19145 9812 21791
rect 9770 19136 9826 19145
rect 9770 19071 9826 19080
rect 9692 18924 9812 18952
rect 9680 18828 9732 18834
rect 9680 18770 9732 18776
rect 9692 18426 9720 18770
rect 9784 18698 9812 18924
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9588 18284 9640 18290
rect 9588 18226 9640 18232
rect 9496 18148 9548 18154
rect 9496 18090 9548 18096
rect 9508 17921 9536 18090
rect 9494 17912 9550 17921
rect 9494 17847 9550 17856
rect 9324 17700 9444 17728
rect 9220 17128 9272 17134
rect 9324 17105 9352 17700
rect 9680 17672 9732 17678
rect 9586 17640 9642 17649
rect 9404 17604 9456 17610
rect 9404 17546 9456 17552
rect 9508 17598 9586 17626
rect 9416 17338 9444 17546
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9220 17070 9272 17076
rect 9310 17096 9366 17105
rect 9310 17031 9366 17040
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9218 16824 9274 16833
rect 9218 16759 9274 16768
rect 9126 15736 9182 15745
rect 9126 15671 9182 15680
rect 9140 15065 9168 15671
rect 9126 15056 9182 15065
rect 9126 14991 9182 15000
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 9036 13864 9088 13870
rect 9034 13832 9036 13841
rect 9088 13832 9090 13841
rect 9140 13802 9168 14758
rect 9034 13767 9090 13776
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9232 13682 9260 16759
rect 9324 15881 9352 16934
rect 9404 15972 9456 15978
rect 9404 15914 9456 15920
rect 9310 15872 9366 15881
rect 9310 15807 9366 15816
rect 9310 15736 9366 15745
rect 9310 15671 9366 15680
rect 9324 15502 9352 15671
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9416 14550 9444 15914
rect 9404 14544 9456 14550
rect 9404 14486 9456 14492
rect 9508 14090 9536 17598
rect 9680 17614 9732 17620
rect 9586 17575 9642 17584
rect 9692 17202 9720 17614
rect 9772 17332 9824 17338
rect 9772 17274 9824 17280
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9784 17116 9812 17274
rect 9876 17241 9904 22607
rect 9968 21486 9996 23140
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10140 22704 10192 22710
rect 10140 22646 10192 22652
rect 10152 21962 10180 22646
rect 10244 22522 10272 22714
rect 10336 22642 10364 23287
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10244 22494 10364 22522
rect 10230 21992 10286 22001
rect 10140 21956 10192 21962
rect 10230 21927 10232 21936
rect 10140 21898 10192 21904
rect 10284 21927 10286 21936
rect 10232 21898 10284 21904
rect 9956 21480 10008 21486
rect 9956 21422 10008 21428
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 10138 21448 10194 21457
rect 9956 21344 10008 21350
rect 9956 21286 10008 21292
rect 9968 20641 9996 21286
rect 9954 20632 10010 20641
rect 9954 20567 10010 20576
rect 9956 20256 10008 20262
rect 9956 20198 10008 20204
rect 9968 19310 9996 20198
rect 10060 19854 10088 21422
rect 10138 21383 10194 21392
rect 10152 20924 10180 21383
rect 10244 21049 10272 21898
rect 10230 21040 10286 21049
rect 10230 20975 10286 20984
rect 10152 20896 10272 20924
rect 10138 20768 10194 20777
rect 10138 20703 10194 20712
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10060 19718 10088 19790
rect 10048 19712 10100 19718
rect 10048 19654 10100 19660
rect 9956 19304 10008 19310
rect 9956 19246 10008 19252
rect 9954 19136 10010 19145
rect 9954 19071 10010 19080
rect 9968 18222 9996 19071
rect 10060 18873 10088 19654
rect 10046 18864 10102 18873
rect 10046 18799 10102 18808
rect 10048 18692 10100 18698
rect 10048 18634 10100 18640
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 9956 18080 10008 18086
rect 9956 18022 10008 18028
rect 9968 17270 9996 18022
rect 10060 17610 10088 18634
rect 10048 17604 10100 17610
rect 10048 17546 10100 17552
rect 9956 17264 10008 17270
rect 9862 17232 9918 17241
rect 9956 17206 10008 17212
rect 9862 17167 9918 17176
rect 9784 17088 9904 17116
rect 9770 16960 9826 16969
rect 9770 16895 9826 16904
rect 9784 16674 9812 16895
rect 9876 16833 9904 17088
rect 9954 17096 10010 17105
rect 9954 17031 10010 17040
rect 9862 16824 9918 16833
rect 9968 16794 9996 17031
rect 9862 16759 9918 16768
rect 9956 16788 10008 16794
rect 9956 16730 10008 16736
rect 9692 16646 9812 16674
rect 9692 16289 9720 16646
rect 10060 16522 10088 17546
rect 10152 17377 10180 20703
rect 10244 19825 10272 20896
rect 10230 19816 10286 19825
rect 10230 19751 10286 19760
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10244 19514 10272 19654
rect 10232 19508 10284 19514
rect 10232 19450 10284 19456
rect 10232 18692 10284 18698
rect 10232 18634 10284 18640
rect 10244 17678 10272 18634
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10138 17368 10194 17377
rect 10138 17303 10194 17312
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 9864 16516 9916 16522
rect 9864 16458 9916 16464
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 9772 16448 9824 16454
rect 9772 16390 9824 16396
rect 9678 16280 9734 16289
rect 9678 16215 9734 16224
rect 9784 16114 9812 16390
rect 9772 16108 9824 16114
rect 9772 16050 9824 16056
rect 9876 15994 9904 16458
rect 10060 16250 10088 16458
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10152 16130 10180 16594
rect 10244 16522 10272 17614
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 9784 15966 9904 15994
rect 9968 16102 10180 16130
rect 9588 15428 9640 15434
rect 9588 15370 9640 15376
rect 9600 15337 9628 15370
rect 9586 15328 9642 15337
rect 9586 15263 9642 15272
rect 9680 14408 9732 14414
rect 9048 13654 9260 13682
rect 9324 14062 9536 14090
rect 9600 14356 9680 14362
rect 9600 14350 9732 14356
rect 9600 14334 9720 14350
rect 9048 11762 9076 13654
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9140 10554 9168 13262
rect 9232 12306 9260 13398
rect 9324 12918 9352 14062
rect 9496 14000 9548 14006
rect 9496 13942 9548 13948
rect 9404 13796 9456 13802
rect 9404 13738 9456 13744
rect 9416 13462 9444 13738
rect 9404 13456 9456 13462
rect 9404 13398 9456 13404
rect 9404 13252 9456 13258
rect 9404 13194 9456 13200
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9220 12300 9272 12306
rect 9324 12288 9352 12854
rect 9416 12442 9444 13194
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9324 12260 9444 12288
rect 9220 12242 9272 12248
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 9232 11257 9260 11698
rect 9218 11248 9274 11257
rect 9218 11183 9274 11192
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9048 10526 9168 10554
rect 9048 7410 9076 10526
rect 9126 10432 9182 10441
rect 9126 10367 9182 10376
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 5545 9076 7142
rect 9034 5536 9090 5545
rect 9034 5471 9090 5480
rect 9048 5234 9076 5471
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 9048 3369 9076 3878
rect 9140 3534 9168 10367
rect 9232 8090 9260 11086
rect 9324 10742 9352 12106
rect 9416 11830 9444 12260
rect 9404 11824 9456 11830
rect 9404 11766 9456 11772
rect 9404 11144 9456 11150
rect 9508 11132 9536 13942
rect 9600 13530 9628 14334
rect 9678 13832 9734 13841
rect 9678 13767 9734 13776
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9586 13424 9642 13433
rect 9586 13359 9642 13368
rect 9600 12442 9628 13359
rect 9692 13326 9720 13767
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9600 11218 9628 12378
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9456 11104 9536 11132
rect 9404 11086 9456 11092
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 10266 9352 10542
rect 9312 10260 9364 10266
rect 9312 10202 9364 10208
rect 9324 9654 9352 10202
rect 9416 10198 9444 10950
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 9416 9518 9444 9862
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9324 8430 9352 9386
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9416 8634 9444 8842
rect 9508 8634 9536 10950
rect 9692 10146 9720 13262
rect 9784 11801 9812 15966
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 9876 14890 9904 15846
rect 9968 15706 9996 16102
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10048 15904 10100 15910
rect 10048 15846 10100 15852
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9954 15328 10010 15337
rect 9954 15263 10010 15272
rect 9864 14884 9916 14890
rect 9864 14826 9916 14832
rect 9864 14544 9916 14550
rect 9862 14512 9864 14521
rect 9916 14512 9918 14521
rect 9862 14447 9918 14456
rect 9968 14226 9996 15263
rect 9876 14198 9996 14226
rect 9876 13938 9904 14198
rect 9954 14104 10010 14113
rect 9954 14039 10010 14048
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9876 12374 9904 13874
rect 9864 12368 9916 12374
rect 9864 12310 9916 12316
rect 9864 12096 9916 12102
rect 9864 12038 9916 12044
rect 9770 11792 9826 11801
rect 9770 11727 9826 11736
rect 9876 11676 9904 12038
rect 9784 11648 9904 11676
rect 9784 10554 9812 11648
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9876 10674 9904 11290
rect 9864 10668 9916 10674
rect 9864 10610 9916 10616
rect 9784 10526 9904 10554
rect 9772 10464 9824 10470
rect 9772 10406 9824 10412
rect 9784 10266 9812 10406
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9770 10160 9826 10169
rect 9600 10130 9770 10146
rect 9588 10124 9770 10130
rect 9640 10118 9770 10124
rect 9770 10095 9826 10104
rect 9588 10066 9640 10072
rect 9600 9654 9628 10066
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9772 10056 9824 10062
rect 9772 9998 9824 10004
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9692 9042 9720 9998
rect 9784 9926 9812 9998
rect 9772 9920 9824 9926
rect 9772 9862 9824 9868
rect 9784 9518 9812 9862
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 9772 9036 9824 9042
rect 9772 8978 9824 8984
rect 9784 8922 9812 8978
rect 9692 8894 9812 8922
rect 9876 8906 9904 10526
rect 9968 10130 9996 14039
rect 10060 12424 10088 15846
rect 10152 15706 10180 15982
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10140 15564 10192 15570
rect 10140 15506 10192 15512
rect 10152 13920 10180 15506
rect 10336 15194 10364 22494
rect 10428 21865 10456 24783
rect 10520 24274 10548 24822
rect 10508 24268 10560 24274
rect 10508 24210 10560 24216
rect 10508 24132 10560 24138
rect 10508 24074 10560 24080
rect 10520 23050 10548 24074
rect 10508 23044 10560 23050
rect 10508 22986 10560 22992
rect 10612 22930 10640 24890
rect 10520 22902 10640 22930
rect 10520 22778 10548 22902
rect 10598 22808 10654 22817
rect 10508 22772 10560 22778
rect 10598 22743 10654 22752
rect 10508 22714 10560 22720
rect 10508 22432 10560 22438
rect 10508 22374 10560 22380
rect 10520 22273 10548 22374
rect 10506 22264 10562 22273
rect 10506 22199 10562 22208
rect 10508 22024 10560 22030
rect 10508 21966 10560 21972
rect 10414 21856 10470 21865
rect 10414 21791 10470 21800
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10428 19281 10456 21626
rect 10520 21078 10548 21966
rect 10508 21072 10560 21078
rect 10508 21014 10560 21020
rect 10520 19553 10548 21014
rect 10612 21010 10640 22743
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10600 20392 10652 20398
rect 10600 20334 10652 20340
rect 10612 19854 10640 20334
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10600 19712 10652 19718
rect 10600 19654 10652 19660
rect 10506 19544 10562 19553
rect 10506 19479 10562 19488
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10414 19272 10470 19281
rect 10414 19207 10470 19216
rect 10520 18873 10548 19314
rect 10506 18864 10562 18873
rect 10506 18799 10562 18808
rect 10416 18692 10468 18698
rect 10416 18634 10468 18640
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 10428 18426 10456 18634
rect 10416 18420 10468 18426
rect 10416 18362 10468 18368
rect 10520 18086 10548 18634
rect 10612 18272 10640 19654
rect 10704 19281 10732 25638
rect 10796 25294 10824 25758
rect 11334 25735 11390 25744
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 11244 25220 11296 25226
rect 11244 25162 11296 25168
rect 10839 25052 11147 25061
rect 10839 25050 10845 25052
rect 10901 25050 10925 25052
rect 10981 25050 11005 25052
rect 11061 25050 11085 25052
rect 11141 25050 11147 25052
rect 10901 24998 10903 25050
rect 11083 24998 11085 25050
rect 10839 24996 10845 24998
rect 10901 24996 10925 24998
rect 10981 24996 11005 24998
rect 11061 24996 11085 24998
rect 11141 24996 11147 24998
rect 10839 24987 11147 24996
rect 11058 24848 11114 24857
rect 10784 24812 10836 24818
rect 11058 24783 11114 24792
rect 10784 24754 10836 24760
rect 10796 24410 10824 24754
rect 10784 24404 10836 24410
rect 10784 24346 10836 24352
rect 11072 24313 11100 24783
rect 11058 24304 11114 24313
rect 10784 24268 10836 24274
rect 11058 24239 11114 24248
rect 10784 24210 10836 24216
rect 10796 24052 10824 24210
rect 10876 24064 10928 24070
rect 10796 24024 10876 24052
rect 10876 24006 10928 24012
rect 10839 23964 11147 23973
rect 10839 23962 10845 23964
rect 10901 23962 10925 23964
rect 10981 23962 11005 23964
rect 11061 23962 11085 23964
rect 11141 23962 11147 23964
rect 10901 23910 10903 23962
rect 11083 23910 11085 23962
rect 10839 23908 10845 23910
rect 10901 23908 10925 23910
rect 10981 23908 11005 23910
rect 11061 23908 11085 23910
rect 11141 23908 11147 23910
rect 10839 23899 11147 23908
rect 11256 23866 11284 25162
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11256 23594 11284 23802
rect 11244 23588 11296 23594
rect 11244 23530 11296 23536
rect 10784 23520 10836 23526
rect 10784 23462 10836 23468
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 11242 23488 11298 23497
rect 10796 23089 10824 23462
rect 10782 23080 10838 23089
rect 11164 23050 11192 23462
rect 11242 23423 11298 23432
rect 10782 23015 10838 23024
rect 11152 23044 11204 23050
rect 11204 22992 11217 23032
rect 11152 22986 11217 22992
rect 10839 22876 11147 22885
rect 10839 22874 10845 22876
rect 10901 22874 10925 22876
rect 10981 22874 11005 22876
rect 11061 22874 11085 22876
rect 11141 22874 11147 22876
rect 10901 22822 10903 22874
rect 11083 22822 11085 22874
rect 10839 22820 10845 22822
rect 10901 22820 10925 22822
rect 10981 22820 11005 22822
rect 11061 22820 11085 22822
rect 11141 22820 11147 22822
rect 10839 22811 11147 22820
rect 11189 22760 11217 22986
rect 11164 22732 11217 22760
rect 11164 22574 11192 22732
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11060 22432 11112 22438
rect 11060 22374 11112 22380
rect 11072 22094 11100 22374
rect 11072 22066 11192 22094
rect 11164 22030 11192 22066
rect 11152 22024 11204 22030
rect 11152 21966 11204 21972
rect 10839 21788 11147 21797
rect 10839 21786 10845 21788
rect 10901 21786 10925 21788
rect 10981 21786 11005 21788
rect 11061 21786 11085 21788
rect 11141 21786 11147 21788
rect 10901 21734 10903 21786
rect 11083 21734 11085 21786
rect 10839 21732 10845 21734
rect 10901 21732 10925 21734
rect 10981 21732 11005 21734
rect 11061 21732 11085 21734
rect 11141 21732 11147 21734
rect 10839 21723 11147 21732
rect 11060 20936 11112 20942
rect 10980 20884 11060 20890
rect 10980 20878 11112 20884
rect 10980 20862 11100 20878
rect 10980 20806 11008 20862
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10839 20700 11147 20709
rect 10839 20698 10845 20700
rect 10901 20698 10925 20700
rect 10981 20698 11005 20700
rect 11061 20698 11085 20700
rect 11141 20698 11147 20700
rect 10901 20646 10903 20698
rect 11083 20646 11085 20698
rect 10839 20644 10845 20646
rect 10901 20644 10925 20646
rect 10981 20644 11005 20646
rect 11061 20644 11085 20646
rect 11141 20644 11147 20646
rect 10839 20635 11147 20644
rect 10876 20528 10928 20534
rect 10876 20470 10928 20476
rect 10784 20460 10836 20466
rect 10784 20402 10836 20408
rect 10796 19854 10824 20402
rect 10784 19848 10836 19854
rect 10888 19825 10916 20470
rect 10784 19790 10836 19796
rect 10874 19816 10930 19825
rect 10874 19751 10930 19760
rect 10839 19612 11147 19621
rect 10839 19610 10845 19612
rect 10901 19610 10925 19612
rect 10981 19610 11005 19612
rect 11061 19610 11085 19612
rect 11141 19610 11147 19612
rect 10901 19558 10903 19610
rect 11083 19558 11085 19610
rect 10839 19556 10845 19558
rect 10901 19556 10925 19558
rect 10981 19556 11005 19558
rect 11061 19556 11085 19558
rect 11141 19556 11147 19558
rect 10839 19547 11147 19556
rect 11256 19496 11284 23423
rect 11348 22642 11376 25735
rect 11518 25528 11574 25537
rect 11518 25463 11574 25472
rect 11428 25356 11480 25362
rect 11428 25298 11480 25304
rect 11440 24954 11468 25298
rect 11428 24948 11480 24954
rect 11428 24890 11480 24896
rect 11426 24304 11482 24313
rect 11426 24239 11428 24248
rect 11480 24239 11482 24248
rect 11428 24210 11480 24216
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11440 23798 11468 24006
rect 11428 23792 11480 23798
rect 11428 23734 11480 23740
rect 11440 23662 11468 23734
rect 11428 23656 11480 23662
rect 11428 23598 11480 23604
rect 11336 22636 11388 22642
rect 11336 22578 11388 22584
rect 11440 22438 11468 23598
rect 11532 23322 11560 25463
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11428 22432 11480 22438
rect 11428 22374 11480 22380
rect 11440 22030 11468 22374
rect 11428 22024 11480 22030
rect 11428 21966 11480 21972
rect 11440 21690 11468 21966
rect 11428 21684 11480 21690
rect 11428 21626 11480 21632
rect 11336 21140 11388 21146
rect 11624 21128 11652 25894
rect 11716 21593 11744 25996
rect 11796 25696 11848 25702
rect 11796 25638 11848 25644
rect 11808 24750 11836 25638
rect 11900 24993 11928 26182
rect 11886 24984 11942 24993
rect 11886 24919 11942 24928
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11796 24744 11848 24750
rect 11796 24686 11848 24692
rect 11808 23526 11836 24686
rect 11900 24449 11928 24822
rect 11886 24440 11942 24449
rect 11886 24375 11942 24384
rect 11886 23624 11942 23633
rect 11886 23559 11888 23568
rect 11940 23559 11942 23568
rect 11888 23530 11940 23536
rect 11796 23520 11848 23526
rect 11796 23462 11848 23468
rect 11888 23044 11940 23050
rect 11888 22986 11940 22992
rect 11702 21584 11758 21593
rect 11702 21519 11758 21528
rect 11796 21344 11848 21350
rect 11796 21286 11848 21292
rect 11336 21082 11388 21088
rect 11440 21100 11652 21128
rect 11072 19468 11284 19496
rect 10690 19272 10746 19281
rect 11072 19242 11100 19468
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 10690 19207 10746 19216
rect 11060 19236 11112 19242
rect 11060 19178 11112 19184
rect 11072 18698 11100 19178
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 11164 18630 11192 19314
rect 11348 18630 11376 21082
rect 11440 21010 11468 21100
rect 11428 21004 11480 21010
rect 11428 20946 11480 20952
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11532 20058 11560 20946
rect 11808 20942 11836 21286
rect 11796 20936 11848 20942
rect 11796 20878 11848 20884
rect 11612 20596 11664 20602
rect 11612 20538 11664 20544
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11532 18834 11560 19858
rect 11520 18828 11572 18834
rect 11520 18770 11572 18776
rect 11152 18624 11204 18630
rect 11336 18624 11388 18630
rect 11204 18584 11284 18612
rect 11152 18566 11204 18572
rect 10839 18524 11147 18533
rect 10839 18522 10845 18524
rect 10901 18522 10925 18524
rect 10981 18522 11005 18524
rect 11061 18522 11085 18524
rect 11141 18522 11147 18524
rect 10901 18470 10903 18522
rect 11083 18470 11085 18522
rect 10839 18468 10845 18470
rect 10901 18468 10925 18470
rect 10981 18468 11005 18470
rect 11061 18468 11085 18470
rect 11141 18468 11147 18470
rect 10839 18459 11147 18468
rect 10612 18244 10916 18272
rect 10690 18184 10746 18193
rect 10690 18119 10746 18128
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10508 17604 10560 17610
rect 10508 17546 10560 17552
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 10428 17105 10456 17274
rect 10414 17096 10470 17105
rect 10414 17031 10470 17040
rect 10416 16584 10468 16590
rect 10416 16526 10468 16532
rect 10244 15166 10364 15194
rect 10244 14074 10272 15166
rect 10428 15076 10456 16526
rect 10520 15706 10548 17546
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10612 17202 10640 17478
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10508 15700 10560 15706
rect 10508 15642 10560 15648
rect 10336 15048 10456 15076
rect 10336 14482 10364 15048
rect 10612 15008 10640 16934
rect 10428 14980 10640 15008
rect 10324 14476 10376 14482
rect 10324 14418 10376 14424
rect 10428 14362 10456 14980
rect 10612 14929 10640 14980
rect 10598 14920 10654 14929
rect 10598 14855 10654 14864
rect 10336 14334 10456 14362
rect 10508 14408 10560 14414
rect 10508 14350 10560 14356
rect 10232 14068 10284 14074
rect 10232 14010 10284 14016
rect 10152 13892 10272 13920
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10152 13161 10180 13738
rect 10138 13152 10194 13161
rect 10138 13087 10194 13096
rect 10140 12640 10192 12646
rect 10244 12628 10272 13892
rect 10192 12600 10272 12628
rect 10140 12582 10192 12588
rect 10060 12396 10272 12424
rect 10048 12300 10100 12306
rect 10048 12242 10100 12248
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10060 10810 10088 12242
rect 10152 10810 10180 12242
rect 10244 12220 10272 12396
rect 10336 12288 10364 14334
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10428 13161 10456 13466
rect 10414 13152 10470 13161
rect 10414 13087 10470 13096
rect 10520 12986 10548 14350
rect 10704 14113 10732 18119
rect 10784 18080 10836 18086
rect 10784 18022 10836 18028
rect 10796 17610 10824 18022
rect 10784 17604 10836 17610
rect 10888 17592 10916 18244
rect 10968 17604 11020 17610
rect 10888 17564 10968 17592
rect 10784 17546 10836 17552
rect 10968 17546 11020 17552
rect 11256 17542 11284 18584
rect 11336 18566 11388 18572
rect 11244 17536 11296 17542
rect 11244 17478 11296 17484
rect 10839 17436 11147 17445
rect 10839 17434 10845 17436
rect 10901 17434 10925 17436
rect 10981 17434 11005 17436
rect 11061 17434 11085 17436
rect 11141 17434 11147 17436
rect 10901 17382 10903 17434
rect 11083 17382 11085 17434
rect 10839 17380 10845 17382
rect 10901 17380 10925 17382
rect 10981 17380 11005 17382
rect 11061 17380 11085 17382
rect 11141 17380 11147 17382
rect 10839 17371 11147 17380
rect 11256 17202 11284 17478
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 10796 16522 10824 17138
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 11256 16454 11284 17138
rect 11348 16794 11376 18566
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11532 17746 11560 18158
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11348 16658 11376 16730
rect 11336 16652 11388 16658
rect 11336 16594 11388 16600
rect 11428 16584 11480 16590
rect 11428 16526 11480 16532
rect 11440 16454 11468 16526
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 10839 16348 11147 16357
rect 10839 16346 10845 16348
rect 10901 16346 10925 16348
rect 10981 16346 11005 16348
rect 11061 16346 11085 16348
rect 11141 16346 11147 16348
rect 10901 16294 10903 16346
rect 11083 16294 11085 16346
rect 10839 16292 10845 16294
rect 10901 16292 10925 16294
rect 10981 16292 11005 16294
rect 11061 16292 11085 16294
rect 11141 16292 11147 16294
rect 10839 16283 11147 16292
rect 11058 16144 11114 16153
rect 11256 16130 11284 16390
rect 11114 16102 11284 16130
rect 11058 16079 11114 16088
rect 11244 15360 11296 15366
rect 11244 15302 11296 15308
rect 10839 15260 11147 15269
rect 10839 15258 10845 15260
rect 10901 15258 10925 15260
rect 10981 15258 11005 15260
rect 11061 15258 11085 15260
rect 11141 15258 11147 15260
rect 10901 15206 10903 15258
rect 11083 15206 11085 15258
rect 10839 15204 10845 15206
rect 10901 15204 10925 15206
rect 10981 15204 11005 15206
rect 11061 15204 11085 15206
rect 11141 15204 11147 15206
rect 10839 15195 11147 15204
rect 10968 15088 11020 15094
rect 10968 15030 11020 15036
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10980 14958 11008 15030
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10980 14260 11008 14894
rect 11072 14793 11100 15030
rect 11058 14784 11114 14793
rect 11058 14719 11114 14728
rect 11256 14414 11284 15302
rect 11348 15162 11376 16390
rect 11336 15156 11388 15162
rect 11336 15098 11388 15104
rect 11244 14408 11296 14414
rect 11244 14350 11296 14356
rect 10980 14232 11284 14260
rect 10839 14172 11147 14181
rect 10839 14170 10845 14172
rect 10901 14170 10925 14172
rect 10981 14170 11005 14172
rect 11061 14170 11085 14172
rect 11141 14170 11147 14172
rect 10901 14118 10903 14170
rect 11083 14118 11085 14170
rect 10839 14116 10845 14118
rect 10901 14116 10925 14118
rect 10981 14116 11005 14118
rect 11061 14116 11085 14118
rect 11141 14116 11147 14118
rect 10690 14104 10746 14113
rect 10839 14107 11147 14116
rect 10600 14068 10652 14074
rect 10690 14039 10746 14048
rect 10600 14010 10652 14016
rect 10612 13938 10640 14010
rect 10600 13932 10652 13938
rect 10600 13874 10652 13880
rect 10692 13864 10744 13870
rect 10598 13832 10654 13841
rect 10692 13806 10744 13812
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10598 13767 10654 13776
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10612 12481 10640 13767
rect 10598 12472 10654 12481
rect 10598 12407 10654 12416
rect 10416 12300 10468 12306
rect 10336 12260 10416 12288
rect 10416 12242 10468 12248
rect 10600 12232 10652 12238
rect 10244 12192 10364 12220
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 10244 11665 10272 11834
rect 10230 11656 10286 11665
rect 10230 11591 10286 11600
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 11082 10272 11494
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 10336 10962 10364 12192
rect 10600 12174 10652 12180
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 10428 11121 10456 12038
rect 10414 11112 10470 11121
rect 10414 11047 10470 11056
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10244 10934 10364 10962
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10140 10804 10192 10810
rect 10140 10746 10192 10752
rect 10046 10704 10102 10713
rect 10046 10639 10102 10648
rect 10060 10146 10088 10639
rect 9956 10124 10008 10130
rect 10060 10118 10180 10146
rect 9956 10066 10008 10072
rect 10048 9920 10100 9926
rect 10152 9897 10180 10118
rect 10048 9862 10100 9868
rect 10138 9888 10194 9897
rect 9954 9344 10010 9353
rect 9954 9279 10010 9288
rect 9968 9110 9996 9279
rect 9956 9104 10008 9110
rect 9956 9046 10008 9052
rect 9864 8900 9916 8906
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9312 8424 9364 8430
rect 9600 8378 9628 8774
rect 9312 8366 9364 8372
rect 9508 8350 9628 8378
rect 9220 8084 9272 8090
rect 9220 8026 9272 8032
rect 9232 7857 9260 8026
rect 9312 7880 9364 7886
rect 9218 7848 9274 7857
rect 9364 7840 9444 7868
rect 9312 7822 9364 7828
rect 9218 7783 9274 7792
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9232 7410 9260 7686
rect 9220 7404 9272 7410
rect 9220 7346 9272 7352
rect 9416 7002 9444 7840
rect 9312 6996 9364 7002
rect 9312 6938 9364 6944
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9232 6390 9260 6734
rect 9324 6390 9352 6938
rect 9508 6730 9536 8350
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9404 6248 9456 6254
rect 9310 6216 9366 6225
rect 9404 6190 9456 6196
rect 9310 6151 9366 6160
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9232 5817 9260 5850
rect 9218 5808 9274 5817
rect 9218 5743 9274 5752
rect 9220 5704 9272 5710
rect 9218 5672 9220 5681
rect 9272 5672 9274 5681
rect 9218 5607 9274 5616
rect 9220 5364 9272 5370
rect 9220 5306 9272 5312
rect 9232 5234 9260 5306
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9324 5137 9352 6151
rect 9416 5370 9444 6190
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9402 5264 9458 5273
rect 9402 5199 9458 5208
rect 9310 5128 9366 5137
rect 9310 5063 9366 5072
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9128 3528 9180 3534
rect 9128 3470 9180 3476
rect 9034 3360 9090 3369
rect 9034 3295 9090 3304
rect 9232 3233 9260 3878
rect 9416 3534 9444 5199
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9404 3528 9456 3534
rect 9310 3496 9366 3505
rect 9404 3470 9456 3476
rect 9310 3431 9366 3440
rect 9324 3398 9352 3431
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9218 3224 9274 3233
rect 9218 3159 9274 3168
rect 9128 3052 9180 3058
rect 8956 3012 9128 3040
rect 8852 2994 8904 3000
rect 9128 2994 9180 3000
rect 9220 2984 9272 2990
rect 9048 2932 9220 2938
rect 9048 2926 9272 2932
rect 9310 2952 9366 2961
rect 9048 2910 9260 2926
rect 8944 2848 8996 2854
rect 8864 2808 8944 2836
rect 8864 1834 8892 2808
rect 8944 2790 8996 2796
rect 9048 2650 9076 2910
rect 9416 2938 9444 3334
rect 9366 2910 9444 2938
rect 9310 2887 9366 2896
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9128 2440 9180 2446
rect 9034 2408 9090 2417
rect 9128 2382 9180 2388
rect 9034 2343 9090 2352
rect 9048 2310 9076 2343
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 9036 2304 9088 2310
rect 9140 2281 9168 2382
rect 9036 2246 9088 2252
rect 9126 2272 9182 2281
rect 8852 1828 8904 1834
rect 8852 1770 8904 1776
rect 8956 1578 8984 2246
rect 9126 2207 9182 2216
rect 9232 1714 9260 2790
rect 9324 2582 9352 2887
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 9508 2446 9536 4694
rect 9496 2440 9548 2446
rect 9496 2382 9548 2388
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9324 2106 9352 2246
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 9324 1873 9352 1906
rect 9310 1864 9366 1873
rect 9310 1799 9366 1808
rect 9404 1760 9456 1766
rect 9232 1686 9352 1714
rect 9404 1702 9456 1708
rect 8772 1550 8892 1578
rect 8956 1550 9260 1578
rect 9324 1562 9352 1686
rect 8114 1527 8170 1536
rect 8036 1414 8524 1442
rect 8114 1320 8170 1329
rect 8114 1255 8170 1264
rect 8128 160 8156 1255
rect 8206 1184 8262 1193
rect 8262 1142 8340 1170
rect 8206 1119 8262 1128
rect 8312 160 8340 1142
rect 8496 160 8524 1414
rect 8864 160 8892 1550
rect 9036 1216 9088 1222
rect 9036 1158 9088 1164
rect 9128 1216 9180 1222
rect 9128 1158 9180 1164
rect 9048 160 9076 1158
rect 9140 610 9168 1158
rect 9128 604 9180 610
rect 9128 546 9180 552
rect 9232 160 9260 1550
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9310 1456 9366 1465
rect 9310 1391 9366 1400
rect 9324 1018 9352 1391
rect 9312 1012 9364 1018
rect 9312 954 9364 960
rect 9416 160 9444 1702
rect 9508 1290 9536 2246
rect 9600 1970 9628 8230
rect 9692 8090 9720 8894
rect 9864 8842 9916 8848
rect 10060 8786 10088 9862
rect 10138 9823 10194 9832
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 9876 8758 10088 8786
rect 9772 8288 9824 8294
rect 9772 8230 9824 8236
rect 9680 8084 9732 8090
rect 9680 8026 9732 8032
rect 9784 7954 9812 8230
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 9692 7721 9720 7754
rect 9678 7712 9734 7721
rect 9678 7647 9734 7656
rect 9784 7342 9812 7890
rect 9876 7585 9904 8758
rect 10046 8664 10102 8673
rect 10046 8599 10102 8608
rect 9956 8084 10008 8090
rect 9956 8026 10008 8032
rect 9862 7576 9918 7585
rect 9862 7511 9918 7520
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9864 7200 9916 7206
rect 9678 7168 9734 7177
rect 9864 7142 9916 7148
rect 9678 7103 9734 7112
rect 9692 6769 9720 7103
rect 9772 6928 9824 6934
rect 9772 6870 9824 6876
rect 9678 6760 9734 6769
rect 9678 6695 9734 6704
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 3058 9720 6598
rect 9784 6440 9812 6870
rect 9876 6662 9904 7142
rect 9968 6866 9996 8026
rect 9956 6860 10008 6866
rect 9956 6802 10008 6808
rect 10060 6746 10088 8599
rect 9968 6718 10088 6746
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9864 6452 9916 6458
rect 9784 6412 9864 6440
rect 9864 6394 9916 6400
rect 9770 6352 9826 6361
rect 9968 6338 9996 6718
rect 10048 6656 10100 6662
rect 10048 6598 10100 6604
rect 9770 6287 9826 6296
rect 9876 6310 9996 6338
rect 9784 5846 9812 6287
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9784 5545 9812 5646
rect 9770 5536 9826 5545
rect 9770 5471 9826 5480
rect 9876 5114 9904 6310
rect 9956 6248 10008 6254
rect 9956 6190 10008 6196
rect 9968 5914 9996 6190
rect 9956 5908 10008 5914
rect 9956 5850 10008 5856
rect 10060 5794 10088 6598
rect 10152 6458 10180 9046
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10244 6322 10272 10934
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10336 9761 10364 10474
rect 10428 10146 10456 10746
rect 10520 10248 10548 11018
rect 10612 10810 10640 12174
rect 10704 11898 10732 13806
rect 10784 13320 10836 13326
rect 10888 13308 10916 13806
rect 11256 13716 11284 14232
rect 11440 14074 11468 16390
rect 11532 15620 11560 17682
rect 11624 15745 11652 20538
rect 11796 20528 11848 20534
rect 11900 20516 11928 22986
rect 11992 21486 12020 26182
rect 12176 25974 12204 26551
rect 12164 25968 12216 25974
rect 12164 25910 12216 25916
rect 12164 25696 12216 25702
rect 12070 25664 12126 25673
rect 12164 25638 12216 25644
rect 12070 25599 12126 25608
rect 12084 25294 12112 25599
rect 12176 25498 12204 25638
rect 12164 25492 12216 25498
rect 12164 25434 12216 25440
rect 12268 25378 12296 26710
rect 12346 26687 12402 26696
rect 12544 26382 12572 27406
rect 12532 26376 12584 26382
rect 12532 26318 12584 26324
rect 12636 26234 12664 33798
rect 12728 31346 12756 34342
rect 12716 31340 12768 31346
rect 12716 31282 12768 31288
rect 12716 29504 12768 29510
rect 12716 29446 12768 29452
rect 12728 29345 12756 29446
rect 12714 29336 12770 29345
rect 12714 29271 12770 29280
rect 12728 29102 12756 29271
rect 12716 29096 12768 29102
rect 12716 29038 12768 29044
rect 12714 28928 12770 28937
rect 12714 28863 12770 28872
rect 12728 28558 12756 28863
rect 12716 28552 12768 28558
rect 12716 28494 12768 28500
rect 12716 28416 12768 28422
rect 12716 28358 12768 28364
rect 12728 28082 12756 28358
rect 12716 28076 12768 28082
rect 12716 28018 12768 28024
rect 12716 27600 12768 27606
rect 12716 27542 12768 27548
rect 12728 27062 12756 27542
rect 12716 27056 12768 27062
rect 12716 26998 12768 27004
rect 12452 26206 12664 26234
rect 12716 26240 12768 26246
rect 12348 26036 12400 26042
rect 12348 25978 12400 25984
rect 12176 25350 12296 25378
rect 12072 25288 12124 25294
rect 12072 25230 12124 25236
rect 12072 24268 12124 24274
rect 12072 24210 12124 24216
rect 12084 23526 12112 24210
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 12084 23322 12112 23462
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 12070 23080 12126 23089
rect 12070 23015 12126 23024
rect 12084 22030 12112 23015
rect 12072 22024 12124 22030
rect 12072 21966 12124 21972
rect 12070 21584 12126 21593
rect 12070 21519 12072 21528
rect 12124 21519 12126 21528
rect 12072 21490 12124 21496
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 12084 20942 12112 21354
rect 12072 20936 12124 20942
rect 11978 20904 12034 20913
rect 12072 20878 12124 20884
rect 11978 20839 12034 20848
rect 11848 20488 11928 20516
rect 11796 20470 11848 20476
rect 11808 18358 11836 20470
rect 11992 19718 12020 20839
rect 12176 20806 12204 25350
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12268 24954 12296 25230
rect 12256 24948 12308 24954
rect 12256 24890 12308 24896
rect 12360 24206 12388 25978
rect 12348 24200 12400 24206
rect 12268 24160 12348 24188
rect 12268 22642 12296 24160
rect 12348 24142 12400 24148
rect 12346 24032 12402 24041
rect 12346 23967 12402 23976
rect 12256 22636 12308 22642
rect 12256 22578 12308 22584
rect 12256 22500 12308 22506
rect 12256 22442 12308 22448
rect 12268 22166 12296 22442
rect 12256 22160 12308 22166
rect 12256 22102 12308 22108
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12070 20496 12126 20505
rect 12070 20431 12072 20440
rect 12124 20431 12126 20440
rect 12072 20402 12124 20408
rect 12164 20256 12216 20262
rect 12268 20244 12296 21966
rect 12216 20216 12296 20244
rect 12164 20198 12216 20204
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 11980 19712 12032 19718
rect 11980 19654 12032 19660
rect 12164 19712 12216 19718
rect 12164 19654 12216 19660
rect 11886 19544 11942 19553
rect 11886 19479 11888 19488
rect 11940 19479 11942 19488
rect 11888 19450 11940 19456
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11716 16114 11744 17546
rect 11808 17105 11836 18294
rect 11794 17096 11850 17105
rect 11794 17031 11850 17040
rect 11794 16824 11850 16833
rect 11794 16759 11850 16768
rect 11808 16590 11836 16759
rect 11796 16584 11848 16590
rect 11796 16526 11848 16532
rect 11704 16108 11756 16114
rect 11704 16050 11756 16056
rect 11716 15858 11744 16050
rect 11808 16046 11836 16526
rect 11796 16040 11848 16046
rect 11796 15982 11848 15988
rect 11716 15830 11836 15858
rect 11610 15736 11666 15745
rect 11666 15694 11744 15722
rect 11610 15671 11666 15680
rect 11532 15592 11652 15620
rect 11520 15496 11572 15502
rect 11520 15438 11572 15444
rect 11532 15094 11560 15438
rect 11520 15088 11572 15094
rect 11520 15030 11572 15036
rect 11624 14958 11652 15592
rect 11716 15162 11744 15694
rect 11808 15638 11836 15830
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11612 14952 11664 14958
rect 11612 14894 11664 14900
rect 11612 14816 11664 14822
rect 11612 14758 11664 14764
rect 11704 14816 11756 14822
rect 11704 14758 11756 14764
rect 11518 14512 11574 14521
rect 11624 14482 11652 14758
rect 11716 14618 11744 14758
rect 11704 14612 11756 14618
rect 11704 14554 11756 14560
rect 11518 14447 11574 14456
rect 11612 14476 11664 14482
rect 11428 14068 11480 14074
rect 11428 14010 11480 14016
rect 11428 13728 11480 13734
rect 11256 13688 11428 13716
rect 11428 13670 11480 13676
rect 10836 13280 10916 13308
rect 10968 13320 11020 13326
rect 10784 13262 10836 13268
rect 11020 13280 11376 13308
rect 10968 13262 11020 13268
rect 11242 13152 11298 13161
rect 10839 13084 11147 13093
rect 11242 13087 11298 13096
rect 10839 13082 10845 13084
rect 10901 13082 10925 13084
rect 10981 13082 11005 13084
rect 11061 13082 11085 13084
rect 11141 13082 11147 13084
rect 10901 13030 10903 13082
rect 11083 13030 11085 13082
rect 10839 13028 10845 13030
rect 10901 13028 10925 13030
rect 10981 13028 11005 13030
rect 11061 13028 11085 13030
rect 11141 13028 11147 13030
rect 10839 13019 11147 13028
rect 11256 12594 11284 13087
rect 11072 12566 11284 12594
rect 11072 12209 11100 12566
rect 11244 12436 11296 12442
rect 11244 12378 11296 12384
rect 11256 12209 11284 12378
rect 11058 12200 11114 12209
rect 11058 12135 11114 12144
rect 11242 12200 11298 12209
rect 11242 12135 11298 12144
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 10839 11996 11147 12005
rect 10839 11994 10845 11996
rect 10901 11994 10925 11996
rect 10981 11994 11005 11996
rect 11061 11994 11085 11996
rect 11141 11994 11147 11996
rect 10901 11942 10903 11994
rect 11083 11942 11085 11994
rect 10839 11940 10845 11942
rect 10901 11940 10925 11942
rect 10981 11940 11005 11942
rect 11061 11940 11085 11942
rect 11141 11940 11147 11942
rect 10839 11931 11147 11940
rect 10692 11892 10744 11898
rect 10692 11834 10744 11840
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10704 10849 10732 11222
rect 11060 11144 11112 11150
rect 11060 11086 11112 11092
rect 11072 10996 11100 11086
rect 11072 10968 11217 10996
rect 10839 10908 11147 10917
rect 10839 10906 10845 10908
rect 10901 10906 10925 10908
rect 10981 10906 11005 10908
rect 11061 10906 11085 10908
rect 11141 10906 11147 10908
rect 10901 10854 10903 10906
rect 11083 10854 11085 10906
rect 10839 10852 10845 10854
rect 10901 10852 10925 10854
rect 10981 10852 11005 10854
rect 11061 10852 11085 10854
rect 11141 10852 11147 10854
rect 10690 10840 10746 10849
rect 10839 10843 11147 10852
rect 10600 10804 10652 10810
rect 11189 10810 11217 10968
rect 10690 10775 10746 10784
rect 11152 10804 11217 10810
rect 10600 10746 10652 10752
rect 11204 10764 11217 10804
rect 11152 10746 11204 10752
rect 11256 10577 11284 12038
rect 11348 11354 11376 13280
rect 11440 12753 11468 13670
rect 11532 13394 11560 14447
rect 11612 14418 11664 14424
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11426 12744 11482 12753
rect 11426 12679 11482 12688
rect 11440 11694 11468 12679
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11336 11348 11388 11354
rect 11532 11336 11560 13330
rect 11624 13025 11652 13466
rect 11610 13016 11666 13025
rect 11610 12951 11666 12960
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11336 11290 11388 11296
rect 11440 11308 11560 11336
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11242 10568 11298 10577
rect 10968 10532 11020 10538
rect 11242 10503 11298 10512
rect 10968 10474 11020 10480
rect 10520 10220 10640 10248
rect 10428 10130 10548 10146
rect 10612 10130 10640 10220
rect 10980 10130 11008 10474
rect 11242 10432 11298 10441
rect 11242 10367 11298 10376
rect 10428 10124 10560 10130
rect 10428 10118 10508 10124
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 10428 9586 10456 10118
rect 10508 10066 10560 10072
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10506 9616 10562 9625
rect 10416 9580 10468 9586
rect 10612 9586 10640 10066
rect 10784 10056 10836 10062
rect 10704 10004 10784 10010
rect 10704 9998 10836 10004
rect 10704 9982 10824 9998
rect 10506 9551 10562 9560
rect 10600 9580 10652 9586
rect 10416 9522 10468 9528
rect 10520 9353 10548 9551
rect 10600 9522 10652 9528
rect 10506 9344 10562 9353
rect 10506 9279 10562 9288
rect 10600 9036 10652 9042
rect 10600 8978 10652 8984
rect 10416 8968 10468 8974
rect 10468 8916 10548 8922
rect 10416 8910 10548 8916
rect 10428 8894 10548 8910
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10428 8634 10456 8774
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10140 6112 10192 6118
rect 10140 6054 10192 6060
rect 9784 5086 9904 5114
rect 9968 5766 10088 5794
rect 9784 5001 9812 5086
rect 9864 5024 9916 5030
rect 9770 4992 9826 5001
rect 9864 4966 9916 4972
rect 9770 4927 9826 4936
rect 9770 4856 9826 4865
rect 9876 4826 9904 4966
rect 9770 4791 9826 4800
rect 9864 4820 9916 4826
rect 9784 3738 9812 4791
rect 9864 4762 9916 4768
rect 9876 3738 9904 4762
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9862 3632 9918 3641
rect 9862 3567 9918 3576
rect 9876 3534 9904 3567
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9968 3058 9996 5766
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 10060 5370 10088 5510
rect 10048 5364 10100 5370
rect 10048 5306 10100 5312
rect 10060 4690 10088 5306
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 10046 4584 10102 4593
rect 10046 4519 10102 4528
rect 10060 4486 10088 4519
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 10060 4026 10088 4422
rect 10152 4214 10180 6054
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10244 4282 10272 5578
rect 10336 5302 10364 8502
rect 10414 7848 10470 7857
rect 10414 7783 10470 7792
rect 10428 5953 10456 7783
rect 10520 7041 10548 8894
rect 10612 7546 10640 8978
rect 10704 8634 10732 9982
rect 11256 9897 11284 10367
rect 11242 9888 11298 9897
rect 10839 9820 11147 9829
rect 11242 9823 11298 9832
rect 10839 9818 10845 9820
rect 10901 9818 10925 9820
rect 10981 9818 11005 9820
rect 11061 9818 11085 9820
rect 11141 9818 11147 9820
rect 10901 9766 10903 9818
rect 11083 9766 11085 9818
rect 10839 9764 10845 9766
rect 10901 9764 10925 9766
rect 10981 9764 11005 9766
rect 11061 9764 11085 9766
rect 11141 9764 11147 9766
rect 10839 9755 11147 9764
rect 10966 9616 11022 9625
rect 10796 9574 10966 9602
rect 10796 9042 10824 9574
rect 10966 9551 11022 9560
rect 11348 9466 11376 11086
rect 10888 9438 11376 9466
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10888 8838 10916 9438
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 10980 8838 11008 8910
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10839 8732 11147 8741
rect 10839 8730 10845 8732
rect 10901 8730 10925 8732
rect 10981 8730 11005 8732
rect 11061 8730 11085 8732
rect 11141 8730 11147 8732
rect 10901 8678 10903 8730
rect 11083 8678 11085 8730
rect 10839 8676 10845 8678
rect 10901 8676 10925 8678
rect 10981 8676 11005 8678
rect 11061 8676 11085 8678
rect 11141 8676 11147 8678
rect 10839 8667 11147 8676
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 10692 8424 10744 8430
rect 10692 8366 10744 8372
rect 10704 7886 10732 8366
rect 10874 8256 10930 8265
rect 10874 8191 10930 8200
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 10796 7732 10824 8026
rect 10888 7857 10916 8191
rect 10874 7848 10930 7857
rect 10874 7783 10930 7792
rect 11072 7750 11100 8570
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 10704 7704 10824 7732
rect 11060 7744 11112 7750
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10704 7188 10732 7704
rect 11164 7732 11192 8298
rect 11256 8090 11284 8910
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11242 7848 11298 7857
rect 11242 7783 11298 7792
rect 11164 7704 11217 7732
rect 11060 7686 11112 7692
rect 10839 7644 11147 7653
rect 10839 7642 10845 7644
rect 10901 7642 10925 7644
rect 10981 7642 11005 7644
rect 11061 7642 11085 7644
rect 11141 7642 11147 7644
rect 10901 7590 10903 7642
rect 11083 7590 11085 7642
rect 10839 7588 10845 7590
rect 10901 7588 10925 7590
rect 10981 7588 11005 7590
rect 11061 7588 11085 7590
rect 11141 7588 11147 7590
rect 10839 7579 11147 7588
rect 11189 7528 11217 7704
rect 10888 7500 11217 7528
rect 10612 7160 10732 7188
rect 10784 7200 10836 7206
rect 10506 7032 10562 7041
rect 10506 6967 10562 6976
rect 10520 6866 10548 6967
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10520 6361 10548 6598
rect 10506 6352 10562 6361
rect 10506 6287 10562 6296
rect 10612 6202 10640 7160
rect 10888 7177 10916 7500
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 10784 7142 10836 7148
rect 10874 7168 10930 7177
rect 10796 6984 10824 7142
rect 10874 7103 10930 7112
rect 10796 6956 10916 6984
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10520 6174 10640 6202
rect 10414 5944 10470 5953
rect 10414 5879 10470 5888
rect 10414 5808 10470 5817
rect 10414 5743 10470 5752
rect 10324 5296 10376 5302
rect 10324 5238 10376 5244
rect 10322 4992 10378 5001
rect 10322 4927 10378 4936
rect 10232 4276 10284 4282
rect 10232 4218 10284 4224
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10060 3998 10180 4026
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10060 3777 10088 3878
rect 10046 3768 10102 3777
rect 10046 3703 10102 3712
rect 10152 3482 10180 3998
rect 10244 3913 10272 4082
rect 10230 3904 10286 3913
rect 10230 3839 10286 3848
rect 10336 3618 10364 4927
rect 10428 4758 10456 5743
rect 10520 4826 10548 6174
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10508 4820 10560 4826
rect 10508 4762 10560 4768
rect 10416 4752 10468 4758
rect 10416 4694 10468 4700
rect 10506 4720 10562 4729
rect 10428 4282 10456 4694
rect 10506 4655 10562 4664
rect 10416 4276 10468 4282
rect 10416 4218 10468 4224
rect 10520 4128 10548 4655
rect 10612 4282 10640 6054
rect 10704 5370 10732 6802
rect 10888 6644 10916 6956
rect 10980 6905 11008 7278
rect 11152 7268 11204 7274
rect 11152 7210 11204 7216
rect 11058 7168 11114 7177
rect 11058 7103 11114 7112
rect 10966 6896 11022 6905
rect 10966 6831 11022 6840
rect 11072 6798 11100 7103
rect 11164 6798 11192 7210
rect 11060 6792 11112 6798
rect 11060 6734 11112 6740
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10888 6616 11217 6644
rect 10839 6556 11147 6565
rect 10839 6554 10845 6556
rect 10901 6554 10925 6556
rect 10981 6554 11005 6556
rect 11061 6554 11085 6556
rect 11141 6554 11147 6556
rect 10901 6502 10903 6554
rect 11083 6502 11085 6554
rect 10839 6500 10845 6502
rect 10901 6500 10925 6502
rect 10981 6500 11005 6502
rect 11061 6500 11085 6502
rect 11141 6500 11147 6502
rect 10839 6491 11147 6500
rect 11189 6440 11217 6616
rect 10980 6412 11217 6440
rect 10782 5944 10838 5953
rect 10782 5879 10838 5888
rect 10796 5574 10824 5879
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10980 5534 11008 6412
rect 11150 6352 11206 6361
rect 11060 6316 11112 6322
rect 11150 6287 11152 6296
rect 11060 6258 11112 6264
rect 11204 6287 11206 6296
rect 11152 6258 11204 6264
rect 11072 6225 11100 6258
rect 11058 6216 11114 6225
rect 11058 6151 11114 6160
rect 11058 6080 11114 6089
rect 11058 6015 11114 6024
rect 11072 5681 11100 6015
rect 11256 5794 11284 7783
rect 11348 7313 11376 9318
rect 11440 9042 11468 11308
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11532 10606 11560 11154
rect 11624 11150 11652 11698
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11610 10840 11666 10849
rect 11610 10775 11666 10784
rect 11520 10600 11572 10606
rect 11520 10542 11572 10548
rect 11532 10130 11560 10542
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11520 9512 11572 9518
rect 11520 9454 11572 9460
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11440 8650 11468 8978
rect 11532 8809 11560 9454
rect 11518 8800 11574 8809
rect 11518 8735 11574 8744
rect 11440 8622 11560 8650
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11334 7304 11390 7313
rect 11334 7239 11390 7248
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11348 5914 11376 6734
rect 11440 6254 11468 8502
rect 11532 7954 11560 8622
rect 11624 8430 11652 10775
rect 11716 9722 11744 12786
rect 11808 11014 11836 14962
rect 11900 14362 11928 19450
rect 11992 15026 12020 19654
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12084 18630 12112 18702
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12072 18352 12124 18358
rect 12072 18294 12124 18300
rect 12084 17678 12112 18294
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12084 17270 12112 17614
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 12070 17096 12126 17105
rect 12070 17031 12126 17040
rect 12084 16998 12112 17031
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12176 16522 12204 19654
rect 12268 17626 12296 19994
rect 12360 19009 12388 23967
rect 12452 23769 12480 26206
rect 12716 26182 12768 26188
rect 12728 25956 12756 26182
rect 12636 25945 12756 25956
rect 12636 25936 12770 25945
rect 12636 25928 12714 25936
rect 12532 25900 12584 25906
rect 12532 25842 12584 25848
rect 12544 25498 12572 25842
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12636 25294 12664 25928
rect 12714 25871 12770 25880
rect 12716 25764 12768 25770
rect 12716 25706 12768 25712
rect 12728 25673 12756 25706
rect 12714 25664 12770 25673
rect 12714 25599 12770 25608
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12636 23848 12664 25230
rect 12820 24698 12848 34711
rect 12912 28762 12940 36518
rect 13004 34406 13032 37606
rect 12992 34400 13044 34406
rect 12992 34342 13044 34348
rect 12992 33516 13044 33522
rect 12992 33458 13044 33464
rect 13004 32774 13032 33458
rect 12992 32768 13044 32774
rect 12992 32710 13044 32716
rect 13096 32609 13124 38898
rect 13188 36582 13216 41534
rect 13312 40828 13620 40837
rect 13312 40826 13318 40828
rect 13374 40826 13398 40828
rect 13454 40826 13478 40828
rect 13534 40826 13558 40828
rect 13614 40826 13620 40828
rect 13374 40774 13376 40826
rect 13556 40774 13558 40826
rect 13312 40772 13318 40774
rect 13374 40772 13398 40774
rect 13454 40772 13478 40774
rect 13534 40772 13558 40774
rect 13614 40772 13620 40774
rect 13312 40763 13620 40772
rect 13648 40526 13676 41550
rect 13544 40520 13596 40526
rect 13544 40462 13596 40468
rect 13636 40520 13688 40526
rect 13636 40462 13688 40468
rect 13556 40089 13584 40462
rect 13542 40080 13598 40089
rect 13542 40015 13598 40024
rect 13312 39740 13620 39749
rect 13312 39738 13318 39740
rect 13374 39738 13398 39740
rect 13454 39738 13478 39740
rect 13534 39738 13558 39740
rect 13614 39738 13620 39740
rect 13374 39686 13376 39738
rect 13556 39686 13558 39738
rect 13312 39684 13318 39686
rect 13374 39684 13398 39686
rect 13454 39684 13478 39686
rect 13534 39684 13558 39686
rect 13614 39684 13620 39686
rect 13312 39675 13620 39684
rect 13740 39642 13768 41670
rect 13728 39636 13780 39642
rect 13728 39578 13780 39584
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 13312 38652 13620 38661
rect 13312 38650 13318 38652
rect 13374 38650 13398 38652
rect 13454 38650 13478 38652
rect 13534 38650 13558 38652
rect 13614 38650 13620 38652
rect 13374 38598 13376 38650
rect 13556 38598 13558 38650
rect 13312 38596 13318 38598
rect 13374 38596 13398 38598
rect 13454 38596 13478 38598
rect 13534 38596 13558 38598
rect 13614 38596 13620 38598
rect 13312 38587 13620 38596
rect 13832 38350 13860 38694
rect 13820 38344 13872 38350
rect 13820 38286 13872 38292
rect 13728 38208 13780 38214
rect 13728 38150 13780 38156
rect 13740 38010 13768 38150
rect 13728 38004 13780 38010
rect 13728 37946 13780 37952
rect 13924 37806 13952 41958
rect 13912 37800 13964 37806
rect 13912 37742 13964 37748
rect 13312 37564 13620 37573
rect 13312 37562 13318 37564
rect 13374 37562 13398 37564
rect 13454 37562 13478 37564
rect 13534 37562 13558 37564
rect 13614 37562 13620 37564
rect 13374 37510 13376 37562
rect 13556 37510 13558 37562
rect 13312 37508 13318 37510
rect 13374 37508 13398 37510
rect 13454 37508 13478 37510
rect 13534 37508 13558 37510
rect 13614 37508 13620 37510
rect 13312 37499 13620 37508
rect 14016 37466 14044 42502
rect 14108 41818 14136 42894
rect 14292 42906 14320 43046
rect 14186 42871 14242 42880
rect 14280 42900 14332 42906
rect 14280 42842 14332 42848
rect 14370 42392 14426 42401
rect 14370 42327 14426 42336
rect 14384 42022 14412 42327
rect 14476 42226 14504 43046
rect 14464 42220 14516 42226
rect 14464 42162 14516 42168
rect 14280 42016 14332 42022
rect 14280 41958 14332 41964
rect 14372 42016 14424 42022
rect 14372 41958 14424 41964
rect 14462 41984 14518 41993
rect 14096 41812 14148 41818
rect 14096 41754 14148 41760
rect 14188 41744 14240 41750
rect 14186 41712 14188 41721
rect 14240 41712 14242 41721
rect 14186 41647 14242 41656
rect 14292 41414 14320 41958
rect 14462 41919 14518 41928
rect 14476 41834 14504 41919
rect 14200 41386 14320 41414
rect 14384 41806 14504 41834
rect 14200 40168 14228 41386
rect 14384 41274 14412 41806
rect 14464 41472 14516 41478
rect 14464 41414 14516 41420
rect 14372 41268 14424 41274
rect 14372 41210 14424 41216
rect 14200 40140 14412 40168
rect 14188 40044 14240 40050
rect 14188 39986 14240 39992
rect 14096 38888 14148 38894
rect 14096 38830 14148 38836
rect 14108 38350 14136 38830
rect 14096 38344 14148 38350
rect 14096 38286 14148 38292
rect 14004 37460 14056 37466
rect 14004 37402 14056 37408
rect 13636 37324 13688 37330
rect 13636 37266 13688 37272
rect 13452 37188 13504 37194
rect 13452 37130 13504 37136
rect 13464 36718 13492 37130
rect 13452 36712 13504 36718
rect 13452 36654 13504 36660
rect 13176 36576 13228 36582
rect 13176 36518 13228 36524
rect 13312 36476 13620 36485
rect 13312 36474 13318 36476
rect 13374 36474 13398 36476
rect 13454 36474 13478 36476
rect 13534 36474 13558 36476
rect 13614 36474 13620 36476
rect 13374 36422 13376 36474
rect 13556 36422 13558 36474
rect 13312 36420 13318 36422
rect 13374 36420 13398 36422
rect 13454 36420 13478 36422
rect 13534 36420 13558 36422
rect 13614 36420 13620 36422
rect 13312 36411 13620 36420
rect 13542 36272 13598 36281
rect 13542 36207 13598 36216
rect 13556 35562 13584 36207
rect 13544 35556 13596 35562
rect 13544 35498 13596 35504
rect 13176 35488 13228 35494
rect 13176 35430 13228 35436
rect 13188 33862 13216 35430
rect 13312 35388 13620 35397
rect 13312 35386 13318 35388
rect 13374 35386 13398 35388
rect 13454 35386 13478 35388
rect 13534 35386 13558 35388
rect 13614 35386 13620 35388
rect 13374 35334 13376 35386
rect 13556 35334 13558 35386
rect 13312 35332 13318 35334
rect 13374 35332 13398 35334
rect 13454 35332 13478 35334
rect 13534 35332 13558 35334
rect 13614 35332 13620 35334
rect 13312 35323 13620 35332
rect 13312 34300 13620 34309
rect 13312 34298 13318 34300
rect 13374 34298 13398 34300
rect 13454 34298 13478 34300
rect 13534 34298 13558 34300
rect 13614 34298 13620 34300
rect 13374 34246 13376 34298
rect 13556 34246 13558 34298
rect 13312 34244 13318 34246
rect 13374 34244 13398 34246
rect 13454 34244 13478 34246
rect 13534 34244 13558 34246
rect 13614 34244 13620 34246
rect 13312 34235 13620 34244
rect 13176 33856 13228 33862
rect 13176 33798 13228 33804
rect 13176 33312 13228 33318
rect 13176 33254 13228 33260
rect 13188 33017 13216 33254
rect 13312 33212 13620 33221
rect 13312 33210 13318 33212
rect 13374 33210 13398 33212
rect 13454 33210 13478 33212
rect 13534 33210 13558 33212
rect 13614 33210 13620 33212
rect 13374 33158 13376 33210
rect 13556 33158 13558 33210
rect 13312 33156 13318 33158
rect 13374 33156 13398 33158
rect 13454 33156 13478 33158
rect 13534 33156 13558 33158
rect 13614 33156 13620 33158
rect 13312 33147 13620 33156
rect 13174 33008 13230 33017
rect 13174 32943 13230 32952
rect 13082 32600 13138 32609
rect 13082 32535 13138 32544
rect 13188 32434 13216 32943
rect 13176 32428 13228 32434
rect 13176 32370 13228 32376
rect 13084 32224 13136 32230
rect 13084 32166 13136 32172
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 13096 32026 13124 32166
rect 13084 32020 13136 32026
rect 13084 31962 13136 31968
rect 13084 31680 13136 31686
rect 13188 31657 13216 32166
rect 13312 32124 13620 32133
rect 13312 32122 13318 32124
rect 13374 32122 13398 32124
rect 13454 32122 13478 32124
rect 13534 32122 13558 32124
rect 13614 32122 13620 32124
rect 13374 32070 13376 32122
rect 13556 32070 13558 32122
rect 13312 32068 13318 32070
rect 13374 32068 13398 32070
rect 13454 32068 13478 32070
rect 13534 32068 13558 32070
rect 13614 32068 13620 32070
rect 13312 32059 13620 32068
rect 13084 31622 13136 31628
rect 13174 31648 13230 31657
rect 12992 31272 13044 31278
rect 12992 31214 13044 31220
rect 13004 30274 13032 31214
rect 13096 30598 13124 31622
rect 13174 31583 13230 31592
rect 13188 31278 13216 31583
rect 13176 31272 13228 31278
rect 13176 31214 13228 31220
rect 13312 31036 13620 31045
rect 13312 31034 13318 31036
rect 13374 31034 13398 31036
rect 13454 31034 13478 31036
rect 13534 31034 13558 31036
rect 13614 31034 13620 31036
rect 13374 30982 13376 31034
rect 13556 30982 13558 31034
rect 13312 30980 13318 30982
rect 13374 30980 13398 30982
rect 13454 30980 13478 30982
rect 13534 30980 13558 30982
rect 13614 30980 13620 30982
rect 13312 30971 13620 30980
rect 13360 30932 13412 30938
rect 13360 30874 13412 30880
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 13004 30246 13216 30274
rect 13372 30258 13400 30874
rect 13648 30716 13676 37266
rect 14002 37088 14058 37097
rect 14002 37023 14058 37032
rect 14016 36854 14044 37023
rect 13728 36848 13780 36854
rect 13728 36790 13780 36796
rect 14004 36848 14056 36854
rect 14004 36790 14056 36796
rect 13740 36281 13768 36790
rect 13912 36304 13964 36310
rect 13726 36272 13782 36281
rect 13912 36246 13964 36252
rect 13726 36207 13782 36216
rect 13728 36032 13780 36038
rect 13728 35974 13780 35980
rect 13820 36032 13872 36038
rect 13820 35974 13872 35980
rect 13740 35834 13768 35974
rect 13728 35828 13780 35834
rect 13728 35770 13780 35776
rect 13832 35290 13860 35974
rect 13820 35284 13872 35290
rect 13820 35226 13872 35232
rect 13820 35012 13872 35018
rect 13820 34954 13872 34960
rect 13832 34610 13860 34954
rect 13820 34604 13872 34610
rect 13820 34546 13872 34552
rect 13924 34490 13952 36246
rect 14108 36242 14136 38286
rect 14096 36236 14148 36242
rect 14096 36178 14148 36184
rect 14200 35986 14228 39986
rect 14384 38010 14412 40140
rect 14476 39817 14504 41414
rect 14568 41274 14596 44540
rect 14646 43072 14702 43081
rect 14646 43007 14702 43016
rect 14660 42838 14688 43007
rect 14648 42832 14700 42838
rect 14648 42774 14700 42780
rect 14648 42560 14700 42566
rect 14648 42502 14700 42508
rect 14660 42362 14688 42502
rect 14648 42356 14700 42362
rect 14648 42298 14700 42304
rect 14648 42220 14700 42226
rect 14648 42162 14700 42168
rect 14660 41274 14688 42162
rect 14752 41274 14780 44540
rect 14936 44010 14964 44540
rect 14936 43982 15056 44010
rect 14924 43920 14976 43926
rect 14924 43862 14976 43868
rect 14832 43648 14884 43654
rect 14832 43590 14884 43596
rect 14844 43314 14872 43590
rect 14936 43314 14964 43862
rect 14832 43308 14884 43314
rect 14832 43250 14884 43256
rect 14924 43308 14976 43314
rect 14924 43250 14976 43256
rect 14924 43104 14976 43110
rect 14924 43046 14976 43052
rect 14936 42770 14964 43046
rect 15028 42922 15056 43982
rect 15120 43314 15148 44540
rect 15304 43738 15332 44540
rect 15474 44540 15530 45000
rect 15658 44540 15714 45000
rect 15842 44540 15898 45000
rect 16026 44540 16082 45000
rect 16210 44540 16266 45000
rect 16394 44540 16450 45000
rect 16578 44540 16634 45000
rect 16762 44540 16818 45000
rect 16946 44540 17002 45000
rect 17130 44540 17186 45000
rect 17314 44540 17370 45000
rect 17498 44540 17554 45000
rect 17682 44540 17738 45000
rect 17866 44540 17922 45000
rect 18050 44540 18106 45000
rect 18234 44540 18290 45000
rect 18418 44540 18474 45000
rect 18602 44540 18658 45000
rect 18786 44540 18842 45000
rect 18970 44540 19026 45000
rect 19154 44540 19210 45000
rect 19338 44540 19394 45000
rect 15382 44503 15438 44512
rect 15396 44418 15424 44503
rect 15488 44418 15516 44540
rect 15396 44390 15516 44418
rect 15474 43888 15530 43897
rect 15474 43823 15530 43832
rect 15212 43722 15332 43738
rect 15200 43716 15332 43722
rect 15252 43710 15332 43716
rect 15200 43658 15252 43664
rect 15488 43314 15516 43823
rect 15672 43761 15700 44540
rect 15856 43874 15884 44540
rect 16040 44010 16068 44540
rect 16224 44146 16252 44540
rect 16224 44118 16344 44146
rect 16040 43982 16252 44010
rect 15856 43846 16160 43874
rect 15658 43752 15714 43761
rect 15658 43687 15714 43696
rect 15784 43548 16092 43557
rect 15784 43546 15790 43548
rect 15846 43546 15870 43548
rect 15926 43546 15950 43548
rect 16006 43546 16030 43548
rect 16086 43546 16092 43548
rect 15846 43494 15848 43546
rect 16028 43494 16030 43546
rect 15784 43492 15790 43494
rect 15846 43492 15870 43494
rect 15926 43492 15950 43494
rect 16006 43492 16030 43494
rect 16086 43492 16092 43494
rect 15784 43483 16092 43492
rect 16132 43450 16160 43846
rect 16224 43450 16252 43982
rect 16316 43466 16344 44118
rect 16408 43602 16436 44540
rect 16408 43574 16528 43602
rect 16120 43444 16172 43450
rect 16120 43386 16172 43392
rect 16212 43444 16264 43450
rect 16316 43438 16436 43466
rect 16212 43386 16264 43392
rect 16408 43382 16436 43438
rect 16304 43376 16356 43382
rect 16304 43318 16356 43324
rect 16396 43376 16448 43382
rect 16396 43318 16448 43324
rect 15108 43308 15160 43314
rect 15108 43250 15160 43256
rect 15476 43308 15528 43314
rect 15476 43250 15528 43256
rect 15660 43308 15712 43314
rect 15660 43250 15712 43256
rect 16120 43308 16172 43314
rect 16120 43250 16172 43256
rect 15028 42894 15240 42922
rect 15108 42832 15160 42838
rect 15108 42774 15160 42780
rect 14924 42764 14976 42770
rect 14924 42706 14976 42712
rect 14924 42560 14976 42566
rect 14924 42502 14976 42508
rect 15016 42560 15068 42566
rect 15016 42502 15068 42508
rect 14830 42392 14886 42401
rect 14830 42327 14886 42336
rect 14844 42106 14872 42327
rect 14936 42226 14964 42502
rect 14924 42220 14976 42226
rect 14924 42162 14976 42168
rect 14844 42078 14964 42106
rect 14832 42016 14884 42022
rect 14832 41958 14884 41964
rect 14844 41585 14872 41958
rect 14936 41750 14964 42078
rect 15028 41818 15056 42502
rect 15016 41812 15068 41818
rect 15016 41754 15068 41760
rect 14924 41744 14976 41750
rect 15120 41698 15148 42774
rect 14924 41686 14976 41692
rect 15028 41670 15148 41698
rect 14830 41576 14886 41585
rect 14830 41511 14886 41520
rect 14832 41472 14884 41478
rect 14832 41414 14884 41420
rect 14556 41268 14608 41274
rect 14556 41210 14608 41216
rect 14648 41268 14700 41274
rect 14648 41210 14700 41216
rect 14740 41268 14792 41274
rect 14740 41210 14792 41216
rect 14844 41177 14872 41414
rect 15028 41274 15056 41670
rect 15212 41596 15240 42894
rect 15304 42758 15516 42786
rect 15304 42362 15332 42758
rect 15488 42702 15516 42758
rect 15384 42696 15436 42702
rect 15384 42638 15436 42644
rect 15476 42696 15528 42702
rect 15476 42638 15528 42644
rect 15292 42356 15344 42362
rect 15292 42298 15344 42304
rect 15396 42242 15424 42638
rect 15476 42560 15528 42566
rect 15476 42502 15528 42508
rect 15488 42362 15516 42502
rect 15566 42392 15622 42401
rect 15476 42356 15528 42362
rect 15566 42327 15622 42336
rect 15476 42298 15528 42304
rect 15304 42214 15424 42242
rect 15304 42022 15332 42214
rect 15580 42140 15608 42327
rect 15396 42112 15608 42140
rect 15396 42022 15424 42112
rect 15292 42016 15344 42022
rect 15292 41958 15344 41964
rect 15384 42016 15436 42022
rect 15384 41958 15436 41964
rect 15476 42016 15528 42022
rect 15476 41958 15528 41964
rect 15488 41857 15516 41958
rect 15474 41848 15530 41857
rect 15474 41783 15530 41792
rect 15672 41732 15700 43250
rect 16132 43217 16160 43250
rect 16118 43208 16174 43217
rect 16118 43143 16174 43152
rect 16212 42696 16264 42702
rect 16210 42664 16212 42673
rect 16264 42664 16266 42673
rect 16210 42599 16266 42608
rect 16120 42560 16172 42566
rect 16120 42502 16172 42508
rect 16212 42560 16264 42566
rect 16212 42502 16264 42508
rect 15784 42460 16092 42469
rect 15784 42458 15790 42460
rect 15846 42458 15870 42460
rect 15926 42458 15950 42460
rect 16006 42458 16030 42460
rect 16086 42458 16092 42460
rect 15846 42406 15848 42458
rect 16028 42406 16030 42458
rect 15784 42404 15790 42406
rect 15846 42404 15870 42406
rect 15926 42404 15950 42406
rect 16006 42404 16030 42406
rect 16086 42404 16092 42406
rect 15784 42395 16092 42404
rect 16132 42362 16160 42502
rect 16224 42362 16252 42502
rect 16120 42356 16172 42362
rect 16120 42298 16172 42304
rect 16212 42356 16264 42362
rect 16212 42298 16264 42304
rect 16316 42226 16344 43318
rect 16396 43104 16448 43110
rect 16396 43046 16448 43052
rect 16408 42786 16436 43046
rect 16500 42906 16528 43574
rect 16592 43110 16620 44540
rect 16580 43104 16632 43110
rect 16580 43046 16632 43052
rect 16488 42900 16540 42906
rect 16488 42842 16540 42848
rect 16578 42800 16634 42809
rect 16408 42758 16528 42786
rect 16396 42628 16448 42634
rect 16396 42570 16448 42576
rect 16408 42265 16436 42570
rect 16500 42294 16528 42758
rect 16776 42770 16804 44540
rect 16960 43178 16988 44540
rect 17144 43602 17172 44540
rect 17328 43874 17356 44540
rect 17328 43846 17448 43874
rect 17144 43574 17356 43602
rect 17224 43308 17276 43314
rect 17224 43250 17276 43256
rect 16948 43172 17000 43178
rect 16948 43114 17000 43120
rect 16578 42735 16634 42744
rect 16764 42764 16816 42770
rect 16488 42288 16540 42294
rect 16394 42256 16450 42265
rect 16304 42220 16356 42226
rect 16488 42230 16540 42236
rect 16592 42226 16620 42735
rect 16764 42706 16816 42712
rect 16856 42696 16908 42702
rect 16856 42638 16908 42644
rect 16394 42191 16450 42200
rect 16580 42220 16632 42226
rect 16304 42162 16356 42168
rect 16580 42162 16632 42168
rect 16302 42120 16358 42129
rect 16358 42078 16528 42106
rect 16302 42055 16358 42064
rect 15844 42016 15896 42022
rect 15844 41958 15896 41964
rect 15750 41848 15806 41857
rect 15750 41783 15806 41792
rect 15764 41750 15792 41783
rect 15580 41704 15700 41732
rect 15752 41744 15804 41750
rect 15212 41568 15332 41596
rect 15304 41562 15332 41568
rect 15304 41534 15404 41562
rect 15376 41460 15404 41534
rect 15198 41440 15254 41449
rect 15376 41432 15424 41460
rect 15198 41375 15254 41384
rect 15212 41274 15240 41375
rect 15016 41268 15068 41274
rect 15016 41210 15068 41216
rect 15200 41268 15252 41274
rect 15200 41210 15252 41216
rect 14554 41168 14610 41177
rect 14554 41103 14556 41112
rect 14608 41103 14610 41112
rect 14830 41168 14886 41177
rect 14830 41103 14886 41112
rect 15198 41168 15254 41177
rect 15396 41138 15424 41432
rect 15580 41274 15608 41704
rect 15752 41686 15804 41692
rect 15660 41608 15712 41614
rect 15856 41596 15884 41958
rect 16500 41614 16528 42078
rect 16580 41744 16632 41750
rect 16580 41686 16632 41692
rect 15712 41568 15884 41596
rect 15936 41608 15988 41614
rect 15660 41550 15712 41556
rect 16304 41608 16356 41614
rect 15936 41550 15988 41556
rect 16026 41576 16082 41585
rect 15948 41460 15976 41550
rect 16026 41511 16082 41520
rect 16224 41568 16304 41596
rect 16040 41478 16068 41511
rect 15672 41432 15976 41460
rect 16028 41472 16080 41478
rect 15568 41268 15620 41274
rect 15568 41210 15620 41216
rect 15198 41103 15254 41112
rect 15384 41132 15436 41138
rect 14556 41074 14608 41080
rect 14924 40928 14976 40934
rect 14922 40896 14924 40905
rect 14976 40896 14978 40905
rect 14922 40831 14978 40840
rect 15212 40730 15240 41103
rect 15384 41074 15436 41080
rect 15568 41132 15620 41138
rect 15568 41074 15620 41080
rect 15476 41064 15528 41070
rect 15476 41006 15528 41012
rect 15384 40928 15436 40934
rect 15384 40870 15436 40876
rect 15200 40724 15252 40730
rect 15200 40666 15252 40672
rect 15396 40526 15424 40870
rect 15488 40730 15516 41006
rect 15476 40724 15528 40730
rect 15476 40666 15528 40672
rect 15384 40520 15436 40526
rect 15384 40462 15436 40468
rect 15292 40452 15344 40458
rect 15292 40394 15344 40400
rect 14924 40384 14976 40390
rect 14924 40326 14976 40332
rect 15106 40352 15162 40361
rect 14648 40044 14700 40050
rect 14648 39986 14700 39992
rect 14462 39808 14518 39817
rect 14462 39743 14518 39752
rect 14556 39092 14608 39098
rect 14556 39034 14608 39040
rect 14372 38004 14424 38010
rect 14372 37946 14424 37952
rect 14278 37768 14334 37777
rect 14278 37703 14334 37712
rect 14108 35958 14228 35986
rect 14004 35080 14056 35086
rect 14004 35022 14056 35028
rect 13832 34462 13952 34490
rect 13726 34232 13782 34241
rect 13726 34167 13782 34176
rect 13740 34066 13768 34167
rect 13832 34134 13860 34462
rect 13820 34128 13872 34134
rect 13820 34070 13872 34076
rect 13728 34060 13780 34066
rect 13728 34002 13780 34008
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 13820 33924 13872 33930
rect 13820 33866 13872 33872
rect 13832 33833 13860 33866
rect 13818 33824 13874 33833
rect 13818 33759 13874 33768
rect 13818 33688 13874 33697
rect 13818 33623 13874 33632
rect 13832 33590 13860 33623
rect 13820 33584 13872 33590
rect 13820 33526 13872 33532
rect 13924 33454 13952 34002
rect 13912 33448 13964 33454
rect 13912 33390 13964 33396
rect 14016 32978 14044 35022
rect 14004 32972 14056 32978
rect 14004 32914 14056 32920
rect 13820 32836 13872 32842
rect 13820 32778 13872 32784
rect 13728 32768 13780 32774
rect 13728 32710 13780 32716
rect 13740 30938 13768 32710
rect 13832 32570 13860 32778
rect 14016 32774 14044 32914
rect 14004 32768 14056 32774
rect 14004 32710 14056 32716
rect 13820 32564 13872 32570
rect 13820 32506 13872 32512
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 13832 31482 13860 32370
rect 14004 32224 14056 32230
rect 14004 32166 14056 32172
rect 13912 31816 13964 31822
rect 14016 31804 14044 32166
rect 13964 31776 14044 31804
rect 13912 31758 13964 31764
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13820 31272 13872 31278
rect 13820 31214 13872 31220
rect 13832 30938 13860 31214
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13820 30932 13872 30938
rect 13820 30874 13872 30880
rect 13818 30832 13874 30841
rect 13818 30767 13874 30776
rect 13648 30688 13768 30716
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 13004 28558 13032 30246
rect 13188 30190 13216 30246
rect 13360 30252 13412 30258
rect 13360 30194 13412 30200
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 13176 30184 13228 30190
rect 13176 30126 13228 30132
rect 13096 28558 13124 30126
rect 13636 30116 13688 30122
rect 13636 30058 13688 30064
rect 13312 29948 13620 29957
rect 13312 29946 13318 29948
rect 13374 29946 13398 29948
rect 13454 29946 13478 29948
rect 13534 29946 13558 29948
rect 13614 29946 13620 29948
rect 13374 29894 13376 29946
rect 13556 29894 13558 29946
rect 13312 29892 13318 29894
rect 13374 29892 13398 29894
rect 13454 29892 13478 29894
rect 13534 29892 13558 29894
rect 13614 29892 13620 29894
rect 13312 29883 13620 29892
rect 13648 29850 13676 30058
rect 13636 29844 13688 29850
rect 13636 29786 13688 29792
rect 13544 29776 13596 29782
rect 13596 29724 13676 29730
rect 13544 29718 13676 29724
rect 13556 29702 13676 29718
rect 13176 29640 13228 29646
rect 13176 29582 13228 29588
rect 13188 29306 13216 29582
rect 13176 29300 13228 29306
rect 13176 29242 13228 29248
rect 13174 28928 13230 28937
rect 13174 28863 13230 28872
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 13084 28552 13136 28558
rect 13084 28494 13136 28500
rect 12900 28008 12952 28014
rect 12898 27976 12900 27985
rect 12952 27976 12954 27985
rect 12898 27911 12954 27920
rect 12898 26616 12954 26625
rect 12898 26551 12954 26560
rect 12912 26382 12940 26551
rect 12900 26376 12952 26382
rect 12900 26318 12952 26324
rect 12900 26036 12952 26042
rect 12900 25978 12952 25984
rect 12912 24818 12940 25978
rect 12900 24812 12952 24818
rect 12900 24754 12952 24760
rect 13004 24721 13032 28494
rect 13096 27878 13124 28494
rect 13188 27946 13216 28863
rect 13312 28860 13620 28869
rect 13312 28858 13318 28860
rect 13374 28858 13398 28860
rect 13454 28858 13478 28860
rect 13534 28858 13558 28860
rect 13614 28858 13620 28860
rect 13374 28806 13376 28858
rect 13556 28806 13558 28858
rect 13312 28804 13318 28806
rect 13374 28804 13398 28806
rect 13454 28804 13478 28806
rect 13534 28804 13558 28806
rect 13614 28804 13620 28806
rect 13312 28795 13620 28804
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 13556 28393 13584 28698
rect 13542 28384 13598 28393
rect 13542 28319 13598 28328
rect 13176 27940 13228 27946
rect 13176 27882 13228 27888
rect 13084 27872 13136 27878
rect 13084 27814 13136 27820
rect 13312 27772 13620 27781
rect 13312 27770 13318 27772
rect 13374 27770 13398 27772
rect 13454 27770 13478 27772
rect 13534 27770 13558 27772
rect 13614 27770 13620 27772
rect 13374 27718 13376 27770
rect 13556 27718 13558 27770
rect 13312 27716 13318 27718
rect 13374 27716 13398 27718
rect 13454 27716 13478 27718
rect 13534 27716 13558 27718
rect 13614 27716 13620 27718
rect 13082 27704 13138 27713
rect 13312 27707 13620 27716
rect 13082 27639 13138 27648
rect 13176 27668 13228 27674
rect 13096 26314 13124 27639
rect 13176 27610 13228 27616
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 13188 26246 13216 27610
rect 13648 27538 13676 29702
rect 13636 27532 13688 27538
rect 13636 27474 13688 27480
rect 13636 26852 13688 26858
rect 13636 26794 13688 26800
rect 13312 26684 13620 26693
rect 13312 26682 13318 26684
rect 13374 26682 13398 26684
rect 13454 26682 13478 26684
rect 13534 26682 13558 26684
rect 13614 26682 13620 26684
rect 13374 26630 13376 26682
rect 13556 26630 13558 26682
rect 13312 26628 13318 26630
rect 13374 26628 13398 26630
rect 13454 26628 13478 26630
rect 13534 26628 13558 26630
rect 13614 26628 13620 26630
rect 13312 26619 13620 26628
rect 13648 26586 13676 26794
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13176 26240 13228 26246
rect 13176 26182 13228 26188
rect 13740 25974 13768 30688
rect 13832 29481 13860 30767
rect 13924 30190 13952 31758
rect 14004 31272 14056 31278
rect 14004 31214 14056 31220
rect 14016 30394 14044 31214
rect 14108 30841 14136 35958
rect 14188 35012 14240 35018
rect 14188 34954 14240 34960
rect 14200 32026 14228 34954
rect 14292 34785 14320 37703
rect 14372 35488 14424 35494
rect 14372 35430 14424 35436
rect 14384 35086 14412 35430
rect 14568 35193 14596 39034
rect 14660 38894 14688 39986
rect 14936 39846 14964 40326
rect 15106 40287 15162 40296
rect 14924 39840 14976 39846
rect 14924 39782 14976 39788
rect 14648 38888 14700 38894
rect 14648 38830 14700 38836
rect 15120 38536 15148 40287
rect 15304 39438 15332 40394
rect 15580 40186 15608 41074
rect 15672 40730 15700 41432
rect 16028 41414 16080 41420
rect 15784 41372 16092 41381
rect 15784 41370 15790 41372
rect 15846 41370 15870 41372
rect 15926 41370 15950 41372
rect 16006 41370 16030 41372
rect 16086 41370 16092 41372
rect 15846 41318 15848 41370
rect 16028 41318 16030 41370
rect 15784 41316 15790 41318
rect 15846 41316 15870 41318
rect 15926 41316 15950 41318
rect 16006 41316 16030 41318
rect 16086 41316 16092 41318
rect 15784 41307 16092 41316
rect 16224 41138 16252 41568
rect 16304 41550 16356 41556
rect 16396 41608 16448 41614
rect 16396 41550 16448 41556
rect 16488 41608 16540 41614
rect 16488 41550 16540 41556
rect 16408 41274 16436 41550
rect 16592 41414 16620 41686
rect 16764 41608 16816 41614
rect 16764 41550 16816 41556
rect 16500 41386 16620 41414
rect 16396 41268 16448 41274
rect 16396 41210 16448 41216
rect 16500 41154 16528 41386
rect 16578 41304 16634 41313
rect 16578 41239 16634 41248
rect 16212 41132 16264 41138
rect 16212 41074 16264 41080
rect 16304 41132 16356 41138
rect 16304 41074 16356 41080
rect 16408 41126 16528 41154
rect 16210 40760 16266 40769
rect 15660 40724 15712 40730
rect 16210 40695 16212 40704
rect 15660 40666 15712 40672
rect 16264 40695 16266 40704
rect 16212 40666 16264 40672
rect 15660 40520 15712 40526
rect 15660 40462 15712 40468
rect 16120 40520 16172 40526
rect 16120 40462 16172 40468
rect 15568 40180 15620 40186
rect 15568 40122 15620 40128
rect 15672 39642 15700 40462
rect 15784 40284 16092 40293
rect 15784 40282 15790 40284
rect 15846 40282 15870 40284
rect 15926 40282 15950 40284
rect 16006 40282 16030 40284
rect 16086 40282 16092 40284
rect 15846 40230 15848 40282
rect 16028 40230 16030 40282
rect 15784 40228 15790 40230
rect 15846 40228 15870 40230
rect 15926 40228 15950 40230
rect 16006 40228 16030 40230
rect 16086 40228 16092 40230
rect 15784 40219 16092 40228
rect 16132 40186 16160 40462
rect 16212 40384 16264 40390
rect 16212 40326 16264 40332
rect 16120 40180 16172 40186
rect 16120 40122 16172 40128
rect 15660 39636 15712 39642
rect 15660 39578 15712 39584
rect 16224 39574 16252 40326
rect 16212 39568 16264 39574
rect 16212 39510 16264 39516
rect 15292 39432 15344 39438
rect 15292 39374 15344 39380
rect 15476 39432 15528 39438
rect 15476 39374 15528 39380
rect 15200 38956 15252 38962
rect 15200 38898 15252 38904
rect 14844 38508 15148 38536
rect 14740 36712 14792 36718
rect 14740 36654 14792 36660
rect 14752 36582 14780 36654
rect 14740 36576 14792 36582
rect 14740 36518 14792 36524
rect 14752 35630 14780 36518
rect 14648 35624 14700 35630
rect 14648 35566 14700 35572
rect 14740 35624 14792 35630
rect 14740 35566 14792 35572
rect 14554 35184 14610 35193
rect 14554 35119 14610 35128
rect 14372 35080 14424 35086
rect 14372 35022 14424 35028
rect 14556 35080 14608 35086
rect 14556 35022 14608 35028
rect 14372 34944 14424 34950
rect 14372 34886 14424 34892
rect 14278 34776 14334 34785
rect 14278 34711 14334 34720
rect 14280 34604 14332 34610
rect 14384 34592 14412 34886
rect 14332 34564 14412 34592
rect 14280 34546 14332 34552
rect 14384 34513 14412 34564
rect 14370 34504 14426 34513
rect 14370 34439 14426 34448
rect 14280 34400 14332 34406
rect 14280 34342 14332 34348
rect 14292 32502 14320 34342
rect 14462 34232 14518 34241
rect 14462 34167 14518 34176
rect 14372 33380 14424 33386
rect 14372 33322 14424 33328
rect 14280 32496 14332 32502
rect 14280 32438 14332 32444
rect 14280 32360 14332 32366
rect 14280 32302 14332 32308
rect 14292 32026 14320 32302
rect 14188 32020 14240 32026
rect 14188 31962 14240 31968
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14200 31142 14228 31962
rect 14278 31784 14334 31793
rect 14278 31719 14334 31728
rect 14188 31136 14240 31142
rect 14188 31078 14240 31084
rect 14094 30832 14150 30841
rect 14292 30818 14320 31719
rect 14094 30767 14150 30776
rect 14200 30790 14320 30818
rect 14200 30734 14228 30790
rect 14188 30728 14240 30734
rect 14094 30696 14150 30705
rect 14188 30670 14240 30676
rect 14094 30631 14150 30640
rect 14004 30388 14056 30394
rect 14004 30330 14056 30336
rect 14016 30258 14044 30330
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 13912 30184 13964 30190
rect 13912 30126 13964 30132
rect 13818 29472 13874 29481
rect 13818 29407 13874 29416
rect 13832 28665 13860 29407
rect 13818 28656 13874 28665
rect 13818 28591 13874 28600
rect 13818 28112 13874 28121
rect 13818 28047 13874 28056
rect 13832 27130 13860 28047
rect 13924 27996 13952 30126
rect 14108 29170 14136 30631
rect 14096 29164 14148 29170
rect 14096 29106 14148 29112
rect 14108 28529 14136 29106
rect 14188 28960 14240 28966
rect 14188 28902 14240 28908
rect 14200 28762 14228 28902
rect 14188 28756 14240 28762
rect 14188 28698 14240 28704
rect 14094 28520 14150 28529
rect 14292 28490 14320 30790
rect 14094 28455 14150 28464
rect 14280 28484 14332 28490
rect 14280 28426 14332 28432
rect 14292 28082 14320 28426
rect 14188 28076 14240 28082
rect 14188 28018 14240 28024
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 13924 27968 14044 27996
rect 13912 27872 13964 27878
rect 13912 27814 13964 27820
rect 13924 27577 13952 27814
rect 13910 27568 13966 27577
rect 13910 27503 13966 27512
rect 13820 27124 13872 27130
rect 13820 27066 13872 27072
rect 13912 27124 13964 27130
rect 13912 27066 13964 27072
rect 13728 25968 13780 25974
rect 13542 25936 13598 25945
rect 13598 25894 13676 25922
rect 13728 25910 13780 25916
rect 13542 25871 13598 25880
rect 13360 25832 13412 25838
rect 13648 25820 13676 25894
rect 13728 25832 13780 25838
rect 13542 25800 13598 25809
rect 13412 25780 13542 25786
rect 13360 25774 13542 25780
rect 13372 25758 13542 25774
rect 13648 25792 13728 25820
rect 13728 25774 13780 25780
rect 13542 25735 13598 25744
rect 13728 25696 13780 25702
rect 13728 25638 13780 25644
rect 13312 25596 13620 25605
rect 13312 25594 13318 25596
rect 13374 25594 13398 25596
rect 13454 25594 13478 25596
rect 13534 25594 13558 25596
rect 13614 25594 13620 25596
rect 13374 25542 13376 25594
rect 13556 25542 13558 25594
rect 13312 25540 13318 25542
rect 13374 25540 13398 25542
rect 13454 25540 13478 25542
rect 13534 25540 13558 25542
rect 13614 25540 13620 25542
rect 13312 25531 13620 25540
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13268 25288 13320 25294
rect 13268 25230 13320 25236
rect 13280 24936 13308 25230
rect 13121 24908 13308 24936
rect 13121 24868 13149 24908
rect 13096 24840 13149 24868
rect 12990 24712 13046 24721
rect 12820 24670 12940 24698
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12820 24274 12848 24550
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12634 23820 12664 23848
rect 12438 23760 12494 23769
rect 12438 23695 12494 23704
rect 12634 23712 12662 23820
rect 12820 23769 12848 24210
rect 12806 23760 12862 23769
rect 12634 23684 12664 23712
rect 12806 23695 12862 23704
rect 12440 23656 12492 23662
rect 12532 23656 12584 23662
rect 12440 23598 12492 23604
rect 12530 23624 12532 23633
rect 12636 23644 12664 23684
rect 12584 23624 12586 23633
rect 12452 23526 12480 23598
rect 12530 23559 12586 23568
rect 12634 23616 12664 23644
rect 12634 23576 12662 23616
rect 12912 23576 12940 24670
rect 12990 24647 13046 24656
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 13004 23866 13032 24550
rect 12992 23860 13044 23866
rect 12992 23802 13044 23808
rect 12634 23548 12664 23576
rect 12440 23520 12492 23526
rect 12440 23462 12492 23468
rect 12452 21350 12480 23462
rect 12636 22094 12664 23548
rect 12544 22066 12664 22094
rect 12820 23548 12940 23576
rect 12544 21962 12572 22066
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 12716 21412 12768 21418
rect 12716 21354 12768 21360
rect 12440 21344 12492 21350
rect 12440 21286 12492 21292
rect 12452 21146 12480 21286
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12544 19530 12572 20198
rect 12452 19502 12572 19530
rect 12346 19000 12402 19009
rect 12346 18935 12402 18944
rect 12346 18728 12402 18737
rect 12346 18663 12402 18672
rect 12360 18057 12388 18663
rect 12452 18358 12480 19502
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12544 18970 12572 19314
rect 12532 18964 12584 18970
rect 12532 18906 12584 18912
rect 12532 18760 12584 18766
rect 12636 18748 12664 20742
rect 12728 20602 12756 21354
rect 12716 20596 12768 20602
rect 12716 20538 12768 20544
rect 12714 20224 12770 20233
rect 12714 20159 12770 20168
rect 12584 18720 12664 18748
rect 12532 18702 12584 18708
rect 12440 18352 12492 18358
rect 12440 18294 12492 18300
rect 12440 18216 12492 18222
rect 12440 18158 12492 18164
rect 12346 18048 12402 18057
rect 12346 17983 12402 17992
rect 12268 17598 12388 17626
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12164 16516 12216 16522
rect 12164 16458 12216 16464
rect 12162 16416 12218 16425
rect 12162 16351 12218 16360
rect 12176 15201 12204 16351
rect 12162 15192 12218 15201
rect 12072 15156 12124 15162
rect 12268 15162 12296 17478
rect 12360 15609 12388 17598
rect 12452 16114 12480 18158
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12346 15600 12402 15609
rect 12346 15535 12402 15544
rect 12452 15502 12480 16050
rect 12440 15496 12492 15502
rect 12360 15444 12440 15450
rect 12360 15438 12492 15444
rect 12360 15422 12480 15438
rect 12162 15127 12218 15136
rect 12256 15156 12308 15162
rect 12072 15098 12124 15104
rect 12256 15098 12308 15104
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 12084 14657 12112 15098
rect 12162 15056 12218 15065
rect 12162 14991 12164 15000
rect 12216 14991 12218 15000
rect 12164 14962 12216 14968
rect 12070 14648 12126 14657
rect 12070 14583 12126 14592
rect 12072 14408 12124 14414
rect 11900 14334 12020 14362
rect 12176 14396 12204 14962
rect 12124 14368 12204 14396
rect 12072 14350 12124 14356
rect 11992 14278 12020 14334
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11900 12986 11928 13330
rect 11992 13190 12020 14214
rect 12070 14104 12126 14113
rect 12070 14039 12126 14048
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11992 12918 12020 13126
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11888 12640 11940 12646
rect 11888 12582 11940 12588
rect 11900 11937 11928 12582
rect 11992 12102 12020 12854
rect 11980 12096 12032 12102
rect 11980 12038 12032 12044
rect 11886 11928 11942 11937
rect 11886 11863 11942 11872
rect 11900 11762 11928 11863
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11886 11656 11942 11665
rect 11886 11591 11942 11600
rect 11796 11008 11848 11014
rect 11796 10950 11848 10956
rect 11808 10713 11836 10950
rect 11794 10704 11850 10713
rect 11794 10639 11850 10648
rect 11808 10062 11836 10639
rect 11796 10056 11848 10062
rect 11796 9998 11848 10004
rect 11704 9716 11756 9722
rect 11704 9658 11756 9664
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11716 7664 11744 9658
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11808 7818 11836 9318
rect 11900 9217 11928 11591
rect 11886 9208 11942 9217
rect 11886 9143 11942 9152
rect 11992 9042 12020 12038
rect 12084 11286 12112 14039
rect 12176 13326 12204 14368
rect 12268 13870 12296 15098
rect 12256 13864 12308 13870
rect 12256 13806 12308 13812
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12176 12918 12204 13262
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 12176 12238 12204 12854
rect 12164 12232 12216 12238
rect 12164 12174 12216 12180
rect 12256 12164 12308 12170
rect 12256 12106 12308 12112
rect 12268 11898 12296 12106
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12070 11112 12126 11121
rect 12070 11047 12126 11056
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11888 8968 11940 8974
rect 11888 8910 11940 8916
rect 11900 8362 11928 8910
rect 11978 8800 12034 8809
rect 11978 8735 12034 8744
rect 11888 8356 11940 8362
rect 11992 8344 12020 8735
rect 12084 8498 12112 11047
rect 12176 8498 12204 11766
rect 12256 11756 12308 11762
rect 12256 11698 12308 11704
rect 12268 11354 12296 11698
rect 12256 11348 12308 11354
rect 12256 11290 12308 11296
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12268 9042 12296 10950
rect 12360 10810 12388 15422
rect 12440 14952 12492 14958
rect 12440 14894 12492 14900
rect 12452 14346 12480 14894
rect 12440 14340 12492 14346
rect 12440 14282 12492 14288
rect 12452 13308 12480 14282
rect 12544 14006 12572 18702
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12636 17105 12664 18022
rect 12622 17096 12678 17105
rect 12622 17031 12678 17040
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12636 14958 12664 15098
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12622 14648 12678 14657
rect 12622 14583 12678 14592
rect 12636 14346 12664 14583
rect 12624 14340 12676 14346
rect 12624 14282 12676 14288
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12728 13569 12756 20159
rect 12714 13560 12770 13569
rect 12714 13495 12770 13504
rect 12532 13320 12584 13326
rect 12452 13280 12532 13308
rect 12532 13262 12584 13268
rect 12716 13252 12768 13258
rect 12716 13194 12768 13200
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12452 11354 12480 12786
rect 12532 12776 12584 12782
rect 12532 12718 12584 12724
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12544 10810 12572 12718
rect 12624 12300 12676 12306
rect 12624 12242 12676 12248
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12532 10804 12584 10810
rect 12532 10746 12584 10752
rect 12360 10062 12388 10746
rect 12440 10668 12492 10674
rect 12440 10610 12492 10616
rect 12348 10056 12400 10062
rect 12348 9998 12400 10004
rect 12348 9716 12400 9722
rect 12348 9658 12400 9664
rect 12360 9353 12388 9658
rect 12346 9344 12402 9353
rect 12346 9279 12402 9288
rect 12346 9208 12402 9217
rect 12346 9143 12402 9152
rect 12256 9036 12308 9042
rect 12256 8978 12308 8984
rect 12254 8528 12310 8537
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12164 8492 12216 8498
rect 12254 8463 12310 8472
rect 12164 8434 12216 8440
rect 12072 8356 12124 8362
rect 11992 8316 12072 8344
rect 11888 8298 11940 8304
rect 12072 8298 12124 8304
rect 11888 7948 11940 7954
rect 11888 7890 11940 7896
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11532 7636 11744 7664
rect 11532 7410 11560 7636
rect 11808 7562 11836 7754
rect 11624 7534 11836 7562
rect 11520 7404 11572 7410
rect 11520 7346 11572 7352
rect 11624 7342 11652 7534
rect 11900 7410 11928 7890
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11612 7336 11664 7342
rect 11518 7304 11574 7313
rect 11612 7278 11664 7284
rect 11518 7239 11574 7248
rect 11532 7206 11560 7239
rect 11520 7200 11572 7206
rect 11520 7142 11572 7148
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11518 7032 11574 7041
rect 11518 6967 11574 6976
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11532 6100 11560 6967
rect 11624 6225 11652 7142
rect 11716 6984 11744 7346
rect 11992 7290 12020 7686
rect 11900 7262 12020 7290
rect 11716 6956 11836 6984
rect 11808 6934 11836 6956
rect 11808 6928 11866 6934
rect 11702 6896 11758 6905
rect 11808 6888 11814 6928
rect 11814 6870 11866 6876
rect 11702 6831 11758 6840
rect 11610 6216 11666 6225
rect 11610 6151 11666 6160
rect 11426 6080 11482 6089
rect 11532 6072 11652 6100
rect 11426 6015 11482 6024
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11256 5766 11376 5794
rect 11058 5672 11114 5681
rect 11058 5607 11114 5616
rect 10980 5506 11284 5534
rect 10839 5468 11147 5477
rect 10839 5466 10845 5468
rect 10901 5466 10925 5468
rect 10981 5466 11005 5468
rect 11061 5466 11085 5468
rect 11141 5466 11147 5468
rect 10901 5414 10903 5466
rect 11083 5414 11085 5466
rect 10839 5412 10845 5414
rect 10901 5412 10925 5414
rect 10981 5412 11005 5414
rect 11061 5412 11085 5414
rect 11141 5412 11147 5414
rect 10839 5403 11147 5412
rect 11256 5370 11284 5506
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 10782 5264 10838 5273
rect 11348 5250 11376 5766
rect 10782 5199 10838 5208
rect 11256 5222 11376 5250
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10704 4622 10732 5034
rect 10796 4690 10824 5199
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 11058 5128 11114 5137
rect 10874 4992 10930 5001
rect 10874 4927 10930 4936
rect 10888 4826 10916 4927
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10874 4720 10930 4729
rect 10784 4684 10836 4690
rect 10874 4655 10930 4664
rect 10784 4626 10836 4632
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10888 4468 10916 4655
rect 10980 4622 11008 5102
rect 11058 5063 11114 5072
rect 10968 4616 11020 4622
rect 11072 4593 11100 5063
rect 11152 4684 11204 4690
rect 11152 4626 11204 4632
rect 10968 4558 11020 4564
rect 11058 4584 11114 4593
rect 11058 4519 11114 4528
rect 10704 4440 10916 4468
rect 11164 4468 11192 4626
rect 11164 4440 11217 4468
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10600 4140 10652 4146
rect 10520 4100 10600 4128
rect 10600 4082 10652 4088
rect 10704 4026 10732 4440
rect 10839 4380 11147 4389
rect 10839 4378 10845 4380
rect 10901 4378 10925 4380
rect 10981 4378 11005 4380
rect 11061 4378 11085 4380
rect 11141 4378 11147 4380
rect 10901 4326 10903 4378
rect 11083 4326 11085 4378
rect 10839 4324 10845 4326
rect 10901 4324 10925 4326
rect 10981 4324 11005 4326
rect 11061 4324 11085 4326
rect 11141 4324 11147 4326
rect 10839 4315 11147 4324
rect 11189 4282 11217 4440
rect 11152 4276 11217 4282
rect 11204 4236 11217 4276
rect 11152 4218 11204 4224
rect 11150 4040 11206 4049
rect 10600 4004 10652 4010
rect 10704 3998 10824 4026
rect 10600 3946 10652 3952
rect 10506 3632 10562 3641
rect 10336 3590 10506 3618
rect 10506 3567 10562 3576
rect 10612 3534 10640 3946
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10600 3528 10652 3534
rect 10152 3454 10548 3482
rect 10600 3470 10652 3476
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9956 3052 10008 3058
rect 9956 2994 10008 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10048 2916 10100 2922
rect 10048 2858 10100 2864
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9772 2848 9824 2854
rect 9772 2790 9824 2796
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9692 1834 9720 2790
rect 9680 1828 9732 1834
rect 9680 1770 9732 1776
rect 9588 1760 9640 1766
rect 9588 1702 9640 1708
rect 9496 1284 9548 1290
rect 9496 1226 9548 1232
rect 9600 160 9628 1702
rect 9784 1562 9812 2790
rect 9864 2304 9916 2310
rect 9864 2246 9916 2252
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9772 1556 9824 1562
rect 9772 1498 9824 1504
rect 9876 1494 9904 2246
rect 9968 2106 9996 2246
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 9864 1488 9916 1494
rect 9864 1430 9916 1436
rect 10060 1412 10088 2858
rect 10138 2544 10194 2553
rect 10138 2479 10194 2488
rect 10152 2446 10180 2479
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10244 2394 10272 2994
rect 10336 2632 10364 3334
rect 10416 2984 10468 2990
rect 10414 2952 10416 2961
rect 10468 2952 10470 2961
rect 10414 2887 10470 2896
rect 10416 2848 10468 2854
rect 10414 2816 10416 2825
rect 10468 2816 10470 2825
rect 10414 2751 10470 2760
rect 10520 2774 10548 3454
rect 10600 3392 10652 3398
rect 10704 3369 10732 3878
rect 10796 3738 10824 3998
rect 11072 3998 11150 4026
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 11072 3602 11100 3998
rect 11150 3975 11206 3984
rect 11256 3924 11284 5222
rect 11334 5128 11390 5137
rect 11334 5063 11390 5072
rect 11348 4146 11376 5063
rect 11440 4826 11468 6015
rect 11518 5536 11574 5545
rect 11518 5471 11574 5480
rect 11532 5166 11560 5471
rect 11520 5160 11572 5166
rect 11624 5137 11652 6072
rect 11716 5534 11744 6831
rect 11796 6452 11848 6458
rect 11796 6394 11848 6400
rect 11808 6322 11836 6394
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11794 6216 11850 6225
rect 11794 6151 11850 6160
rect 11808 5710 11836 6151
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11716 5506 11836 5534
rect 11702 5400 11758 5409
rect 11808 5370 11836 5506
rect 11702 5335 11704 5344
rect 11756 5335 11758 5344
rect 11796 5364 11848 5370
rect 11704 5306 11756 5312
rect 11796 5306 11848 5312
rect 11900 5250 11928 7262
rect 12084 6798 12112 8298
rect 12176 7886 12204 8434
rect 12164 7880 12216 7886
rect 12164 7822 12216 7828
rect 12162 7576 12218 7585
rect 12162 7511 12218 7520
rect 12176 7002 12204 7511
rect 12268 7313 12296 8463
rect 12360 8265 12388 9143
rect 12346 8256 12402 8265
rect 12346 8191 12402 8200
rect 12452 7954 12480 10610
rect 12636 10266 12664 12242
rect 12728 11558 12756 13194
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12820 10441 12848 23548
rect 13096 23118 13124 24840
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13188 23866 13216 24754
rect 13372 24682 13400 25434
rect 13740 25294 13768 25638
rect 13728 25288 13780 25294
rect 13728 25230 13780 25236
rect 13832 24993 13860 27066
rect 13924 26994 13952 27066
rect 13912 26988 13964 26994
rect 13912 26930 13964 26936
rect 13910 25936 13966 25945
rect 13910 25871 13966 25880
rect 13924 25498 13952 25871
rect 13912 25492 13964 25498
rect 13912 25434 13964 25440
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13818 24984 13874 24993
rect 13818 24919 13874 24928
rect 13636 24812 13688 24818
rect 13636 24754 13688 24760
rect 13728 24812 13780 24818
rect 13728 24754 13780 24760
rect 13360 24676 13412 24682
rect 13360 24618 13412 24624
rect 13312 24508 13620 24517
rect 13312 24506 13318 24508
rect 13374 24506 13398 24508
rect 13454 24506 13478 24508
rect 13534 24506 13558 24508
rect 13614 24506 13620 24508
rect 13374 24454 13376 24506
rect 13556 24454 13558 24506
rect 13312 24452 13318 24454
rect 13374 24452 13398 24454
rect 13454 24452 13478 24454
rect 13534 24452 13558 24454
rect 13614 24452 13620 24454
rect 13312 24443 13620 24452
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13556 24290 13584 24346
rect 13648 24290 13676 24754
rect 13556 24262 13676 24290
rect 13740 24206 13768 24754
rect 13924 24698 13952 25230
rect 13832 24670 13952 24698
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 13174 23760 13230 23769
rect 13174 23695 13230 23704
rect 13188 23594 13216 23695
rect 13176 23588 13228 23594
rect 13176 23530 13228 23536
rect 13312 23420 13620 23429
rect 13312 23418 13318 23420
rect 13374 23418 13398 23420
rect 13454 23418 13478 23420
rect 13534 23418 13558 23420
rect 13614 23418 13620 23420
rect 13374 23366 13376 23418
rect 13556 23366 13558 23418
rect 13312 23364 13318 23366
rect 13374 23364 13398 23366
rect 13454 23364 13478 23366
rect 13534 23364 13558 23366
rect 13614 23364 13620 23366
rect 13312 23355 13620 23364
rect 12900 23112 12952 23118
rect 12900 23054 12952 23060
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 12912 18630 12940 23054
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 12990 22536 13046 22545
rect 12990 22471 13046 22480
rect 13004 21690 13032 22471
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 13096 21554 13124 22578
rect 13312 22332 13620 22341
rect 13312 22330 13318 22332
rect 13374 22330 13398 22332
rect 13454 22330 13478 22332
rect 13534 22330 13558 22332
rect 13614 22330 13620 22332
rect 13374 22278 13376 22330
rect 13556 22278 13558 22330
rect 13312 22276 13318 22278
rect 13374 22276 13398 22278
rect 13454 22276 13478 22278
rect 13534 22276 13558 22278
rect 13614 22276 13620 22278
rect 13312 22267 13620 22276
rect 13648 22216 13676 24142
rect 13832 23730 13860 24670
rect 13912 24608 13964 24614
rect 13912 24550 13964 24556
rect 13924 24206 13952 24550
rect 13912 24200 13964 24206
rect 13912 24142 13964 24148
rect 13912 24064 13964 24070
rect 13912 24006 13964 24012
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13924 23322 13952 24006
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 13728 23248 13780 23254
rect 13728 23190 13780 23196
rect 13910 23216 13966 23225
rect 13556 22188 13676 22216
rect 13268 22160 13320 22166
rect 13174 22128 13230 22137
rect 13268 22102 13320 22108
rect 13174 22063 13230 22072
rect 13084 21548 13136 21554
rect 13084 21490 13136 21496
rect 12992 21480 13044 21486
rect 12992 21422 13044 21428
rect 13004 21146 13032 21422
rect 12992 21140 13044 21146
rect 12992 21082 13044 21088
rect 12990 21040 13046 21049
rect 12990 20975 13046 20984
rect 13004 19802 13032 20975
rect 13096 20806 13124 21490
rect 13084 20800 13136 20806
rect 13084 20742 13136 20748
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13096 20262 13124 20538
rect 13188 20398 13216 22063
rect 13280 21554 13308 22102
rect 13556 22094 13584 22188
rect 13556 22066 13676 22094
rect 13648 22001 13676 22066
rect 13634 21992 13690 22001
rect 13634 21927 13690 21936
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13312 21244 13620 21253
rect 13312 21242 13318 21244
rect 13374 21242 13398 21244
rect 13454 21242 13478 21244
rect 13534 21242 13558 21244
rect 13614 21242 13620 21244
rect 13374 21190 13376 21242
rect 13556 21190 13558 21242
rect 13312 21188 13318 21190
rect 13374 21188 13398 21190
rect 13454 21188 13478 21190
rect 13534 21188 13558 21190
rect 13614 21188 13620 21190
rect 13312 21179 13620 21188
rect 13544 21072 13596 21078
rect 13542 21040 13544 21049
rect 13596 21040 13598 21049
rect 13542 20975 13598 20984
rect 13544 20936 13596 20942
rect 13544 20878 13596 20884
rect 13556 20777 13584 20878
rect 13542 20768 13598 20777
rect 13542 20703 13598 20712
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13084 20256 13136 20262
rect 13084 20198 13136 20204
rect 13188 20058 13216 20334
rect 13312 20156 13620 20165
rect 13312 20154 13318 20156
rect 13374 20154 13398 20156
rect 13454 20154 13478 20156
rect 13534 20154 13558 20156
rect 13614 20154 13620 20156
rect 13374 20102 13376 20154
rect 13556 20102 13558 20154
rect 13312 20100 13318 20102
rect 13374 20100 13398 20102
rect 13454 20100 13478 20102
rect 13534 20100 13558 20102
rect 13614 20100 13620 20102
rect 13312 20091 13620 20100
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13544 19848 13596 19854
rect 13004 19774 13308 19802
rect 13544 19790 13596 19796
rect 12992 19712 13044 19718
rect 12992 19654 13044 19660
rect 13004 19310 13032 19654
rect 13084 19440 13136 19446
rect 13084 19382 13136 19388
rect 12992 19304 13044 19310
rect 12992 19246 13044 19252
rect 13096 19122 13124 19382
rect 13280 19156 13308 19774
rect 13358 19544 13414 19553
rect 13556 19514 13584 19790
rect 13358 19479 13414 19488
rect 13544 19508 13596 19514
rect 13372 19446 13400 19479
rect 13544 19450 13596 19456
rect 13360 19440 13412 19446
rect 13360 19382 13412 19388
rect 13004 19094 13124 19122
rect 13188 19128 13308 19156
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12912 18358 12940 18566
rect 12900 18352 12952 18358
rect 12900 18294 12952 18300
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12912 15008 12940 18158
rect 13004 17082 13032 19094
rect 13188 17678 13216 19128
rect 13312 19068 13620 19077
rect 13312 19066 13318 19068
rect 13374 19066 13398 19068
rect 13454 19066 13478 19068
rect 13534 19066 13558 19068
rect 13614 19066 13620 19068
rect 13374 19014 13376 19066
rect 13556 19014 13558 19066
rect 13312 19012 13318 19014
rect 13374 19012 13398 19014
rect 13454 19012 13478 19014
rect 13534 19012 13558 19014
rect 13614 19012 13620 19014
rect 13312 19003 13620 19012
rect 13648 18952 13676 21927
rect 13740 21434 13768 23190
rect 13910 23151 13912 23160
rect 13964 23151 13966 23160
rect 13912 23122 13964 23128
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13832 22778 13860 23054
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 13832 21690 13860 22714
rect 13924 22642 13952 23122
rect 13912 22636 13964 22642
rect 13912 22578 13964 22584
rect 13910 22400 13966 22409
rect 13910 22335 13966 22344
rect 13924 22030 13952 22335
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 13740 21406 13860 21434
rect 13728 21344 13780 21350
rect 13832 21321 13860 21406
rect 13728 21286 13780 21292
rect 13818 21312 13874 21321
rect 13740 21128 13768 21286
rect 13818 21247 13874 21256
rect 13740 21100 13860 21128
rect 13832 20992 13860 21100
rect 13556 18924 13676 18952
rect 13740 20964 13860 20992
rect 13556 18222 13584 18924
rect 13634 18320 13690 18329
rect 13634 18255 13690 18264
rect 13544 18216 13596 18222
rect 13544 18158 13596 18164
rect 13312 17980 13620 17989
rect 13312 17978 13318 17980
rect 13374 17978 13398 17980
rect 13454 17978 13478 17980
rect 13534 17978 13558 17980
rect 13614 17978 13620 17980
rect 13374 17926 13376 17978
rect 13556 17926 13558 17978
rect 13312 17924 13318 17926
rect 13374 17924 13398 17926
rect 13454 17924 13478 17926
rect 13534 17924 13558 17926
rect 13614 17924 13620 17926
rect 13312 17915 13620 17924
rect 13176 17672 13228 17678
rect 13176 17614 13228 17620
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17202 13124 17478
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 13004 17054 13124 17082
rect 12992 16992 13044 16998
rect 12992 16934 13044 16940
rect 13004 16522 13032 16934
rect 12992 16516 13044 16522
rect 12992 16458 13044 16464
rect 12992 15020 13044 15026
rect 12912 14980 12992 15008
rect 12912 14929 12940 14980
rect 12992 14962 13044 14968
rect 12898 14920 12954 14929
rect 12898 14855 12954 14864
rect 12992 14272 13044 14278
rect 13096 14260 13124 17054
rect 13176 16992 13228 16998
rect 13176 16934 13228 16940
rect 13188 16590 13216 16934
rect 13312 16892 13620 16901
rect 13312 16890 13318 16892
rect 13374 16890 13398 16892
rect 13454 16890 13478 16892
rect 13534 16890 13558 16892
rect 13614 16890 13620 16892
rect 13374 16838 13376 16890
rect 13556 16838 13558 16890
rect 13312 16836 13318 16838
rect 13374 16836 13398 16838
rect 13454 16836 13478 16838
rect 13534 16836 13558 16838
rect 13614 16836 13620 16838
rect 13312 16827 13620 16836
rect 13176 16584 13228 16590
rect 13176 16526 13228 16532
rect 13174 15872 13230 15881
rect 13174 15807 13230 15816
rect 13188 15570 13216 15807
rect 13312 15804 13620 15813
rect 13312 15802 13318 15804
rect 13374 15802 13398 15804
rect 13454 15802 13478 15804
rect 13534 15802 13558 15804
rect 13614 15802 13620 15804
rect 13374 15750 13376 15802
rect 13556 15750 13558 15802
rect 13312 15748 13318 15750
rect 13374 15748 13398 15750
rect 13454 15748 13478 15750
rect 13534 15748 13558 15750
rect 13614 15748 13620 15750
rect 13312 15739 13620 15748
rect 13176 15564 13228 15570
rect 13176 15506 13228 15512
rect 13648 14958 13676 18255
rect 13740 17882 13768 20964
rect 13820 20800 13872 20806
rect 13820 20742 13872 20748
rect 13832 18766 13860 20742
rect 14016 20346 14044 27968
rect 14200 27962 14228 28018
rect 14384 28014 14412 33322
rect 14476 32042 14504 34167
rect 14568 33930 14596 35022
rect 14556 33924 14608 33930
rect 14556 33866 14608 33872
rect 14556 32768 14608 32774
rect 14556 32710 14608 32716
rect 14568 32298 14596 32710
rect 14556 32292 14608 32298
rect 14556 32234 14608 32240
rect 14476 32014 14596 32042
rect 14464 31952 14516 31958
rect 14464 31894 14516 31900
rect 14372 28008 14424 28014
rect 14200 27934 14320 27962
rect 14372 27950 14424 27956
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14200 27418 14228 27610
rect 14108 27390 14228 27418
rect 14108 27130 14136 27390
rect 14188 27328 14240 27334
rect 14188 27270 14240 27276
rect 14096 27124 14148 27130
rect 14096 27066 14148 27072
rect 14200 26994 14228 27270
rect 14188 26988 14240 26994
rect 14188 26930 14240 26936
rect 14186 25936 14242 25945
rect 14186 25871 14242 25880
rect 14096 25424 14148 25430
rect 14200 25412 14228 25871
rect 14148 25384 14228 25412
rect 14096 25366 14148 25372
rect 14292 25158 14320 27934
rect 14476 27878 14504 31894
rect 14568 30376 14596 32014
rect 14660 30977 14688 35566
rect 14738 34232 14794 34241
rect 14738 34167 14794 34176
rect 14752 33998 14780 34167
rect 14740 33992 14792 33998
rect 14740 33934 14792 33940
rect 14740 33856 14792 33862
rect 14740 33798 14792 33804
rect 14752 33658 14780 33798
rect 14740 33652 14792 33658
rect 14740 33594 14792 33600
rect 14740 33448 14792 33454
rect 14740 33390 14792 33396
rect 14752 32065 14780 33390
rect 14844 32881 14872 38508
rect 15212 38486 15240 38898
rect 15200 38480 15252 38486
rect 15200 38422 15252 38428
rect 15016 38276 15068 38282
rect 15016 38218 15068 38224
rect 15028 34542 15056 38218
rect 15108 37868 15160 37874
rect 15108 37810 15160 37816
rect 15120 37466 15148 37810
rect 15108 37460 15160 37466
rect 15108 37402 15160 37408
rect 15212 36666 15240 38422
rect 15488 38214 15516 39374
rect 16224 39273 16252 39510
rect 16210 39264 16266 39273
rect 15784 39196 16092 39205
rect 16210 39199 16266 39208
rect 15784 39194 15790 39196
rect 15846 39194 15870 39196
rect 15926 39194 15950 39196
rect 16006 39194 16030 39196
rect 16086 39194 16092 39196
rect 15846 39142 15848 39194
rect 16028 39142 16030 39194
rect 15784 39140 15790 39142
rect 15846 39140 15870 39142
rect 15926 39140 15950 39142
rect 16006 39140 16030 39142
rect 16086 39140 16092 39142
rect 15784 39131 16092 39140
rect 15476 38208 15528 38214
rect 15476 38150 15528 38156
rect 15568 38208 15620 38214
rect 15568 38150 15620 38156
rect 15580 38010 15608 38150
rect 15784 38108 16092 38117
rect 15784 38106 15790 38108
rect 15846 38106 15870 38108
rect 15926 38106 15950 38108
rect 16006 38106 16030 38108
rect 16086 38106 16092 38108
rect 15846 38054 15848 38106
rect 16028 38054 16030 38106
rect 15784 38052 15790 38054
rect 15846 38052 15870 38054
rect 15926 38052 15950 38054
rect 16006 38052 16030 38054
rect 16086 38052 16092 38054
rect 15658 38040 15714 38049
rect 15784 38043 16092 38052
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15568 38004 15620 38010
rect 15714 37984 15884 37992
rect 15658 37975 15884 37984
rect 15672 37964 15884 37975
rect 15568 37946 15620 37952
rect 15488 37890 15516 37946
rect 15292 37868 15344 37874
rect 15488 37862 15792 37890
rect 15856 37874 15884 37964
rect 15292 37810 15344 37816
rect 15304 37777 15332 37810
rect 15290 37768 15346 37777
rect 15290 37703 15346 37712
rect 15568 37256 15620 37262
rect 15568 37198 15620 37204
rect 15580 36786 15608 37198
rect 15764 37108 15792 37862
rect 15844 37868 15896 37874
rect 15844 37810 15896 37816
rect 15844 37120 15896 37126
rect 15764 37080 15844 37108
rect 15844 37062 15896 37068
rect 15784 37020 16092 37029
rect 15784 37018 15790 37020
rect 15846 37018 15870 37020
rect 15926 37018 15950 37020
rect 16006 37018 16030 37020
rect 16086 37018 16092 37020
rect 15846 36966 15848 37018
rect 16028 36966 16030 37018
rect 15784 36964 15790 36966
rect 15846 36964 15870 36966
rect 15926 36964 15950 36966
rect 16006 36964 16030 36966
rect 16086 36964 16092 36966
rect 15784 36955 16092 36964
rect 15384 36780 15436 36786
rect 15384 36722 15436 36728
rect 15568 36780 15620 36786
rect 15568 36722 15620 36728
rect 15120 36638 15240 36666
rect 15120 35873 15148 36638
rect 15200 36576 15252 36582
rect 15200 36518 15252 36524
rect 15106 35864 15162 35873
rect 15106 35799 15162 35808
rect 15212 35766 15240 36518
rect 15292 36372 15344 36378
rect 15292 36314 15344 36320
rect 15304 36106 15332 36314
rect 15292 36100 15344 36106
rect 15292 36042 15344 36048
rect 15396 35834 15424 36722
rect 15476 36576 15528 36582
rect 15476 36518 15528 36524
rect 15488 36378 15516 36518
rect 15476 36372 15528 36378
rect 15476 36314 15528 36320
rect 15476 36032 15528 36038
rect 15580 36009 15608 36722
rect 16212 36100 16264 36106
rect 16212 36042 16264 36048
rect 15476 35974 15528 35980
rect 15566 36000 15622 36009
rect 15488 35834 15516 35974
rect 15566 35935 15622 35944
rect 15384 35828 15436 35834
rect 15384 35770 15436 35776
rect 15476 35828 15528 35834
rect 15476 35770 15528 35776
rect 15200 35760 15252 35766
rect 15200 35702 15252 35708
rect 15382 35728 15438 35737
rect 15580 35714 15608 35935
rect 15784 35932 16092 35941
rect 15784 35930 15790 35932
rect 15846 35930 15870 35932
rect 15926 35930 15950 35932
rect 16006 35930 16030 35932
rect 16086 35930 16092 35932
rect 15846 35878 15848 35930
rect 16028 35878 16030 35930
rect 15784 35876 15790 35878
rect 15846 35876 15870 35878
rect 15926 35876 15950 35878
rect 16006 35876 16030 35878
rect 16086 35876 16092 35878
rect 15784 35867 16092 35876
rect 16224 35766 16252 36042
rect 16212 35760 16264 35766
rect 15382 35663 15438 35672
rect 15488 35686 15608 35714
rect 15842 35728 15898 35737
rect 15200 35624 15252 35630
rect 15200 35566 15252 35572
rect 15016 34536 15068 34542
rect 15016 34478 15068 34484
rect 15016 34400 15068 34406
rect 15016 34342 15068 34348
rect 15028 33833 15056 34342
rect 15212 34241 15240 35566
rect 15292 34944 15344 34950
rect 15292 34886 15344 34892
rect 15198 34232 15254 34241
rect 15198 34167 15254 34176
rect 15200 33856 15252 33862
rect 15014 33824 15070 33833
rect 15200 33798 15252 33804
rect 15014 33759 15070 33768
rect 15028 33658 15056 33759
rect 15016 33652 15068 33658
rect 15016 33594 15068 33600
rect 15212 33522 15240 33798
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15016 33448 15068 33454
rect 15016 33390 15068 33396
rect 14830 32872 14886 32881
rect 14830 32807 14886 32816
rect 14832 32768 14884 32774
rect 14832 32710 14884 32716
rect 14844 32298 14872 32710
rect 14832 32292 14884 32298
rect 14832 32234 14884 32240
rect 14738 32056 14794 32065
rect 14738 31991 14794 32000
rect 14740 31952 14792 31958
rect 14740 31894 14792 31900
rect 14752 31657 14780 31894
rect 14738 31648 14794 31657
rect 14738 31583 14794 31592
rect 14844 31396 14872 32234
rect 15028 31793 15056 33390
rect 15304 32434 15332 34886
rect 15396 34649 15424 35663
rect 15488 34785 15516 35686
rect 16212 35702 16264 35708
rect 15842 35663 15898 35672
rect 15856 35222 15884 35663
rect 15844 35216 15896 35222
rect 15658 35184 15714 35193
rect 15580 35142 15658 35170
rect 15474 34776 15530 34785
rect 15474 34711 15530 34720
rect 15382 34640 15438 34649
rect 15382 34575 15438 34584
rect 15384 34196 15436 34202
rect 15384 34138 15436 34144
rect 15396 33114 15424 34138
rect 15580 33538 15608 35142
rect 15844 35158 15896 35164
rect 15658 35119 15714 35128
rect 16212 35012 16264 35018
rect 16212 34954 16264 34960
rect 15784 34844 16092 34853
rect 15784 34842 15790 34844
rect 15846 34842 15870 34844
rect 15926 34842 15950 34844
rect 16006 34842 16030 34844
rect 16086 34842 16092 34844
rect 15846 34790 15848 34842
rect 16028 34790 16030 34842
rect 15784 34788 15790 34790
rect 15846 34788 15870 34790
rect 15926 34788 15950 34790
rect 16006 34788 16030 34790
rect 16086 34788 16092 34790
rect 15784 34779 16092 34788
rect 15660 33992 15712 33998
rect 15660 33934 15712 33940
rect 15672 33697 15700 33934
rect 15784 33756 16092 33765
rect 15784 33754 15790 33756
rect 15846 33754 15870 33756
rect 15926 33754 15950 33756
rect 16006 33754 16030 33756
rect 16086 33754 16092 33756
rect 15846 33702 15848 33754
rect 16028 33702 16030 33754
rect 15784 33700 15790 33702
rect 15846 33700 15870 33702
rect 15926 33700 15950 33702
rect 16006 33700 16030 33702
rect 16086 33700 16092 33702
rect 15658 33688 15714 33697
rect 15784 33691 16092 33700
rect 15658 33623 15714 33632
rect 15488 33510 15608 33538
rect 16120 33516 16172 33522
rect 15384 33108 15436 33114
rect 15384 33050 15436 33056
rect 15292 32428 15344 32434
rect 15292 32370 15344 32376
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 15120 31929 15148 32302
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 15106 31920 15162 31929
rect 15106 31855 15108 31864
rect 15160 31855 15162 31864
rect 15108 31826 15160 31832
rect 15014 31784 15070 31793
rect 15014 31719 15070 31728
rect 14924 31680 14976 31686
rect 14924 31622 14976 31628
rect 14936 31414 14964 31622
rect 14752 31368 14872 31396
rect 14924 31408 14976 31414
rect 14646 30968 14702 30977
rect 14646 30903 14702 30912
rect 14752 30870 14780 31368
rect 14924 31350 14976 31356
rect 15212 31260 15240 31962
rect 14844 31232 15240 31260
rect 14740 30864 14792 30870
rect 14740 30806 14792 30812
rect 14648 30388 14700 30394
rect 14568 30348 14648 30376
rect 14568 29850 14596 30348
rect 14648 30330 14700 30336
rect 14844 30054 14872 31232
rect 15016 30932 15068 30938
rect 15016 30874 15068 30880
rect 15028 30734 15056 30874
rect 15304 30802 15332 32370
rect 15488 32280 15516 33510
rect 16120 33458 16172 33464
rect 16132 33114 16160 33458
rect 16120 33108 16172 33114
rect 16120 33050 16172 33056
rect 16224 33017 16252 34954
rect 16210 33008 16266 33017
rect 16210 32943 16266 32952
rect 15660 32904 15712 32910
rect 15660 32846 15712 32852
rect 15396 32252 15516 32280
rect 15292 30796 15344 30802
rect 15292 30738 15344 30744
rect 15016 30728 15068 30734
rect 15016 30670 15068 30676
rect 15108 30728 15160 30734
rect 15160 30676 15332 30682
rect 15108 30670 15332 30676
rect 14832 30048 14884 30054
rect 14832 29990 14884 29996
rect 14556 29844 14608 29850
rect 14556 29786 14608 29792
rect 14556 29640 14608 29646
rect 14556 29582 14608 29588
rect 14568 29510 14596 29582
rect 14648 29572 14700 29578
rect 14648 29514 14700 29520
rect 14556 29504 14608 29510
rect 14556 29446 14608 29452
rect 14556 29096 14608 29102
rect 14660 29084 14688 29514
rect 14740 29300 14792 29306
rect 14740 29242 14792 29248
rect 14608 29056 14688 29084
rect 14556 29038 14608 29044
rect 14752 28994 14780 29242
rect 14568 28966 14780 28994
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14372 26308 14424 26314
rect 14372 26250 14424 26256
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14280 25152 14332 25158
rect 14280 25094 14332 25100
rect 14108 24274 14136 25094
rect 14280 24744 14332 24750
rect 14280 24686 14332 24692
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14108 23633 14136 24006
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14094 23624 14150 23633
rect 14094 23559 14150 23568
rect 14200 22658 14228 23802
rect 14292 23526 14320 24686
rect 14384 23746 14412 26250
rect 14476 25129 14504 27814
rect 14568 26874 14596 28966
rect 14844 28914 14872 29990
rect 15028 29594 15056 30670
rect 15120 30654 15332 30670
rect 15108 30252 15160 30258
rect 15108 30194 15160 30200
rect 15120 29753 15148 30194
rect 15106 29744 15162 29753
rect 15106 29679 15162 29688
rect 14752 28886 14872 28914
rect 14936 29566 15056 29594
rect 14648 28416 14700 28422
rect 14648 28358 14700 28364
rect 14660 28014 14688 28358
rect 14648 28008 14700 28014
rect 14648 27950 14700 27956
rect 14752 27614 14780 28886
rect 14832 28620 14884 28626
rect 14936 28608 14964 29566
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 14884 28580 14964 28608
rect 14832 28562 14884 28568
rect 14752 27586 14872 27614
rect 14568 26846 14688 26874
rect 14556 26784 14608 26790
rect 14556 26726 14608 26732
rect 14568 26382 14596 26726
rect 14556 26376 14608 26382
rect 14556 26318 14608 26324
rect 14660 25838 14688 26846
rect 14738 26752 14794 26761
rect 14738 26687 14794 26696
rect 14752 26042 14780 26687
rect 14844 26586 14872 27586
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14740 26036 14792 26042
rect 14740 25978 14792 25984
rect 14648 25832 14700 25838
rect 14648 25774 14700 25780
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14462 25120 14518 25129
rect 14462 25055 14518 25064
rect 14462 24304 14518 24313
rect 14518 24262 14596 24290
rect 14462 24239 14518 24248
rect 14568 24206 14596 24262
rect 14752 24206 14780 25638
rect 14832 25152 14884 25158
rect 14832 25094 14884 25100
rect 14844 24818 14872 25094
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14740 24200 14792 24206
rect 14740 24142 14792 24148
rect 14568 23866 14596 24142
rect 14844 24052 14872 24754
rect 14660 24024 14872 24052
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14384 23718 14596 23746
rect 14280 23520 14332 23526
rect 14280 23462 14332 23468
rect 14108 22630 14228 22658
rect 14108 20942 14136 22630
rect 14188 22432 14240 22438
rect 14188 22374 14240 22380
rect 14200 21554 14228 22374
rect 14188 21548 14240 21554
rect 14240 21508 14320 21536
rect 14188 21490 14240 21496
rect 14096 20936 14148 20942
rect 14096 20878 14148 20884
rect 14108 20466 14136 20878
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14096 20460 14148 20466
rect 14096 20402 14148 20408
rect 13924 20318 14044 20346
rect 14096 20324 14148 20330
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 13820 18352 13872 18358
rect 13820 18294 13872 18300
rect 13728 17876 13780 17882
rect 13728 17818 13780 17824
rect 13832 17678 13860 18294
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13740 16590 13768 17614
rect 13924 17202 13952 20318
rect 14096 20266 14148 20272
rect 14002 20224 14058 20233
rect 14002 20159 14058 20168
rect 14016 19378 14044 20159
rect 14108 20058 14136 20266
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14096 19848 14148 19854
rect 14096 19790 14148 19796
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 14002 19272 14058 19281
rect 14108 19258 14136 19790
rect 14058 19230 14136 19258
rect 14002 19207 14058 19216
rect 14108 18630 14136 19230
rect 14096 18624 14148 18630
rect 14096 18566 14148 18572
rect 14108 18222 14136 18566
rect 14096 18216 14148 18222
rect 14096 18158 14148 18164
rect 14108 17746 14136 18158
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13912 17196 13964 17202
rect 13912 17138 13964 17144
rect 13728 16584 13780 16590
rect 13728 16526 13780 16532
rect 13268 14952 13320 14958
rect 13044 14232 13124 14260
rect 13188 14912 13268 14940
rect 12992 14214 13044 14220
rect 12900 14000 12952 14006
rect 12900 13942 12952 13948
rect 12912 11830 12940 13942
rect 13004 13190 13032 14214
rect 13188 14074 13216 14912
rect 13268 14894 13320 14900
rect 13636 14952 13688 14958
rect 13636 14894 13688 14900
rect 13740 14770 13768 16526
rect 13820 15904 13872 15910
rect 13820 15846 13872 15852
rect 13832 15094 13860 15846
rect 13924 15638 13952 17138
rect 14016 16250 14044 17478
rect 14200 17134 14228 20810
rect 14292 18834 14320 21508
rect 14464 21344 14516 21350
rect 14464 21286 14516 21292
rect 14476 20942 14504 21286
rect 14464 20936 14516 20942
rect 14464 20878 14516 20884
rect 14476 20602 14504 20878
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14384 19718 14412 19790
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14280 18828 14332 18834
rect 14280 18770 14332 18776
rect 14278 18456 14334 18465
rect 14278 18391 14334 18400
rect 14292 18358 14320 18391
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14384 17762 14412 19450
rect 14292 17734 14412 17762
rect 14188 17128 14240 17134
rect 14188 17070 14240 17076
rect 14096 17060 14148 17066
rect 14096 17002 14148 17008
rect 14108 16794 14136 17002
rect 14200 16794 14228 17070
rect 14096 16788 14148 16794
rect 14096 16730 14148 16736
rect 14188 16788 14240 16794
rect 14188 16730 14240 16736
rect 14004 16244 14056 16250
rect 14004 16186 14056 16192
rect 14292 16130 14320 17734
rect 14372 17672 14424 17678
rect 14372 17614 14424 17620
rect 14200 16102 14320 16130
rect 14096 15972 14148 15978
rect 14096 15914 14148 15920
rect 13912 15632 13964 15638
rect 13912 15574 13964 15580
rect 14108 15502 14136 15914
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13820 15088 13872 15094
rect 13820 15030 13872 15036
rect 13820 14952 13872 14958
rect 13820 14894 13872 14900
rect 13648 14742 13768 14770
rect 13312 14716 13620 14725
rect 13312 14714 13318 14716
rect 13374 14714 13398 14716
rect 13454 14714 13478 14716
rect 13534 14714 13558 14716
rect 13614 14714 13620 14716
rect 13374 14662 13376 14714
rect 13556 14662 13558 14714
rect 13312 14660 13318 14662
rect 13374 14660 13398 14662
rect 13454 14660 13478 14662
rect 13534 14660 13558 14662
rect 13614 14660 13620 14662
rect 13312 14651 13620 14660
rect 13648 14618 13676 14742
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13312 13628 13620 13637
rect 13312 13626 13318 13628
rect 13374 13626 13398 13628
rect 13454 13626 13478 13628
rect 13534 13626 13558 13628
rect 13614 13626 13620 13628
rect 13374 13574 13376 13626
rect 13556 13574 13558 13626
rect 13312 13572 13318 13574
rect 13374 13572 13398 13574
rect 13454 13572 13478 13574
rect 13534 13572 13558 13574
rect 13614 13572 13620 13574
rect 13312 13563 13620 13572
rect 13648 13308 13676 14554
rect 13832 14006 13860 14894
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13648 13280 13860 13308
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13004 12850 13032 13126
rect 13096 12918 13124 13194
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13004 12102 13032 12786
rect 13096 12238 13124 12854
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12900 11824 12952 11830
rect 12900 11766 12952 11772
rect 12912 10606 12940 11766
rect 13004 11014 13032 12038
rect 13096 11393 13124 12038
rect 13082 11384 13138 11393
rect 13082 11319 13138 11328
rect 13084 11280 13136 11286
rect 13084 11222 13136 11228
rect 12992 11008 13044 11014
rect 12992 10950 13044 10956
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12806 10432 12862 10441
rect 12806 10367 12862 10376
rect 12624 10260 12676 10266
rect 13096 10248 13124 11222
rect 13188 10742 13216 12718
rect 13312 12540 13620 12549
rect 13312 12538 13318 12540
rect 13374 12538 13398 12540
rect 13454 12538 13478 12540
rect 13534 12538 13558 12540
rect 13614 12538 13620 12540
rect 13374 12486 13376 12538
rect 13556 12486 13558 12538
rect 13312 12484 13318 12486
rect 13374 12484 13398 12486
rect 13454 12484 13478 12486
rect 13534 12484 13558 12486
rect 13614 12484 13620 12486
rect 13312 12475 13620 12484
rect 13740 12238 13768 12922
rect 13832 12481 13860 13280
rect 13924 13274 13952 15438
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14016 14482 14044 14962
rect 14108 14770 14136 15438
rect 14200 14872 14228 16102
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 14292 15201 14320 15982
rect 14278 15192 14334 15201
rect 14278 15127 14334 15136
rect 14200 14844 14320 14872
rect 14108 14742 14228 14770
rect 14004 14476 14056 14482
rect 14004 14418 14056 14424
rect 14016 13870 14044 14418
rect 14200 14090 14228 14742
rect 14292 14385 14320 14844
rect 14384 14414 14412 17614
rect 14476 17610 14504 20402
rect 14568 17814 14596 23718
rect 14660 22681 14688 24024
rect 14832 23724 14884 23730
rect 14832 23666 14884 23672
rect 14738 23624 14794 23633
rect 14844 23610 14872 23666
rect 14794 23582 14872 23610
rect 14738 23559 14794 23568
rect 14844 23118 14872 23582
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14646 22672 14702 22681
rect 14646 22607 14702 22616
rect 14648 22432 14700 22438
rect 14648 22374 14700 22380
rect 14660 22001 14688 22374
rect 14740 22228 14792 22234
rect 14740 22170 14792 22176
rect 14752 22137 14780 22170
rect 14738 22128 14794 22137
rect 14738 22063 14794 22072
rect 14646 21992 14702 22001
rect 14936 21978 14964 28580
rect 15028 28422 15056 29446
rect 15198 29064 15254 29073
rect 15198 28999 15254 29008
rect 15212 28914 15240 28999
rect 15120 28886 15240 28914
rect 15016 28416 15068 28422
rect 15016 28358 15068 28364
rect 15016 26308 15068 26314
rect 15016 26250 15068 26256
rect 15028 26042 15056 26250
rect 15016 26036 15068 26042
rect 15016 25978 15068 25984
rect 15120 25974 15148 28886
rect 15198 28656 15254 28665
rect 15198 28591 15254 28600
rect 15212 28558 15240 28591
rect 15200 28552 15252 28558
rect 15200 28494 15252 28500
rect 15200 28416 15252 28422
rect 15200 28358 15252 28364
rect 15212 26994 15240 28358
rect 15304 28218 15332 30654
rect 15292 28212 15344 28218
rect 15292 28154 15344 28160
rect 15304 28082 15332 28154
rect 15292 28076 15344 28082
rect 15292 28018 15344 28024
rect 15200 26988 15252 26994
rect 15200 26930 15252 26936
rect 15212 26382 15240 26930
rect 15292 26784 15344 26790
rect 15292 26726 15344 26732
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 15304 26234 15332 26726
rect 15212 26206 15332 26234
rect 15108 25968 15160 25974
rect 15108 25910 15160 25916
rect 15108 25832 15160 25838
rect 15108 25774 15160 25780
rect 15014 24168 15070 24177
rect 15014 24103 15070 24112
rect 15028 23866 15056 24103
rect 15016 23860 15068 23866
rect 15016 23802 15068 23808
rect 15028 22030 15056 23802
rect 15120 23066 15148 25774
rect 15212 23633 15240 26206
rect 15292 25832 15344 25838
rect 15292 25774 15344 25780
rect 15304 25362 15332 25774
rect 15292 25356 15344 25362
rect 15292 25298 15344 25304
rect 15292 25152 15344 25158
rect 15292 25094 15344 25100
rect 15304 24614 15332 25094
rect 15292 24608 15344 24614
rect 15292 24550 15344 24556
rect 15396 24177 15424 32252
rect 15672 32026 15700 32846
rect 16224 32774 16252 32943
rect 16212 32768 16264 32774
rect 16212 32710 16264 32716
rect 15784 32668 16092 32677
rect 15784 32666 15790 32668
rect 15846 32666 15870 32668
rect 15926 32666 15950 32668
rect 16006 32666 16030 32668
rect 16086 32666 16092 32668
rect 15846 32614 15848 32666
rect 16028 32614 16030 32666
rect 15784 32612 15790 32614
rect 15846 32612 15870 32614
rect 15926 32612 15950 32614
rect 16006 32612 16030 32614
rect 16086 32612 16092 32614
rect 15784 32603 16092 32612
rect 16316 32552 16344 41074
rect 16408 40934 16436 41126
rect 16396 40928 16448 40934
rect 16396 40870 16448 40876
rect 16488 40928 16540 40934
rect 16488 40870 16540 40876
rect 16500 40458 16528 40870
rect 16488 40452 16540 40458
rect 16488 40394 16540 40400
rect 16592 39982 16620 41239
rect 16776 41206 16804 41550
rect 16868 41478 16896 42638
rect 16948 42628 17000 42634
rect 16948 42570 17000 42576
rect 16960 41698 16988 42570
rect 17132 42220 17184 42226
rect 17132 42162 17184 42168
rect 16960 41670 17080 41698
rect 16948 41608 17000 41614
rect 16948 41550 17000 41556
rect 16856 41472 16908 41478
rect 16856 41414 16908 41420
rect 16960 41274 16988 41550
rect 16948 41268 17000 41274
rect 16948 41210 17000 41216
rect 16764 41200 16816 41206
rect 17052 41177 17080 41670
rect 16764 41142 16816 41148
rect 17038 41168 17094 41177
rect 16672 41132 16724 41138
rect 16672 41074 16724 41080
rect 16856 41132 16908 41138
rect 16856 41074 16908 41080
rect 16948 41132 17000 41138
rect 17038 41103 17094 41112
rect 16948 41074 17000 41080
rect 16684 40186 16712 41074
rect 16764 40996 16816 41002
rect 16764 40938 16816 40944
rect 16776 40730 16804 40938
rect 16764 40724 16816 40730
rect 16764 40666 16816 40672
rect 16764 40520 16816 40526
rect 16764 40462 16816 40468
rect 16672 40180 16724 40186
rect 16672 40122 16724 40128
rect 16488 39976 16540 39982
rect 16488 39918 16540 39924
rect 16580 39976 16632 39982
rect 16580 39918 16632 39924
rect 16672 39976 16724 39982
rect 16672 39918 16724 39924
rect 16500 39273 16528 39918
rect 16684 39658 16712 39918
rect 16592 39630 16712 39658
rect 16592 39574 16620 39630
rect 16580 39568 16632 39574
rect 16580 39510 16632 39516
rect 16486 39264 16542 39273
rect 16486 39199 16542 39208
rect 16396 39092 16448 39098
rect 16396 39034 16448 39040
rect 16408 38554 16436 39034
rect 16776 38654 16804 40462
rect 16868 39522 16896 41074
rect 16960 40390 16988 41074
rect 17040 41064 17092 41070
rect 17040 41006 17092 41012
rect 17052 40662 17080 41006
rect 17040 40656 17092 40662
rect 17040 40598 17092 40604
rect 16948 40384 17000 40390
rect 16948 40326 17000 40332
rect 17040 40384 17092 40390
rect 17040 40326 17092 40332
rect 16948 40112 17000 40118
rect 16946 40080 16948 40089
rect 17000 40080 17002 40089
rect 16946 40015 17002 40024
rect 16868 39494 16988 39522
rect 16856 39432 16908 39438
rect 16856 39374 16908 39380
rect 16868 39302 16896 39374
rect 16856 39296 16908 39302
rect 16856 39238 16908 39244
rect 16856 38956 16908 38962
rect 16856 38898 16908 38904
rect 16592 38626 16804 38654
rect 16396 38548 16448 38554
rect 16396 38490 16448 38496
rect 16488 37800 16540 37806
rect 16488 37742 16540 37748
rect 16500 37262 16528 37742
rect 16488 37256 16540 37262
rect 16488 37198 16540 37204
rect 16500 35086 16528 37198
rect 16592 35494 16620 38626
rect 16672 37800 16724 37806
rect 16868 37788 16896 38898
rect 16724 37760 16896 37788
rect 16672 37742 16724 37748
rect 16672 36712 16724 36718
rect 16672 36654 16724 36660
rect 16684 36174 16712 36654
rect 16672 36168 16724 36174
rect 16672 36110 16724 36116
rect 16580 35488 16632 35494
rect 16580 35430 16632 35436
rect 16488 35080 16540 35086
rect 16408 35028 16488 35034
rect 16408 35022 16540 35028
rect 16408 35006 16528 35022
rect 16408 34950 16436 35006
rect 16396 34944 16448 34950
rect 16396 34886 16448 34892
rect 16394 34640 16450 34649
rect 16684 34610 16712 36110
rect 16960 35329 16988 39494
rect 17052 36825 17080 40326
rect 17144 39522 17172 42162
rect 17236 41750 17264 43250
rect 17328 42770 17356 43574
rect 17420 43466 17448 43846
rect 17512 43602 17540 44540
rect 17696 44010 17724 44540
rect 17696 43994 17816 44010
rect 17696 43988 17828 43994
rect 17696 43982 17776 43988
rect 17776 43930 17828 43936
rect 17512 43574 17632 43602
rect 17420 43450 17540 43466
rect 17420 43444 17552 43450
rect 17420 43438 17500 43444
rect 17500 43386 17552 43392
rect 17500 43308 17552 43314
rect 17500 43250 17552 43256
rect 17512 42838 17540 43250
rect 17500 42832 17552 42838
rect 17500 42774 17552 42780
rect 17316 42764 17368 42770
rect 17316 42706 17368 42712
rect 17604 42650 17632 43574
rect 17880 42770 17908 44540
rect 17960 43308 18012 43314
rect 17960 43250 18012 43256
rect 17972 42906 18000 43250
rect 18064 43110 18092 44540
rect 18144 43308 18196 43314
rect 18144 43250 18196 43256
rect 18052 43104 18104 43110
rect 18052 43046 18104 43052
rect 17960 42900 18012 42906
rect 17960 42842 18012 42848
rect 17868 42764 17920 42770
rect 17868 42706 17920 42712
rect 17774 42664 17830 42673
rect 17500 42628 17552 42634
rect 17604 42622 17774 42650
rect 17774 42599 17830 42608
rect 17500 42570 17552 42576
rect 17316 42220 17368 42226
rect 17316 42162 17368 42168
rect 17224 41744 17276 41750
rect 17224 41686 17276 41692
rect 17224 41608 17276 41614
rect 17224 41550 17276 41556
rect 17236 41274 17264 41550
rect 17224 41268 17276 41274
rect 17224 41210 17276 41216
rect 17224 41132 17276 41138
rect 17224 41074 17276 41080
rect 17236 40730 17264 41074
rect 17224 40724 17276 40730
rect 17224 40666 17276 40672
rect 17328 40186 17356 42162
rect 17406 41712 17462 41721
rect 17406 41647 17462 41656
rect 17420 41478 17448 41647
rect 17408 41472 17460 41478
rect 17408 41414 17460 41420
rect 17512 41274 17540 42570
rect 17776 42560 17828 42566
rect 17776 42502 17828 42508
rect 17682 42120 17738 42129
rect 17682 42055 17738 42064
rect 17696 41614 17724 42055
rect 17592 41608 17644 41614
rect 17592 41550 17644 41556
rect 17684 41608 17736 41614
rect 17684 41550 17736 41556
rect 17500 41268 17552 41274
rect 17500 41210 17552 41216
rect 17408 41200 17460 41206
rect 17408 41142 17460 41148
rect 17420 40526 17448 41142
rect 17500 41132 17552 41138
rect 17500 41074 17552 41080
rect 17408 40520 17460 40526
rect 17408 40462 17460 40468
rect 17316 40180 17368 40186
rect 17316 40122 17368 40128
rect 17144 39494 17264 39522
rect 17132 39432 17184 39438
rect 17132 39374 17184 39380
rect 17144 38729 17172 39374
rect 17236 39137 17264 39494
rect 17408 39432 17460 39438
rect 17408 39374 17460 39380
rect 17316 39296 17368 39302
rect 17316 39238 17368 39244
rect 17222 39128 17278 39137
rect 17222 39063 17278 39072
rect 17130 38720 17186 38729
rect 17130 38655 17186 38664
rect 17328 37505 17356 39238
rect 17420 39098 17448 39374
rect 17408 39092 17460 39098
rect 17408 39034 17460 39040
rect 17314 37496 17370 37505
rect 17314 37431 17370 37440
rect 17316 37120 17368 37126
rect 17316 37062 17368 37068
rect 17038 36816 17094 36825
rect 17038 36751 17094 36760
rect 17052 36650 17080 36751
rect 17040 36644 17092 36650
rect 17040 36586 17092 36592
rect 17224 36032 17276 36038
rect 17224 35974 17276 35980
rect 17040 35692 17092 35698
rect 17040 35634 17092 35640
rect 16946 35320 17002 35329
rect 17052 35290 17080 35634
rect 17236 35630 17264 35974
rect 17328 35873 17356 37062
rect 17408 36168 17460 36174
rect 17408 36110 17460 36116
rect 17314 35864 17370 35873
rect 17420 35834 17448 36110
rect 17314 35799 17370 35808
rect 17408 35828 17460 35834
rect 17408 35770 17460 35776
rect 17224 35624 17276 35630
rect 17224 35566 17276 35572
rect 17132 35488 17184 35494
rect 17132 35430 17184 35436
rect 17224 35488 17276 35494
rect 17224 35430 17276 35436
rect 16946 35255 17002 35264
rect 17040 35284 17092 35290
rect 17040 35226 17092 35232
rect 16394 34575 16450 34584
rect 16672 34604 16724 34610
rect 16132 32524 16344 32552
rect 15752 32292 15804 32298
rect 15752 32234 15804 32240
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 15488 31482 15516 31826
rect 15764 31686 15792 32234
rect 15844 32224 15896 32230
rect 15844 32166 15896 32172
rect 15936 32224 15988 32230
rect 15936 32166 15988 32172
rect 15856 31890 15884 32166
rect 15844 31884 15896 31890
rect 15844 31826 15896 31832
rect 15948 31686 15976 32166
rect 15752 31680 15804 31686
rect 15672 31640 15752 31668
rect 15476 31476 15528 31482
rect 15476 31418 15528 31424
rect 15672 31385 15700 31640
rect 15752 31622 15804 31628
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 15784 31580 16092 31589
rect 15784 31578 15790 31580
rect 15846 31578 15870 31580
rect 15926 31578 15950 31580
rect 16006 31578 16030 31580
rect 16086 31578 16092 31580
rect 15846 31526 15848 31578
rect 16028 31526 16030 31578
rect 15784 31524 15790 31526
rect 15846 31524 15870 31526
rect 15926 31524 15950 31526
rect 16006 31524 16030 31526
rect 16086 31524 16092 31526
rect 15784 31515 16092 31524
rect 15474 31376 15530 31385
rect 15474 31311 15530 31320
rect 15658 31376 15714 31385
rect 15658 31311 15714 31320
rect 15488 31192 15516 31311
rect 15568 31204 15620 31210
rect 15488 31164 15568 31192
rect 15568 31146 15620 31152
rect 16132 30802 16160 32524
rect 16212 32428 16264 32434
rect 16212 32370 16264 32376
rect 16224 30938 16252 32370
rect 16408 32314 16436 34575
rect 16672 34546 16724 34552
rect 16948 34604 17000 34610
rect 16948 34546 17000 34552
rect 16580 34468 16632 34474
rect 16580 34410 16632 34416
rect 16592 34202 16620 34410
rect 16580 34196 16632 34202
rect 16580 34138 16632 34144
rect 16580 33924 16632 33930
rect 16580 33866 16632 33872
rect 16592 33658 16620 33866
rect 16580 33652 16632 33658
rect 16580 33594 16632 33600
rect 16684 32570 16712 34546
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16764 34060 16816 34066
rect 16764 34002 16816 34008
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 16580 32428 16632 32434
rect 16580 32370 16632 32376
rect 16408 32286 16528 32314
rect 16592 32298 16620 32370
rect 16396 32224 16448 32230
rect 16396 32166 16448 32172
rect 16304 31680 16356 31686
rect 16304 31622 16356 31628
rect 16316 31346 16344 31622
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16302 31104 16358 31113
rect 16302 31039 16358 31048
rect 16212 30932 16264 30938
rect 16212 30874 16264 30880
rect 15660 30796 15712 30802
rect 15580 30756 15660 30784
rect 15474 30152 15530 30161
rect 15474 30087 15530 30096
rect 15488 29510 15516 30087
rect 15580 29714 15608 30756
rect 15660 30738 15712 30744
rect 16120 30796 16172 30802
rect 16316 30784 16344 31039
rect 16120 30738 16172 30744
rect 16224 30756 16344 30784
rect 15658 30696 15714 30705
rect 16224 30648 16252 30756
rect 16408 30734 16436 32166
rect 16396 30728 16448 30734
rect 16396 30670 16448 30676
rect 15658 30631 15714 30640
rect 15568 29708 15620 29714
rect 15568 29650 15620 29656
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15476 28960 15528 28966
rect 15476 28902 15528 28908
rect 15488 28626 15516 28902
rect 15476 28620 15528 28626
rect 15476 28562 15528 28568
rect 15476 28008 15528 28014
rect 15476 27950 15528 27956
rect 15488 27674 15516 27950
rect 15476 27668 15528 27674
rect 15476 27610 15528 27616
rect 15476 27532 15528 27538
rect 15580 27520 15608 29650
rect 15672 27713 15700 30631
rect 16132 30620 16252 30648
rect 16304 30660 16356 30666
rect 15784 30492 16092 30501
rect 15784 30490 15790 30492
rect 15846 30490 15870 30492
rect 15926 30490 15950 30492
rect 16006 30490 16030 30492
rect 16086 30490 16092 30492
rect 15846 30438 15848 30490
rect 16028 30438 16030 30490
rect 15784 30436 15790 30438
rect 15846 30436 15870 30438
rect 15926 30436 15950 30438
rect 16006 30436 16030 30438
rect 16086 30436 16092 30438
rect 15784 30427 16092 30436
rect 15784 29404 16092 29413
rect 15784 29402 15790 29404
rect 15846 29402 15870 29404
rect 15926 29402 15950 29404
rect 16006 29402 16030 29404
rect 16086 29402 16092 29404
rect 15846 29350 15848 29402
rect 16028 29350 16030 29402
rect 15784 29348 15790 29350
rect 15846 29348 15870 29350
rect 15926 29348 15950 29350
rect 16006 29348 16030 29350
rect 16086 29348 16092 29350
rect 15784 29339 16092 29348
rect 15784 28316 16092 28325
rect 15784 28314 15790 28316
rect 15846 28314 15870 28316
rect 15926 28314 15950 28316
rect 16006 28314 16030 28316
rect 16086 28314 16092 28316
rect 15846 28262 15848 28314
rect 16028 28262 16030 28314
rect 15784 28260 15790 28262
rect 15846 28260 15870 28262
rect 15926 28260 15950 28262
rect 16006 28260 16030 28262
rect 16086 28260 16092 28262
rect 15784 28251 16092 28260
rect 15658 27704 15714 27713
rect 15658 27639 15714 27648
rect 15528 27492 15608 27520
rect 15476 27474 15528 27480
rect 15476 25968 15528 25974
rect 15476 25910 15528 25916
rect 15382 24168 15438 24177
rect 15382 24103 15438 24112
rect 15198 23624 15254 23633
rect 15198 23559 15254 23568
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23322 15240 23462
rect 15200 23316 15252 23322
rect 15200 23258 15252 23264
rect 15200 23180 15252 23186
rect 15384 23180 15436 23186
rect 15252 23140 15384 23168
rect 15200 23122 15252 23128
rect 15384 23122 15436 23128
rect 15120 23038 15332 23066
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15108 22500 15160 22506
rect 15108 22442 15160 22448
rect 15120 22234 15148 22442
rect 15108 22228 15160 22234
rect 15108 22170 15160 22176
rect 14646 21927 14702 21936
rect 14752 21950 14964 21978
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 14660 21078 14688 21927
rect 14648 21072 14700 21078
rect 14648 21014 14700 21020
rect 14648 19712 14700 19718
rect 14648 19654 14700 19660
rect 14660 19310 14688 19654
rect 14648 19304 14700 19310
rect 14648 19246 14700 19252
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14464 17604 14516 17610
rect 14464 17546 14516 17552
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14476 16153 14504 17274
rect 14752 16250 14780 21950
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14844 20448 14872 21830
rect 15028 21729 15056 21966
rect 15014 21720 15070 21729
rect 15014 21655 15070 21664
rect 15212 21570 15240 22918
rect 15304 21978 15332 23038
rect 15488 22094 15516 25910
rect 15580 25838 15608 27492
rect 15784 27228 16092 27237
rect 15784 27226 15790 27228
rect 15846 27226 15870 27228
rect 15926 27226 15950 27228
rect 16006 27226 16030 27228
rect 16086 27226 16092 27228
rect 15846 27174 15848 27226
rect 16028 27174 16030 27226
rect 15784 27172 15790 27174
rect 15846 27172 15870 27174
rect 15926 27172 15950 27174
rect 16006 27172 16030 27174
rect 16086 27172 16092 27174
rect 15784 27163 16092 27172
rect 15660 26240 15712 26246
rect 15660 26182 15712 26188
rect 15568 25832 15620 25838
rect 15568 25774 15620 25780
rect 15568 25152 15620 25158
rect 15566 25120 15568 25129
rect 15620 25120 15622 25129
rect 15566 25055 15622 25064
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15580 24410 15608 24550
rect 15568 24404 15620 24410
rect 15568 24346 15620 24352
rect 15672 24070 15700 26182
rect 15784 26140 16092 26149
rect 15784 26138 15790 26140
rect 15846 26138 15870 26140
rect 15926 26138 15950 26140
rect 16006 26138 16030 26140
rect 16086 26138 16092 26140
rect 15846 26086 15848 26138
rect 16028 26086 16030 26138
rect 15784 26084 15790 26086
rect 15846 26084 15870 26086
rect 15926 26084 15950 26086
rect 16006 26084 16030 26086
rect 16086 26084 16092 26086
rect 15784 26075 16092 26084
rect 16132 25922 16160 30620
rect 16304 30602 16356 30608
rect 16210 30424 16266 30433
rect 16316 30394 16344 30602
rect 16210 30359 16266 30368
rect 16304 30388 16356 30394
rect 16224 26450 16252 30359
rect 16304 30330 16356 30336
rect 16500 30274 16528 32286
rect 16580 32292 16632 32298
rect 16580 32234 16632 32240
rect 16580 31680 16632 31686
rect 16580 31622 16632 31628
rect 16592 31278 16620 31622
rect 16580 31272 16632 31278
rect 16580 31214 16632 31220
rect 16592 30802 16620 31214
rect 16580 30796 16632 30802
rect 16580 30738 16632 30744
rect 16500 30246 16620 30274
rect 16684 30258 16712 32506
rect 16776 31736 16804 34002
rect 16868 32892 16896 34138
rect 16960 33998 16988 34546
rect 16948 33992 17000 33998
rect 16948 33934 17000 33940
rect 17144 33862 17172 35430
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 17130 33416 17186 33425
rect 17130 33351 17186 33360
rect 16868 32864 17080 32892
rect 16856 32768 16908 32774
rect 16856 32710 16908 32716
rect 16868 31890 16896 32710
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16856 31748 16908 31754
rect 16776 31708 16856 31736
rect 16856 31690 16908 31696
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16776 30938 16804 31078
rect 16764 30932 16816 30938
rect 16764 30874 16816 30880
rect 16764 30592 16816 30598
rect 16764 30534 16816 30540
rect 16304 28484 16356 28490
rect 16304 28426 16356 28432
rect 16316 28082 16344 28426
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16304 27396 16356 27402
rect 16304 27338 16356 27344
rect 16316 27130 16344 27338
rect 16304 27124 16356 27130
rect 16304 27066 16356 27072
rect 16592 26874 16620 30246
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16684 28558 16712 30194
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16776 28370 16804 30534
rect 16316 26846 16620 26874
rect 16684 28342 16804 28370
rect 16212 26444 16264 26450
rect 16212 26386 16264 26392
rect 16210 26208 16266 26217
rect 16210 26143 16266 26152
rect 16224 26042 16252 26143
rect 16212 26036 16264 26042
rect 16212 25978 16264 25984
rect 16132 25894 16252 25922
rect 16224 25430 16252 25894
rect 16212 25424 16264 25430
rect 16212 25366 16264 25372
rect 16210 25256 16266 25265
rect 16210 25191 16266 25200
rect 15784 25052 16092 25061
rect 15784 25050 15790 25052
rect 15846 25050 15870 25052
rect 15926 25050 15950 25052
rect 16006 25050 16030 25052
rect 16086 25050 16092 25052
rect 15846 24998 15848 25050
rect 16028 24998 16030 25050
rect 15784 24996 15790 24998
rect 15846 24996 15870 24998
rect 15926 24996 15950 24998
rect 16006 24996 16030 24998
rect 16086 24996 16092 24998
rect 15784 24987 16092 24996
rect 16120 24676 16172 24682
rect 16120 24618 16172 24624
rect 15660 24064 15712 24070
rect 15660 24006 15712 24012
rect 15784 23964 16092 23973
rect 15784 23962 15790 23964
rect 15846 23962 15870 23964
rect 15926 23962 15950 23964
rect 16006 23962 16030 23964
rect 16086 23962 16092 23964
rect 15846 23910 15848 23962
rect 16028 23910 16030 23962
rect 15784 23908 15790 23910
rect 15846 23908 15870 23910
rect 15926 23908 15950 23910
rect 16006 23908 16030 23910
rect 16086 23908 16092 23910
rect 15784 23899 16092 23908
rect 16132 23866 16160 24618
rect 16120 23860 16172 23866
rect 16120 23802 16172 23808
rect 15750 23624 15806 23633
rect 15750 23559 15806 23568
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15672 23118 15700 23462
rect 15660 23112 15712 23118
rect 15660 23054 15712 23060
rect 15764 22964 15792 23559
rect 16120 23316 16172 23322
rect 16120 23258 16172 23264
rect 15672 22936 15792 22964
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15580 22574 15608 22714
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 15488 22066 15608 22094
rect 15304 21950 15516 21978
rect 15292 21888 15344 21894
rect 15292 21830 15344 21836
rect 15028 21554 15240 21570
rect 15016 21548 15240 21554
rect 15068 21542 15240 21548
rect 15016 21490 15068 21496
rect 14924 21344 14976 21350
rect 15304 21298 15332 21830
rect 15384 21480 15436 21486
rect 15384 21422 15436 21428
rect 14924 21286 14976 21292
rect 14936 20913 14964 21286
rect 15120 21270 15332 21298
rect 15016 20936 15068 20942
rect 14922 20904 14978 20913
rect 15016 20878 15068 20884
rect 14922 20839 14978 20848
rect 15028 20806 15056 20878
rect 15016 20800 15068 20806
rect 15016 20742 15068 20748
rect 14924 20460 14976 20466
rect 14844 20420 14924 20448
rect 14924 20402 14976 20408
rect 14936 19961 14964 20402
rect 14922 19952 14978 19961
rect 14922 19887 14978 19896
rect 14832 19780 14884 19786
rect 14832 19722 14884 19728
rect 14844 19378 14872 19722
rect 15028 19394 15056 20742
rect 15120 19514 15148 21270
rect 15292 20936 15344 20942
rect 15396 20924 15424 21422
rect 15344 20896 15424 20924
rect 15292 20878 15344 20884
rect 15304 20602 15332 20878
rect 15292 20596 15344 20602
rect 15292 20538 15344 20544
rect 15384 19916 15436 19922
rect 15488 19904 15516 21950
rect 15436 19876 15516 19904
rect 15384 19858 15436 19864
rect 15290 19816 15346 19825
rect 15474 19816 15530 19825
rect 15346 19774 15424 19802
rect 15290 19751 15346 19760
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14936 19366 15056 19394
rect 14936 18986 14964 19366
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15028 19174 15056 19246
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14936 18958 15056 18986
rect 14922 18864 14978 18873
rect 14922 18799 14924 18808
rect 14976 18799 14978 18808
rect 14924 18770 14976 18776
rect 14924 18692 14976 18698
rect 14924 18634 14976 18640
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14844 17202 14872 17546
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14832 16992 14884 16998
rect 14832 16934 14884 16940
rect 14740 16244 14792 16250
rect 14660 16204 14740 16232
rect 14462 16144 14518 16153
rect 14462 16079 14518 16088
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14372 14408 14424 14414
rect 14278 14376 14334 14385
rect 14372 14350 14424 14356
rect 14278 14311 14334 14320
rect 14108 14062 14228 14090
rect 14004 13864 14056 13870
rect 14004 13806 14056 13812
rect 14108 13530 14136 14062
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 14096 13524 14148 13530
rect 14096 13466 14148 13472
rect 14200 13462 14228 13942
rect 14188 13456 14240 13462
rect 14188 13398 14240 13404
rect 14188 13320 14240 13326
rect 13924 13246 14044 13274
rect 14188 13262 14240 13268
rect 13912 13184 13964 13190
rect 13912 13126 13964 13132
rect 13818 12472 13874 12481
rect 13924 12442 13952 13126
rect 14016 12850 14044 13246
rect 14004 12844 14056 12850
rect 14004 12786 14056 12792
rect 13818 12407 13874 12416
rect 13912 12436 13964 12442
rect 13912 12378 13964 12384
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 14094 12336 14150 12345
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13636 12164 13688 12170
rect 13636 12106 13688 12112
rect 13266 11928 13322 11937
rect 13266 11863 13322 11872
rect 13280 11762 13308 11863
rect 13268 11756 13320 11762
rect 13268 11698 13320 11704
rect 13312 11452 13620 11461
rect 13312 11450 13318 11452
rect 13374 11450 13398 11452
rect 13454 11450 13478 11452
rect 13534 11450 13558 11452
rect 13614 11450 13620 11452
rect 13374 11398 13376 11450
rect 13556 11398 13558 11450
rect 13312 11396 13318 11398
rect 13374 11396 13398 11398
rect 13454 11396 13478 11398
rect 13534 11396 13558 11398
rect 13614 11396 13620 11398
rect 13312 11387 13620 11396
rect 13176 10736 13228 10742
rect 13176 10678 13228 10684
rect 13176 10600 13228 10606
rect 13176 10542 13228 10548
rect 12624 10202 12676 10208
rect 12820 10220 13124 10248
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 12544 9897 12572 9930
rect 12820 9897 12848 10220
rect 13188 10130 13216 10542
rect 13312 10364 13620 10373
rect 13312 10362 13318 10364
rect 13374 10362 13398 10364
rect 13454 10362 13478 10364
rect 13534 10362 13558 10364
rect 13614 10362 13620 10364
rect 13374 10310 13376 10362
rect 13556 10310 13558 10362
rect 13312 10308 13318 10310
rect 13374 10308 13398 10310
rect 13454 10308 13478 10310
rect 13534 10308 13558 10310
rect 13614 10308 13620 10310
rect 13312 10299 13620 10308
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 12530 9888 12586 9897
rect 12530 9823 12586 9832
rect 12806 9888 12862 9897
rect 12806 9823 12862 9832
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12532 9172 12584 9178
rect 12532 9114 12584 9120
rect 12544 8129 12572 9114
rect 12636 8922 12664 9454
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12808 9376 12860 9382
rect 12808 9318 12860 9324
rect 12728 9110 12756 9318
rect 12716 9104 12768 9110
rect 12716 9046 12768 9052
rect 12636 8894 12756 8922
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8498 12664 8774
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12530 8120 12586 8129
rect 12530 8055 12586 8064
rect 12440 7948 12492 7954
rect 12440 7890 12492 7896
rect 12636 7868 12664 8434
rect 12728 8022 12756 8894
rect 12820 8537 12848 9318
rect 12912 9042 12940 10066
rect 13082 9888 13138 9897
rect 13082 9823 13138 9832
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12992 8968 13044 8974
rect 12898 8936 12954 8945
rect 12954 8916 12992 8922
rect 12954 8910 13044 8916
rect 12954 8894 13032 8910
rect 12898 8871 12954 8880
rect 12806 8528 12862 8537
rect 12990 8528 13046 8537
rect 12806 8463 12862 8472
rect 12912 8486 12990 8514
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12530 7848 12586 7857
rect 12636 7840 12756 7868
rect 12530 7783 12586 7792
rect 12254 7304 12310 7313
rect 12254 7239 12310 7248
rect 12440 7268 12492 7274
rect 12440 7210 12492 7216
rect 12164 6996 12216 7002
rect 12348 6996 12400 7002
rect 12164 6938 12216 6944
rect 12268 6956 12348 6984
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12084 6458 12112 6734
rect 12072 6452 12124 6458
rect 12072 6394 12124 6400
rect 12268 6338 12296 6956
rect 12348 6938 12400 6944
rect 12452 6712 12480 7210
rect 12360 6684 12480 6712
rect 12360 6458 12388 6684
rect 12544 6610 12572 7783
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12636 7041 12664 7482
rect 12728 7410 12756 7840
rect 12820 7410 12848 7890
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12728 7177 12756 7346
rect 12714 7168 12770 7177
rect 12714 7103 12770 7112
rect 12622 7032 12678 7041
rect 12622 6967 12678 6976
rect 12716 6792 12768 6798
rect 12714 6760 12716 6769
rect 12768 6760 12770 6769
rect 12624 6724 12676 6730
rect 12714 6695 12770 6704
rect 12624 6666 12676 6672
rect 12452 6582 12572 6610
rect 12348 6452 12400 6458
rect 12348 6394 12400 6400
rect 12084 6310 12296 6338
rect 12346 6352 12402 6361
rect 12084 5794 12112 6310
rect 12346 6287 12348 6296
rect 12400 6287 12402 6296
rect 12348 6258 12400 6264
rect 12346 6216 12402 6225
rect 11808 5222 11928 5250
rect 11992 5766 12112 5794
rect 12176 6174 12346 6202
rect 12176 5778 12204 6174
rect 12346 6151 12402 6160
rect 12452 6118 12480 6582
rect 12636 6474 12664 6666
rect 12544 6446 12664 6474
rect 12806 6488 12862 6497
rect 12716 6452 12768 6458
rect 12544 6186 12572 6446
rect 12806 6423 12862 6432
rect 12716 6394 12768 6400
rect 12532 6180 12584 6186
rect 12532 6122 12584 6128
rect 12440 6112 12492 6118
rect 12440 6054 12492 6060
rect 12624 6112 12676 6118
rect 12624 6054 12676 6060
rect 12346 5944 12402 5953
rect 12256 5908 12308 5914
rect 12346 5879 12402 5888
rect 12256 5850 12308 5856
rect 12164 5772 12216 5778
rect 11520 5102 11572 5108
rect 11610 5128 11666 5137
rect 11610 5063 11666 5072
rect 11702 4856 11758 4865
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11612 4820 11664 4826
rect 11702 4791 11758 4800
rect 11612 4762 11664 4768
rect 11428 4684 11480 4690
rect 11428 4626 11480 4632
rect 11440 4593 11468 4626
rect 11624 4593 11652 4762
rect 11426 4584 11482 4593
rect 11426 4519 11482 4528
rect 11610 4584 11666 4593
rect 11610 4519 11666 4528
rect 11716 4282 11744 4791
rect 11704 4276 11756 4282
rect 11440 4236 11652 4264
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11164 3896 11284 3924
rect 11336 3936 11388 3942
rect 11164 3670 11192 3896
rect 11336 3878 11388 3884
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 11242 3632 11298 3641
rect 11060 3596 11112 3602
rect 11242 3567 11298 3576
rect 11060 3538 11112 3544
rect 10600 3334 10652 3340
rect 10690 3360 10746 3369
rect 10612 2938 10640 3334
rect 10690 3295 10746 3304
rect 10839 3292 11147 3301
rect 10839 3290 10845 3292
rect 10901 3290 10925 3292
rect 10981 3290 11005 3292
rect 11061 3290 11085 3292
rect 11141 3290 11147 3292
rect 10901 3238 10903 3290
rect 11083 3238 11085 3290
rect 10839 3236 10845 3238
rect 10901 3236 10925 3238
rect 10981 3236 11005 3238
rect 11061 3236 11085 3238
rect 11141 3236 11147 3238
rect 10839 3227 11147 3236
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 10782 3088 10838 3097
rect 10782 3023 10784 3032
rect 10836 3023 10838 3032
rect 10784 2994 10836 3000
rect 10612 2910 10824 2938
rect 10692 2848 10744 2854
rect 10690 2816 10692 2825
rect 10744 2816 10746 2825
rect 10520 2746 10640 2774
rect 10690 2751 10746 2760
rect 10612 2666 10640 2746
rect 10612 2638 10732 2666
rect 10336 2604 10548 2632
rect 10520 2530 10548 2604
rect 10520 2502 10640 2530
rect 10244 2366 10364 2394
rect 10336 2360 10364 2366
rect 10336 2332 10456 2360
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10140 1760 10192 1766
rect 10140 1702 10192 1708
rect 10048 1406 10100 1412
rect 9772 1352 9824 1358
rect 10048 1348 10100 1354
rect 10152 1306 10180 1702
rect 9824 1300 9904 1306
rect 9772 1294 9904 1300
rect 9784 1278 9904 1294
rect 9680 1216 9732 1222
rect 9680 1158 9732 1164
rect 9772 1216 9824 1222
rect 9772 1158 9824 1164
rect 9692 678 9720 1158
rect 9680 672 9732 678
rect 9680 614 9732 620
rect 9784 160 9812 1158
rect 9876 728 9904 1278
rect 10060 1278 10180 1306
rect 10060 1193 10088 1278
rect 10244 1193 10272 2246
rect 10324 1488 10376 1494
rect 10324 1430 10376 1436
rect 10046 1184 10102 1193
rect 10046 1119 10102 1128
rect 10230 1184 10286 1193
rect 10230 1119 10286 1128
rect 10046 1048 10102 1057
rect 10230 1048 10286 1057
rect 10102 1006 10180 1034
rect 10046 983 10102 992
rect 10046 912 10102 921
rect 10046 847 10102 856
rect 10060 814 10088 847
rect 10048 808 10100 814
rect 10048 750 10100 756
rect 9876 700 9996 728
rect 9968 160 9996 700
rect 10152 160 10180 1006
rect 10230 983 10286 992
rect 10244 882 10272 983
rect 10232 876 10284 882
rect 10232 818 10284 824
rect 10230 776 10286 785
rect 10230 711 10232 720
rect 10284 711 10286 720
rect 10232 682 10284 688
rect 10336 160 10364 1430
rect 10428 202 10456 2332
rect 10508 1760 10560 1766
rect 10508 1702 10560 1708
rect 10416 196 10468 202
rect 7470 96 7526 105
rect 7470 31 7526 40
rect 7562 -300 7618 160
rect 7746 -300 7802 160
rect 7930 -300 7986 160
rect 8114 -300 8170 160
rect 8298 -300 8354 160
rect 8482 -300 8538 160
rect 8574 96 8630 105
rect 8666 82 8722 160
rect 8630 54 8722 82
rect 8574 31 8630 40
rect 8666 -300 8722 54
rect 8850 -300 8906 160
rect 9034 -300 9090 160
rect 9218 -300 9274 160
rect 9402 -300 9458 160
rect 9586 -300 9642 160
rect 9770 -300 9826 160
rect 9954 -300 10010 160
rect 10138 -300 10194 160
rect 10322 -300 10378 160
rect 10520 160 10548 1702
rect 10612 1562 10640 2502
rect 10704 2446 10732 2638
rect 10796 2530 10824 2910
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10888 2689 10916 2790
rect 10874 2680 10930 2689
rect 10874 2615 10930 2624
rect 10980 2530 11008 3130
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11072 2961 11100 2994
rect 11058 2952 11114 2961
rect 11058 2887 11114 2896
rect 11164 2825 11192 2994
rect 11150 2816 11206 2825
rect 11150 2751 11206 2760
rect 10796 2502 11008 2530
rect 11256 2446 11284 3567
rect 10692 2440 10744 2446
rect 11152 2440 11204 2446
rect 10692 2382 10744 2388
rect 11150 2408 11152 2417
rect 11244 2440 11296 2446
rect 11204 2408 11206 2417
rect 11244 2382 11296 2388
rect 11150 2343 11206 2352
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 10839 2204 11147 2213
rect 10839 2202 10845 2204
rect 10901 2202 10925 2204
rect 10981 2202 11005 2204
rect 11061 2202 11085 2204
rect 11141 2202 11147 2204
rect 10901 2150 10903 2202
rect 11083 2150 11085 2202
rect 10839 2148 10845 2150
rect 10901 2148 10925 2150
rect 10981 2148 11005 2150
rect 11061 2148 11085 2150
rect 11141 2148 11147 2150
rect 10839 2139 11147 2148
rect 11152 1896 11204 1902
rect 11152 1838 11204 1844
rect 10876 1828 10928 1834
rect 10876 1770 10928 1776
rect 10692 1760 10744 1766
rect 10692 1702 10744 1708
rect 10600 1556 10652 1562
rect 10600 1498 10652 1504
rect 10600 1216 10652 1222
rect 10600 1158 10652 1164
rect 10612 1018 10640 1158
rect 10600 1012 10652 1018
rect 10600 954 10652 960
rect 10600 604 10652 610
rect 10600 546 10652 552
rect 10416 138 10468 144
rect 10506 -300 10562 160
rect 10612 82 10640 546
rect 10704 252 10732 1702
rect 10888 1601 10916 1770
rect 10874 1592 10930 1601
rect 10874 1527 10930 1536
rect 11060 1352 11112 1358
rect 11164 1306 11192 1838
rect 11256 1358 11284 2246
rect 11348 2038 11376 3878
rect 11440 3738 11468 4236
rect 11624 4162 11652 4236
rect 11704 4218 11756 4224
rect 11624 4146 11744 4162
rect 11520 4140 11572 4146
rect 11624 4140 11756 4146
rect 11624 4134 11704 4140
rect 11520 4082 11572 4088
rect 11704 4082 11756 4088
rect 11532 3738 11560 4082
rect 11808 4010 11836 5222
rect 11886 5128 11942 5137
rect 11886 5063 11942 5072
rect 11900 4690 11928 5063
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11992 4622 12020 5766
rect 12164 5714 12216 5720
rect 12176 5302 12204 5714
rect 12268 5370 12296 5850
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 12360 5114 12388 5879
rect 12440 5704 12492 5710
rect 12530 5672 12586 5681
rect 12492 5652 12530 5658
rect 12440 5646 12530 5652
rect 12452 5630 12530 5646
rect 12530 5607 12586 5616
rect 12636 5284 12664 6054
rect 12728 5914 12756 6394
rect 12716 5908 12768 5914
rect 12716 5850 12768 5856
rect 12714 5808 12770 5817
rect 12714 5743 12770 5752
rect 12176 5086 12388 5114
rect 12452 5256 12664 5284
rect 12070 4856 12126 4865
rect 12070 4791 12126 4800
rect 11980 4616 12032 4622
rect 11980 4558 12032 4564
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11978 4448 12034 4457
rect 11900 4321 11928 4422
rect 11978 4383 12034 4392
rect 11886 4312 11942 4321
rect 11886 4247 11942 4256
rect 11796 4004 11848 4010
rect 11796 3946 11848 3952
rect 11612 3936 11664 3942
rect 11888 3936 11940 3942
rect 11794 3904 11850 3913
rect 11612 3878 11664 3884
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11520 3732 11572 3738
rect 11520 3674 11572 3680
rect 11624 3641 11652 3878
rect 11716 3862 11794 3890
rect 11610 3632 11666 3641
rect 11610 3567 11666 3576
rect 11518 3360 11574 3369
rect 11518 3295 11574 3304
rect 11532 3176 11560 3295
rect 11440 3148 11560 3176
rect 11440 2854 11468 3148
rect 11716 3058 11744 3862
rect 11888 3878 11940 3884
rect 11794 3839 11850 3848
rect 11796 3528 11848 3534
rect 11796 3470 11848 3476
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11612 2984 11664 2990
rect 11702 2952 11758 2961
rect 11664 2932 11702 2938
rect 11612 2926 11702 2932
rect 11624 2910 11702 2926
rect 11702 2887 11758 2896
rect 11428 2848 11480 2854
rect 11428 2790 11480 2796
rect 11428 2644 11480 2650
rect 11428 2586 11480 2592
rect 11520 2644 11572 2650
rect 11520 2586 11572 2592
rect 11440 2446 11468 2586
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11428 2304 11480 2310
rect 11426 2272 11428 2281
rect 11480 2272 11482 2281
rect 11426 2207 11482 2216
rect 11336 2032 11388 2038
rect 11336 1974 11388 1980
rect 11532 1358 11560 2586
rect 11704 2576 11756 2582
rect 11808 2553 11836 3470
rect 11900 3233 11928 3878
rect 11992 3618 12020 4383
rect 12084 4146 12112 4791
rect 12176 4729 12204 5086
rect 12452 4978 12480 5256
rect 12728 5234 12756 5743
rect 12716 5228 12768 5234
rect 12716 5170 12768 5176
rect 12532 5160 12584 5166
rect 12820 5137 12848 6423
rect 12912 6089 12940 8486
rect 12990 8463 13046 8472
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13004 7886 13032 8366
rect 12992 7880 13044 7886
rect 12992 7822 13044 7828
rect 12992 7404 13044 7410
rect 12992 7346 13044 7352
rect 13004 7002 13032 7346
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 12990 6760 13046 6769
rect 12990 6695 13046 6704
rect 13004 6118 13032 6695
rect 13096 6361 13124 9823
rect 13176 9512 13228 9518
rect 13176 9454 13228 9460
rect 13188 9160 13216 9454
rect 13312 9276 13620 9285
rect 13312 9274 13318 9276
rect 13374 9274 13398 9276
rect 13454 9274 13478 9276
rect 13534 9274 13558 9276
rect 13614 9274 13620 9276
rect 13374 9222 13376 9274
rect 13556 9222 13558 9274
rect 13312 9220 13318 9222
rect 13374 9220 13398 9222
rect 13454 9220 13478 9222
rect 13534 9220 13558 9222
rect 13614 9220 13620 9222
rect 13312 9211 13620 9220
rect 13188 9132 13492 9160
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13188 8430 13216 8910
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13280 8276 13308 8774
rect 13464 8294 13492 9132
rect 13544 8492 13596 8498
rect 13648 8480 13676 12106
rect 13910 11928 13966 11937
rect 13910 11863 13966 11872
rect 13728 11756 13780 11762
rect 13728 11698 13780 11704
rect 13740 11529 13768 11698
rect 13820 11552 13872 11558
rect 13726 11520 13782 11529
rect 13820 11494 13872 11500
rect 13726 11455 13782 11464
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13740 10606 13768 11290
rect 13728 10600 13780 10606
rect 13728 10542 13780 10548
rect 13726 10432 13782 10441
rect 13726 10367 13782 10376
rect 13740 9178 13768 10367
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 13728 8900 13780 8906
rect 13728 8842 13780 8848
rect 13596 8452 13676 8480
rect 13544 8434 13596 8440
rect 13636 8356 13688 8362
rect 13740 8344 13768 8842
rect 13832 8498 13860 11494
rect 13924 11150 13952 11863
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 13912 11008 13964 11014
rect 13912 10950 13964 10956
rect 13924 10674 13952 10950
rect 14016 10674 14044 12310
rect 14094 12271 14096 12280
rect 14148 12271 14150 12280
rect 14096 12242 14148 12248
rect 14200 12238 14228 13262
rect 14280 12912 14332 12918
rect 14280 12854 14332 12860
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14096 11756 14148 11762
rect 14096 11698 14148 11704
rect 14108 11393 14136 11698
rect 14094 11384 14150 11393
rect 14094 11319 14150 11328
rect 14096 11280 14148 11286
rect 14096 11222 14148 11228
rect 14108 10985 14136 11222
rect 14094 10976 14150 10985
rect 14094 10911 14150 10920
rect 14094 10840 14150 10849
rect 14094 10775 14150 10784
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 14004 10668 14056 10674
rect 14004 10610 14056 10616
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 13924 9450 13952 10202
rect 14004 10056 14056 10062
rect 14108 10044 14136 10775
rect 14200 10062 14228 12174
rect 14292 10130 14320 12854
rect 14384 11540 14412 14350
rect 14476 12442 14504 15438
rect 14568 15337 14596 15574
rect 14554 15328 14610 15337
rect 14554 15263 14610 15272
rect 14556 13456 14608 13462
rect 14556 13398 14608 13404
rect 14464 12436 14516 12442
rect 14464 12378 14516 12384
rect 14568 12238 14596 13398
rect 14660 13394 14688 16204
rect 14740 16186 14792 16192
rect 14740 15972 14792 15978
rect 14740 15914 14792 15920
rect 14752 15162 14780 15914
rect 14740 15156 14792 15162
rect 14740 15098 14792 15104
rect 14844 14906 14872 16934
rect 14936 15552 14964 18634
rect 15028 16114 15056 18958
rect 15120 18426 15148 19246
rect 15396 18426 15424 19774
rect 15474 19751 15530 19760
rect 15488 19174 15516 19751
rect 15476 19168 15528 19174
rect 15476 19110 15528 19116
rect 15580 18986 15608 22066
rect 15672 21536 15700 22936
rect 15784 22876 16092 22885
rect 15784 22874 15790 22876
rect 15846 22874 15870 22876
rect 15926 22874 15950 22876
rect 16006 22874 16030 22876
rect 16086 22874 16092 22876
rect 15846 22822 15848 22874
rect 16028 22822 16030 22874
rect 15784 22820 15790 22822
rect 15846 22820 15870 22822
rect 15926 22820 15950 22822
rect 16006 22820 16030 22822
rect 16086 22820 16092 22822
rect 15784 22811 16092 22820
rect 15784 21788 16092 21797
rect 15784 21786 15790 21788
rect 15846 21786 15870 21788
rect 15926 21786 15950 21788
rect 16006 21786 16030 21788
rect 16086 21786 16092 21788
rect 15846 21734 15848 21786
rect 16028 21734 16030 21786
rect 15784 21732 15790 21734
rect 15846 21732 15870 21734
rect 15926 21732 15950 21734
rect 16006 21732 16030 21734
rect 16086 21732 16092 21734
rect 15784 21723 16092 21732
rect 15672 21508 15792 21536
rect 15764 20788 15792 21508
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15948 21146 15976 21286
rect 15936 21140 15988 21146
rect 15936 21082 15988 21088
rect 16132 20890 16160 23258
rect 16224 23254 16252 25191
rect 16212 23248 16264 23254
rect 16212 23190 16264 23196
rect 16316 21894 16344 26846
rect 16580 26444 16632 26450
rect 16580 26386 16632 26392
rect 16396 26308 16448 26314
rect 16396 26250 16448 26256
rect 16408 25838 16436 26250
rect 16488 26240 16540 26246
rect 16488 26182 16540 26188
rect 16396 25832 16448 25838
rect 16396 25774 16448 25780
rect 16396 25492 16448 25498
rect 16396 25434 16448 25440
rect 16408 23610 16436 25434
rect 16500 25294 16528 26182
rect 16592 25362 16620 26386
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16488 25288 16540 25294
rect 16488 25230 16540 25236
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24818 16620 25094
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16408 23582 16620 23610
rect 16592 23361 16620 23582
rect 16578 23352 16634 23361
rect 16578 23287 16634 23296
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16500 22094 16528 22578
rect 16684 22094 16712 28342
rect 16868 28082 16896 31690
rect 16946 31376 17002 31385
rect 16946 31311 17002 31320
rect 16960 31210 16988 31311
rect 16948 31204 17000 31210
rect 16948 31146 17000 31152
rect 16960 29646 16988 31146
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 17052 29209 17080 32864
rect 17144 32570 17172 33351
rect 17236 33114 17264 35430
rect 17408 35080 17460 35086
rect 17314 35048 17370 35057
rect 17408 35022 17460 35028
rect 17314 34983 17370 34992
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17328 32774 17356 34983
rect 17420 32910 17448 35022
rect 17408 32904 17460 32910
rect 17408 32846 17460 32852
rect 17316 32768 17368 32774
rect 17316 32710 17368 32716
rect 17132 32564 17184 32570
rect 17132 32506 17184 32512
rect 17130 32464 17186 32473
rect 17130 32399 17186 32408
rect 17144 30841 17172 32399
rect 17420 31929 17448 32846
rect 17406 31920 17462 31929
rect 17406 31855 17462 31864
rect 17130 30832 17186 30841
rect 17130 30767 17186 30776
rect 17316 30592 17368 30598
rect 17316 30534 17368 30540
rect 17132 30388 17184 30394
rect 17132 30330 17184 30336
rect 17144 29850 17172 30330
rect 17328 30258 17356 30534
rect 17420 30394 17448 31855
rect 17408 30388 17460 30394
rect 17408 30330 17460 30336
rect 17316 30252 17368 30258
rect 17316 30194 17368 30200
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 17038 29200 17094 29209
rect 17038 29135 17094 29144
rect 16856 28076 16908 28082
rect 16856 28018 16908 28024
rect 17144 27878 17172 29786
rect 17316 29232 17368 29238
rect 17316 29174 17368 29180
rect 17132 27872 17184 27878
rect 17132 27814 17184 27820
rect 16948 27464 17000 27470
rect 16948 27406 17000 27412
rect 16960 27130 16988 27406
rect 17040 27328 17092 27334
rect 17040 27270 17092 27276
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 17052 27062 17080 27270
rect 17040 27056 17092 27062
rect 17040 26998 17092 27004
rect 16948 26920 17000 26926
rect 17144 26874 17172 27814
rect 17328 26976 17356 29174
rect 17406 29064 17462 29073
rect 17406 28999 17462 29008
rect 17000 26868 17172 26874
rect 16948 26862 17172 26868
rect 16960 26846 17172 26862
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 16854 26616 16910 26625
rect 16854 26551 16910 26560
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 16776 26042 16804 26318
rect 16764 26036 16816 26042
rect 16764 25978 16816 25984
rect 16868 25910 16896 26551
rect 17052 26382 17080 26726
rect 16948 26376 17000 26382
rect 16948 26318 17000 26324
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 16856 25904 16908 25910
rect 16856 25846 16908 25852
rect 16764 25696 16816 25702
rect 16816 25656 16896 25684
rect 16764 25638 16816 25644
rect 16868 25362 16896 25656
rect 16960 25498 16988 26318
rect 16948 25492 17000 25498
rect 16948 25434 17000 25440
rect 17040 25424 17092 25430
rect 17040 25366 17092 25372
rect 16856 25356 16908 25362
rect 16856 25298 16908 25304
rect 16762 25256 16818 25265
rect 16762 25191 16818 25200
rect 16776 22794 16804 25191
rect 16868 24750 16896 25298
rect 16946 24848 17002 24857
rect 16946 24783 17002 24792
rect 16856 24744 16908 24750
rect 16856 24686 16908 24692
rect 16776 22766 16896 22794
rect 16764 22704 16816 22710
rect 16764 22646 16816 22652
rect 16408 22066 16528 22094
rect 16592 22066 16712 22094
rect 16776 22094 16804 22646
rect 16868 22273 16896 22766
rect 16854 22264 16910 22273
rect 16960 22234 16988 24783
rect 16854 22199 16910 22208
rect 16948 22228 17000 22234
rect 16948 22170 17000 22176
rect 16776 22066 16896 22094
rect 16408 21962 16436 22066
rect 16396 21956 16448 21962
rect 16396 21898 16448 21904
rect 16304 21888 16356 21894
rect 16304 21830 16356 21836
rect 16486 21448 16542 21457
rect 16592 21434 16620 22066
rect 16764 22024 16816 22030
rect 16542 21406 16620 21434
rect 16684 21984 16764 22012
rect 16486 21383 16542 21392
rect 16302 21040 16358 21049
rect 16302 20975 16358 20984
rect 16132 20862 16252 20890
rect 15672 20760 15792 20788
rect 16120 20800 16172 20806
rect 15672 19718 15700 20760
rect 16120 20742 16172 20748
rect 15784 20700 16092 20709
rect 15784 20698 15790 20700
rect 15846 20698 15870 20700
rect 15926 20698 15950 20700
rect 16006 20698 16030 20700
rect 16086 20698 16092 20700
rect 15846 20646 15848 20698
rect 16028 20646 16030 20698
rect 15784 20644 15790 20646
rect 15846 20644 15870 20646
rect 15926 20644 15950 20646
rect 16006 20644 16030 20646
rect 16086 20644 16092 20646
rect 15784 20635 16092 20644
rect 16132 20602 16160 20742
rect 16120 20596 16172 20602
rect 16120 20538 16172 20544
rect 16028 20528 16080 20534
rect 16224 20482 16252 20862
rect 16080 20476 16252 20482
rect 16028 20470 16252 20476
rect 16040 20454 16252 20470
rect 15660 19712 15712 19718
rect 15660 19654 15712 19660
rect 16212 19712 16264 19718
rect 16212 19654 16264 19660
rect 15784 19612 16092 19621
rect 15784 19610 15790 19612
rect 15846 19610 15870 19612
rect 15926 19610 15950 19612
rect 16006 19610 16030 19612
rect 16086 19610 16092 19612
rect 15846 19558 15848 19610
rect 16028 19558 16030 19610
rect 15784 19556 15790 19558
rect 15846 19556 15870 19558
rect 15926 19556 15950 19558
rect 16006 19556 16030 19558
rect 16086 19556 16092 19558
rect 15784 19547 16092 19556
rect 15660 19508 15712 19514
rect 15660 19450 15712 19456
rect 15488 18958 15608 18986
rect 15108 18420 15160 18426
rect 15108 18362 15160 18368
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15384 18284 15436 18290
rect 15384 18226 15436 18232
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15120 16998 15148 18158
rect 15200 17536 15252 17542
rect 15200 17478 15252 17484
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15212 17134 15240 17478
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 15108 16992 15160 16998
rect 15108 16934 15160 16940
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15198 16552 15254 16561
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15016 15564 15068 15570
rect 14936 15524 15016 15552
rect 15016 15506 15068 15512
rect 14922 15328 14978 15337
rect 14922 15263 14978 15272
rect 14752 14878 14872 14906
rect 14752 14414 14780 14878
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14740 14408 14792 14414
rect 14844 14385 14872 14758
rect 14936 14618 14964 15263
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 15028 14521 15056 15506
rect 15014 14512 15070 14521
rect 15014 14447 15070 14456
rect 15016 14408 15068 14414
rect 14740 14350 14792 14356
rect 14830 14376 14886 14385
rect 15120 14385 15148 16526
rect 15198 16487 15254 16496
rect 15212 16250 15240 16487
rect 15200 16244 15252 16250
rect 15200 16186 15252 16192
rect 15304 16114 15332 17478
rect 15396 17320 15424 18226
rect 15488 18193 15516 18958
rect 15568 18828 15620 18834
rect 15568 18770 15620 18776
rect 15474 18184 15530 18193
rect 15474 18119 15530 18128
rect 15580 17882 15608 18770
rect 15672 18170 15700 19450
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15856 18766 15884 19110
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15784 18524 16092 18533
rect 15784 18522 15790 18524
rect 15846 18522 15870 18524
rect 15926 18522 15950 18524
rect 16006 18522 16030 18524
rect 16086 18522 16092 18524
rect 15846 18470 15848 18522
rect 16028 18470 16030 18522
rect 15784 18468 15790 18470
rect 15846 18468 15870 18470
rect 15926 18468 15950 18470
rect 16006 18468 16030 18470
rect 16086 18468 16092 18470
rect 15784 18459 16092 18468
rect 15672 18142 15792 18170
rect 15764 17954 15792 18142
rect 15672 17926 15792 17954
rect 15568 17876 15620 17882
rect 15568 17818 15620 17824
rect 15476 17332 15528 17338
rect 15396 17292 15476 17320
rect 15476 17274 15528 17280
rect 15384 17128 15436 17134
rect 15382 17096 15384 17105
rect 15436 17096 15438 17105
rect 15382 17031 15438 17040
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15394 16584 15446 16590
rect 15394 16526 15446 16532
rect 15292 16108 15344 16114
rect 15292 16050 15344 16056
rect 15396 15706 15424 16526
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15212 15570 15240 15642
rect 15200 15564 15252 15570
rect 15200 15506 15252 15512
rect 15292 15496 15344 15502
rect 15292 15438 15344 15444
rect 15198 15192 15254 15201
rect 15198 15127 15254 15136
rect 15212 14822 15240 15127
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15016 14350 15068 14356
rect 15106 14376 15162 14385
rect 14830 14311 14886 14320
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 13462 14780 14214
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14660 12850 14688 13330
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14738 12608 14794 12617
rect 14660 12374 14688 12582
rect 14738 12543 14794 12552
rect 14648 12368 14700 12374
rect 14648 12310 14700 12316
rect 14556 12232 14608 12238
rect 14556 12174 14608 12180
rect 14464 11552 14516 11558
rect 14384 11512 14464 11540
rect 14384 11150 14412 11512
rect 14464 11494 14516 11500
rect 14568 11370 14596 12174
rect 14646 11792 14702 11801
rect 14646 11727 14702 11736
rect 14476 11342 14596 11370
rect 14372 11144 14424 11150
rect 14372 11086 14424 11092
rect 14280 10124 14332 10130
rect 14280 10066 14332 10072
rect 14056 10016 14136 10044
rect 14004 9998 14056 10004
rect 13912 9444 13964 9450
rect 13912 9386 13964 9392
rect 13924 9217 13952 9386
rect 14002 9344 14058 9353
rect 14002 9279 14058 9288
rect 13910 9208 13966 9217
rect 13910 9143 13966 9152
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13688 8316 13768 8344
rect 13636 8298 13688 8304
rect 13188 8248 13308 8276
rect 13452 8288 13504 8294
rect 13188 6984 13216 8248
rect 13452 8230 13504 8236
rect 13312 8188 13620 8197
rect 13312 8186 13318 8188
rect 13374 8186 13398 8188
rect 13454 8186 13478 8188
rect 13534 8186 13558 8188
rect 13614 8186 13620 8188
rect 13374 8134 13376 8186
rect 13556 8134 13558 8186
rect 13312 8132 13318 8134
rect 13374 8132 13398 8134
rect 13454 8132 13478 8134
rect 13534 8132 13558 8134
rect 13614 8132 13620 8134
rect 13312 8123 13620 8132
rect 13740 7936 13768 8316
rect 13924 8090 13952 8774
rect 14016 8265 14044 9279
rect 14002 8256 14058 8265
rect 14002 8191 14058 8200
rect 14002 8120 14058 8129
rect 13912 8084 13964 8090
rect 14002 8055 14058 8064
rect 13912 8026 13964 8032
rect 13820 7948 13872 7954
rect 13740 7908 13820 7936
rect 13820 7890 13872 7896
rect 14016 7834 14044 8055
rect 13832 7806 14044 7834
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13312 7100 13620 7109
rect 13312 7098 13318 7100
rect 13374 7098 13398 7100
rect 13454 7098 13478 7100
rect 13534 7098 13558 7100
rect 13614 7098 13620 7100
rect 13374 7046 13376 7098
rect 13556 7046 13558 7098
rect 13312 7044 13318 7046
rect 13374 7044 13398 7046
rect 13454 7044 13478 7046
rect 13534 7044 13558 7046
rect 13614 7044 13620 7046
rect 13312 7035 13620 7044
rect 13188 6956 13492 6984
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13268 6792 13320 6798
rect 13268 6734 13320 6740
rect 13082 6352 13138 6361
rect 13082 6287 13138 6296
rect 13280 6236 13308 6734
rect 13372 6322 13400 6802
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13096 6208 13308 6236
rect 12992 6112 13044 6118
rect 12898 6080 12954 6089
rect 12992 6054 13044 6060
rect 12898 6015 12954 6024
rect 13096 5846 13124 6208
rect 13464 6100 13492 6956
rect 13648 6798 13676 7142
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6390 13768 6734
rect 13728 6384 13780 6390
rect 13634 6352 13690 6361
rect 13728 6326 13780 6332
rect 13634 6287 13690 6296
rect 13188 6072 13492 6100
rect 13084 5840 13136 5846
rect 13084 5782 13136 5788
rect 12900 5704 12952 5710
rect 13188 5702 13216 6072
rect 13312 6012 13620 6021
rect 13312 6010 13318 6012
rect 13374 6010 13398 6012
rect 13454 6010 13478 6012
rect 13534 6010 13558 6012
rect 13614 6010 13620 6012
rect 13374 5958 13376 6010
rect 13556 5958 13558 6010
rect 13312 5956 13318 5958
rect 13374 5956 13398 5958
rect 13454 5956 13478 5958
rect 13534 5956 13558 5958
rect 13614 5956 13620 5958
rect 13312 5947 13620 5956
rect 13648 5896 13676 6287
rect 13751 6180 13803 6186
rect 12900 5646 12952 5652
rect 13096 5674 13216 5702
rect 13372 5868 13676 5896
rect 13740 6128 13751 6168
rect 13740 6122 13803 6128
rect 12912 5409 12940 5646
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12898 5400 12954 5409
rect 12898 5335 12954 5344
rect 12532 5102 12584 5108
rect 12806 5128 12862 5137
rect 12360 4950 12480 4978
rect 12360 4808 12388 4950
rect 12266 4780 12388 4808
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 12162 4720 12218 4729
rect 12266 4706 12294 4780
rect 12263 4690 12294 4706
rect 12346 4720 12402 4729
rect 12162 4655 12218 4664
rect 12256 4684 12308 4690
rect 12346 4655 12402 4664
rect 12256 4626 12308 4632
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 12176 3670 12204 4422
rect 12254 4312 12310 4321
rect 12254 4247 12310 4256
rect 12268 3738 12296 4247
rect 12360 4146 12388 4655
rect 12452 4554 12480 4791
rect 12544 4570 12572 5102
rect 12716 5092 12768 5098
rect 12636 5052 12716 5080
rect 12636 4690 12664 5052
rect 12806 5063 12862 5072
rect 12716 5034 12768 5040
rect 12714 4856 12770 4865
rect 12714 4791 12770 4800
rect 12624 4684 12676 4690
rect 12624 4626 12676 4632
rect 12728 4570 12756 4791
rect 13004 4758 13032 5510
rect 13096 5234 13124 5674
rect 13372 5534 13400 5868
rect 13740 5778 13768 6122
rect 13728 5772 13780 5778
rect 13728 5714 13780 5720
rect 13636 5636 13688 5642
rect 13636 5578 13688 5584
rect 13188 5506 13400 5534
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13188 5114 13216 5506
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13372 5234 13400 5306
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13360 5228 13412 5234
rect 13360 5170 13412 5176
rect 13096 5098 13216 5114
rect 13084 5092 13216 5098
rect 13136 5086 13216 5092
rect 13280 5080 13308 5170
rect 13280 5052 13400 5080
rect 13084 5034 13136 5040
rect 13372 5012 13400 5052
rect 13464 5030 13492 5510
rect 13542 5400 13598 5409
rect 13648 5370 13676 5578
rect 13728 5568 13780 5574
rect 13832 5556 13860 7806
rect 14004 7744 14056 7750
rect 14004 7686 14056 7692
rect 14016 7478 14044 7686
rect 14004 7472 14056 7478
rect 13910 7440 13966 7449
rect 14004 7414 14056 7420
rect 13910 7375 13966 7384
rect 13924 7274 13952 7375
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14004 7268 14056 7274
rect 14004 7210 14056 7216
rect 13910 7168 13966 7177
rect 13910 7103 13966 7112
rect 13924 6934 13952 7103
rect 13912 6928 13964 6934
rect 13912 6870 13964 6876
rect 14016 6798 14044 7210
rect 14108 6934 14136 10016
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9518 14228 9998
rect 14188 9512 14240 9518
rect 14186 9480 14188 9489
rect 14240 9480 14242 9489
rect 14292 9450 14320 10066
rect 14186 9415 14242 9424
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14292 9353 14320 9386
rect 14278 9344 14334 9353
rect 14278 9279 14334 9288
rect 14384 8974 14412 11086
rect 14476 10266 14504 11342
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14556 10192 14608 10198
rect 14462 10160 14518 10169
rect 14660 10169 14688 11727
rect 14556 10134 14608 10140
rect 14646 10160 14702 10169
rect 14462 10095 14518 10104
rect 14476 10062 14504 10095
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14568 9518 14596 10134
rect 14646 10095 14702 10104
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14476 9178 14504 9386
rect 14554 9208 14610 9217
rect 14464 9172 14516 9178
rect 14554 9143 14610 9152
rect 14464 9114 14516 9120
rect 14372 8968 14424 8974
rect 14200 8928 14372 8956
rect 14200 7478 14228 8928
rect 14372 8910 14424 8916
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14278 7984 14334 7993
rect 14278 7919 14334 7928
rect 14188 7472 14240 7478
rect 14188 7414 14240 7420
rect 14186 7032 14242 7041
rect 14186 6967 14242 6976
rect 14096 6928 14148 6934
rect 14096 6870 14148 6876
rect 14004 6792 14056 6798
rect 14200 6780 14228 6967
rect 14004 6734 14056 6740
rect 14108 6752 14228 6780
rect 14016 6662 14044 6734
rect 14004 6656 14056 6662
rect 14108 6633 14136 6752
rect 14004 6598 14056 6604
rect 14094 6624 14150 6633
rect 14016 6118 14044 6598
rect 14094 6559 14150 6568
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14004 6112 14056 6118
rect 13910 6080 13966 6089
rect 14004 6054 14056 6060
rect 13910 6015 13966 6024
rect 13924 5778 13952 6015
rect 14016 5953 14044 6054
rect 14200 5953 14228 6258
rect 14002 5944 14058 5953
rect 14002 5879 14058 5888
rect 14186 5944 14242 5953
rect 14186 5879 14242 5888
rect 14016 5846 14044 5879
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13912 5772 13964 5778
rect 13912 5714 13964 5720
rect 14292 5702 14320 7919
rect 14384 5710 14412 8434
rect 14568 7664 14596 9143
rect 14752 7886 14780 12543
rect 14844 11762 14872 14311
rect 15028 13326 15056 14350
rect 15106 14311 15162 14320
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15016 13320 15068 13326
rect 14936 13280 15016 13308
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14832 11280 14884 11286
rect 14832 11222 14884 11228
rect 14844 10792 14872 11222
rect 14936 11014 14964 13280
rect 15016 13262 15068 13268
rect 15106 13152 15162 13161
rect 15106 13087 15162 13096
rect 15016 12776 15068 12782
rect 15120 12764 15148 13087
rect 15068 12736 15148 12764
rect 15016 12718 15068 12724
rect 15106 11792 15162 11801
rect 15028 11750 15106 11778
rect 15028 11286 15056 11750
rect 15106 11727 15162 11736
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15016 11280 15068 11286
rect 15016 11222 15068 11228
rect 15120 11014 15148 11630
rect 14924 11008 14976 11014
rect 15108 11008 15160 11014
rect 14976 10956 15056 10962
rect 14924 10950 15056 10956
rect 15108 10950 15160 10956
rect 14936 10934 15056 10950
rect 14924 10804 14976 10810
rect 14844 10764 14924 10792
rect 14924 10746 14976 10752
rect 14832 10464 14884 10470
rect 14832 10406 14884 10412
rect 14844 9110 14872 10406
rect 15028 10112 15056 10934
rect 15120 10674 15148 10950
rect 15212 10674 15240 13874
rect 15304 13870 15332 15438
rect 15384 14408 15436 14414
rect 15384 14350 15436 14356
rect 15396 13870 15424 14350
rect 15488 14113 15516 16934
rect 15672 16046 15700 17926
rect 15784 17436 16092 17445
rect 15784 17434 15790 17436
rect 15846 17434 15870 17436
rect 15926 17434 15950 17436
rect 16006 17434 16030 17436
rect 16086 17434 16092 17436
rect 15846 17382 15848 17434
rect 16028 17382 16030 17434
rect 15784 17380 15790 17382
rect 15846 17380 15870 17382
rect 15926 17380 15950 17382
rect 16006 17380 16030 17382
rect 16086 17380 16092 17382
rect 15784 17371 16092 17380
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15764 16658 15792 17274
rect 16026 16688 16082 16697
rect 15752 16652 15804 16658
rect 16026 16623 16028 16632
rect 15752 16594 15804 16600
rect 16080 16623 16082 16632
rect 16028 16594 16080 16600
rect 15784 16348 16092 16357
rect 15784 16346 15790 16348
rect 15846 16346 15870 16348
rect 15926 16346 15950 16348
rect 16006 16346 16030 16348
rect 16086 16346 16092 16348
rect 15846 16294 15848 16346
rect 16028 16294 16030 16346
rect 15784 16292 15790 16294
rect 15846 16292 15870 16294
rect 15926 16292 15950 16294
rect 16006 16292 16030 16294
rect 16086 16292 16092 16294
rect 15784 16283 16092 16292
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15660 15564 15712 15570
rect 15660 15506 15712 15512
rect 15566 15464 15622 15473
rect 15566 15399 15622 15408
rect 15474 14104 15530 14113
rect 15474 14039 15530 14048
rect 15292 13864 15344 13870
rect 15292 13806 15344 13812
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15580 13802 15608 15399
rect 15672 15094 15700 15506
rect 15784 15260 16092 15269
rect 15784 15258 15790 15260
rect 15846 15258 15870 15260
rect 15926 15258 15950 15260
rect 16006 15258 16030 15260
rect 16086 15258 16092 15260
rect 15846 15206 15848 15258
rect 16028 15206 16030 15258
rect 15784 15204 15790 15206
rect 15846 15204 15870 15206
rect 15926 15204 15950 15206
rect 16006 15204 16030 15206
rect 16086 15204 16092 15206
rect 15784 15195 16092 15204
rect 16132 15162 16160 19178
rect 16224 18290 16252 19654
rect 16212 18284 16264 18290
rect 16212 18226 16264 18232
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16224 16794 16252 16934
rect 16212 16788 16264 16794
rect 16212 16730 16264 16736
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16224 15502 16252 15982
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 15660 15088 15712 15094
rect 15660 15030 15712 15036
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15936 14816 15988 14822
rect 15936 14758 15988 14764
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 15672 14074 15700 14758
rect 15948 14618 15976 14758
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15784 14172 16092 14181
rect 15784 14170 15790 14172
rect 15846 14170 15870 14172
rect 15926 14170 15950 14172
rect 16006 14170 16030 14172
rect 16086 14170 16092 14172
rect 15846 14118 15848 14170
rect 16028 14118 16030 14170
rect 15784 14116 15790 14118
rect 15846 14116 15870 14118
rect 15926 14116 15950 14118
rect 16006 14116 16030 14118
rect 16086 14116 16092 14118
rect 15784 14107 16092 14116
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15660 13932 15712 13938
rect 15660 13874 15712 13880
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15672 13682 15700 13874
rect 15752 13796 15804 13802
rect 15752 13738 15804 13744
rect 15488 13654 15700 13682
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 15304 12850 15332 13466
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15290 12472 15346 12481
rect 15290 12407 15346 12416
rect 15304 12306 15332 12407
rect 15292 12300 15344 12306
rect 15292 12242 15344 12248
rect 15290 12064 15346 12073
rect 15290 11999 15346 12008
rect 15304 11676 15332 11999
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15396 11801 15424 11834
rect 15382 11792 15438 11801
rect 15488 11762 15516 13654
rect 15764 13172 15792 13738
rect 15934 13288 15990 13297
rect 15934 13223 15936 13232
rect 15988 13223 15990 13232
rect 15936 13194 15988 13200
rect 15672 13144 15792 13172
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15580 11898 15608 12582
rect 15672 12481 15700 13144
rect 15784 13084 16092 13093
rect 15784 13082 15790 13084
rect 15846 13082 15870 13084
rect 15926 13082 15950 13084
rect 16006 13082 16030 13084
rect 16086 13082 16092 13084
rect 15846 13030 15848 13082
rect 16028 13030 16030 13082
rect 15784 13028 15790 13030
rect 15846 13028 15870 13030
rect 15926 13028 15950 13030
rect 16006 13028 16030 13030
rect 16086 13028 16092 13030
rect 15784 13019 16092 13028
rect 16132 12968 16160 14758
rect 16224 14657 16252 15438
rect 16210 14648 16266 14657
rect 16210 14583 16266 14592
rect 16316 14385 16344 20975
rect 16396 20936 16448 20942
rect 16396 20878 16448 20884
rect 16408 20602 16436 20878
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16580 20868 16632 20874
rect 16580 20810 16632 20816
rect 16500 20777 16528 20810
rect 16486 20768 16542 20777
rect 16486 20703 16542 20712
rect 16486 20632 16542 20641
rect 16396 20596 16448 20602
rect 16592 20602 16620 20810
rect 16486 20567 16542 20576
rect 16580 20596 16632 20602
rect 16396 20538 16448 20544
rect 16408 20058 16436 20538
rect 16396 20052 16448 20058
rect 16396 19994 16448 20000
rect 16396 19916 16448 19922
rect 16396 19858 16448 19864
rect 16408 18086 16436 19858
rect 16396 18080 16448 18086
rect 16396 18022 16448 18028
rect 16408 17678 16436 18022
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16302 14376 16358 14385
rect 16212 14340 16264 14346
rect 16302 14311 16358 14320
rect 16212 14282 16264 14288
rect 16224 13938 16252 14282
rect 16212 13932 16264 13938
rect 16212 13874 16264 13880
rect 16408 13818 16436 17614
rect 16500 16833 16528 20567
rect 16580 20538 16632 20544
rect 16684 20398 16712 21984
rect 16764 21966 16816 21972
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16672 20392 16724 20398
rect 16672 20334 16724 20340
rect 16580 20256 16632 20262
rect 16580 20198 16632 20204
rect 16592 18193 16620 20198
rect 16776 19922 16804 21626
rect 16868 20602 16896 22066
rect 17052 21146 17080 25366
rect 17144 25362 17172 26846
rect 17236 26948 17356 26976
rect 17236 25498 17264 26948
rect 17316 26784 17368 26790
rect 17314 26752 17316 26761
rect 17368 26752 17370 26761
rect 17314 26687 17370 26696
rect 17316 26580 17368 26586
rect 17316 26522 17368 26528
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 17132 25356 17184 25362
rect 17132 25298 17184 25304
rect 17132 25220 17184 25226
rect 17132 25162 17184 25168
rect 17144 23798 17172 25162
rect 17132 23792 17184 23798
rect 17132 23734 17184 23740
rect 17144 22545 17172 23734
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17130 22536 17186 22545
rect 17130 22471 17186 22480
rect 17130 21992 17186 22001
rect 17130 21927 17186 21936
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17144 20890 17172 21927
rect 17236 21690 17264 22646
rect 17224 21684 17276 21690
rect 17224 21626 17276 21632
rect 17052 20862 17172 20890
rect 16856 20596 16908 20602
rect 16856 20538 16908 20544
rect 16868 20058 16896 20538
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16764 19916 16816 19922
rect 16764 19858 16816 19864
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 16764 18624 16816 18630
rect 16764 18566 16816 18572
rect 16578 18184 16634 18193
rect 16578 18119 16634 18128
rect 16580 17876 16632 17882
rect 16580 17818 16632 17824
rect 16486 16824 16542 16833
rect 16486 16759 16542 16768
rect 16486 16552 16542 16561
rect 16592 16522 16620 17818
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16684 17134 16712 17546
rect 16672 17128 16724 17134
rect 16672 17070 16724 17076
rect 16486 16487 16542 16496
rect 16580 16516 16632 16522
rect 16500 15162 16528 16487
rect 16580 16458 16632 16464
rect 16684 16232 16712 17070
rect 16592 16204 16712 16232
rect 16592 15434 16620 16204
rect 16672 16108 16724 16114
rect 16672 16050 16724 16056
rect 16684 15745 16712 16050
rect 16670 15736 16726 15745
rect 16670 15671 16726 15680
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16580 15156 16632 15162
rect 16580 15098 16632 15104
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16500 13954 16528 14350
rect 16592 14346 16620 15098
rect 16580 14340 16632 14346
rect 16580 14282 16632 14288
rect 16500 13926 16620 13954
rect 16212 13796 16264 13802
rect 16212 13738 16264 13744
rect 16316 13790 16436 13818
rect 16224 13326 16252 13738
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 15948 12940 16160 12968
rect 15658 12472 15714 12481
rect 15658 12407 15714 12416
rect 15948 12170 15976 12940
rect 16224 12782 16252 13262
rect 16212 12776 16264 12782
rect 16118 12744 16174 12753
rect 16212 12718 16264 12724
rect 16118 12679 16120 12688
rect 16172 12679 16174 12688
rect 16120 12650 16172 12656
rect 16028 12232 16080 12238
rect 16080 12192 16160 12220
rect 16028 12174 16080 12180
rect 15936 12164 15988 12170
rect 15672 12124 15936 12152
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15672 11778 15700 12124
rect 15936 12106 15988 12112
rect 15784 11996 16092 12005
rect 15784 11994 15790 11996
rect 15846 11994 15870 11996
rect 15926 11994 15950 11996
rect 16006 11994 16030 11996
rect 16086 11994 16092 11996
rect 15846 11942 15848 11994
rect 16028 11942 16030 11994
rect 15784 11940 15790 11942
rect 15846 11940 15870 11942
rect 15926 11940 15950 11942
rect 16006 11940 16030 11942
rect 16086 11940 16092 11942
rect 15784 11931 16092 11940
rect 15382 11727 15438 11736
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15580 11750 15700 11778
rect 15304 11648 15424 11676
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15304 10849 15332 11290
rect 15290 10840 15346 10849
rect 15290 10775 15346 10784
rect 15396 10742 15424 11648
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15108 10668 15160 10674
rect 15108 10610 15160 10616
rect 15200 10668 15252 10674
rect 15200 10610 15252 10616
rect 15108 10124 15160 10130
rect 14936 10084 15108 10112
rect 14936 9586 14964 10084
rect 15108 10066 15160 10072
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14922 9208 14978 9217
rect 14922 9143 14978 9152
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14568 7636 14780 7664
rect 14646 7576 14702 7585
rect 14646 7511 14702 7520
rect 14556 7472 14608 7478
rect 14556 7414 14608 7420
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14476 6458 14504 7346
rect 14568 7002 14596 7414
rect 14660 7002 14688 7511
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14752 6458 14780 7636
rect 14830 7440 14886 7449
rect 14830 7375 14886 7384
rect 14844 6769 14872 7375
rect 14936 6798 14964 9143
rect 15212 8974 15240 10610
rect 15290 9616 15346 9625
rect 15488 9602 15516 11698
rect 15580 11082 15608 11750
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15346 9574 15516 9602
rect 15580 9976 15608 11018
rect 15672 10985 15700 11086
rect 16132 11082 16160 12192
rect 16120 11076 16172 11082
rect 16120 11018 16172 11024
rect 16224 11014 16252 12718
rect 16316 12617 16344 13790
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16408 12850 16436 13670
rect 16488 13252 16540 13258
rect 16488 13194 16540 13200
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16302 12608 16358 12617
rect 16302 12543 16358 12552
rect 16302 12472 16358 12481
rect 16358 12430 16436 12458
rect 16302 12407 16358 12416
rect 16302 12064 16358 12073
rect 16302 11999 16358 12008
rect 16316 11830 16344 11999
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16212 11008 16264 11014
rect 15658 10976 15714 10985
rect 16212 10950 16264 10956
rect 15658 10911 15714 10920
rect 15784 10908 16092 10917
rect 15784 10906 15790 10908
rect 15846 10906 15870 10908
rect 15926 10906 15950 10908
rect 16006 10906 16030 10908
rect 16086 10906 16092 10908
rect 15846 10854 15848 10906
rect 16028 10854 16030 10906
rect 15784 10852 15790 10854
rect 15846 10852 15870 10854
rect 15926 10852 15950 10854
rect 16006 10852 16030 10854
rect 16086 10852 16092 10854
rect 15784 10843 16092 10852
rect 16224 10849 16252 10950
rect 16210 10840 16266 10849
rect 16408 10810 16436 12430
rect 16210 10775 16266 10784
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16396 10804 16448 10810
rect 16396 10746 16448 10752
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 16316 10690 16344 10746
rect 16500 10690 16528 13194
rect 15844 10532 15896 10538
rect 15844 10474 15896 10480
rect 15856 10266 15884 10474
rect 15844 10260 15896 10266
rect 15844 10202 15896 10208
rect 15948 10062 15976 10678
rect 16120 10668 16172 10674
rect 16316 10662 16528 10690
rect 16592 10674 16620 13926
rect 16684 13546 16712 15671
rect 16776 13682 16804 18566
rect 16856 18420 16908 18426
rect 16856 18362 16908 18368
rect 16868 14482 16896 18362
rect 16960 18329 16988 18634
rect 16946 18320 17002 18329
rect 16946 18255 17002 18264
rect 16948 16176 17000 16182
rect 16946 16144 16948 16153
rect 17000 16144 17002 16153
rect 16946 16079 17002 16088
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16960 15473 16988 15846
rect 16946 15464 17002 15473
rect 16946 15399 17002 15408
rect 16948 15360 17000 15366
rect 16948 15302 17000 15308
rect 16856 14476 16908 14482
rect 16856 14418 16908 14424
rect 16960 13705 16988 15302
rect 16946 13696 17002 13705
rect 16776 13654 16896 13682
rect 16684 13518 16804 13546
rect 16672 13320 16724 13326
rect 16670 13288 16672 13297
rect 16724 13288 16726 13297
rect 16670 13223 16726 13232
rect 16670 12744 16726 12753
rect 16670 12679 16726 12688
rect 16684 11880 16712 12679
rect 16776 12170 16804 13518
rect 16868 12238 16896 13654
rect 16946 13631 17002 13640
rect 17052 13258 17080 20862
rect 17132 20800 17184 20806
rect 17132 20742 17184 20748
rect 17040 13252 17092 13258
rect 17040 13194 17092 13200
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16960 12617 16988 12786
rect 16946 12608 17002 12617
rect 16946 12543 17002 12552
rect 16856 12232 16908 12238
rect 16856 12174 16908 12180
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 16684 11852 16804 11880
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16580 10668 16632 10674
rect 16120 10610 16172 10616
rect 16580 10610 16632 10616
rect 16028 10600 16080 10606
rect 16028 10542 16080 10548
rect 16040 10062 16068 10542
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 15580 9948 15884 9976
rect 15290 9551 15346 9560
rect 15476 9376 15528 9382
rect 15304 9336 15476 9364
rect 15200 8968 15252 8974
rect 15200 8910 15252 8916
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15028 7721 15056 7890
rect 15014 7712 15070 7721
rect 15014 7647 15070 7656
rect 15120 7596 15148 8570
rect 15212 8498 15240 8910
rect 15304 8673 15332 9336
rect 15476 9318 15528 9324
rect 15580 9178 15608 9948
rect 15856 9908 15884 9948
rect 16040 9908 16068 9998
rect 16132 9926 16160 10610
rect 16302 10568 16358 10577
rect 16224 10526 16302 10554
rect 15658 9888 15714 9897
rect 15856 9880 16068 9908
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 15658 9823 15714 9832
rect 15672 9674 15700 9823
rect 15784 9820 16092 9829
rect 15784 9818 15790 9820
rect 15846 9818 15870 9820
rect 15926 9818 15950 9820
rect 16006 9818 16030 9820
rect 16086 9818 16092 9820
rect 15846 9766 15848 9818
rect 16028 9766 16030 9818
rect 15784 9764 15790 9766
rect 15846 9764 15870 9766
rect 15926 9764 15950 9766
rect 16006 9764 16030 9766
rect 16086 9764 16092 9766
rect 15784 9755 16092 9764
rect 16224 9704 16252 10526
rect 16302 10503 16358 10512
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 9897 16344 10406
rect 16396 9920 16448 9926
rect 16302 9888 16358 9897
rect 16396 9862 16448 9868
rect 16302 9823 16358 9832
rect 16304 9716 16356 9722
rect 16224 9676 16304 9704
rect 15672 9646 15792 9674
rect 16408 9674 16436 9862
rect 16304 9658 16356 9664
rect 15660 9580 15712 9586
rect 15660 9522 15712 9528
rect 15672 9489 15700 9522
rect 15658 9480 15714 9489
rect 15658 9415 15714 9424
rect 15764 9217 15792 9646
rect 16406 9646 16436 9674
rect 16684 9654 16712 11698
rect 16776 11150 16804 11852
rect 16868 11762 16896 12174
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16764 11144 16816 11150
rect 16816 11104 16896 11132
rect 16764 11086 16816 11092
rect 16764 10192 16816 10198
rect 16764 10134 16816 10140
rect 16672 9648 16724 9654
rect 16028 9580 16080 9586
rect 16028 9522 16080 9528
rect 16304 9580 16356 9586
rect 16406 9568 16434 9646
rect 16672 9590 16724 9596
rect 16356 9540 16434 9568
rect 16304 9522 16356 9528
rect 15750 9208 15806 9217
rect 15568 9172 15620 9178
rect 15750 9143 15806 9152
rect 15568 9114 15620 9120
rect 15384 9104 15436 9110
rect 15384 9046 15436 9052
rect 15290 8664 15346 8673
rect 15290 8599 15346 8608
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15028 7568 15148 7596
rect 14924 6792 14976 6798
rect 14830 6760 14886 6769
rect 14924 6734 14976 6740
rect 14830 6695 14886 6704
rect 15028 6644 15056 7568
rect 15396 7274 15424 9046
rect 15474 8936 15530 8945
rect 15936 8900 15988 8906
rect 15474 8871 15530 8880
rect 15488 8634 15516 8871
rect 15672 8860 15936 8888
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15488 8498 15516 8570
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15672 8294 15700 8860
rect 15936 8842 15988 8848
rect 16040 8838 16068 9522
rect 16684 9518 16712 9590
rect 16120 9512 16172 9518
rect 16672 9512 16724 9518
rect 16120 9454 16172 9460
rect 16500 9472 16672 9500
rect 16132 9160 16160 9454
rect 16212 9172 16264 9178
rect 16132 9132 16212 9160
rect 16212 9114 16264 9120
rect 16120 8968 16172 8974
rect 16396 8968 16448 8974
rect 16120 8910 16172 8916
rect 16394 8936 16396 8945
rect 16448 8936 16450 8945
rect 16028 8832 16080 8838
rect 16132 8820 16160 8910
rect 16394 8871 16450 8880
rect 16132 8792 16344 8820
rect 16028 8774 16080 8780
rect 15784 8732 16092 8741
rect 15784 8730 15790 8732
rect 15846 8730 15870 8732
rect 15926 8730 15950 8732
rect 16006 8730 16030 8732
rect 16086 8730 16092 8732
rect 15846 8678 15848 8730
rect 16028 8678 16030 8730
rect 15784 8676 15790 8678
rect 15846 8676 15870 8678
rect 15926 8676 15950 8678
rect 16006 8676 16030 8678
rect 16086 8676 16092 8678
rect 15784 8667 16092 8676
rect 16210 8664 16266 8673
rect 16210 8599 16212 8608
rect 16264 8599 16266 8608
rect 16212 8570 16264 8576
rect 15844 8560 15896 8566
rect 15764 8520 15844 8548
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15488 7342 15516 7822
rect 15764 7750 15792 8520
rect 15844 8502 15896 8508
rect 16120 8560 16172 8566
rect 16120 8502 16172 8508
rect 15844 8424 15896 8430
rect 15844 8366 15896 8372
rect 15856 8090 15884 8366
rect 16132 8090 16160 8502
rect 16316 8498 16344 8792
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16210 8120 16266 8129
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 16120 8084 16172 8090
rect 16210 8055 16266 8064
rect 16120 8026 16172 8032
rect 15936 7880 15988 7886
rect 15988 7840 16160 7868
rect 15936 7822 15988 7828
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15752 7744 15804 7750
rect 15752 7686 15804 7692
rect 15672 7460 15700 7686
rect 15784 7644 16092 7653
rect 15784 7642 15790 7644
rect 15846 7642 15870 7644
rect 15926 7642 15950 7644
rect 16006 7642 16030 7644
rect 16086 7642 16092 7644
rect 15846 7590 15848 7642
rect 16028 7590 16030 7642
rect 15784 7588 15790 7590
rect 15846 7588 15870 7590
rect 15926 7588 15950 7590
rect 16006 7588 16030 7590
rect 16086 7588 16092 7590
rect 15784 7579 16092 7588
rect 16132 7546 16160 7840
rect 16224 7721 16252 8055
rect 16394 7984 16450 7993
rect 16500 7954 16528 9472
rect 16672 9454 16724 9460
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8974 16620 9318
rect 16776 9024 16804 10134
rect 16684 8996 16804 9024
rect 16580 8968 16632 8974
rect 16580 8910 16632 8916
rect 16684 8634 16712 8996
rect 16672 8628 16724 8634
rect 16672 8570 16724 8576
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16670 8120 16726 8129
rect 16776 8090 16804 8434
rect 16670 8055 16672 8064
rect 16724 8055 16726 8064
rect 16764 8084 16816 8090
rect 16672 8026 16724 8032
rect 16764 8026 16816 8032
rect 16394 7919 16450 7928
rect 16488 7948 16540 7954
rect 16304 7744 16356 7750
rect 16210 7712 16266 7721
rect 16408 7721 16436 7919
rect 16488 7890 16540 7896
rect 16304 7686 16356 7692
rect 16394 7712 16450 7721
rect 16210 7647 16266 7656
rect 16120 7540 16172 7546
rect 16120 7482 16172 7488
rect 16212 7540 16264 7546
rect 16316 7528 16344 7686
rect 16394 7647 16450 7656
rect 16316 7500 16436 7528
rect 16212 7482 16264 7488
rect 15752 7472 15804 7478
rect 15672 7432 15752 7460
rect 15752 7414 15804 7420
rect 15476 7336 15528 7342
rect 15476 7278 15528 7284
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15752 7268 15804 7274
rect 15752 7210 15804 7216
rect 15304 6956 15608 6984
rect 15304 6769 15332 6956
rect 15384 6860 15436 6866
rect 15384 6802 15436 6808
rect 15290 6760 15346 6769
rect 15290 6695 15346 6704
rect 14936 6616 15056 6644
rect 15200 6656 15252 6662
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14016 5674 14320 5702
rect 14372 5704 14424 5710
rect 13912 5636 13964 5642
rect 13912 5578 13964 5584
rect 13780 5528 13860 5556
rect 13728 5510 13780 5516
rect 13924 5386 13952 5578
rect 13542 5335 13598 5344
rect 13636 5364 13688 5370
rect 13556 5098 13584 5335
rect 13636 5306 13688 5312
rect 13728 5364 13780 5370
rect 13728 5306 13780 5312
rect 13832 5358 13952 5386
rect 13740 5234 13768 5306
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13188 4984 13400 5012
rect 13452 5024 13504 5030
rect 13188 4865 13216 4984
rect 13452 4966 13504 4972
rect 13312 4924 13620 4933
rect 13312 4922 13318 4924
rect 13374 4922 13398 4924
rect 13454 4922 13478 4924
rect 13534 4922 13558 4924
rect 13614 4922 13620 4924
rect 13374 4870 13376 4922
rect 13556 4870 13558 4922
rect 13312 4868 13318 4870
rect 13374 4868 13398 4870
rect 13454 4868 13478 4870
rect 13534 4868 13558 4870
rect 13614 4868 13620 4870
rect 13174 4856 13230 4865
rect 13312 4859 13620 4868
rect 13084 4820 13136 4826
rect 13648 4808 13676 5170
rect 13728 5024 13780 5030
rect 13728 4966 13780 4972
rect 13174 4791 13230 4800
rect 13084 4762 13136 4768
rect 13372 4780 13676 4808
rect 12992 4752 13044 4758
rect 12992 4694 13044 4700
rect 12440 4548 12492 4554
rect 12544 4542 12756 4570
rect 12440 4490 12492 4496
rect 12992 4480 13044 4486
rect 12438 4448 12494 4457
rect 12898 4448 12954 4457
rect 12494 4406 12898 4434
rect 12438 4383 12494 4392
rect 12992 4422 13044 4428
rect 12898 4383 12954 4392
rect 13004 4298 13032 4422
rect 12452 4270 13032 4298
rect 12348 4140 12400 4146
rect 12348 4082 12400 4088
rect 12452 4049 12480 4270
rect 13096 4146 13124 4762
rect 13268 4752 13320 4758
rect 13174 4720 13230 4729
rect 13268 4694 13320 4700
rect 13174 4655 13176 4664
rect 13228 4655 13230 4664
rect 13176 4626 13228 4632
rect 13280 4536 13308 4694
rect 13372 4622 13400 4780
rect 13452 4684 13504 4690
rect 13452 4626 13504 4632
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13188 4508 13308 4536
rect 13188 4185 13216 4508
rect 13464 4434 13492 4626
rect 13544 4616 13596 4622
rect 13280 4406 13492 4434
rect 13522 4564 13544 4604
rect 13740 4570 13768 4966
rect 13832 4826 13860 5358
rect 14016 5080 14044 5674
rect 14372 5646 14424 5652
rect 14096 5636 14148 5642
rect 14096 5578 14148 5584
rect 13924 5052 14044 5080
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13522 4558 13596 4564
rect 13174 4176 13230 4185
rect 13084 4140 13136 4146
rect 13174 4111 13230 4120
rect 13084 4082 13136 4088
rect 12532 4072 12584 4078
rect 12438 4040 12494 4049
rect 12348 4004 12400 4010
rect 12992 4072 13044 4078
rect 12584 4032 12992 4060
rect 12532 4014 12584 4020
rect 13280 4049 13308 4406
rect 13522 4298 13550 4558
rect 13360 4276 13412 4282
rect 13360 4218 13412 4224
rect 13464 4270 13550 4298
rect 13648 4542 13768 4570
rect 13372 4185 13400 4218
rect 13358 4176 13414 4185
rect 13358 4111 13414 4120
rect 13360 4072 13412 4078
rect 12992 4014 13044 4020
rect 13266 4040 13322 4049
rect 12438 3975 12494 3984
rect 13176 4004 13228 4010
rect 12348 3946 12400 3952
rect 13464 4049 13492 4270
rect 13544 4208 13596 4214
rect 13648 4196 13676 4542
rect 13924 4434 13952 5052
rect 14108 4978 14136 5578
rect 14476 5386 14504 6054
rect 14554 5944 14610 5953
rect 14554 5879 14610 5888
rect 14200 5370 14504 5386
rect 14188 5364 14504 5370
rect 14240 5358 14504 5364
rect 14188 5306 14240 5312
rect 14280 5296 14332 5302
rect 14186 5264 14242 5273
rect 14280 5238 14332 5244
rect 14186 5199 14242 5208
rect 14200 5001 14228 5199
rect 14016 4950 14136 4978
rect 14186 4992 14242 5001
rect 14016 4554 14044 4950
rect 14186 4927 14242 4936
rect 14292 4842 14320 5238
rect 14568 5137 14596 5879
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14554 5128 14610 5137
rect 14554 5063 14610 5072
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14554 4992 14610 5001
rect 14384 4865 14412 4966
rect 14096 4820 14148 4826
rect 14096 4762 14148 4768
rect 14200 4814 14320 4842
rect 14370 4856 14426 4865
rect 14108 4729 14136 4762
rect 14094 4720 14150 4729
rect 14094 4655 14150 4664
rect 14200 4604 14228 4814
rect 14370 4791 14426 4800
rect 14476 4740 14504 4966
rect 14554 4927 14610 4936
rect 14568 4758 14596 4927
rect 14292 4712 14504 4740
rect 14556 4752 14608 4758
rect 14292 4622 14320 4712
rect 14556 4694 14608 4700
rect 14660 4690 14688 5510
rect 14752 5370 14780 6258
rect 14830 5808 14886 5817
rect 14830 5743 14886 5752
rect 14844 5642 14872 5743
rect 14936 5702 14964 6616
rect 15200 6598 15252 6604
rect 15108 6384 15160 6390
rect 15108 6326 15160 6332
rect 15014 6216 15070 6225
rect 15014 6151 15070 6160
rect 15028 5817 15056 6151
rect 15014 5808 15070 5817
rect 15014 5743 15070 5752
rect 14936 5674 15056 5702
rect 14832 5636 14884 5642
rect 14832 5578 14884 5584
rect 14740 5364 14792 5370
rect 14740 5306 14792 5312
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14936 5234 14964 5306
rect 15028 5302 15056 5674
rect 15120 5370 15148 6326
rect 15212 6322 15240 6598
rect 15290 6488 15346 6497
rect 15290 6423 15346 6432
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15304 6089 15332 6423
rect 15396 6118 15424 6802
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15580 6746 15608 6956
rect 15660 6860 15712 6866
rect 15764 6848 15792 7210
rect 16224 7206 16252 7482
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16212 7200 16264 7206
rect 16212 7142 16264 7148
rect 15712 6820 15792 6848
rect 15660 6802 15712 6808
rect 15488 6474 15516 6734
rect 15580 6718 16252 6746
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15566 6488 15622 6497
rect 15488 6446 15566 6474
rect 15384 6112 15436 6118
rect 15290 6080 15346 6089
rect 15384 6054 15436 6060
rect 15290 6015 15346 6024
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15016 5296 15068 5302
rect 15212 5250 15240 5510
rect 15016 5238 15068 5244
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 15120 5222 15240 5250
rect 14738 5128 14794 5137
rect 15120 5098 15148 5222
rect 15200 5160 15252 5166
rect 15198 5128 15200 5137
rect 15252 5128 15254 5137
rect 14738 5063 14794 5072
rect 15108 5092 15160 5098
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14752 4622 14780 5063
rect 15198 5063 15254 5072
rect 15108 5034 15160 5040
rect 15304 4826 15332 6015
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 15396 5710 15424 5850
rect 15488 5778 15516 6446
rect 15566 6423 15622 6432
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5846 15608 6054
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15672 5624 15700 6598
rect 15784 6556 16092 6565
rect 15784 6554 15790 6556
rect 15846 6554 15870 6556
rect 15926 6554 15950 6556
rect 16006 6554 16030 6556
rect 16086 6554 16092 6556
rect 15846 6502 15848 6554
rect 16028 6502 16030 6554
rect 15784 6500 15790 6502
rect 15846 6500 15870 6502
rect 15926 6500 15950 6502
rect 16006 6500 16030 6502
rect 16086 6500 16092 6502
rect 15784 6491 16092 6500
rect 16224 6497 16252 6718
rect 16210 6488 16266 6497
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15844 6452 15896 6458
rect 16028 6452 16080 6458
rect 15896 6412 16028 6440
rect 15844 6394 15896 6400
rect 16316 6458 16344 7346
rect 16408 7206 16436 7500
rect 16500 7342 16528 7890
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16684 7342 16712 7686
rect 16868 7528 16896 11104
rect 16960 9194 16988 12106
rect 17144 11354 17172 20742
rect 17222 20360 17278 20369
rect 17222 20295 17278 20304
rect 17236 19378 17264 20295
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17328 18222 17356 26522
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17420 15688 17448 28999
rect 17512 20806 17540 41074
rect 17604 41002 17632 41550
rect 17788 41120 17816 42502
rect 17868 42152 17920 42158
rect 17868 42094 17920 42100
rect 17696 41092 17816 41120
rect 17592 40996 17644 41002
rect 17592 40938 17644 40944
rect 17696 40186 17724 41092
rect 17776 40996 17828 41002
rect 17776 40938 17828 40944
rect 17788 40526 17816 40938
rect 17880 40934 17908 42094
rect 17958 41848 18014 41857
rect 17958 41783 18014 41792
rect 17972 41478 18000 41783
rect 18156 41698 18184 43250
rect 18248 43194 18276 44540
rect 18432 44010 18460 44540
rect 18432 43982 18552 44010
rect 18524 43926 18552 43982
rect 18512 43920 18564 43926
rect 18512 43862 18564 43868
rect 18616 43314 18644 44540
rect 18694 43344 18750 43353
rect 18604 43308 18656 43314
rect 18694 43279 18696 43288
rect 18604 43250 18656 43256
rect 18748 43279 18750 43288
rect 18696 43250 18748 43256
rect 18248 43166 18736 43194
rect 18604 43104 18656 43110
rect 18604 43046 18656 43052
rect 18257 43004 18565 43013
rect 18257 43002 18263 43004
rect 18319 43002 18343 43004
rect 18399 43002 18423 43004
rect 18479 43002 18503 43004
rect 18559 43002 18565 43004
rect 18319 42950 18321 43002
rect 18501 42950 18503 43002
rect 18257 42948 18263 42950
rect 18319 42948 18343 42950
rect 18399 42948 18423 42950
rect 18479 42948 18503 42950
rect 18559 42948 18565 42950
rect 18257 42939 18565 42948
rect 18326 42664 18382 42673
rect 18326 42599 18382 42608
rect 18340 42566 18368 42599
rect 18328 42560 18380 42566
rect 18328 42502 18380 42508
rect 18616 42294 18644 43046
rect 18708 42566 18736 43166
rect 18696 42560 18748 42566
rect 18696 42502 18748 42508
rect 18236 42288 18288 42294
rect 18236 42230 18288 42236
rect 18604 42288 18656 42294
rect 18604 42230 18656 42236
rect 18248 42129 18276 42230
rect 18234 42120 18290 42129
rect 18234 42055 18290 42064
rect 18257 41916 18565 41925
rect 18257 41914 18263 41916
rect 18319 41914 18343 41916
rect 18399 41914 18423 41916
rect 18479 41914 18503 41916
rect 18559 41914 18565 41916
rect 18319 41862 18321 41914
rect 18501 41862 18503 41914
rect 18257 41860 18263 41862
rect 18319 41860 18343 41862
rect 18399 41860 18423 41862
rect 18479 41860 18503 41862
rect 18559 41860 18565 41862
rect 18257 41851 18565 41860
rect 18800 41818 18828 44540
rect 18878 43208 18934 43217
rect 18878 43143 18934 43152
rect 18892 42634 18920 43143
rect 18880 42628 18932 42634
rect 18880 42570 18932 42576
rect 18984 42362 19012 44540
rect 19064 43716 19116 43722
rect 19064 43658 19116 43664
rect 19076 43314 19104 43658
rect 19064 43308 19116 43314
rect 19064 43250 19116 43256
rect 19062 42800 19118 42809
rect 19062 42735 19064 42744
rect 19116 42735 19118 42744
rect 19064 42706 19116 42712
rect 18972 42356 19024 42362
rect 18972 42298 19024 42304
rect 19168 42158 19196 44540
rect 19248 43920 19300 43926
rect 19248 43862 19300 43868
rect 19156 42152 19208 42158
rect 19156 42094 19208 42100
rect 18788 41812 18840 41818
rect 18788 41754 18840 41760
rect 18064 41670 18184 41698
rect 18236 41744 18288 41750
rect 18236 41686 18288 41692
rect 18064 41614 18092 41670
rect 18052 41608 18104 41614
rect 18052 41550 18104 41556
rect 18144 41540 18196 41546
rect 18144 41482 18196 41488
rect 17960 41472 18012 41478
rect 17960 41414 18012 41420
rect 18156 41414 18184 41482
rect 18064 41386 18184 41414
rect 18064 41018 18092 41386
rect 18248 41274 18276 41686
rect 18788 41540 18840 41546
rect 18788 41482 18840 41488
rect 18236 41268 18288 41274
rect 18236 41210 18288 41216
rect 18694 41168 18750 41177
rect 18236 41132 18288 41138
rect 18288 41092 18644 41120
rect 18694 41103 18750 41112
rect 18236 41074 18288 41080
rect 17972 40990 18092 41018
rect 17868 40928 17920 40934
rect 17868 40870 17920 40876
rect 17776 40520 17828 40526
rect 17776 40462 17828 40468
rect 17776 40384 17828 40390
rect 17776 40326 17828 40332
rect 17684 40180 17736 40186
rect 17684 40122 17736 40128
rect 17592 40044 17644 40050
rect 17592 39986 17644 39992
rect 17604 39642 17632 39986
rect 17682 39808 17738 39817
rect 17682 39743 17738 39752
rect 17696 39642 17724 39743
rect 17592 39636 17644 39642
rect 17592 39578 17644 39584
rect 17684 39636 17736 39642
rect 17684 39578 17736 39584
rect 17592 39500 17644 39506
rect 17592 39442 17644 39448
rect 17604 37482 17632 39442
rect 17788 39030 17816 40326
rect 17868 40044 17920 40050
rect 17868 39986 17920 39992
rect 17880 39642 17908 39986
rect 17972 39642 18000 40990
rect 18052 40928 18104 40934
rect 18052 40870 18104 40876
rect 18064 40118 18092 40870
rect 18257 40828 18565 40837
rect 18257 40826 18263 40828
rect 18319 40826 18343 40828
rect 18399 40826 18423 40828
rect 18479 40826 18503 40828
rect 18559 40826 18565 40828
rect 18319 40774 18321 40826
rect 18501 40774 18503 40826
rect 18257 40772 18263 40774
rect 18319 40772 18343 40774
rect 18399 40772 18423 40774
rect 18479 40772 18503 40774
rect 18559 40772 18565 40774
rect 18257 40763 18565 40772
rect 18326 40624 18382 40633
rect 18326 40559 18382 40568
rect 18144 40520 18196 40526
rect 18144 40462 18196 40468
rect 18234 40488 18290 40497
rect 18052 40112 18104 40118
rect 18156 40089 18184 40462
rect 18234 40423 18290 40432
rect 18248 40118 18276 40423
rect 18236 40112 18288 40118
rect 18052 40054 18104 40060
rect 18142 40080 18198 40089
rect 18236 40054 18288 40060
rect 18340 40050 18368 40559
rect 18420 40384 18472 40390
rect 18420 40326 18472 40332
rect 18432 40225 18460 40326
rect 18418 40216 18474 40225
rect 18418 40151 18474 40160
rect 18616 40089 18644 41092
rect 18602 40080 18658 40089
rect 18142 40015 18198 40024
rect 18328 40044 18380 40050
rect 18602 40015 18658 40024
rect 18328 39986 18380 39992
rect 18052 39908 18104 39914
rect 18052 39850 18104 39856
rect 17868 39636 17920 39642
rect 17868 39578 17920 39584
rect 17960 39636 18012 39642
rect 17960 39578 18012 39584
rect 18064 39370 18092 39850
rect 18708 39846 18736 41103
rect 18144 39840 18196 39846
rect 18144 39782 18196 39788
rect 18696 39840 18748 39846
rect 18696 39782 18748 39788
rect 18156 39624 18184 39782
rect 18257 39740 18565 39749
rect 18257 39738 18263 39740
rect 18319 39738 18343 39740
rect 18399 39738 18423 39740
rect 18479 39738 18503 39740
rect 18559 39738 18565 39740
rect 18319 39686 18321 39738
rect 18501 39686 18503 39738
rect 18257 39684 18263 39686
rect 18319 39684 18343 39686
rect 18399 39684 18423 39686
rect 18479 39684 18503 39686
rect 18559 39684 18565 39686
rect 18257 39675 18565 39684
rect 18694 39672 18750 39681
rect 18156 39596 18460 39624
rect 18236 39432 18288 39438
rect 18236 39374 18288 39380
rect 18326 39400 18382 39409
rect 18052 39364 18104 39370
rect 18052 39306 18104 39312
rect 18144 39364 18196 39370
rect 18144 39306 18196 39312
rect 17958 39264 18014 39273
rect 18156 39250 18184 39306
rect 18014 39222 18184 39250
rect 17958 39199 18014 39208
rect 18248 39098 18276 39374
rect 18326 39335 18328 39344
rect 18380 39335 18382 39344
rect 18328 39306 18380 39312
rect 18326 39128 18382 39137
rect 18236 39092 18288 39098
rect 18326 39063 18328 39072
rect 18236 39034 18288 39040
rect 18380 39063 18382 39072
rect 18328 39034 18380 39040
rect 17776 39024 17828 39030
rect 17776 38966 17828 38972
rect 18050 38992 18106 39001
rect 18432 38962 18460 39596
rect 18616 39616 18694 39624
rect 18616 39607 18750 39616
rect 18616 39596 18736 39607
rect 18512 39568 18564 39574
rect 18616 39556 18644 39596
rect 18564 39528 18644 39556
rect 18512 39510 18564 39516
rect 18800 39302 18828 41482
rect 19064 41472 19116 41478
rect 19064 41414 19116 41420
rect 19076 41138 19104 41414
rect 19260 41274 19288 43862
rect 19352 42106 19380 44540
rect 19982 44024 20038 44033
rect 19432 43988 19484 43994
rect 19982 43959 20038 43968
rect 19432 43930 19484 43936
rect 19444 43450 19472 43930
rect 19708 43852 19760 43858
rect 19708 43794 19760 43800
rect 19432 43444 19484 43450
rect 19432 43386 19484 43392
rect 19524 42832 19576 42838
rect 19524 42774 19576 42780
rect 19352 42078 19472 42106
rect 19340 42016 19392 42022
rect 19338 41984 19340 41993
rect 19392 41984 19394 41993
rect 19338 41919 19394 41928
rect 19444 41818 19472 42078
rect 19432 41812 19484 41818
rect 19432 41754 19484 41760
rect 19432 41540 19484 41546
rect 19432 41482 19484 41488
rect 19340 41472 19392 41478
rect 19340 41414 19392 41420
rect 19248 41268 19300 41274
rect 19248 41210 19300 41216
rect 18972 41132 19024 41138
rect 18972 41074 19024 41080
rect 19064 41132 19116 41138
rect 19064 41074 19116 41080
rect 18878 41032 18934 41041
rect 18878 40967 18934 40976
rect 18892 40050 18920 40967
rect 18880 40044 18932 40050
rect 18880 39986 18932 39992
rect 18880 39840 18932 39846
rect 18880 39782 18932 39788
rect 18788 39296 18840 39302
rect 18602 39264 18658 39273
rect 18788 39238 18840 39244
rect 18602 39199 18658 39208
rect 18050 38927 18052 38936
rect 18104 38927 18106 38936
rect 18328 38956 18380 38962
rect 18052 38898 18104 38904
rect 18328 38898 18380 38904
rect 18420 38956 18472 38962
rect 18420 38898 18472 38904
rect 18144 38820 18196 38826
rect 18340 38808 18368 38898
rect 18420 38820 18472 38826
rect 18340 38780 18420 38808
rect 18144 38762 18196 38768
rect 18420 38762 18472 38768
rect 18156 38350 18184 38762
rect 18257 38652 18565 38661
rect 18257 38650 18263 38652
rect 18319 38650 18343 38652
rect 18399 38650 18423 38652
rect 18479 38650 18503 38652
rect 18559 38650 18565 38652
rect 18319 38598 18321 38650
rect 18501 38598 18503 38650
rect 18257 38596 18263 38598
rect 18319 38596 18343 38598
rect 18399 38596 18423 38598
rect 18479 38596 18503 38598
rect 18559 38596 18565 38598
rect 18257 38587 18565 38596
rect 18328 38548 18380 38554
rect 18328 38490 18380 38496
rect 18340 38350 18368 38490
rect 17684 38344 17736 38350
rect 17684 38286 17736 38292
rect 18144 38344 18196 38350
rect 18144 38286 18196 38292
rect 18328 38344 18380 38350
rect 18328 38286 18380 38292
rect 17696 38010 17724 38286
rect 17776 38276 17828 38282
rect 17776 38218 17828 38224
rect 17684 38004 17736 38010
rect 17684 37946 17736 37952
rect 17788 37670 17816 38218
rect 18144 38208 18196 38214
rect 18064 38168 18144 38196
rect 17868 37868 17920 37874
rect 17868 37810 17920 37816
rect 17776 37664 17828 37670
rect 17776 37606 17828 37612
rect 17604 37454 17816 37482
rect 17592 37392 17644 37398
rect 17592 37334 17644 37340
rect 17604 35714 17632 37334
rect 17684 36032 17736 36038
rect 17684 35974 17736 35980
rect 17696 35834 17724 35974
rect 17684 35828 17736 35834
rect 17684 35770 17736 35776
rect 17604 35686 17724 35714
rect 17592 34400 17644 34406
rect 17592 34342 17644 34348
rect 17604 34202 17632 34342
rect 17592 34196 17644 34202
rect 17592 34138 17644 34144
rect 17592 33856 17644 33862
rect 17592 33798 17644 33804
rect 17604 31754 17632 33798
rect 17592 31748 17644 31754
rect 17592 31690 17644 31696
rect 17592 31340 17644 31346
rect 17592 31282 17644 31288
rect 17604 30682 17632 31282
rect 17696 30802 17724 35686
rect 17788 31838 17816 37454
rect 17880 35680 17908 37810
rect 17960 35692 18012 35698
rect 17880 35652 17960 35680
rect 17960 35634 18012 35640
rect 18064 35018 18092 38168
rect 18144 38150 18196 38156
rect 18144 37936 18196 37942
rect 18144 37878 18196 37884
rect 18156 37346 18184 37878
rect 18257 37564 18565 37573
rect 18257 37562 18263 37564
rect 18319 37562 18343 37564
rect 18399 37562 18423 37564
rect 18479 37562 18503 37564
rect 18559 37562 18565 37564
rect 18319 37510 18321 37562
rect 18501 37510 18503 37562
rect 18257 37508 18263 37510
rect 18319 37508 18343 37510
rect 18399 37508 18423 37510
rect 18479 37508 18503 37510
rect 18559 37508 18565 37510
rect 18257 37499 18565 37508
rect 18156 37318 18276 37346
rect 18144 36780 18196 36786
rect 18144 36722 18196 36728
rect 18156 36689 18184 36722
rect 18142 36680 18198 36689
rect 18248 36666 18276 37318
rect 18418 36952 18474 36961
rect 18418 36887 18474 36896
rect 18432 36786 18460 36887
rect 18420 36780 18472 36786
rect 18420 36722 18472 36728
rect 18326 36680 18382 36689
rect 18248 36638 18326 36666
rect 18142 36615 18198 36624
rect 18326 36615 18382 36624
rect 18257 36476 18565 36485
rect 18257 36474 18263 36476
rect 18319 36474 18343 36476
rect 18399 36474 18423 36476
rect 18479 36474 18503 36476
rect 18559 36474 18565 36476
rect 18319 36422 18321 36474
rect 18501 36422 18503 36474
rect 18257 36420 18263 36422
rect 18319 36420 18343 36422
rect 18399 36420 18423 36422
rect 18479 36420 18503 36422
rect 18559 36420 18565 36422
rect 18257 36411 18565 36420
rect 18616 36394 18644 39199
rect 18892 39001 18920 39782
rect 18984 39488 19012 41074
rect 19156 41064 19208 41070
rect 19156 41006 19208 41012
rect 19064 40520 19116 40526
rect 19064 40462 19116 40468
rect 19076 40186 19104 40462
rect 19064 40180 19116 40186
rect 19064 40122 19116 40128
rect 19064 39840 19116 39846
rect 19064 39782 19116 39788
rect 19076 39681 19104 39782
rect 19062 39672 19118 39681
rect 19062 39607 19118 39616
rect 18984 39460 19104 39488
rect 18972 39296 19024 39302
rect 18972 39238 19024 39244
rect 18984 39098 19012 39238
rect 18972 39092 19024 39098
rect 18972 39034 19024 39040
rect 18878 38992 18934 39001
rect 18878 38927 18934 38936
rect 19076 38654 19104 39460
rect 18892 38626 19104 38654
rect 18696 37256 18748 37262
rect 18788 37256 18840 37262
rect 18696 37198 18748 37204
rect 18786 37224 18788 37233
rect 18840 37224 18842 37233
rect 18708 36922 18736 37198
rect 18786 37159 18842 37168
rect 18696 36916 18748 36922
rect 18696 36858 18748 36864
rect 18694 36408 18750 36417
rect 18512 36372 18564 36378
rect 18616 36366 18694 36394
rect 18694 36343 18750 36352
rect 18512 36314 18564 36320
rect 18328 36304 18380 36310
rect 18328 36246 18380 36252
rect 18340 35834 18368 36246
rect 18420 36168 18472 36174
rect 18418 36136 18420 36145
rect 18472 36136 18474 36145
rect 18418 36071 18474 36080
rect 18524 35834 18552 36314
rect 18892 36224 18920 38626
rect 18972 38208 19024 38214
rect 18972 38150 19024 38156
rect 18984 38049 19012 38150
rect 18970 38040 19026 38049
rect 18970 37975 19026 37984
rect 18972 37868 19024 37874
rect 19168 37856 19196 41006
rect 19352 40168 19380 41414
rect 19444 40730 19472 41482
rect 19536 40730 19564 42774
rect 19616 42220 19668 42226
rect 19616 42162 19668 42168
rect 19432 40724 19484 40730
rect 19432 40666 19484 40672
rect 19524 40724 19576 40730
rect 19524 40666 19576 40672
rect 19432 40520 19484 40526
rect 19432 40462 19484 40468
rect 19260 40140 19380 40168
rect 19260 40050 19288 40140
rect 19248 40044 19300 40050
rect 19248 39986 19300 39992
rect 19340 40044 19392 40050
rect 19340 39986 19392 39992
rect 19352 39642 19380 39986
rect 19444 39642 19472 40462
rect 19524 39840 19576 39846
rect 19524 39782 19576 39788
rect 19340 39636 19392 39642
rect 19340 39578 19392 39584
rect 19432 39636 19484 39642
rect 19432 39578 19484 39584
rect 19248 39432 19300 39438
rect 19246 39400 19248 39409
rect 19432 39432 19484 39438
rect 19300 39400 19302 39409
rect 19432 39374 19484 39380
rect 19246 39335 19302 39344
rect 19248 39092 19300 39098
rect 19248 39034 19300 39040
rect 19260 38554 19288 39034
rect 19340 38956 19392 38962
rect 19340 38898 19392 38904
rect 19248 38548 19300 38554
rect 19248 38490 19300 38496
rect 19352 37942 19380 38898
rect 19444 38486 19472 39374
rect 19536 38826 19564 39782
rect 19628 39098 19656 42162
rect 19720 41177 19748 43794
rect 19800 43648 19852 43654
rect 19800 43590 19852 43596
rect 19812 43450 19840 43590
rect 19800 43444 19852 43450
rect 19800 43386 19852 43392
rect 19996 43314 20024 43959
rect 21178 43616 21234 43625
rect 20729 43548 21037 43557
rect 21178 43551 21234 43560
rect 20729 43546 20735 43548
rect 20791 43546 20815 43548
rect 20871 43546 20895 43548
rect 20951 43546 20975 43548
rect 21031 43546 21037 43548
rect 20791 43494 20793 43546
rect 20973 43494 20975 43546
rect 20729 43492 20735 43494
rect 20791 43492 20815 43494
rect 20871 43492 20895 43494
rect 20951 43492 20975 43494
rect 21031 43492 21037 43494
rect 20729 43483 21037 43492
rect 19984 43308 20036 43314
rect 19984 43250 20036 43256
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 19982 43072 20038 43081
rect 19982 43007 20038 43016
rect 19996 42906 20024 43007
rect 19984 42900 20036 42906
rect 19984 42842 20036 42848
rect 19892 42628 19944 42634
rect 19892 42570 19944 42576
rect 19904 42106 19932 42570
rect 19812 42078 19932 42106
rect 19812 41562 19840 42078
rect 19892 42016 19944 42022
rect 19892 41958 19944 41964
rect 19904 41732 19932 41958
rect 19904 41704 20116 41732
rect 19812 41534 19932 41562
rect 19798 41440 19854 41449
rect 19798 41375 19854 41384
rect 19706 41168 19762 41177
rect 19706 41103 19762 41112
rect 19812 40594 19840 41375
rect 19800 40588 19852 40594
rect 19800 40530 19852 40536
rect 19904 40474 19932 41534
rect 19720 40446 19932 40474
rect 19984 40520 20036 40526
rect 19984 40462 20036 40468
rect 19720 39953 19748 40446
rect 19800 40384 19852 40390
rect 19800 40326 19852 40332
rect 19812 40186 19840 40326
rect 19800 40180 19852 40186
rect 19800 40122 19852 40128
rect 19892 40044 19944 40050
rect 19892 39986 19944 39992
rect 19706 39944 19762 39953
rect 19706 39879 19762 39888
rect 19800 39840 19852 39846
rect 19800 39782 19852 39788
rect 19706 39536 19762 39545
rect 19706 39471 19762 39480
rect 19720 39438 19748 39471
rect 19708 39432 19760 39438
rect 19708 39374 19760 39380
rect 19616 39092 19668 39098
rect 19616 39034 19668 39040
rect 19524 38820 19576 38826
rect 19524 38762 19576 38768
rect 19708 38752 19760 38758
rect 19708 38694 19760 38700
rect 19432 38480 19484 38486
rect 19432 38422 19484 38428
rect 19432 38344 19484 38350
rect 19432 38286 19484 38292
rect 19524 38344 19576 38350
rect 19524 38286 19576 38292
rect 19340 37936 19392 37942
rect 19340 37878 19392 37884
rect 18972 37810 19024 37816
rect 19076 37828 19196 37856
rect 19248 37868 19300 37874
rect 18984 37466 19012 37810
rect 18972 37460 19024 37466
rect 18972 37402 19024 37408
rect 18972 37256 19024 37262
rect 18972 37198 19024 37204
rect 18984 36922 19012 37198
rect 18972 36916 19024 36922
rect 18972 36858 19024 36864
rect 18970 36816 19026 36825
rect 18970 36751 19026 36760
rect 18984 36310 19012 36751
rect 18972 36304 19024 36310
rect 18972 36246 19024 36252
rect 18800 36196 18920 36224
rect 18328 35828 18380 35834
rect 18328 35770 18380 35776
rect 18512 35828 18564 35834
rect 18512 35770 18564 35776
rect 18800 35737 18828 36196
rect 18972 36168 19024 36174
rect 18972 36110 19024 36116
rect 18880 36100 18932 36106
rect 18880 36042 18932 36048
rect 18786 35728 18842 35737
rect 18786 35663 18842 35672
rect 18696 35624 18748 35630
rect 18696 35566 18748 35572
rect 18144 35488 18196 35494
rect 18144 35430 18196 35436
rect 18156 35018 18184 35430
rect 18257 35388 18565 35397
rect 18257 35386 18263 35388
rect 18319 35386 18343 35388
rect 18399 35386 18423 35388
rect 18479 35386 18503 35388
rect 18559 35386 18565 35388
rect 18319 35334 18321 35386
rect 18501 35334 18503 35386
rect 18257 35332 18263 35334
rect 18319 35332 18343 35334
rect 18399 35332 18423 35334
rect 18479 35332 18503 35334
rect 18559 35332 18565 35334
rect 18257 35323 18565 35332
rect 18708 35086 18736 35566
rect 18892 35290 18920 36042
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18696 35080 18748 35086
rect 18696 35022 18748 35028
rect 18052 35012 18104 35018
rect 18052 34954 18104 34960
rect 18144 35012 18196 35018
rect 18144 34954 18196 34960
rect 18064 34678 18092 34954
rect 18984 34950 19012 36110
rect 18512 34944 18564 34950
rect 18512 34886 18564 34892
rect 18604 34944 18656 34950
rect 18604 34886 18656 34892
rect 18972 34944 19024 34950
rect 18972 34886 19024 34892
rect 18524 34678 18552 34886
rect 18052 34672 18104 34678
rect 18052 34614 18104 34620
rect 18512 34672 18564 34678
rect 18512 34614 18564 34620
rect 18257 34300 18565 34309
rect 18257 34298 18263 34300
rect 18319 34298 18343 34300
rect 18399 34298 18423 34300
rect 18479 34298 18503 34300
rect 18559 34298 18565 34300
rect 18319 34246 18321 34298
rect 18501 34246 18503 34298
rect 18257 34244 18263 34246
rect 18319 34244 18343 34246
rect 18399 34244 18423 34246
rect 18479 34244 18503 34246
rect 18559 34244 18565 34246
rect 18257 34235 18565 34244
rect 18512 34196 18564 34202
rect 18616 34184 18644 34886
rect 18970 34504 19026 34513
rect 18970 34439 19026 34448
rect 18696 34400 18748 34406
rect 18696 34342 18748 34348
rect 18564 34156 18644 34184
rect 18512 34138 18564 34144
rect 18604 34060 18656 34066
rect 18604 34002 18656 34008
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 18510 33960 18566 33969
rect 18248 33658 18276 33934
rect 18510 33895 18566 33904
rect 18524 33658 18552 33895
rect 18236 33652 18288 33658
rect 18236 33594 18288 33600
rect 18512 33652 18564 33658
rect 18512 33594 18564 33600
rect 18142 33552 18198 33561
rect 18142 33487 18198 33496
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 18064 32473 18092 33050
rect 18050 32464 18106 32473
rect 17960 32428 18012 32434
rect 18050 32399 18106 32408
rect 17960 32370 18012 32376
rect 17972 31958 18000 32370
rect 17960 31952 18012 31958
rect 17960 31894 18012 31900
rect 18156 31906 18184 33487
rect 18257 33212 18565 33221
rect 18257 33210 18263 33212
rect 18319 33210 18343 33212
rect 18399 33210 18423 33212
rect 18479 33210 18503 33212
rect 18559 33210 18565 33212
rect 18319 33158 18321 33210
rect 18501 33158 18503 33210
rect 18257 33156 18263 33158
rect 18319 33156 18343 33158
rect 18399 33156 18423 33158
rect 18479 33156 18503 33158
rect 18559 33156 18565 33158
rect 18257 33147 18565 33156
rect 18616 32910 18644 34002
rect 18708 33998 18736 34342
rect 18786 34096 18842 34105
rect 18786 34031 18842 34040
rect 18696 33992 18748 33998
rect 18696 33934 18748 33940
rect 18800 33980 18828 34031
rect 18880 33992 18932 33998
rect 18800 33952 18880 33980
rect 18694 33552 18750 33561
rect 18694 33487 18750 33496
rect 18708 33017 18736 33487
rect 18694 33008 18750 33017
rect 18694 32943 18750 32952
rect 18604 32904 18656 32910
rect 18604 32846 18656 32852
rect 18694 32872 18750 32881
rect 18800 32842 18828 33952
rect 18880 33934 18932 33940
rect 18984 33522 19012 34439
rect 19076 33561 19104 37828
rect 19248 37810 19300 37816
rect 19154 37768 19210 37777
rect 19154 37703 19210 37712
rect 19168 37466 19196 37703
rect 19156 37460 19208 37466
rect 19156 37402 19208 37408
rect 19156 36916 19208 36922
rect 19156 36858 19208 36864
rect 19168 35698 19196 36858
rect 19260 36854 19288 37810
rect 19340 37664 19392 37670
rect 19340 37606 19392 37612
rect 19352 37330 19380 37606
rect 19340 37324 19392 37330
rect 19340 37266 19392 37272
rect 19444 36922 19472 38286
rect 19536 38010 19564 38286
rect 19616 38208 19668 38214
rect 19616 38150 19668 38156
rect 19524 38004 19576 38010
rect 19524 37946 19576 37952
rect 19524 37868 19576 37874
rect 19524 37810 19576 37816
rect 19432 36916 19484 36922
rect 19432 36858 19484 36864
rect 19248 36848 19300 36854
rect 19248 36790 19300 36796
rect 19340 36100 19392 36106
rect 19340 36042 19392 36048
rect 19156 35692 19208 35698
rect 19156 35634 19208 35640
rect 19248 35556 19300 35562
rect 19248 35498 19300 35504
rect 19156 35488 19208 35494
rect 19156 35430 19208 35436
rect 19168 35086 19196 35430
rect 19260 35329 19288 35498
rect 19246 35320 19302 35329
rect 19246 35255 19302 35264
rect 19352 35204 19380 36042
rect 19536 36038 19564 37810
rect 19524 36032 19576 36038
rect 19524 35974 19576 35980
rect 19628 35834 19656 38150
rect 19720 37194 19748 38694
rect 19812 38554 19840 39782
rect 19904 39114 19932 39986
rect 19996 39302 20024 40462
rect 19984 39296 20036 39302
rect 19984 39238 20036 39244
rect 19904 39086 20024 39114
rect 19892 38956 19944 38962
rect 19892 38898 19944 38904
rect 19800 38548 19852 38554
rect 19800 38490 19852 38496
rect 19904 37806 19932 38898
rect 19996 38486 20024 39086
rect 20088 39030 20116 41704
rect 20180 41414 20208 43250
rect 20729 42460 21037 42469
rect 20729 42458 20735 42460
rect 20791 42458 20815 42460
rect 20871 42458 20895 42460
rect 20951 42458 20975 42460
rect 21031 42458 21037 42460
rect 20791 42406 20793 42458
rect 20973 42406 20975 42458
rect 20729 42404 20735 42406
rect 20791 42404 20815 42406
rect 20871 42404 20895 42406
rect 20951 42404 20975 42406
rect 21031 42404 21037 42406
rect 20729 42395 21037 42404
rect 21192 42362 21220 43551
rect 21272 43104 21324 43110
rect 21272 43046 21324 43052
rect 21284 42537 21312 43046
rect 21270 42528 21326 42537
rect 21270 42463 21326 42472
rect 21180 42356 21232 42362
rect 21180 42298 21232 42304
rect 20628 42220 20680 42226
rect 20628 42162 20680 42168
rect 20444 41608 20496 41614
rect 20444 41550 20496 41556
rect 20180 41386 20300 41414
rect 20168 40928 20220 40934
rect 20168 40870 20220 40876
rect 20180 39642 20208 40870
rect 20272 40186 20300 41386
rect 20352 40452 20404 40458
rect 20352 40394 20404 40400
rect 20260 40180 20312 40186
rect 20260 40122 20312 40128
rect 20260 40044 20312 40050
rect 20260 39986 20312 39992
rect 20168 39636 20220 39642
rect 20168 39578 20220 39584
rect 20076 39024 20128 39030
rect 20076 38966 20128 38972
rect 19984 38480 20036 38486
rect 19984 38422 20036 38428
rect 20076 38412 20128 38418
rect 20076 38354 20128 38360
rect 19984 38208 20036 38214
rect 19984 38150 20036 38156
rect 19892 37800 19944 37806
rect 19892 37742 19944 37748
rect 19800 37664 19852 37670
rect 19800 37606 19852 37612
rect 19892 37664 19944 37670
rect 19892 37606 19944 37612
rect 19812 37398 19840 37606
rect 19800 37392 19852 37398
rect 19800 37334 19852 37340
rect 19708 37188 19760 37194
rect 19708 37130 19760 37136
rect 19800 37188 19852 37194
rect 19800 37130 19852 37136
rect 19812 36553 19840 37130
rect 19904 36582 19932 37606
rect 19892 36576 19944 36582
rect 19798 36544 19854 36553
rect 19892 36518 19944 36524
rect 19798 36479 19854 36488
rect 19892 36168 19944 36174
rect 19892 36110 19944 36116
rect 19524 35828 19576 35834
rect 19524 35770 19576 35776
rect 19616 35828 19668 35834
rect 19616 35770 19668 35776
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 19444 35290 19472 35634
rect 19432 35284 19484 35290
rect 19432 35226 19484 35232
rect 19260 35176 19380 35204
rect 19156 35080 19208 35086
rect 19156 35022 19208 35028
rect 19156 34128 19208 34134
rect 19156 34070 19208 34076
rect 19168 33862 19196 34070
rect 19156 33856 19208 33862
rect 19156 33798 19208 33804
rect 19062 33552 19118 33561
rect 18972 33516 19024 33522
rect 18892 33476 18972 33504
rect 18694 32807 18750 32816
rect 18788 32836 18840 32842
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 18248 32337 18276 32370
rect 18234 32328 18290 32337
rect 18234 32263 18290 32272
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 18257 32124 18565 32133
rect 18257 32122 18263 32124
rect 18319 32122 18343 32124
rect 18399 32122 18423 32124
rect 18479 32122 18503 32124
rect 18559 32122 18565 32124
rect 18319 32070 18321 32122
rect 18501 32070 18503 32122
rect 18257 32068 18263 32070
rect 18319 32068 18343 32070
rect 18399 32068 18423 32070
rect 18479 32068 18503 32070
rect 18559 32068 18565 32070
rect 18257 32059 18565 32068
rect 18616 32026 18644 32166
rect 18604 32020 18656 32026
rect 18604 31962 18656 31968
rect 18156 31878 18276 31906
rect 17788 31810 18092 31838
rect 17868 31748 17920 31754
rect 17868 31690 17920 31696
rect 17684 30796 17736 30802
rect 17684 30738 17736 30744
rect 17776 30728 17828 30734
rect 17604 30654 17724 30682
rect 17776 30670 17828 30676
rect 17696 30598 17724 30654
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17684 30592 17736 30598
rect 17684 30534 17736 30540
rect 17604 30394 17632 30534
rect 17788 30394 17816 30670
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 17776 30388 17828 30394
rect 17776 30330 17828 30336
rect 17592 29776 17644 29782
rect 17592 29718 17644 29724
rect 17604 29306 17632 29718
rect 17592 29300 17644 29306
rect 17592 29242 17644 29248
rect 17776 29164 17828 29170
rect 17776 29106 17828 29112
rect 17590 29064 17646 29073
rect 17646 29022 17724 29050
rect 17590 28999 17646 29008
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17604 27470 17632 27814
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 17696 26874 17724 29022
rect 17788 28121 17816 29106
rect 17880 29034 17908 31690
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17868 29028 17920 29034
rect 17868 28970 17920 28976
rect 17972 28218 18000 30670
rect 18064 28506 18092 31810
rect 18248 31793 18276 31878
rect 18234 31784 18290 31793
rect 18708 31754 18736 32807
rect 18788 32778 18840 32784
rect 18234 31719 18290 31728
rect 18420 31748 18472 31754
rect 18420 31690 18472 31696
rect 18524 31726 18736 31754
rect 18788 31748 18840 31754
rect 18432 31385 18460 31690
rect 18418 31376 18474 31385
rect 18524 31346 18552 31726
rect 18788 31690 18840 31696
rect 18604 31680 18656 31686
rect 18656 31640 18736 31668
rect 18604 31622 18656 31628
rect 18708 31346 18736 31640
rect 18800 31482 18828 31690
rect 18788 31476 18840 31482
rect 18788 31418 18840 31424
rect 18418 31311 18474 31320
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18696 31340 18748 31346
rect 18696 31282 18748 31288
rect 18236 31272 18288 31278
rect 18142 31240 18198 31249
rect 18788 31272 18840 31278
rect 18288 31249 18368 31260
rect 18288 31240 18382 31249
rect 18288 31232 18326 31240
rect 18236 31214 18288 31220
rect 18142 31175 18198 31184
rect 18788 31214 18840 31220
rect 18326 31175 18382 31184
rect 18156 30734 18184 31175
rect 18420 31136 18472 31142
rect 18696 31136 18748 31142
rect 18472 31096 18644 31124
rect 18420 31078 18472 31084
rect 18257 31036 18565 31045
rect 18257 31034 18263 31036
rect 18319 31034 18343 31036
rect 18399 31034 18423 31036
rect 18479 31034 18503 31036
rect 18559 31034 18565 31036
rect 18319 30982 18321 31034
rect 18501 30982 18503 31034
rect 18257 30980 18263 30982
rect 18319 30980 18343 30982
rect 18399 30980 18423 30982
rect 18479 30980 18503 30982
rect 18559 30980 18565 30982
rect 18257 30971 18565 30980
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18236 30660 18288 30666
rect 18236 30602 18288 30608
rect 18144 30252 18196 30258
rect 18144 30194 18196 30200
rect 18156 29850 18184 30194
rect 18248 30161 18276 30602
rect 18234 30152 18290 30161
rect 18234 30087 18290 30096
rect 18257 29948 18565 29957
rect 18257 29946 18263 29948
rect 18319 29946 18343 29948
rect 18399 29946 18423 29948
rect 18479 29946 18503 29948
rect 18559 29946 18565 29948
rect 18319 29894 18321 29946
rect 18501 29894 18503 29946
rect 18257 29892 18263 29894
rect 18319 29892 18343 29894
rect 18399 29892 18423 29894
rect 18479 29892 18503 29894
rect 18559 29892 18565 29894
rect 18257 29883 18565 29892
rect 18144 29844 18196 29850
rect 18144 29786 18196 29792
rect 18616 29714 18644 31096
rect 18694 31104 18696 31113
rect 18748 31104 18750 31113
rect 18694 31039 18750 31048
rect 18800 30977 18828 31214
rect 18786 30968 18842 30977
rect 18786 30903 18842 30912
rect 18788 30728 18840 30734
rect 18788 30670 18840 30676
rect 18800 30394 18828 30670
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 18892 30274 18920 33476
rect 19062 33487 19118 33496
rect 18972 33458 19024 33464
rect 19260 32994 19288 35176
rect 19432 35148 19484 35154
rect 19352 35108 19432 35136
rect 19352 34746 19380 35108
rect 19432 35090 19484 35096
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 19536 34678 19564 35770
rect 19616 35692 19668 35698
rect 19616 35634 19668 35640
rect 19524 34672 19576 34678
rect 19524 34614 19576 34620
rect 19340 34604 19392 34610
rect 19340 34546 19392 34552
rect 19432 34604 19484 34610
rect 19432 34546 19484 34552
rect 19352 34202 19380 34546
rect 19340 34196 19392 34202
rect 19340 34138 19392 34144
rect 19444 34105 19472 34546
rect 19628 34202 19656 35634
rect 19904 35562 19932 36110
rect 19996 35766 20024 38150
rect 20088 36310 20116 38354
rect 20272 38010 20300 39986
rect 20364 38894 20392 40394
rect 20352 38888 20404 38894
rect 20352 38830 20404 38836
rect 20456 38842 20484 41550
rect 20536 41540 20588 41546
rect 20536 41482 20588 41488
rect 20548 40905 20576 41482
rect 20534 40896 20590 40905
rect 20534 40831 20590 40840
rect 20640 39098 20668 42162
rect 21272 41676 21324 41682
rect 21272 41618 21324 41624
rect 21284 41449 21312 41618
rect 21270 41440 21326 41449
rect 20729 41372 21037 41381
rect 21270 41375 21326 41384
rect 20729 41370 20735 41372
rect 20791 41370 20815 41372
rect 20871 41370 20895 41372
rect 20951 41370 20975 41372
rect 21031 41370 21037 41372
rect 20791 41318 20793 41370
rect 20973 41318 20975 41370
rect 20729 41316 20735 41318
rect 20791 41316 20815 41318
rect 20871 41316 20895 41318
rect 20951 41316 20975 41318
rect 21031 41316 21037 41318
rect 20729 41307 21037 41316
rect 21088 41132 21140 41138
rect 21088 41074 21140 41080
rect 20729 40284 21037 40293
rect 20729 40282 20735 40284
rect 20791 40282 20815 40284
rect 20871 40282 20895 40284
rect 20951 40282 20975 40284
rect 21031 40282 21037 40284
rect 20791 40230 20793 40282
rect 20973 40230 20975 40282
rect 20729 40228 20735 40230
rect 20791 40228 20815 40230
rect 20871 40228 20895 40230
rect 20951 40228 20975 40230
rect 21031 40228 21037 40230
rect 20729 40219 21037 40228
rect 20996 39840 21048 39846
rect 20994 39808 20996 39817
rect 21048 39808 21050 39817
rect 20994 39743 21050 39752
rect 20729 39196 21037 39205
rect 20729 39194 20735 39196
rect 20791 39194 20815 39196
rect 20871 39194 20895 39196
rect 20951 39194 20975 39196
rect 21031 39194 21037 39196
rect 20791 39142 20793 39194
rect 20973 39142 20975 39194
rect 20729 39140 20735 39142
rect 20791 39140 20815 39142
rect 20871 39140 20895 39142
rect 20951 39140 20975 39142
rect 21031 39140 21037 39142
rect 20729 39131 21037 39140
rect 20628 39092 20680 39098
rect 20628 39034 20680 39040
rect 20456 38814 20576 38842
rect 20444 38752 20496 38758
rect 20442 38720 20444 38729
rect 20496 38720 20498 38729
rect 20442 38655 20498 38664
rect 20260 38004 20312 38010
rect 20260 37946 20312 37952
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 20180 37262 20208 37810
rect 20444 37664 20496 37670
rect 20442 37632 20444 37641
rect 20496 37632 20498 37641
rect 20442 37567 20498 37576
rect 20260 37324 20312 37330
rect 20260 37266 20312 37272
rect 20168 37256 20220 37262
rect 20272 37233 20300 37266
rect 20168 37198 20220 37204
rect 20258 37224 20314 37233
rect 20258 37159 20314 37168
rect 20168 36780 20220 36786
rect 20168 36722 20220 36728
rect 20180 36378 20208 36722
rect 20168 36372 20220 36378
rect 20168 36314 20220 36320
rect 20076 36304 20128 36310
rect 20076 36246 20128 36252
rect 19984 35760 20036 35766
rect 19984 35702 20036 35708
rect 20088 35698 20116 36246
rect 20548 36174 20576 38814
rect 20729 38108 21037 38117
rect 20729 38106 20735 38108
rect 20791 38106 20815 38108
rect 20871 38106 20895 38108
rect 20951 38106 20975 38108
rect 21031 38106 21037 38108
rect 20791 38054 20793 38106
rect 20973 38054 20975 38106
rect 20729 38052 20735 38054
rect 20791 38052 20815 38054
rect 20871 38052 20895 38054
rect 20951 38052 20975 38054
rect 21031 38052 21037 38054
rect 20729 38043 21037 38052
rect 20729 37020 21037 37029
rect 20729 37018 20735 37020
rect 20791 37018 20815 37020
rect 20871 37018 20895 37020
rect 20951 37018 20975 37020
rect 21031 37018 21037 37020
rect 20791 36966 20793 37018
rect 20973 36966 20975 37018
rect 20729 36964 20735 36966
rect 20791 36964 20815 36966
rect 20871 36964 20895 36966
rect 20951 36964 20975 36966
rect 21031 36964 21037 36966
rect 20729 36955 21037 36964
rect 20536 36168 20588 36174
rect 20536 36110 20588 36116
rect 20729 35932 21037 35941
rect 20729 35930 20735 35932
rect 20791 35930 20815 35932
rect 20871 35930 20895 35932
rect 20951 35930 20975 35932
rect 21031 35930 21037 35932
rect 20791 35878 20793 35930
rect 20973 35878 20975 35930
rect 20729 35876 20735 35878
rect 20791 35876 20815 35878
rect 20871 35876 20895 35878
rect 20951 35876 20975 35878
rect 21031 35876 21037 35878
rect 20729 35867 21037 35876
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 20536 35692 20588 35698
rect 20536 35634 20588 35640
rect 19892 35556 19944 35562
rect 19892 35498 19944 35504
rect 19708 35488 19760 35494
rect 19708 35430 19760 35436
rect 19984 35488 20036 35494
rect 19984 35430 20036 35436
rect 20350 35456 20406 35465
rect 19524 34196 19576 34202
rect 19524 34138 19576 34144
rect 19616 34196 19668 34202
rect 19616 34138 19668 34144
rect 19430 34096 19486 34105
rect 19430 34031 19486 34040
rect 19432 33992 19484 33998
rect 19432 33934 19484 33940
rect 19340 33312 19392 33318
rect 19338 33280 19340 33289
rect 19392 33280 19394 33289
rect 19338 33215 19394 33224
rect 19444 33114 19472 33934
rect 19536 33833 19564 34138
rect 19616 33992 19668 33998
rect 19720 33969 19748 35430
rect 19892 34604 19944 34610
rect 19892 34546 19944 34552
rect 19616 33934 19668 33940
rect 19706 33960 19762 33969
rect 19522 33824 19578 33833
rect 19522 33759 19578 33768
rect 19628 33658 19656 33934
rect 19706 33895 19762 33904
rect 19800 33856 19852 33862
rect 19800 33798 19852 33804
rect 19616 33652 19668 33658
rect 19616 33594 19668 33600
rect 19524 33516 19576 33522
rect 19524 33458 19576 33464
rect 19432 33108 19484 33114
rect 19432 33050 19484 33056
rect 18984 32966 19288 32994
rect 18984 30376 19012 32966
rect 19340 32904 19392 32910
rect 19168 32864 19340 32892
rect 19062 31920 19118 31929
rect 19062 31855 19064 31864
rect 19116 31855 19118 31864
rect 19064 31826 19116 31832
rect 19064 31748 19116 31754
rect 19064 31690 19116 31696
rect 19076 31278 19104 31690
rect 19064 31272 19116 31278
rect 19064 31214 19116 31220
rect 19062 31104 19118 31113
rect 19168 31090 19196 32864
rect 19340 32846 19392 32852
rect 19432 32768 19484 32774
rect 19430 32736 19432 32745
rect 19484 32736 19486 32745
rect 19430 32671 19486 32680
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 19352 31754 19380 32506
rect 19536 32502 19564 33458
rect 19706 33280 19762 33289
rect 19706 33215 19762 33224
rect 19720 33114 19748 33215
rect 19708 33108 19760 33114
rect 19708 33050 19760 33056
rect 19616 32836 19668 32842
rect 19616 32778 19668 32784
rect 19524 32496 19576 32502
rect 19430 32464 19486 32473
rect 19524 32438 19576 32444
rect 19430 32399 19486 32408
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19248 31340 19300 31346
rect 19248 31282 19300 31288
rect 19260 31210 19288 31282
rect 19248 31204 19300 31210
rect 19248 31146 19300 31152
rect 19118 31062 19196 31090
rect 19246 31104 19302 31113
rect 19062 31039 19118 31048
rect 19246 31039 19302 31048
rect 19260 30938 19288 31039
rect 19444 30954 19472 32399
rect 19628 31754 19656 32778
rect 19812 32042 19840 33798
rect 19904 32298 19932 34546
rect 19996 32910 20024 35430
rect 20350 35391 20406 35400
rect 20364 35290 20392 35391
rect 20352 35284 20404 35290
rect 20352 35226 20404 35232
rect 20444 35148 20496 35154
rect 20444 35090 20496 35096
rect 20456 34490 20484 35090
rect 20548 34746 20576 35634
rect 20628 35624 20680 35630
rect 20628 35566 20680 35572
rect 20536 34740 20588 34746
rect 20536 34682 20588 34688
rect 20456 34462 20576 34490
rect 20352 34400 20404 34406
rect 20444 34400 20496 34406
rect 20352 34342 20404 34348
rect 20442 34368 20444 34377
rect 20496 34368 20498 34377
rect 20076 34060 20128 34066
rect 20076 34002 20128 34008
rect 20088 32910 20116 34002
rect 20168 33992 20220 33998
rect 20168 33934 20220 33940
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 20076 32904 20128 32910
rect 20076 32846 20128 32852
rect 20074 32736 20130 32745
rect 20074 32671 20130 32680
rect 19892 32292 19944 32298
rect 19892 32234 19944 32240
rect 19720 32026 19840 32042
rect 19708 32020 19840 32026
rect 19760 32014 19840 32020
rect 19708 31962 19760 31968
rect 19890 31784 19946 31793
rect 19616 31748 19668 31754
rect 19890 31719 19946 31728
rect 19616 31690 19668 31696
rect 19616 31340 19668 31346
rect 19616 31282 19668 31288
rect 19800 31340 19852 31346
rect 19800 31282 19852 31288
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19352 30926 19472 30954
rect 19154 30832 19210 30841
rect 19154 30767 19210 30776
rect 18984 30348 19104 30376
rect 18800 30246 18920 30274
rect 18972 30252 19024 30258
rect 18696 30048 18748 30054
rect 18696 29990 18748 29996
rect 18604 29708 18656 29714
rect 18604 29650 18656 29656
rect 18604 29504 18656 29510
rect 18604 29446 18656 29452
rect 18257 28860 18565 28869
rect 18257 28858 18263 28860
rect 18319 28858 18343 28860
rect 18399 28858 18423 28860
rect 18479 28858 18503 28860
rect 18559 28858 18565 28860
rect 18319 28806 18321 28858
rect 18501 28806 18503 28858
rect 18257 28804 18263 28806
rect 18319 28804 18343 28806
rect 18399 28804 18423 28806
rect 18479 28804 18503 28806
rect 18559 28804 18565 28806
rect 18257 28795 18565 28804
rect 18064 28478 18184 28506
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 17774 28112 17830 28121
rect 17774 28047 17830 28056
rect 17868 28008 17920 28014
rect 17920 27968 18000 27996
rect 17868 27950 17920 27956
rect 17776 27872 17828 27878
rect 17776 27814 17828 27820
rect 17788 27674 17816 27814
rect 17776 27668 17828 27674
rect 17776 27610 17828 27616
rect 17776 27328 17828 27334
rect 17776 27270 17828 27276
rect 17604 26846 17724 26874
rect 17500 20800 17552 20806
rect 17500 20742 17552 20748
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 17512 17338 17540 20402
rect 17604 19802 17632 26846
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17696 26382 17724 26726
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17788 25770 17816 27270
rect 17868 26988 17920 26994
rect 17868 26930 17920 26936
rect 17880 26790 17908 26930
rect 17868 26784 17920 26790
rect 17868 26726 17920 26732
rect 17868 26580 17920 26586
rect 17868 26522 17920 26528
rect 17776 25764 17828 25770
rect 17776 25706 17828 25712
rect 17880 25265 17908 26522
rect 17866 25256 17922 25265
rect 17866 25191 17922 25200
rect 17868 25152 17920 25158
rect 17868 25094 17920 25100
rect 17880 24954 17908 25094
rect 17868 24948 17920 24954
rect 17868 24890 17920 24896
rect 17684 24744 17736 24750
rect 17684 24686 17736 24692
rect 17696 24410 17724 24686
rect 17868 24608 17920 24614
rect 17868 24550 17920 24556
rect 17684 24404 17736 24410
rect 17684 24346 17736 24352
rect 17880 24206 17908 24550
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17774 23352 17830 23361
rect 17774 23287 17830 23296
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 17696 21162 17724 23122
rect 17788 21457 17816 23287
rect 17880 23066 17908 23802
rect 17972 23186 18000 27968
rect 18064 27606 18092 28358
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 18052 27328 18104 27334
rect 18052 27270 18104 27276
rect 18064 26586 18092 27270
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 18156 26466 18184 28478
rect 18257 27772 18565 27781
rect 18257 27770 18263 27772
rect 18319 27770 18343 27772
rect 18399 27770 18423 27772
rect 18479 27770 18503 27772
rect 18559 27770 18565 27772
rect 18319 27718 18321 27770
rect 18501 27718 18503 27770
rect 18257 27716 18263 27718
rect 18319 27716 18343 27718
rect 18399 27716 18423 27718
rect 18479 27716 18503 27718
rect 18559 27716 18565 27718
rect 18257 27707 18565 27716
rect 18616 27033 18644 29446
rect 18602 27024 18658 27033
rect 18602 26959 18658 26968
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 18257 26684 18565 26693
rect 18257 26682 18263 26684
rect 18319 26682 18343 26684
rect 18399 26682 18423 26684
rect 18479 26682 18503 26684
rect 18559 26682 18565 26684
rect 18319 26630 18321 26682
rect 18501 26630 18503 26682
rect 18257 26628 18263 26630
rect 18319 26628 18343 26630
rect 18399 26628 18423 26630
rect 18479 26628 18503 26630
rect 18559 26628 18565 26630
rect 18257 26619 18565 26628
rect 18616 26586 18644 26862
rect 18604 26580 18656 26586
rect 18604 26522 18656 26528
rect 18064 26438 18184 26466
rect 18064 23322 18092 26438
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 18156 25838 18184 26318
rect 18524 25945 18552 26318
rect 18708 26024 18736 29990
rect 18800 28150 18828 30246
rect 18972 30194 19024 30200
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18892 29306 18920 29990
rect 18984 29850 19012 30194
rect 18972 29844 19024 29850
rect 18972 29786 19024 29792
rect 18880 29300 18932 29306
rect 19076 29288 19104 30348
rect 18880 29242 18932 29248
rect 18984 29260 19104 29288
rect 18880 29164 18932 29170
rect 18880 29106 18932 29112
rect 18892 28762 18920 29106
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18788 28144 18840 28150
rect 18788 28086 18840 28092
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18788 27464 18840 27470
rect 18788 27406 18840 27412
rect 18800 27130 18828 27406
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 18892 26976 18920 28018
rect 18984 27130 19012 29260
rect 19062 29200 19118 29209
rect 19168 29170 19196 30767
rect 19246 30152 19302 30161
rect 19246 30087 19302 30096
rect 19260 29209 19288 30087
rect 19246 29200 19302 29209
rect 19062 29135 19118 29144
rect 19156 29164 19208 29170
rect 19076 28150 19104 29135
rect 19246 29135 19302 29144
rect 19156 29106 19208 29112
rect 19248 29096 19300 29102
rect 19248 29038 19300 29044
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19168 28642 19196 28970
rect 19260 28762 19288 29038
rect 19248 28756 19300 28762
rect 19248 28698 19300 28704
rect 19168 28614 19288 28642
rect 19156 28484 19208 28490
rect 19156 28426 19208 28432
rect 19064 28144 19116 28150
rect 19064 28086 19116 28092
rect 19168 27130 19196 28426
rect 19260 28257 19288 28614
rect 19246 28248 19302 28257
rect 19246 28183 19302 28192
rect 19246 28112 19302 28121
rect 19246 28047 19302 28056
rect 18972 27124 19024 27130
rect 18972 27066 19024 27072
rect 19156 27124 19208 27130
rect 19156 27066 19208 27072
rect 18892 26948 19012 26976
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18878 26888 18934 26897
rect 18800 26518 18828 26862
rect 18878 26823 18934 26832
rect 18788 26512 18840 26518
rect 18788 26454 18840 26460
rect 18892 26382 18920 26823
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18880 26376 18932 26382
rect 18880 26318 18932 26324
rect 18800 26042 18828 26318
rect 18616 25996 18736 26024
rect 18788 26036 18840 26042
rect 18510 25936 18566 25945
rect 18510 25871 18566 25880
rect 18144 25832 18196 25838
rect 18144 25774 18196 25780
rect 18156 24750 18184 25774
rect 18257 25596 18565 25605
rect 18257 25594 18263 25596
rect 18319 25594 18343 25596
rect 18399 25594 18423 25596
rect 18479 25594 18503 25596
rect 18559 25594 18565 25596
rect 18319 25542 18321 25594
rect 18501 25542 18503 25594
rect 18257 25540 18263 25542
rect 18319 25540 18343 25542
rect 18399 25540 18423 25542
rect 18479 25540 18503 25542
rect 18559 25540 18565 25542
rect 18257 25531 18565 25540
rect 18616 24886 18644 25996
rect 18788 25978 18840 25984
rect 18892 25922 18920 26318
rect 18708 25906 18920 25922
rect 18696 25900 18920 25906
rect 18748 25894 18920 25900
rect 18696 25842 18748 25848
rect 18984 25786 19012 26948
rect 19064 26852 19116 26858
rect 19064 26794 19116 26800
rect 19076 26217 19104 26794
rect 19062 26208 19118 26217
rect 19062 26143 19118 26152
rect 18800 25758 19012 25786
rect 18604 24880 18656 24886
rect 18604 24822 18656 24828
rect 18144 24744 18196 24750
rect 18144 24686 18196 24692
rect 18052 23316 18104 23322
rect 18052 23258 18104 23264
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17880 23038 18092 23066
rect 17774 21448 17830 21457
rect 17774 21383 17830 21392
rect 17696 21134 17908 21162
rect 17776 20596 17828 20602
rect 17776 20538 17828 20544
rect 17788 20058 17816 20538
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17774 19952 17830 19961
rect 17774 19887 17830 19896
rect 17604 19774 17724 19802
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 19378 17632 19654
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17590 17640 17646 17649
rect 17696 17626 17724 19774
rect 17788 19334 17816 19887
rect 17880 19514 17908 21134
rect 17960 20256 18012 20262
rect 17960 20198 18012 20204
rect 17868 19508 17920 19514
rect 17868 19450 17920 19456
rect 17788 19306 17908 19334
rect 17646 17598 17724 17626
rect 17590 17575 17646 17584
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17776 17264 17828 17270
rect 17776 17206 17828 17212
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17236 15660 17448 15688
rect 17236 11529 17264 15660
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17328 13841 17356 15506
rect 17408 15496 17460 15502
rect 17408 15438 17460 15444
rect 17420 14929 17448 15438
rect 17512 15026 17540 16730
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17696 15416 17724 16390
rect 17788 16017 17816 17206
rect 17880 16998 17908 19306
rect 17972 18290 18000 20198
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17972 17202 18000 18226
rect 18064 17610 18092 23038
rect 18156 22506 18184 24686
rect 18604 24608 18656 24614
rect 18604 24550 18656 24556
rect 18257 24508 18565 24517
rect 18257 24506 18263 24508
rect 18319 24506 18343 24508
rect 18399 24506 18423 24508
rect 18479 24506 18503 24508
rect 18559 24506 18565 24508
rect 18319 24454 18321 24506
rect 18501 24454 18503 24506
rect 18257 24452 18263 24454
rect 18319 24452 18343 24454
rect 18399 24452 18423 24454
rect 18479 24452 18503 24454
rect 18559 24452 18565 24454
rect 18257 24443 18565 24452
rect 18236 24404 18288 24410
rect 18616 24392 18644 24550
rect 18288 24364 18644 24392
rect 18236 24346 18288 24352
rect 18604 24064 18656 24070
rect 18604 24006 18656 24012
rect 18257 23420 18565 23429
rect 18257 23418 18263 23420
rect 18319 23418 18343 23420
rect 18399 23418 18423 23420
rect 18479 23418 18503 23420
rect 18559 23418 18565 23420
rect 18319 23366 18321 23418
rect 18501 23366 18503 23418
rect 18257 23364 18263 23366
rect 18319 23364 18343 23366
rect 18399 23364 18423 23366
rect 18479 23364 18503 23366
rect 18559 23364 18565 23366
rect 18257 23355 18565 23364
rect 18616 23118 18644 24006
rect 18696 23656 18748 23662
rect 18696 23598 18748 23604
rect 18708 23322 18736 23598
rect 18696 23316 18748 23322
rect 18696 23258 18748 23264
rect 18604 23112 18656 23118
rect 18604 23054 18656 23060
rect 18696 22976 18748 22982
rect 18696 22918 18748 22924
rect 18708 22710 18736 22918
rect 18696 22704 18748 22710
rect 18696 22646 18748 22652
rect 18512 22636 18564 22642
rect 18564 22596 18644 22624
rect 18512 22578 18564 22584
rect 18144 22500 18196 22506
rect 18144 22442 18196 22448
rect 18156 22030 18184 22442
rect 18257 22332 18565 22341
rect 18257 22330 18263 22332
rect 18319 22330 18343 22332
rect 18399 22330 18423 22332
rect 18479 22330 18503 22332
rect 18559 22330 18565 22332
rect 18319 22278 18321 22330
rect 18501 22278 18503 22330
rect 18257 22276 18263 22278
rect 18319 22276 18343 22278
rect 18399 22276 18423 22278
rect 18479 22276 18503 22278
rect 18559 22276 18565 22278
rect 18257 22267 18565 22276
rect 18616 22234 18644 22596
rect 18604 22228 18656 22234
rect 18604 22170 18656 22176
rect 18420 22160 18472 22166
rect 18696 22160 18748 22166
rect 18420 22102 18472 22108
rect 18616 22108 18696 22114
rect 18616 22102 18748 22108
rect 18328 22092 18380 22098
rect 18248 22052 18328 22080
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 18144 21344 18196 21350
rect 18248 21332 18276 22052
rect 18328 22034 18380 22040
rect 18432 22030 18460 22102
rect 18616 22086 18736 22102
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18340 21690 18368 21830
rect 18328 21684 18380 21690
rect 18328 21626 18380 21632
rect 18196 21304 18276 21332
rect 18144 21286 18196 21292
rect 18156 19922 18184 21286
rect 18257 21244 18565 21253
rect 18257 21242 18263 21244
rect 18319 21242 18343 21244
rect 18399 21242 18423 21244
rect 18479 21242 18503 21244
rect 18559 21242 18565 21244
rect 18319 21190 18321 21242
rect 18501 21190 18503 21242
rect 18257 21188 18263 21190
rect 18319 21188 18343 21190
rect 18399 21188 18423 21190
rect 18479 21188 18503 21190
rect 18559 21188 18565 21190
rect 18257 21179 18565 21188
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18432 20466 18460 21082
rect 18420 20460 18472 20466
rect 18420 20402 18472 20408
rect 18257 20156 18565 20165
rect 18257 20154 18263 20156
rect 18319 20154 18343 20156
rect 18399 20154 18423 20156
rect 18479 20154 18503 20156
rect 18559 20154 18565 20156
rect 18319 20102 18321 20154
rect 18501 20102 18503 20154
rect 18257 20100 18263 20102
rect 18319 20100 18343 20102
rect 18399 20100 18423 20102
rect 18479 20100 18503 20102
rect 18559 20100 18565 20102
rect 18257 20091 18565 20100
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18156 19242 18184 19858
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18432 19514 18460 19654
rect 18420 19508 18472 19514
rect 18420 19450 18472 19456
rect 18144 19236 18196 19242
rect 18144 19178 18196 19184
rect 18257 19068 18565 19077
rect 18257 19066 18263 19068
rect 18319 19066 18343 19068
rect 18399 19066 18423 19068
rect 18479 19066 18503 19068
rect 18559 19066 18565 19068
rect 18319 19014 18321 19066
rect 18501 19014 18503 19066
rect 18257 19012 18263 19014
rect 18319 19012 18343 19014
rect 18399 19012 18423 19014
rect 18479 19012 18503 19014
rect 18559 19012 18565 19014
rect 18257 19003 18565 19012
rect 18257 17980 18565 17989
rect 18257 17978 18263 17980
rect 18319 17978 18343 17980
rect 18399 17978 18423 17980
rect 18479 17978 18503 17980
rect 18559 17978 18565 17980
rect 18319 17926 18321 17978
rect 18501 17926 18503 17978
rect 18257 17924 18263 17926
rect 18319 17924 18343 17926
rect 18399 17924 18423 17926
rect 18479 17924 18503 17926
rect 18559 17924 18565 17926
rect 18257 17915 18565 17924
rect 18052 17604 18104 17610
rect 18052 17546 18104 17552
rect 17960 17196 18012 17202
rect 17960 17138 18012 17144
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17868 16992 17920 16998
rect 17868 16934 17920 16940
rect 17972 16794 18000 17138
rect 18064 17105 18092 17138
rect 18050 17096 18106 17105
rect 18050 17031 18106 17040
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17960 16788 18012 16794
rect 17960 16730 18012 16736
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17774 16008 17830 16017
rect 17774 15943 17830 15952
rect 17604 15388 17724 15416
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17406 14920 17462 14929
rect 17406 14855 17462 14864
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17314 13832 17370 13841
rect 17314 13767 17370 13776
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 12306 17356 13670
rect 17420 13530 17448 14214
rect 17512 13938 17540 14962
rect 17500 13932 17552 13938
rect 17500 13874 17552 13880
rect 17408 13524 17460 13530
rect 17408 13466 17460 13472
rect 17316 12300 17368 12306
rect 17316 12242 17368 12248
rect 17328 12209 17356 12242
rect 17314 12200 17370 12209
rect 17314 12135 17370 12144
rect 17222 11520 17278 11529
rect 17222 11455 17278 11464
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17420 11082 17448 13466
rect 17512 11762 17540 13874
rect 17604 13734 17632 15388
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 17696 14385 17724 15030
rect 17682 14376 17738 14385
rect 17682 14311 17738 14320
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17590 13560 17646 13569
rect 17590 13495 17646 13504
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11150 17540 11494
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17224 11076 17276 11082
rect 17224 11018 17276 11024
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17132 10736 17184 10742
rect 17038 10704 17094 10713
rect 17132 10678 17184 10684
rect 17038 10639 17040 10648
rect 17092 10639 17094 10648
rect 17040 10610 17092 10616
rect 17038 10296 17094 10305
rect 17038 10231 17094 10240
rect 17052 9353 17080 10231
rect 17038 9344 17094 9353
rect 17038 9279 17094 9288
rect 16960 9166 17080 9194
rect 17144 9178 17172 10678
rect 17236 10130 17264 11018
rect 17408 10532 17460 10538
rect 17408 10474 17460 10480
rect 17420 10130 17448 10474
rect 17224 10124 17276 10130
rect 17224 10066 17276 10072
rect 17408 10124 17460 10130
rect 17408 10066 17460 10072
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 16868 7500 16988 7528
rect 16764 7472 16816 7478
rect 16764 7414 16816 7420
rect 16488 7336 16540 7342
rect 16672 7336 16724 7342
rect 16488 7278 16540 7284
rect 16578 7304 16634 7313
rect 16672 7278 16724 7284
rect 16578 7239 16634 7248
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16394 7032 16450 7041
rect 16394 6967 16450 6976
rect 16210 6423 16266 6432
rect 16304 6452 16356 6458
rect 16028 6394 16080 6400
rect 16304 6394 16356 6400
rect 15764 5846 15792 6394
rect 16408 6338 16436 6967
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16212 6316 16264 6322
rect 16212 6258 16264 6264
rect 16316 6310 16436 6338
rect 16592 6322 16620 7239
rect 16684 6866 16712 7278
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 16684 6322 16712 6802
rect 16776 6440 16804 7414
rect 16960 7410 16988 7500
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16868 6769 16896 7346
rect 17052 6798 17080 9166
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17236 8634 17264 9658
rect 17316 8900 17368 8906
rect 17420 8888 17448 10066
rect 17604 9330 17632 13495
rect 17696 12889 17724 14214
rect 17682 12880 17738 12889
rect 17682 12815 17738 12824
rect 17682 12336 17738 12345
rect 17682 12271 17738 12280
rect 17696 11014 17724 12271
rect 17788 11665 17816 15943
rect 17868 13252 17920 13258
rect 17868 13194 17920 13200
rect 17880 11937 17908 13194
rect 17866 11928 17922 11937
rect 17866 11863 17922 11872
rect 17972 11812 18000 16594
rect 18064 16561 18092 16934
rect 18257 16892 18565 16901
rect 18257 16890 18263 16892
rect 18319 16890 18343 16892
rect 18399 16890 18423 16892
rect 18479 16890 18503 16892
rect 18559 16890 18565 16892
rect 18319 16838 18321 16890
rect 18501 16838 18503 16890
rect 18257 16836 18263 16838
rect 18319 16836 18343 16838
rect 18399 16836 18423 16838
rect 18479 16836 18503 16838
rect 18559 16836 18565 16838
rect 18257 16827 18565 16836
rect 18420 16584 18472 16590
rect 18050 16552 18106 16561
rect 18420 16526 18472 16532
rect 18050 16487 18106 16496
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18064 16250 18092 16390
rect 18432 16250 18460 16526
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18524 16250 18552 16390
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18512 16244 18564 16250
rect 18512 16186 18564 16192
rect 18257 15804 18565 15813
rect 18257 15802 18263 15804
rect 18319 15802 18343 15804
rect 18399 15802 18423 15804
rect 18479 15802 18503 15804
rect 18559 15802 18565 15804
rect 18319 15750 18321 15802
rect 18501 15750 18503 15802
rect 18257 15748 18263 15750
rect 18319 15748 18343 15750
rect 18399 15748 18423 15750
rect 18479 15748 18503 15750
rect 18559 15748 18565 15750
rect 18257 15739 18565 15748
rect 18418 15600 18474 15609
rect 18474 15558 18552 15586
rect 18418 15535 18474 15544
rect 18524 15026 18552 15558
rect 18616 15366 18644 22086
rect 18800 21128 18828 25758
rect 19064 25492 19116 25498
rect 19064 25434 19116 25440
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 18984 24342 19012 25366
rect 18972 24336 19024 24342
rect 18972 24278 19024 24284
rect 18880 23248 18932 23254
rect 18880 23190 18932 23196
rect 18892 21622 18920 23190
rect 18984 22098 19012 24278
rect 19076 24154 19104 25434
rect 19260 25129 19288 28047
rect 19352 27130 19380 30926
rect 19524 30728 19576 30734
rect 19524 30670 19576 30676
rect 19536 29782 19564 30670
rect 19628 30394 19656 31282
rect 19708 31136 19760 31142
rect 19708 31078 19760 31084
rect 19720 30394 19748 31078
rect 19812 30977 19840 31282
rect 19798 30968 19854 30977
rect 19798 30903 19854 30912
rect 19800 30728 19852 30734
rect 19800 30670 19852 30676
rect 19616 30388 19668 30394
rect 19616 30330 19668 30336
rect 19708 30388 19760 30394
rect 19708 30330 19760 30336
rect 19616 30252 19668 30258
rect 19616 30194 19668 30200
rect 19708 30252 19760 30258
rect 19708 30194 19760 30200
rect 19524 29776 19576 29782
rect 19524 29718 19576 29724
rect 19522 29608 19578 29617
rect 19522 29543 19578 29552
rect 19432 28212 19484 28218
rect 19432 28154 19484 28160
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19340 26512 19392 26518
rect 19338 26480 19340 26489
rect 19392 26480 19394 26489
rect 19338 26415 19394 26424
rect 19340 25152 19392 25158
rect 19246 25120 19302 25129
rect 19444 25140 19472 28154
rect 19536 25294 19564 29543
rect 19628 29306 19656 30194
rect 19616 29300 19668 29306
rect 19616 29242 19668 29248
rect 19616 28960 19668 28966
rect 19616 28902 19668 28908
rect 19628 28762 19656 28902
rect 19616 28756 19668 28762
rect 19616 28698 19668 28704
rect 19720 28694 19748 30194
rect 19812 29102 19840 30670
rect 19904 29850 19932 31719
rect 19984 31680 20036 31686
rect 19984 31622 20036 31628
rect 19996 31278 20024 31622
rect 19984 31272 20036 31278
rect 19984 31214 20036 31220
rect 19984 30592 20036 30598
rect 19984 30534 20036 30540
rect 19892 29844 19944 29850
rect 19892 29786 19944 29792
rect 19892 29164 19944 29170
rect 19892 29106 19944 29112
rect 19800 29096 19852 29102
rect 19800 29038 19852 29044
rect 19800 28960 19852 28966
rect 19800 28902 19852 28908
rect 19708 28688 19760 28694
rect 19708 28630 19760 28636
rect 19720 28218 19748 28630
rect 19708 28212 19760 28218
rect 19708 28154 19760 28160
rect 19812 28150 19840 28902
rect 19616 28144 19668 28150
rect 19616 28086 19668 28092
rect 19800 28144 19852 28150
rect 19800 28086 19852 28092
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19444 25112 19564 25140
rect 19340 25094 19392 25100
rect 19246 25055 19302 25064
rect 19076 24126 19196 24154
rect 19064 23520 19116 23526
rect 19064 23462 19116 23468
rect 19076 23322 19104 23462
rect 19168 23338 19196 24126
rect 19352 23730 19380 25094
rect 19432 24608 19484 24614
rect 19432 24550 19484 24556
rect 19444 23866 19472 24550
rect 19432 23860 19484 23866
rect 19432 23802 19484 23808
rect 19340 23724 19392 23730
rect 19340 23666 19392 23672
rect 19340 23588 19392 23594
rect 19340 23530 19392 23536
rect 19352 23474 19380 23530
rect 19352 23446 19472 23474
rect 19338 23352 19394 23361
rect 19064 23316 19116 23322
rect 19168 23310 19288 23338
rect 19064 23258 19116 23264
rect 19156 23248 19208 23254
rect 19156 23190 19208 23196
rect 19064 22432 19116 22438
rect 19064 22374 19116 22380
rect 18972 22092 19024 22098
rect 18972 22034 19024 22040
rect 19076 22030 19104 22374
rect 19168 22166 19196 23190
rect 19156 22160 19208 22166
rect 19156 22102 19208 22108
rect 19064 22024 19116 22030
rect 19260 21978 19288 23310
rect 19338 23287 19394 23296
rect 19064 21966 19116 21972
rect 18972 21956 19024 21962
rect 18972 21898 19024 21904
rect 19168 21950 19288 21978
rect 18880 21616 18932 21622
rect 18880 21558 18932 21564
rect 18708 21100 18828 21128
rect 18708 19334 18736 21100
rect 18892 21026 18920 21558
rect 18984 21049 19012 21898
rect 19062 21448 19118 21457
rect 19062 21383 19118 21392
rect 18800 20998 18920 21026
rect 18970 21040 19026 21049
rect 18800 20602 18828 20998
rect 18970 20975 19026 20984
rect 18880 20936 18932 20942
rect 18880 20878 18932 20884
rect 18972 20936 19024 20942
rect 18972 20878 19024 20884
rect 18788 20596 18840 20602
rect 18788 20538 18840 20544
rect 18892 20262 18920 20878
rect 18880 20256 18932 20262
rect 18880 20198 18932 20204
rect 18984 20058 19012 20878
rect 18972 20052 19024 20058
rect 18972 19994 19024 20000
rect 19076 19938 19104 21383
rect 18892 19910 19104 19938
rect 18708 19306 18828 19334
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 18358 18736 18566
rect 18696 18352 18748 18358
rect 18696 18294 18748 18300
rect 18800 18204 18828 19306
rect 18708 18176 18828 18204
rect 18708 16658 18736 18176
rect 18892 18034 18920 19910
rect 19168 19768 19196 21950
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19260 21554 19288 21830
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19352 21486 19380 23287
rect 19340 21480 19392 21486
rect 19340 21422 19392 21428
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19340 21344 19392 21350
rect 19340 21286 19392 21292
rect 19260 20346 19288 21286
rect 19352 21010 19380 21286
rect 19340 21004 19392 21010
rect 19340 20946 19392 20952
rect 19444 20942 19472 23446
rect 19536 22545 19564 25112
rect 19628 24857 19656 28086
rect 19706 27704 19762 27713
rect 19762 27662 19840 27690
rect 19904 27674 19932 29106
rect 19996 28558 20024 30534
rect 20088 30190 20116 32671
rect 20180 32230 20208 33934
rect 20260 33516 20312 33522
rect 20260 33458 20312 33464
rect 20272 33425 20300 33458
rect 20258 33416 20314 33425
rect 20258 33351 20314 33360
rect 20364 32881 20392 34342
rect 20442 34303 20498 34312
rect 20444 33312 20496 33318
rect 20442 33280 20444 33289
rect 20496 33280 20498 33289
rect 20442 33215 20498 33224
rect 20548 33096 20576 34462
rect 20456 33068 20576 33096
rect 20350 32872 20406 32881
rect 20350 32807 20406 32816
rect 20168 32224 20220 32230
rect 20168 32166 20220 32172
rect 20260 31680 20312 31686
rect 20260 31622 20312 31628
rect 20272 31482 20300 31622
rect 20260 31476 20312 31482
rect 20260 31418 20312 31424
rect 20456 31226 20484 33068
rect 20536 32836 20588 32842
rect 20536 32778 20588 32784
rect 20548 32201 20576 32778
rect 20534 32192 20590 32201
rect 20534 32127 20590 32136
rect 20640 31822 20668 35566
rect 20729 34844 21037 34853
rect 20729 34842 20735 34844
rect 20791 34842 20815 34844
rect 20871 34842 20895 34844
rect 20951 34842 20975 34844
rect 21031 34842 21037 34844
rect 20791 34790 20793 34842
rect 20973 34790 20975 34842
rect 20729 34788 20735 34790
rect 20791 34788 20815 34790
rect 20871 34788 20895 34790
rect 20951 34788 20975 34790
rect 21031 34788 21037 34790
rect 20729 34779 21037 34788
rect 20729 33756 21037 33765
rect 20729 33754 20735 33756
rect 20791 33754 20815 33756
rect 20871 33754 20895 33756
rect 20951 33754 20975 33756
rect 21031 33754 21037 33756
rect 20791 33702 20793 33754
rect 20973 33702 20975 33754
rect 20729 33700 20735 33702
rect 20791 33700 20815 33702
rect 20871 33700 20895 33702
rect 20951 33700 20975 33702
rect 21031 33700 21037 33702
rect 20729 33691 21037 33700
rect 20729 32668 21037 32677
rect 20729 32666 20735 32668
rect 20791 32666 20815 32668
rect 20871 32666 20895 32668
rect 20951 32666 20975 32668
rect 21031 32666 21037 32668
rect 20791 32614 20793 32666
rect 20973 32614 20975 32666
rect 20729 32612 20735 32614
rect 20791 32612 20815 32614
rect 20871 32612 20895 32614
rect 20951 32612 20975 32614
rect 21031 32612 21037 32614
rect 20729 32603 21037 32612
rect 20628 31816 20680 31822
rect 20628 31758 20680 31764
rect 20729 31580 21037 31589
rect 20729 31578 20735 31580
rect 20791 31578 20815 31580
rect 20871 31578 20895 31580
rect 20951 31578 20975 31580
rect 21031 31578 21037 31580
rect 20791 31526 20793 31578
rect 20973 31526 20975 31578
rect 20729 31524 20735 31526
rect 20791 31524 20815 31526
rect 20871 31524 20895 31526
rect 20951 31524 20975 31526
rect 21031 31524 21037 31526
rect 20729 31515 21037 31524
rect 20628 31476 20680 31482
rect 20364 31198 20484 31226
rect 20548 31436 20628 31464
rect 20364 30818 20392 31198
rect 20444 31136 20496 31142
rect 20442 31104 20444 31113
rect 20496 31104 20498 31113
rect 20442 31039 20498 31048
rect 20364 30790 20484 30818
rect 20168 30388 20220 30394
rect 20168 30330 20220 30336
rect 20076 30184 20128 30190
rect 20076 30126 20128 30132
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20088 28762 20116 29990
rect 20180 29238 20208 30330
rect 20456 30138 20484 30790
rect 20272 30110 20484 30138
rect 20168 29232 20220 29238
rect 20168 29174 20220 29180
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 19984 28416 20036 28422
rect 19984 28358 20036 28364
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 19706 27639 19762 27648
rect 19708 26784 19760 26790
rect 19708 26726 19760 26732
rect 19614 24848 19670 24857
rect 19614 24783 19670 24792
rect 19616 24744 19668 24750
rect 19616 24686 19668 24692
rect 19628 24256 19656 24686
rect 19720 24426 19748 26726
rect 19812 24562 19840 27662
rect 19892 27668 19944 27674
rect 19892 27610 19944 27616
rect 19996 27470 20024 28358
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19892 26784 19944 26790
rect 19892 26726 19944 26732
rect 19904 25673 19932 26726
rect 19890 25664 19946 25673
rect 19890 25599 19946 25608
rect 19812 24534 19932 24562
rect 19720 24398 19840 24426
rect 19628 24228 19748 24256
rect 19616 24132 19668 24138
rect 19616 24074 19668 24080
rect 19522 22536 19578 22545
rect 19522 22471 19578 22480
rect 19522 22400 19578 22409
rect 19522 22335 19578 22344
rect 19536 21706 19564 22335
rect 19628 21842 19656 24074
rect 19720 23254 19748 24228
rect 19708 23248 19760 23254
rect 19708 23190 19760 23196
rect 19708 23112 19760 23118
rect 19708 23054 19760 23060
rect 19720 22778 19748 23054
rect 19708 22772 19760 22778
rect 19708 22714 19760 22720
rect 19706 22536 19762 22545
rect 19706 22471 19762 22480
rect 19720 21962 19748 22471
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 19628 21814 19748 21842
rect 19536 21678 19656 21706
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19352 20466 19380 20810
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19260 20318 19472 20346
rect 19340 19780 19392 19786
rect 19168 19740 19340 19768
rect 19340 19722 19392 19728
rect 19064 19712 19116 19718
rect 19064 19654 19116 19660
rect 18872 18006 18920 18034
rect 18872 17898 18900 18006
rect 18800 17870 18900 17898
rect 18800 17762 18828 17870
rect 18800 17734 18920 17762
rect 18788 17196 18840 17202
rect 18788 17138 18840 17144
rect 18696 16652 18748 16658
rect 18696 16594 18748 16600
rect 18800 16590 18828 17138
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18892 16454 18920 17734
rect 19076 17660 19104 19654
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19156 19168 19208 19174
rect 19156 19110 19208 19116
rect 19248 19168 19300 19174
rect 19248 19110 19300 19116
rect 19168 18358 19196 19110
rect 19156 18352 19208 18358
rect 19156 18294 19208 18300
rect 19260 17882 19288 19110
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19156 17672 19208 17678
rect 19076 17632 19156 17660
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18694 16144 18750 16153
rect 18694 16079 18750 16088
rect 18708 16046 18736 16079
rect 18696 16040 18748 16046
rect 19076 16028 19104 17632
rect 19156 17614 19208 17620
rect 18748 16000 19104 16028
rect 18696 15982 18748 15988
rect 18696 15496 18748 15502
rect 18696 15438 18748 15444
rect 18604 15360 18656 15366
rect 18604 15302 18656 15308
rect 18708 15201 18736 15438
rect 18788 15360 18840 15366
rect 18840 15320 18920 15348
rect 18788 15302 18840 15308
rect 18694 15192 18750 15201
rect 18694 15127 18750 15136
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18696 15020 18748 15026
rect 18748 14980 18828 15008
rect 18696 14962 18748 14968
rect 18052 14816 18104 14822
rect 18052 14758 18104 14764
rect 18064 14006 18092 14758
rect 18156 14414 18184 14962
rect 18604 14816 18656 14822
rect 18604 14758 18656 14764
rect 18257 14716 18565 14725
rect 18257 14714 18263 14716
rect 18319 14714 18343 14716
rect 18399 14714 18423 14716
rect 18479 14714 18503 14716
rect 18559 14714 18565 14716
rect 18319 14662 18321 14714
rect 18501 14662 18503 14714
rect 18257 14660 18263 14662
rect 18319 14660 18343 14662
rect 18399 14660 18423 14662
rect 18479 14660 18503 14662
rect 18559 14660 18565 14662
rect 18257 14651 18565 14660
rect 18616 14618 18644 14758
rect 18604 14612 18656 14618
rect 18604 14554 18656 14560
rect 18696 14544 18748 14550
rect 18696 14486 18748 14492
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18234 14376 18290 14385
rect 18234 14311 18290 14320
rect 18052 14000 18104 14006
rect 18052 13942 18104 13948
rect 18144 13864 18196 13870
rect 18144 13806 18196 13812
rect 18156 13530 18184 13806
rect 18248 13734 18276 14311
rect 18708 14006 18736 14486
rect 18800 14482 18828 14980
rect 18788 14476 18840 14482
rect 18788 14418 18840 14424
rect 18696 14000 18748 14006
rect 18696 13942 18748 13948
rect 18604 13932 18656 13938
rect 18604 13874 18656 13880
rect 18616 13818 18644 13874
rect 18616 13790 18736 13818
rect 18236 13728 18288 13734
rect 18236 13670 18288 13676
rect 18604 13728 18656 13734
rect 18604 13670 18656 13676
rect 18257 13628 18565 13637
rect 18257 13626 18263 13628
rect 18319 13626 18343 13628
rect 18399 13626 18423 13628
rect 18479 13626 18503 13628
rect 18559 13626 18565 13628
rect 18319 13574 18321 13626
rect 18501 13574 18503 13626
rect 18257 13572 18263 13574
rect 18319 13572 18343 13574
rect 18399 13572 18423 13574
rect 18479 13572 18503 13574
rect 18559 13572 18565 13574
rect 18257 13563 18565 13572
rect 18144 13524 18196 13530
rect 18144 13466 18196 13472
rect 18156 12986 18184 13466
rect 18616 13410 18644 13670
rect 18340 13382 18644 13410
rect 18052 12980 18104 12986
rect 18052 12922 18104 12928
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18064 12238 18092 12922
rect 18340 12782 18368 13382
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18432 12782 18460 13126
rect 18616 12850 18644 13126
rect 18604 12844 18656 12850
rect 18604 12786 18656 12792
rect 18328 12776 18380 12782
rect 18328 12718 18380 12724
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18156 12442 18184 12582
rect 18257 12540 18565 12549
rect 18257 12538 18263 12540
rect 18319 12538 18343 12540
rect 18399 12538 18423 12540
rect 18479 12538 18503 12540
rect 18559 12538 18565 12540
rect 18319 12486 18321 12538
rect 18501 12486 18503 12538
rect 18257 12484 18263 12486
rect 18319 12484 18343 12486
rect 18399 12484 18423 12486
rect 18479 12484 18503 12486
rect 18559 12484 18565 12486
rect 18257 12475 18565 12484
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 18236 12368 18288 12374
rect 18236 12310 18288 12316
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 17880 11784 18000 11812
rect 17774 11656 17830 11665
rect 17774 11591 17830 11600
rect 17788 11082 17816 11591
rect 17776 11076 17828 11082
rect 17776 11018 17828 11024
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17776 10464 17828 10470
rect 17774 10432 17776 10441
rect 17828 10432 17830 10441
rect 17774 10367 17830 10376
rect 17684 10056 17736 10062
rect 17682 10024 17684 10033
rect 17776 10056 17828 10062
rect 17736 10024 17738 10033
rect 17880 10033 17908 11784
rect 18248 11762 18276 12310
rect 18616 12238 18644 12582
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18340 11762 18368 12038
rect 18236 11756 18288 11762
rect 18236 11698 18288 11704
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18248 11642 18276 11698
rect 18524 11694 18552 12038
rect 18064 11614 18276 11642
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 17958 11384 18014 11393
rect 18064 11354 18092 11614
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 17958 11319 18014 11328
rect 18052 11348 18104 11354
rect 17776 9998 17828 10004
rect 17866 10024 17922 10033
rect 17682 9959 17738 9968
rect 17788 9908 17816 9998
rect 17866 9959 17922 9968
rect 17368 8860 17448 8888
rect 17512 9302 17632 9330
rect 17696 9880 17816 9908
rect 17316 8842 17368 8848
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17420 8430 17448 8570
rect 17512 8548 17540 9302
rect 17510 8520 17540 8548
rect 17592 8560 17644 8566
rect 17510 8480 17538 8520
rect 17592 8502 17644 8508
rect 17510 8452 17540 8480
rect 17132 8424 17184 8430
rect 17408 8424 17460 8430
rect 17184 8384 17264 8412
rect 17132 8366 17184 8372
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17144 7478 17172 8230
rect 17236 7478 17264 8384
rect 17408 8366 17460 8372
rect 17408 8288 17460 8294
rect 17408 8230 17460 8236
rect 17314 8120 17370 8129
rect 17314 8055 17370 8064
rect 17132 7472 17184 7478
rect 17132 7414 17184 7420
rect 17224 7472 17276 7478
rect 17224 7414 17276 7420
rect 17130 7304 17186 7313
rect 17130 7239 17186 7248
rect 17040 6792 17092 6798
rect 16854 6760 16910 6769
rect 17040 6734 17092 6740
rect 16854 6695 16910 6704
rect 16776 6412 17080 6440
rect 16762 6352 16818 6361
rect 16580 6316 16632 6322
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15488 5596 15700 5624
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15396 5370 15424 5510
rect 15384 5364 15436 5370
rect 15384 5306 15436 5312
rect 15382 5264 15438 5273
rect 15488 5234 15516 5596
rect 15856 5534 15884 6258
rect 15580 5506 15884 5534
rect 16040 5534 16068 6258
rect 16224 5794 16252 6258
rect 16132 5766 16252 5794
rect 16132 5642 16160 5766
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 16224 5545 16252 5646
rect 16210 5536 16266 5545
rect 16040 5506 16160 5534
rect 15382 5199 15438 5208
rect 15476 5228 15528 5234
rect 15396 5098 15424 5199
rect 15476 5170 15528 5176
rect 15384 5092 15436 5098
rect 15384 5034 15436 5040
rect 15580 4826 15608 5506
rect 15784 5468 16092 5477
rect 15784 5466 15790 5468
rect 15846 5466 15870 5468
rect 15926 5466 15950 5468
rect 16006 5466 16030 5468
rect 16086 5466 16092 5468
rect 15846 5414 15848 5466
rect 16028 5414 16030 5466
rect 15784 5412 15790 5414
rect 15846 5412 15870 5414
rect 15926 5412 15950 5414
rect 16006 5412 16030 5414
rect 16086 5412 16092 5414
rect 15784 5403 16092 5412
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15764 5273 15792 5306
rect 15750 5264 15806 5273
rect 16132 5216 16160 5506
rect 16210 5471 16266 5480
rect 16212 5364 16264 5370
rect 16316 5352 16344 6310
rect 16580 6258 16632 6264
rect 16672 6316 16724 6322
rect 16818 6310 16988 6338
rect 16762 6287 16818 6296
rect 16672 6258 16724 6264
rect 16396 6248 16448 6254
rect 16448 6208 16528 6236
rect 16396 6190 16448 6196
rect 16500 5710 16528 6208
rect 16764 6180 16816 6186
rect 16764 6122 16816 6128
rect 16580 6112 16632 6118
rect 16580 6054 16632 6060
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16316 5324 16436 5352
rect 16212 5306 16264 5312
rect 15750 5199 15806 5208
rect 15856 5188 16160 5216
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15568 4820 15620 4826
rect 15568 4762 15620 4768
rect 15660 4820 15712 4826
rect 15660 4762 15712 4768
rect 15200 4752 15252 4758
rect 15672 4706 15700 4762
rect 15252 4700 15700 4706
rect 15200 4694 15700 4700
rect 15212 4678 15700 4694
rect 15108 4650 15160 4656
rect 14844 4622 15047 4638
rect 14108 4576 14228 4604
rect 14280 4616 14332 4622
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 13740 4406 13952 4434
rect 13740 4282 13768 4406
rect 14108 4282 14136 4576
rect 14740 4616 14792 4622
rect 14646 4584 14702 4593
rect 14280 4558 14332 4564
rect 14384 4542 14646 4570
rect 14188 4480 14240 4486
rect 14186 4448 14188 4457
rect 14240 4448 14242 4457
rect 14186 4383 14242 4392
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 13596 4168 13676 4196
rect 13820 4208 13872 4214
rect 13544 4150 13596 4156
rect 14384 4162 14412 4542
rect 14740 4558 14792 4564
rect 14832 4616 15047 4622
rect 14884 4610 15047 4616
rect 15019 4604 15047 4610
rect 15019 4598 15108 4604
rect 15019 4592 15160 4598
rect 15019 4576 15148 4592
rect 14832 4558 14884 4564
rect 14646 4519 14702 4528
rect 14924 4548 14976 4554
rect 15752 4548 15804 4554
rect 14924 4490 14976 4496
rect 15672 4508 15752 4536
rect 14464 4480 14516 4486
rect 14936 4434 14964 4490
rect 15672 4457 15700 4508
rect 15752 4490 15804 4496
rect 15856 4468 15884 5188
rect 16120 5092 16172 5098
rect 16224 5080 16252 5306
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16172 5052 16252 5080
rect 16120 5034 16172 5040
rect 16316 4536 16344 5170
rect 16224 4508 16344 4536
rect 14516 4428 14964 4434
rect 14464 4422 14964 4428
rect 14476 4406 14964 4422
rect 15658 4448 15714 4457
rect 15856 4440 16160 4468
rect 15658 4383 15714 4392
rect 15784 4380 16092 4389
rect 15784 4378 15790 4380
rect 15846 4378 15870 4380
rect 15926 4378 15950 4380
rect 16006 4378 16030 4380
rect 16086 4378 16092 4380
rect 15846 4326 15848 4378
rect 16028 4326 16030 4378
rect 15784 4324 15790 4326
rect 15846 4324 15870 4326
rect 15926 4324 15950 4326
rect 16006 4324 16030 4326
rect 16086 4324 16092 4326
rect 15290 4312 15346 4321
rect 15784 4315 16092 4324
rect 14660 4270 14964 4298
rect 14660 4196 14688 4270
rect 14936 4214 14964 4270
rect 15346 4270 15516 4298
rect 15290 4247 15346 4256
rect 13872 4156 14412 4162
rect 13820 4150 14412 4156
rect 13832 4134 14412 4150
rect 14476 4168 14688 4196
rect 14832 4208 14884 4214
rect 14476 4128 14504 4168
rect 14832 4150 14884 4156
rect 14924 4208 14976 4214
rect 14924 4150 14976 4156
rect 14442 4100 14504 4128
rect 13820 4072 13872 4078
rect 13360 4014 13412 4020
rect 13450 4040 13506 4049
rect 13266 3975 13322 3984
rect 13176 3946 13228 3952
rect 12360 3754 12388 3946
rect 12806 3904 12862 3913
rect 12806 3839 12862 3848
rect 13015 3904 13071 3913
rect 13015 3839 13071 3848
rect 12256 3732 12308 3738
rect 12360 3726 12572 3754
rect 12256 3674 12308 3680
rect 12164 3664 12216 3670
rect 11992 3590 12112 3618
rect 12440 3664 12492 3670
rect 12164 3606 12216 3612
rect 12438 3632 12440 3641
rect 12492 3632 12494 3641
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11886 3224 11942 3233
rect 11886 3159 11942 3168
rect 11886 3088 11942 3097
rect 11886 3023 11888 3032
rect 11940 3023 11942 3032
rect 11888 2994 11940 3000
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11704 2518 11756 2524
rect 11794 2544 11850 2553
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 11624 1412 11652 2246
rect 11612 1406 11664 1412
rect 11112 1300 11192 1306
rect 11060 1294 11192 1300
rect 11244 1352 11296 1358
rect 11244 1294 11296 1300
rect 11520 1352 11572 1358
rect 11716 1358 11744 2518
rect 11794 2479 11850 2488
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 11808 1873 11836 2314
rect 11900 1970 11928 2858
rect 11992 2394 12020 3470
rect 12084 3176 12112 3590
rect 12544 3618 12572 3726
rect 12820 3618 12848 3839
rect 12898 3768 12954 3777
rect 13029 3754 13057 3839
rect 12898 3703 12954 3712
rect 13004 3726 13057 3754
rect 12912 3670 12940 3703
rect 12544 3590 12664 3618
rect 12728 3602 12848 3618
rect 12900 3664 12952 3670
rect 13004 3652 13032 3726
rect 13188 3720 13216 3946
rect 13372 3924 13400 4014
rect 13450 3975 13506 3984
rect 13556 4020 13820 4026
rect 14442 4060 14470 4100
rect 13556 4014 13872 4020
rect 14384 4032 14470 4060
rect 14844 4060 14872 4150
rect 14844 4032 14962 4060
rect 13556 3998 13860 4014
rect 13912 4004 13964 4010
rect 13556 3924 13584 3998
rect 13912 3946 13964 3952
rect 14004 4004 14056 4010
rect 14384 3992 14412 4032
rect 14934 4026 14962 4032
rect 14934 3998 15332 4026
rect 14056 3964 14412 3992
rect 14571 3964 14872 3992
rect 14004 3946 14056 3952
rect 13372 3896 13584 3924
rect 13924 3913 13952 3946
rect 14464 3936 14516 3942
rect 13910 3904 13966 3913
rect 14571 3924 14599 3964
rect 14516 3896 14599 3924
rect 14844 3924 14872 3964
rect 15200 3936 15252 3942
rect 14844 3896 14964 3924
rect 14464 3878 14516 3884
rect 13312 3836 13620 3845
rect 13910 3839 13966 3848
rect 13312 3834 13318 3836
rect 13374 3834 13398 3836
rect 13454 3834 13478 3836
rect 13534 3834 13558 3836
rect 13614 3834 13620 3836
rect 13374 3782 13376 3834
rect 13556 3782 13558 3834
rect 13312 3780 13318 3782
rect 13374 3780 13398 3782
rect 13454 3780 13478 3782
rect 13534 3780 13558 3782
rect 13614 3780 13620 3782
rect 13312 3771 13620 3780
rect 14094 3768 14150 3777
rect 13740 3726 14044 3754
rect 13740 3720 13768 3726
rect 13188 3692 13768 3720
rect 13820 3664 13872 3670
rect 13004 3624 13584 3652
rect 12900 3606 12952 3612
rect 12438 3567 12494 3576
rect 12256 3528 12308 3534
rect 12532 3528 12584 3534
rect 12308 3488 12388 3516
rect 12256 3470 12308 3476
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12084 3148 12204 3176
rect 12070 3088 12126 3097
rect 12070 3023 12072 3032
rect 12124 3023 12126 3032
rect 12072 2994 12124 3000
rect 12176 2922 12204 3148
rect 12164 2916 12216 2922
rect 12164 2858 12216 2864
rect 12268 2825 12296 3334
rect 12254 2816 12310 2825
rect 12254 2751 12310 2760
rect 12360 2530 12388 3488
rect 12452 3488 12532 3516
rect 12452 3369 12480 3488
rect 12532 3470 12584 3476
rect 12636 3482 12664 3590
rect 12716 3596 12848 3602
rect 12768 3590 12848 3596
rect 12716 3538 12768 3544
rect 12636 3454 13492 3482
rect 12624 3392 12676 3398
rect 12438 3360 12494 3369
rect 12808 3392 12860 3398
rect 12624 3334 12676 3340
rect 12714 3360 12770 3369
rect 12438 3295 12494 3304
rect 12440 3052 12492 3058
rect 12440 2994 12492 3000
rect 12452 2825 12480 2994
rect 12438 2816 12494 2825
rect 12438 2751 12494 2760
rect 12636 2530 12664 3334
rect 12992 3392 13044 3398
rect 12808 3334 12860 3340
rect 12912 3352 12992 3380
rect 12714 3295 12770 3304
rect 12728 3194 12756 3295
rect 12820 3194 12848 3334
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12820 2961 12848 2994
rect 12806 2952 12862 2961
rect 12806 2887 12862 2896
rect 12912 2836 12940 3352
rect 12992 3334 13044 3340
rect 13358 3392 13410 3398
rect 13358 3334 13410 3340
rect 12990 3224 13046 3233
rect 13046 3182 13308 3210
rect 13372 3194 13400 3334
rect 12990 3159 13046 3168
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 13096 2938 13124 2994
rect 12992 2916 13044 2922
rect 13096 2910 13216 2938
rect 12992 2858 13044 2864
rect 12820 2808 12940 2836
rect 12714 2544 12770 2553
rect 12360 2502 12480 2530
rect 12636 2502 12714 2530
rect 12256 2440 12308 2446
rect 11992 2366 12204 2394
rect 12452 2417 12480 2502
rect 12714 2479 12770 2488
rect 12532 2440 12584 2446
rect 12256 2382 12308 2388
rect 12438 2408 12494 2417
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 11992 1873 12020 2246
rect 11794 1864 11850 1873
rect 11794 1799 11850 1808
rect 11978 1864 12034 1873
rect 11978 1799 12034 1808
rect 11888 1760 11940 1766
rect 11888 1702 11940 1708
rect 11796 1420 11848 1426
rect 11794 1408 11796 1417
rect 11848 1408 11850 1417
rect 11612 1348 11664 1354
rect 11704 1352 11756 1358
rect 11520 1294 11572 1300
rect 11794 1343 11850 1352
rect 11704 1294 11756 1300
rect 11072 1278 11192 1294
rect 11900 1290 11928 1702
rect 11980 1488 12032 1494
rect 11980 1430 12032 1436
rect 11428 1284 11480 1290
rect 11428 1226 11480 1232
rect 11888 1284 11940 1290
rect 11888 1226 11940 1232
rect 10839 1116 11147 1125
rect 10839 1114 10845 1116
rect 10901 1114 10925 1116
rect 10981 1114 11005 1116
rect 11061 1114 11085 1116
rect 11141 1114 11147 1116
rect 10901 1062 10903 1114
rect 11083 1062 11085 1114
rect 10839 1060 10845 1062
rect 10901 1060 10925 1062
rect 10981 1060 11005 1062
rect 11061 1060 11085 1062
rect 11141 1060 11147 1062
rect 10839 1051 11147 1060
rect 11244 1012 11296 1018
rect 11244 954 11296 960
rect 11150 912 11206 921
rect 10968 876 11020 882
rect 11150 847 11206 856
rect 10968 818 11020 824
rect 10704 224 10824 252
rect 10690 82 10746 160
rect 10612 54 10746 82
rect 10796 82 10824 224
rect 10874 82 10930 160
rect 10980 134 11008 818
rect 11060 672 11112 678
rect 11060 614 11112 620
rect 11072 160 11100 614
rect 11164 542 11192 847
rect 11152 536 11204 542
rect 11152 478 11204 484
rect 11256 160 11284 954
rect 11440 160 11468 1226
rect 11520 1216 11572 1222
rect 11520 1158 11572 1164
rect 11704 1216 11756 1222
rect 11704 1158 11756 1164
rect 11532 1018 11560 1158
rect 11520 1012 11572 1018
rect 11520 954 11572 960
rect 11518 776 11574 785
rect 11518 711 11574 720
rect 11532 406 11560 711
rect 11520 400 11572 406
rect 11520 342 11572 348
rect 10796 54 10930 82
rect 10968 128 11020 134
rect 10968 70 11020 76
rect 10690 -300 10746 54
rect 10874 -300 10930 54
rect 11058 -300 11114 160
rect 11242 -300 11298 160
rect 11426 -300 11482 160
rect 11610 82 11666 160
rect 11716 82 11744 1158
rect 11796 1012 11848 1018
rect 11796 954 11848 960
rect 11808 160 11836 954
rect 11992 160 12020 1430
rect 12084 1057 12112 2246
rect 12176 1834 12204 2366
rect 12164 1828 12216 1834
rect 12164 1770 12216 1776
rect 12268 1426 12296 2382
rect 12532 2382 12584 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 12438 2343 12494 2352
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12452 1902 12480 2246
rect 12440 1896 12492 1902
rect 12440 1838 12492 1844
rect 12544 1766 12572 2382
rect 12636 2145 12664 2382
rect 12820 2281 12848 2808
rect 13004 2564 13032 2858
rect 13188 2854 13216 2910
rect 13280 2904 13308 3182
rect 13360 3188 13412 3194
rect 13464 3176 13492 3454
rect 13556 3380 13584 3624
rect 13872 3624 13952 3652
rect 13820 3606 13872 3612
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 13636 3392 13688 3398
rect 13556 3352 13636 3380
rect 13636 3334 13688 3340
rect 13832 3346 13860 3470
rect 13924 3448 13952 3624
rect 14016 3516 14044 3726
rect 14094 3703 14150 3712
rect 14738 3768 14794 3777
rect 14738 3703 14794 3712
rect 14108 3670 14136 3703
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 14016 3488 14688 3516
rect 13924 3420 14228 3448
rect 14200 3380 14228 3420
rect 14200 3352 14504 3380
rect 13832 3318 14026 3346
rect 13998 3210 14026 3318
rect 14186 3224 14242 3233
rect 13912 3188 13964 3194
rect 13464 3148 13912 3176
rect 13360 3130 13412 3136
rect 13998 3182 14044 3210
rect 13912 3130 13964 3136
rect 14016 2990 14044 3182
rect 14370 3224 14426 3233
rect 14186 3159 14242 3168
rect 14280 3188 14332 3194
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 14004 2984 14056 2990
rect 14004 2926 14056 2932
rect 14200 2938 14228 3159
rect 14476 3176 14504 3352
rect 14660 3194 14688 3488
rect 14752 3346 14780 3703
rect 14936 3670 14964 3896
rect 15028 3896 15200 3924
rect 14924 3664 14976 3670
rect 14924 3606 14976 3612
rect 14832 3596 14884 3602
rect 14832 3538 14884 3544
rect 14844 3466 14872 3538
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14752 3318 14964 3346
rect 14830 3224 14886 3233
rect 14370 3159 14372 3168
rect 14280 3130 14332 3136
rect 14424 3159 14426 3168
rect 14372 3130 14424 3136
rect 14458 3148 14504 3176
rect 14648 3188 14700 3194
rect 14300 3040 14328 3130
rect 14363 3052 14415 3058
rect 14300 3012 14363 3040
rect 14458 3040 14486 3148
rect 14830 3159 14886 3168
rect 14648 3130 14700 3136
rect 14844 3126 14872 3159
rect 14832 3120 14884 3126
rect 14832 3062 14884 3068
rect 14648 3052 14700 3058
rect 14458 3012 14648 3040
rect 14363 2994 14415 3000
rect 14648 2994 14700 3000
rect 14936 2990 14964 3318
rect 14924 2984 14976 2990
rect 13360 2916 13412 2922
rect 13280 2876 13360 2904
rect 13360 2858 13412 2864
rect 13176 2848 13228 2854
rect 13740 2825 13768 2926
rect 14200 2910 14412 2938
rect 14924 2926 14976 2932
rect 13820 2848 13872 2854
rect 13176 2790 13228 2796
rect 13726 2816 13782 2825
rect 13820 2790 13872 2796
rect 13912 2848 13964 2854
rect 14280 2848 14332 2854
rect 13912 2790 13964 2796
rect 14200 2808 14280 2836
rect 13312 2748 13620 2757
rect 13726 2751 13782 2760
rect 13312 2746 13318 2748
rect 13374 2746 13398 2748
rect 13454 2746 13478 2748
rect 13534 2746 13558 2748
rect 13614 2746 13620 2748
rect 13374 2694 13376 2746
rect 13556 2694 13558 2746
rect 13312 2692 13318 2694
rect 13374 2692 13398 2694
rect 13454 2692 13478 2694
rect 13534 2692 13558 2694
rect 13614 2692 13620 2694
rect 13312 2683 13620 2692
rect 13832 2689 13860 2790
rect 13818 2680 13874 2689
rect 13924 2666 13952 2790
rect 14002 2680 14058 2689
rect 13924 2638 14002 2666
rect 13818 2615 13874 2624
rect 14002 2615 14058 2624
rect 13004 2536 13492 2564
rect 13464 2462 13492 2536
rect 13726 2544 13782 2553
rect 14002 2544 14058 2553
rect 13912 2508 13964 2514
rect 13726 2479 13782 2488
rect 12900 2440 12952 2446
rect 13360 2440 13412 2446
rect 12900 2382 12952 2388
rect 12990 2408 13046 2417
rect 12806 2272 12862 2281
rect 12806 2207 12862 2216
rect 12912 2145 12940 2382
rect 13464 2434 13584 2462
rect 13556 2428 13584 2434
rect 13636 2440 13688 2446
rect 13556 2400 13636 2428
rect 13360 2382 13412 2388
rect 13636 2382 13688 2388
rect 12990 2343 13046 2352
rect 13004 2310 13032 2343
rect 12992 2304 13044 2310
rect 13372 2281 13400 2382
rect 13740 2310 13768 2479
rect 13832 2468 13912 2496
rect 13728 2304 13780 2310
rect 12992 2246 13044 2252
rect 13358 2272 13414 2281
rect 13728 2246 13780 2252
rect 13358 2207 13414 2216
rect 12622 2136 12678 2145
rect 12622 2071 12678 2080
rect 12898 2136 12954 2145
rect 13832 2122 13860 2468
rect 14200 2530 14228 2808
rect 14384 2825 14412 2910
rect 14280 2790 14332 2796
rect 14370 2816 14426 2825
rect 14660 2808 14918 2836
rect 14660 2802 14688 2808
rect 14370 2751 14426 2760
rect 14476 2774 14688 2802
rect 14890 2802 14918 2808
rect 14890 2774 14964 2802
rect 14372 2576 14424 2582
rect 14002 2479 14058 2488
rect 14108 2502 14228 2530
rect 14292 2536 14372 2564
rect 13912 2450 13964 2456
rect 12898 2071 12954 2080
rect 13464 2094 13860 2122
rect 12624 1964 12676 1970
rect 12676 1924 12756 1952
rect 12624 1906 12676 1912
rect 12532 1760 12584 1766
rect 12532 1702 12584 1708
rect 12622 1728 12678 1737
rect 12622 1663 12678 1672
rect 12440 1556 12492 1562
rect 12360 1516 12440 1544
rect 12256 1420 12308 1426
rect 12256 1362 12308 1368
rect 12256 1284 12308 1290
rect 12256 1226 12308 1232
rect 12164 1216 12216 1222
rect 12164 1158 12216 1164
rect 12070 1048 12126 1057
rect 12070 983 12126 992
rect 12176 160 12204 1158
rect 12268 610 12296 1226
rect 12256 604 12308 610
rect 12256 546 12308 552
rect 12360 160 12388 1516
rect 12440 1498 12492 1504
rect 12636 1494 12664 1663
rect 12624 1488 12676 1494
rect 12624 1430 12676 1436
rect 12728 1358 12756 1924
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 12808 1828 12860 1834
rect 12808 1770 12860 1776
rect 12820 1737 12848 1770
rect 12806 1728 12862 1737
rect 12806 1663 12862 1672
rect 12912 1394 12940 1838
rect 12992 1760 13044 1766
rect 12992 1702 13044 1708
rect 13084 1760 13136 1766
rect 13464 1748 13492 2094
rect 14016 2088 14044 2479
rect 13924 2060 14044 2088
rect 13544 2032 13596 2038
rect 13596 1992 13768 2020
rect 13544 1974 13596 1980
rect 13740 1952 13768 1992
rect 13924 1952 13952 2060
rect 14108 1986 14136 2502
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 13740 1924 13952 1952
rect 14016 1958 14136 1986
rect 13636 1828 13688 1834
rect 13636 1770 13688 1776
rect 13084 1702 13136 1708
rect 13188 1720 13492 1748
rect 12820 1366 12940 1394
rect 12716 1352 12768 1358
rect 12716 1294 12768 1300
rect 12440 1284 12492 1290
rect 12440 1226 12492 1232
rect 12452 338 12480 1226
rect 12716 1216 12768 1222
rect 12530 1184 12586 1193
rect 12530 1119 12586 1128
rect 12636 1164 12716 1170
rect 12636 1158 12768 1164
rect 12636 1142 12756 1158
rect 12544 746 12572 1119
rect 12532 740 12584 746
rect 12532 682 12584 688
rect 12440 332 12492 338
rect 12440 274 12492 280
rect 11610 54 11744 82
rect 11610 -300 11666 54
rect 11794 -300 11850 160
rect 11978 -300 12034 160
rect 12162 -300 12218 160
rect 12346 -300 12402 160
rect 12530 82 12586 160
rect 12636 82 12664 1142
rect 12530 54 12664 82
rect 12714 82 12770 160
rect 12820 82 12848 1366
rect 12900 1284 12952 1290
rect 12900 1226 12952 1232
rect 12912 649 12940 1226
rect 12898 640 12954 649
rect 12898 575 12954 584
rect 12714 54 12848 82
rect 12898 82 12954 160
rect 13004 82 13032 1702
rect 13096 160 13124 1702
rect 12898 54 13032 82
rect 12530 -300 12586 54
rect 12714 -300 12770 54
rect 12898 -300 12954 54
rect 13082 -300 13138 160
rect 13188 82 13216 1720
rect 13312 1660 13620 1669
rect 13312 1658 13318 1660
rect 13374 1658 13398 1660
rect 13454 1658 13478 1660
rect 13534 1658 13558 1660
rect 13614 1658 13620 1660
rect 13374 1606 13376 1658
rect 13556 1606 13558 1658
rect 13312 1604 13318 1606
rect 13374 1604 13398 1606
rect 13454 1604 13478 1606
rect 13534 1604 13558 1606
rect 13614 1604 13620 1606
rect 13312 1595 13620 1604
rect 13648 1494 13676 1770
rect 13728 1760 13780 1766
rect 13728 1702 13780 1708
rect 13360 1488 13412 1494
rect 13360 1430 13412 1436
rect 13636 1488 13688 1494
rect 13636 1430 13688 1436
rect 13268 1420 13320 1426
rect 13268 1362 13320 1368
rect 13280 882 13308 1362
rect 13372 1329 13400 1430
rect 13740 1394 13768 1702
rect 13648 1366 13768 1394
rect 13544 1352 13596 1358
rect 13358 1320 13414 1329
rect 13358 1255 13414 1264
rect 13542 1320 13544 1329
rect 13596 1320 13598 1329
rect 13542 1255 13598 1264
rect 13268 876 13320 882
rect 13268 818 13320 824
rect 13544 808 13596 814
rect 13358 776 13414 785
rect 13358 711 13414 720
rect 13542 776 13544 785
rect 13596 776 13598 785
rect 13542 711 13598 720
rect 13268 672 13320 678
rect 13266 640 13268 649
rect 13320 640 13322 649
rect 13266 575 13322 584
rect 13372 270 13400 711
rect 13360 264 13412 270
rect 13648 218 13676 1366
rect 14016 1306 14044 1958
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 14108 1494 14136 1838
rect 14200 1766 14228 2382
rect 14292 2038 14320 2536
rect 14372 2518 14424 2524
rect 14372 2372 14424 2378
rect 14372 2314 14424 2320
rect 14384 2038 14412 2314
rect 14476 2310 14504 2774
rect 14568 2638 14780 2666
rect 14464 2304 14516 2310
rect 14464 2246 14516 2252
rect 14464 2100 14516 2106
rect 14464 2042 14516 2048
rect 14280 2032 14332 2038
rect 14280 1974 14332 1980
rect 14372 2032 14424 2038
rect 14372 1974 14424 1980
rect 14280 1896 14332 1902
rect 14280 1838 14332 1844
rect 14188 1760 14240 1766
rect 14188 1702 14240 1708
rect 14186 1592 14242 1601
rect 14292 1544 14320 1838
rect 14476 1834 14504 2042
rect 14568 2009 14596 2638
rect 14648 2576 14700 2582
rect 14648 2518 14700 2524
rect 14554 2000 14610 2009
rect 14554 1935 14610 1944
rect 14660 1952 14688 2518
rect 14752 2428 14780 2638
rect 14832 2440 14884 2446
rect 14752 2400 14832 2428
rect 14832 2382 14884 2388
rect 14936 2310 14964 2774
rect 15028 2530 15056 3896
rect 15200 3878 15252 3884
rect 15304 3754 15332 3998
rect 15488 3992 15516 4270
rect 15844 4276 15896 4282
rect 15764 4236 15844 4264
rect 15660 4208 15712 4214
rect 15660 4150 15712 4156
rect 15672 4078 15700 4150
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15488 3964 15608 3992
rect 15580 3890 15608 3964
rect 15764 3913 15792 4236
rect 15844 4218 15896 4224
rect 16132 4146 16160 4440
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 16028 4072 16080 4078
rect 16028 4014 16080 4020
rect 15750 3904 15806 3913
rect 15580 3862 15700 3890
rect 15304 3726 15608 3754
rect 15384 3664 15436 3670
rect 15106 3632 15162 3641
rect 15436 3624 15516 3652
rect 15384 3606 15436 3612
rect 15106 3567 15162 3576
rect 15200 3596 15252 3602
rect 15120 3369 15148 3567
rect 15200 3538 15252 3544
rect 15106 3360 15162 3369
rect 15106 3295 15162 3304
rect 15106 3224 15162 3233
rect 15212 3194 15240 3538
rect 15384 3392 15436 3398
rect 15304 3352 15384 3380
rect 15106 3159 15162 3168
rect 15200 3188 15252 3194
rect 15120 3126 15148 3159
rect 15200 3130 15252 3136
rect 15108 3120 15160 3126
rect 15108 3062 15160 3068
rect 15304 2990 15332 3352
rect 15488 3369 15516 3624
rect 15580 3516 15608 3726
rect 15672 3618 15700 3862
rect 15750 3839 15806 3848
rect 15672 3590 15792 3618
rect 15660 3528 15712 3534
rect 15580 3488 15660 3516
rect 15384 3334 15436 3340
rect 15474 3360 15530 3369
rect 15474 3295 15530 3304
rect 15474 3224 15530 3233
rect 15474 3159 15530 3168
rect 15488 3126 15516 3159
rect 15476 3120 15528 3126
rect 15476 3062 15528 3068
rect 15292 2984 15344 2990
rect 15580 2972 15608 3488
rect 15660 3470 15712 3476
rect 15764 3380 15792 3590
rect 15844 3528 15896 3534
rect 15842 3496 15844 3505
rect 16040 3505 16068 4014
rect 16224 3670 16252 4508
rect 16302 4448 16358 4457
rect 16302 4383 16358 4392
rect 16212 3664 16264 3670
rect 16212 3606 16264 3612
rect 16316 3534 16344 4383
rect 16408 4282 16436 5324
rect 16486 5264 16542 5273
rect 16486 5199 16488 5208
rect 16540 5199 16542 5208
rect 16488 5170 16540 5176
rect 16488 5024 16540 5030
rect 16488 4966 16540 4972
rect 16500 4486 16528 4966
rect 16592 4622 16620 6054
rect 16670 5808 16726 5817
rect 16776 5794 16804 6122
rect 16854 5808 16910 5817
rect 16776 5766 16854 5794
rect 16670 5743 16726 5752
rect 16854 5743 16910 5752
rect 16684 5642 16712 5743
rect 16672 5636 16724 5642
rect 16672 5578 16724 5584
rect 16960 5574 16988 6310
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16948 5568 17000 5574
rect 16948 5510 17000 5516
rect 16764 5296 16816 5302
rect 16868 5273 16896 5510
rect 16764 5238 16816 5244
rect 16854 5264 16910 5273
rect 16776 5030 16804 5238
rect 16854 5199 16910 5208
rect 16764 5024 16816 5030
rect 16764 4966 16816 4972
rect 16854 4720 16910 4729
rect 16672 4684 16724 4690
rect 16960 4690 16988 5510
rect 17052 5409 17080 6412
rect 17144 6322 17172 7239
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 17132 5840 17184 5846
rect 17184 5800 17264 5828
rect 17132 5782 17184 5788
rect 17038 5400 17094 5409
rect 17038 5335 17094 5344
rect 17040 5228 17092 5234
rect 17040 5170 17092 5176
rect 17052 5001 17080 5170
rect 17038 4992 17094 5001
rect 17038 4927 17094 4936
rect 16854 4655 16910 4664
rect 16948 4684 17000 4690
rect 16672 4626 16724 4632
rect 16580 4616 16632 4622
rect 16580 4558 16632 4564
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16396 4276 16448 4282
rect 16396 4218 16448 4224
rect 16486 4176 16542 4185
rect 16396 4140 16448 4146
rect 16486 4111 16542 4120
rect 16396 4082 16448 4088
rect 16304 3528 16356 3534
rect 15896 3496 15898 3505
rect 15842 3431 15898 3440
rect 16026 3496 16082 3505
rect 16304 3470 16356 3476
rect 16026 3431 16082 3440
rect 16408 3448 16436 4082
rect 16500 3913 16528 4111
rect 16486 3904 16542 3913
rect 16486 3839 16542 3848
rect 16408 3420 16528 3448
rect 15672 3352 15792 3380
rect 16120 3392 16172 3398
rect 15672 3233 15700 3352
rect 16120 3334 16172 3340
rect 16394 3360 16450 3369
rect 15784 3292 16092 3301
rect 15784 3290 15790 3292
rect 15846 3290 15870 3292
rect 15926 3290 15950 3292
rect 16006 3290 16030 3292
rect 16086 3290 16092 3292
rect 15846 3238 15848 3290
rect 16028 3238 16030 3290
rect 15784 3236 15790 3238
rect 15846 3236 15870 3238
rect 15926 3236 15950 3238
rect 16006 3236 16030 3238
rect 16086 3236 16092 3238
rect 15658 3224 15714 3233
rect 15784 3227 16092 3236
rect 15658 3159 15714 3168
rect 16132 3074 16160 3334
rect 16394 3295 16450 3304
rect 16304 3120 16356 3126
rect 15292 2926 15344 2932
rect 15396 2944 15608 2972
rect 15672 3046 16160 3074
rect 16302 3088 16304 3097
rect 16356 3088 16358 3097
rect 15292 2848 15344 2854
rect 15212 2808 15292 2836
rect 15028 2502 15148 2530
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14924 2304 14976 2310
rect 14924 2246 14976 2252
rect 14752 2122 14780 2246
rect 14752 2094 15056 2122
rect 14924 2032 14976 2038
rect 14922 2000 14924 2009
rect 14976 2000 14978 2009
rect 14660 1924 14872 1952
rect 14922 1935 14978 1944
rect 14464 1828 14516 1834
rect 14740 1828 14792 1834
rect 14464 1770 14516 1776
rect 14568 1788 14740 1816
rect 14242 1536 14320 1544
rect 14186 1527 14320 1536
rect 14200 1516 14320 1527
rect 14096 1488 14148 1494
rect 14096 1430 14148 1436
rect 14188 1420 14240 1426
rect 14568 1408 14596 1788
rect 14740 1770 14792 1776
rect 14648 1556 14700 1562
rect 14648 1498 14700 1504
rect 14188 1362 14240 1368
rect 14476 1380 14596 1408
rect 13820 1284 13872 1290
rect 14016 1278 14136 1306
rect 13820 1226 13872 1232
rect 13832 864 13860 1226
rect 14004 1012 14056 1018
rect 14004 954 14056 960
rect 13912 876 13964 882
rect 13832 836 13912 864
rect 13912 818 13964 824
rect 13912 740 13964 746
rect 13912 682 13964 688
rect 13728 604 13780 610
rect 13924 592 13952 682
rect 14016 660 14044 954
rect 13780 564 13952 592
rect 13985 632 14044 660
rect 13728 546 13780 552
rect 13985 524 14013 632
rect 13924 496 14013 524
rect 13924 456 13952 496
rect 14108 456 14136 1278
rect 14200 796 14228 1362
rect 14476 1018 14504 1380
rect 14660 1306 14688 1498
rect 14566 1278 14688 1306
rect 14738 1320 14794 1329
rect 14566 1204 14594 1278
rect 14732 1264 14738 1272
rect 14732 1255 14794 1264
rect 14732 1244 14780 1255
rect 14732 1204 14760 1244
rect 14566 1176 14596 1204
rect 14568 1018 14596 1176
rect 14660 1176 14760 1204
rect 14464 1012 14516 1018
rect 14464 954 14516 960
rect 14556 1012 14608 1018
rect 14556 954 14608 960
rect 14200 768 14596 796
rect 14280 672 14332 678
rect 14280 614 14332 620
rect 14292 474 14320 614
rect 13924 428 13960 456
rect 13728 332 13780 338
rect 13728 274 13780 280
rect 13360 206 13412 212
rect 13556 190 13676 218
rect 13266 82 13322 160
rect 13188 54 13322 82
rect 13266 -300 13322 54
rect 13450 82 13506 160
rect 13556 82 13584 190
rect 13450 54 13584 82
rect 13634 82 13690 160
rect 13740 82 13768 274
rect 13932 252 13960 428
rect 13832 224 13960 252
rect 14016 428 14136 456
rect 14280 468 14332 474
rect 13832 160 13860 224
rect 14016 160 14044 428
rect 14280 410 14332 416
rect 14372 468 14424 474
rect 14372 410 14424 416
rect 14188 400 14240 406
rect 14188 342 14240 348
rect 14200 160 14228 342
rect 14384 160 14412 410
rect 14568 160 14596 768
rect 14660 377 14688 1176
rect 14844 1018 14872 1924
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 14832 1012 14884 1018
rect 14832 954 14884 960
rect 14740 808 14792 814
rect 14936 796 14964 1838
rect 15028 1562 15056 2094
rect 15016 1556 15068 1562
rect 15016 1498 15068 1504
rect 15016 1420 15068 1426
rect 15016 1362 15068 1368
rect 15028 1222 15056 1362
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 15016 1012 15068 1018
rect 15016 954 15068 960
rect 15028 796 15056 954
rect 14792 768 14964 796
rect 14994 768 15056 796
rect 14740 750 14792 756
rect 14994 728 15022 768
rect 15120 728 15148 2502
rect 14844 700 15022 728
rect 15053 700 15148 728
rect 14844 474 14872 700
rect 15053 626 15081 700
rect 15212 660 15240 2808
rect 15396 2825 15424 2944
rect 15476 2848 15528 2854
rect 15292 2790 15344 2796
rect 15382 2816 15438 2825
rect 15476 2790 15528 2796
rect 15382 2751 15438 2760
rect 15292 2100 15344 2106
rect 15292 2042 15344 2048
rect 15304 1902 15332 2042
rect 15292 1896 15344 1902
rect 15292 1838 15344 1844
rect 15488 1714 15516 2790
rect 15672 2496 15700 3046
rect 16302 3023 16358 3032
rect 15844 2984 15896 2990
rect 15844 2926 15896 2932
rect 15583 2468 15700 2496
rect 15583 2394 15611 2468
rect 15028 598 15081 626
rect 15120 632 15240 660
rect 15304 1686 15516 1714
rect 15580 2366 15611 2394
rect 15856 2378 15884 2926
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 15948 2378 15976 2858
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15660 2372 15712 2378
rect 14832 468 14884 474
rect 14832 410 14884 416
rect 14924 468 14976 474
rect 14924 410 14976 416
rect 14646 368 14702 377
rect 14936 354 14964 410
rect 14646 303 14702 312
rect 14752 326 14964 354
rect 14752 160 14780 326
rect 15028 252 15056 598
rect 15120 474 15148 632
rect 15304 592 15332 1686
rect 15384 1556 15436 1562
rect 15384 1498 15436 1504
rect 15476 1556 15528 1562
rect 15476 1498 15528 1504
rect 15396 746 15424 1498
rect 15384 740 15436 746
rect 15384 682 15436 688
rect 15212 564 15332 592
rect 15108 468 15160 474
rect 15108 410 15160 416
rect 15212 354 15240 564
rect 15292 468 15344 474
rect 15292 410 15344 416
rect 15304 377 15332 410
rect 15488 388 15516 1498
rect 14936 224 15056 252
rect 15120 326 15240 354
rect 15290 368 15346 377
rect 14936 160 14964 224
rect 15120 160 15148 326
rect 15290 303 15346 312
rect 15396 360 15516 388
rect 15396 184 15424 360
rect 15580 320 15608 2366
rect 15660 2314 15712 2320
rect 15844 2372 15896 2378
rect 15844 2314 15896 2320
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15304 160 15424 184
rect 15488 292 15608 320
rect 15488 160 15516 292
rect 15672 160 15700 2314
rect 15784 2204 16092 2213
rect 15784 2202 15790 2204
rect 15846 2202 15870 2204
rect 15926 2202 15950 2204
rect 16006 2202 16030 2204
rect 16086 2202 16092 2204
rect 15846 2150 15848 2202
rect 16028 2150 16030 2202
rect 15784 2148 15790 2150
rect 15846 2148 15870 2150
rect 15926 2148 15950 2150
rect 16006 2148 16030 2150
rect 16086 2148 16092 2150
rect 15784 2139 16092 2148
rect 16028 1896 16080 1902
rect 16132 1884 16160 2790
rect 16408 2650 16436 3295
rect 16500 3233 16528 3420
rect 16684 3233 16712 4626
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 16776 3777 16804 4422
rect 16868 4214 16896 4655
rect 16948 4626 17000 4632
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 16856 4208 16908 4214
rect 16856 4150 16908 4156
rect 16946 4040 17002 4049
rect 16946 3975 17002 3984
rect 16960 3942 16988 3975
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 16762 3768 16818 3777
rect 16762 3703 16818 3712
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16762 3360 16818 3369
rect 16762 3295 16818 3304
rect 16486 3224 16542 3233
rect 16486 3159 16542 3168
rect 16670 3224 16726 3233
rect 16776 3194 16804 3295
rect 16670 3159 16726 3168
rect 16764 3188 16816 3194
rect 16488 3052 16540 3058
rect 16488 2994 16540 3000
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16500 2836 16528 2994
rect 16592 2961 16620 2994
rect 16684 2990 16712 3159
rect 16764 3130 16816 3136
rect 16672 2984 16724 2990
rect 16578 2952 16634 2961
rect 16672 2926 16724 2932
rect 16578 2887 16634 2896
rect 16868 2854 16896 3402
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16856 2848 16908 2854
rect 16500 2808 16620 2836
rect 16592 2802 16620 2808
rect 16592 2774 16804 2802
rect 16856 2790 16908 2796
rect 16396 2644 16448 2650
rect 16396 2586 16448 2592
rect 16580 2644 16632 2650
rect 16580 2586 16632 2592
rect 16488 2576 16540 2582
rect 16486 2544 16488 2553
rect 16540 2544 16542 2553
rect 16486 2479 16542 2488
rect 16488 2440 16540 2446
rect 16486 2408 16488 2417
rect 16540 2408 16542 2417
rect 16486 2343 16542 2352
rect 16488 2304 16540 2310
rect 16210 2272 16266 2281
rect 16488 2246 16540 2252
rect 16210 2207 16266 2216
rect 16224 2106 16252 2207
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16396 2100 16448 2106
rect 16396 2042 16448 2048
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16080 1856 16160 1884
rect 16028 1838 16080 1844
rect 15934 1456 15990 1465
rect 16316 1442 16344 1906
rect 16408 1766 16436 2042
rect 16500 1850 16528 2246
rect 16592 2106 16620 2586
rect 16672 2440 16724 2446
rect 16776 2417 16804 2774
rect 16672 2382 16724 2388
rect 16762 2408 16818 2417
rect 16580 2100 16632 2106
rect 16580 2042 16632 2048
rect 16500 1822 16620 1850
rect 16396 1760 16448 1766
rect 16396 1702 16448 1708
rect 16488 1760 16540 1766
rect 16488 1702 16540 1708
rect 16500 1494 16528 1702
rect 16592 1562 16620 1822
rect 16580 1556 16632 1562
rect 16580 1498 16632 1504
rect 16488 1488 16540 1494
rect 15990 1414 16252 1442
rect 16316 1414 16436 1442
rect 16488 1430 16540 1436
rect 15934 1391 15990 1400
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 15784 1116 16092 1125
rect 15784 1114 15790 1116
rect 15846 1114 15870 1116
rect 15926 1114 15950 1116
rect 16006 1114 16030 1116
rect 16086 1114 16092 1116
rect 15846 1062 15848 1114
rect 16028 1062 16030 1114
rect 15784 1060 15790 1062
rect 15846 1060 15870 1062
rect 15926 1060 15950 1062
rect 16006 1060 16030 1062
rect 16086 1060 16092 1062
rect 15784 1051 16092 1060
rect 15752 876 15804 882
rect 15752 818 15804 824
rect 15844 876 15896 882
rect 15844 818 15896 824
rect 15764 377 15792 818
rect 15856 746 15884 818
rect 15844 740 15896 746
rect 15844 682 15896 688
rect 16028 740 16080 746
rect 16028 682 16080 688
rect 16040 490 16068 682
rect 15948 462 16068 490
rect 15750 368 15806 377
rect 15750 303 15806 312
rect 13634 54 13768 82
rect 13450 -300 13506 54
rect 13634 -300 13690 54
rect 13818 -300 13874 160
rect 14002 -300 14058 160
rect 14186 -300 14242 160
rect 14370 -300 14426 160
rect 14554 -300 14610 160
rect 14738 -300 14794 160
rect 14922 -300 14978 160
rect 15106 -300 15162 160
rect 15290 156 15424 160
rect 15290 -300 15346 156
rect 15474 -300 15530 160
rect 15658 -300 15714 160
rect 15842 82 15898 160
rect 15948 82 15976 462
rect 16132 388 16160 1294
rect 16224 1057 16252 1414
rect 16304 1352 16356 1358
rect 16302 1320 16304 1329
rect 16356 1320 16358 1329
rect 16302 1255 16358 1264
rect 16304 1216 16356 1222
rect 16302 1184 16304 1193
rect 16356 1184 16358 1193
rect 16302 1119 16358 1128
rect 16210 1048 16266 1057
rect 16210 983 16266 992
rect 16408 932 16436 1414
rect 16580 1352 16632 1358
rect 16580 1294 16632 1300
rect 16488 1216 16540 1222
rect 16488 1158 16540 1164
rect 16040 360 16160 388
rect 16224 904 16436 932
rect 16040 160 16068 360
rect 16224 160 16252 904
rect 16500 728 16528 1158
rect 16592 746 16620 1294
rect 16408 700 16528 728
rect 16580 740 16632 746
rect 16408 160 16436 700
rect 16580 682 16632 688
rect 15842 54 15976 82
rect 15842 -300 15898 54
rect 16026 -300 16082 160
rect 16210 -300 16266 160
rect 16394 -300 16450 160
rect 16578 82 16634 160
rect 16684 82 16712 2382
rect 16762 2343 16818 2352
rect 16960 2281 16988 3130
rect 17052 2310 17080 4422
rect 17040 2304 17092 2310
rect 16946 2272 17002 2281
rect 17040 2246 17092 2252
rect 16946 2207 17002 2216
rect 17040 1964 17092 1970
rect 17040 1906 17092 1912
rect 16946 1592 17002 1601
rect 16946 1527 17002 1536
rect 16856 1488 16908 1494
rect 16856 1430 16908 1436
rect 16762 776 16818 785
rect 16762 711 16764 720
rect 16816 711 16818 720
rect 16764 682 16816 688
rect 16578 54 16712 82
rect 16762 82 16818 160
rect 16868 82 16896 1430
rect 16960 1426 16988 1527
rect 16948 1420 17000 1426
rect 16948 1362 17000 1368
rect 16762 54 16896 82
rect 16946 82 17002 160
rect 17052 82 17080 1906
rect 17144 1494 17172 4490
rect 17236 4486 17264 5800
rect 17328 4758 17356 8055
rect 17316 4752 17368 4758
rect 17316 4694 17368 4700
rect 17224 4480 17276 4486
rect 17224 4422 17276 4428
rect 17224 4276 17276 4282
rect 17224 4218 17276 4224
rect 17236 3670 17264 4218
rect 17420 4146 17448 8230
rect 17512 5234 17540 8452
rect 17604 7954 17632 8502
rect 17696 8294 17724 9880
rect 17868 9648 17920 9654
rect 17868 9590 17920 9596
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17788 8498 17816 8842
rect 17880 8566 17908 9590
rect 17972 8974 18000 11319
rect 18052 11290 18104 11296
rect 18156 10062 18184 11494
rect 18257 11452 18565 11461
rect 18257 11450 18263 11452
rect 18319 11450 18343 11452
rect 18399 11450 18423 11452
rect 18479 11450 18503 11452
rect 18559 11450 18565 11452
rect 18319 11398 18321 11450
rect 18501 11398 18503 11450
rect 18257 11396 18263 11398
rect 18319 11396 18343 11398
rect 18399 11396 18423 11398
rect 18479 11396 18503 11398
rect 18559 11396 18565 11398
rect 18257 11387 18565 11396
rect 18708 11354 18736 13790
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18800 11898 18828 12786
rect 18892 12102 18920 15320
rect 18984 14482 19012 16000
rect 19352 15570 19380 19246
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19248 15496 19300 15502
rect 19248 15438 19300 15444
rect 19076 14822 19104 15438
rect 19156 15428 19208 15434
rect 19156 15370 19208 15376
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18972 14476 19024 14482
rect 18972 14418 19024 14424
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18984 13530 19012 13874
rect 19064 13796 19116 13802
rect 19064 13738 19116 13744
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 19076 12900 19104 13738
rect 18984 12872 19104 12900
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18984 11778 19012 12872
rect 19062 12608 19118 12617
rect 19062 12543 19118 12552
rect 19076 12442 19104 12543
rect 19064 12436 19116 12442
rect 19064 12378 19116 12384
rect 19168 12374 19196 15370
rect 19260 14618 19288 15438
rect 19340 15360 19392 15366
rect 19340 15302 19392 15308
rect 19248 14612 19300 14618
rect 19248 14554 19300 14560
rect 19248 14476 19300 14482
rect 19248 14418 19300 14424
rect 19260 13394 19288 14418
rect 19352 13802 19380 15302
rect 19444 15094 19472 20318
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19628 19666 19656 21678
rect 19720 21146 19748 21814
rect 19708 21140 19760 21146
rect 19708 21082 19760 21088
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 19720 20398 19748 20742
rect 19708 20392 19760 20398
rect 19708 20334 19760 20340
rect 19536 16017 19564 19654
rect 19628 19638 19748 19666
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19628 18426 19656 19314
rect 19616 18420 19668 18426
rect 19616 18362 19668 18368
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19628 17270 19656 17614
rect 19720 17338 19748 19638
rect 19708 17332 19760 17338
rect 19708 17274 19760 17280
rect 19616 17264 19668 17270
rect 19616 17206 19668 17212
rect 19812 17105 19840 24398
rect 19904 23322 19932 24534
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19904 22778 19932 23122
rect 19996 22930 20024 27066
rect 20088 26518 20116 28358
rect 20272 26874 20300 30110
rect 20352 30048 20404 30054
rect 20444 30048 20496 30054
rect 20352 29990 20404 29996
rect 20442 30016 20444 30025
rect 20496 30016 20498 30025
rect 20180 26846 20300 26874
rect 20076 26512 20128 26518
rect 20076 26454 20128 26460
rect 20076 26240 20128 26246
rect 20076 26182 20128 26188
rect 20088 23594 20116 26182
rect 20076 23588 20128 23594
rect 20076 23530 20128 23536
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 20088 23050 20116 23258
rect 20076 23044 20128 23050
rect 20076 22986 20128 22992
rect 19996 22902 20116 22930
rect 19892 22772 19944 22778
rect 19892 22714 19944 22720
rect 20088 22094 20116 22902
rect 19996 22066 20116 22094
rect 19892 21344 19944 21350
rect 19890 21312 19892 21321
rect 19944 21312 19946 21321
rect 19890 21247 19946 21256
rect 19892 21072 19944 21078
rect 19892 21014 19944 21020
rect 19798 17096 19854 17105
rect 19798 17031 19854 17040
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19616 16720 19668 16726
rect 19616 16662 19668 16668
rect 19522 16008 19578 16017
rect 19522 15943 19578 15952
rect 19628 15706 19656 16662
rect 19708 16584 19760 16590
rect 19708 16526 19760 16532
rect 19720 16250 19748 16526
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 19720 15706 19748 16186
rect 19812 15706 19840 16934
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19708 15700 19760 15706
rect 19708 15642 19760 15648
rect 19800 15700 19852 15706
rect 19800 15642 19852 15648
rect 19524 15632 19576 15638
rect 19524 15574 19576 15580
rect 19432 15088 19484 15094
rect 19432 15030 19484 15036
rect 19536 14906 19564 15574
rect 19536 14878 19840 14906
rect 19708 14816 19760 14822
rect 19708 14758 19760 14764
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19616 14272 19668 14278
rect 19616 14214 19668 14220
rect 19340 13796 19392 13802
rect 19340 13738 19392 13744
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19260 12374 19288 13330
rect 19444 12918 19472 14214
rect 19524 13864 19576 13870
rect 19524 13806 19576 13812
rect 19536 13705 19564 13806
rect 19522 13696 19578 13705
rect 19522 13631 19578 13640
rect 19432 12912 19484 12918
rect 19432 12854 19484 12860
rect 19524 12708 19576 12714
rect 19524 12650 19576 12656
rect 19340 12640 19392 12646
rect 19340 12582 19392 12588
rect 19352 12434 19380 12582
rect 19352 12406 19472 12434
rect 19156 12368 19208 12374
rect 19156 12310 19208 12316
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 19338 12200 19394 12209
rect 19338 12135 19394 12144
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 18892 11750 19012 11778
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 18800 11082 18828 11222
rect 18892 11150 18920 11750
rect 18970 11248 19026 11257
rect 18970 11183 19026 11192
rect 19156 11212 19208 11218
rect 18880 11144 18932 11150
rect 18880 11086 18932 11092
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 18788 11076 18840 11082
rect 18788 11018 18840 11024
rect 18257 10364 18565 10373
rect 18257 10362 18263 10364
rect 18319 10362 18343 10364
rect 18399 10362 18423 10364
rect 18479 10362 18503 10364
rect 18559 10362 18565 10364
rect 18319 10310 18321 10362
rect 18501 10310 18503 10362
rect 18257 10308 18263 10310
rect 18319 10308 18343 10310
rect 18399 10308 18423 10310
rect 18479 10308 18503 10310
rect 18559 10308 18565 10310
rect 18257 10299 18565 10308
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18510 10024 18566 10033
rect 18510 9959 18566 9968
rect 18524 9586 18552 9959
rect 18616 9722 18644 11018
rect 18786 10976 18842 10985
rect 18786 10911 18842 10920
rect 18696 10668 18748 10674
rect 18696 10610 18748 10616
rect 18708 10266 18736 10610
rect 18800 10266 18828 10911
rect 18880 10804 18932 10810
rect 18880 10746 18932 10752
rect 18892 10266 18920 10746
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18880 10260 18932 10266
rect 18880 10202 18932 10208
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18694 10024 18750 10033
rect 18694 9959 18750 9968
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18708 9518 18736 9959
rect 18800 9518 18828 10066
rect 18880 9716 18932 9722
rect 18880 9658 18932 9664
rect 18696 9512 18748 9518
rect 18696 9454 18748 9460
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18050 9208 18106 9217
rect 18030 9152 18050 9194
rect 18030 9143 18106 9152
rect 18030 9132 18092 9143
rect 18064 8974 18092 9132
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17868 8560 17920 8566
rect 17920 8520 18000 8548
rect 17868 8502 17920 8508
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17684 8288 17736 8294
rect 17684 8230 17736 8236
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17684 7880 17736 7886
rect 17684 7822 17736 7828
rect 17696 7546 17724 7822
rect 17788 7750 17816 8434
rect 17776 7744 17828 7750
rect 17828 7704 17908 7732
rect 17776 7686 17828 7692
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17682 7440 17738 7449
rect 17682 7375 17738 7384
rect 17590 7304 17646 7313
rect 17590 7239 17646 7248
rect 17604 5370 17632 7239
rect 17696 6322 17724 7375
rect 17776 6656 17828 6662
rect 17776 6598 17828 6604
rect 17684 6316 17736 6322
rect 17684 6258 17736 6264
rect 17684 6180 17736 6186
rect 17684 6122 17736 6128
rect 17696 6089 17724 6122
rect 17682 6080 17738 6089
rect 17682 6015 17738 6024
rect 17682 5808 17738 5817
rect 17682 5743 17738 5752
rect 17696 5370 17724 5743
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17696 5234 17724 5306
rect 17500 5228 17552 5234
rect 17500 5170 17552 5176
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17498 4856 17554 4865
rect 17498 4791 17554 4800
rect 17512 4214 17540 4791
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17408 4140 17460 4146
rect 17408 4082 17460 4088
rect 17328 4026 17356 4082
rect 17696 4026 17724 5170
rect 17788 4758 17816 6598
rect 17880 6254 17908 7704
rect 17972 7410 18000 8520
rect 18156 8294 18184 9318
rect 18257 9276 18565 9285
rect 18257 9274 18263 9276
rect 18319 9274 18343 9276
rect 18399 9274 18423 9276
rect 18479 9274 18503 9276
rect 18559 9274 18565 9276
rect 18319 9222 18321 9274
rect 18501 9222 18503 9274
rect 18257 9220 18263 9222
rect 18319 9220 18343 9222
rect 18399 9220 18423 9222
rect 18479 9220 18503 9222
rect 18559 9220 18565 9222
rect 18257 9211 18565 9220
rect 18694 9208 18750 9217
rect 18432 9152 18694 9160
rect 18892 9194 18920 9658
rect 18432 9143 18750 9152
rect 18800 9166 18920 9194
rect 18432 9132 18736 9143
rect 18326 8936 18382 8945
rect 18326 8871 18328 8880
rect 18380 8871 18382 8880
rect 18328 8842 18380 8848
rect 18432 8294 18460 9132
rect 18800 9058 18828 9166
rect 18616 9030 18828 9058
rect 18878 9072 18934 9081
rect 18512 8832 18564 8838
rect 18512 8774 18564 8780
rect 18524 8430 18552 8774
rect 18616 8498 18644 9030
rect 18878 9007 18934 9016
rect 18788 8968 18840 8974
rect 18788 8910 18840 8916
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18708 8537 18736 8842
rect 18694 8528 18750 8537
rect 18604 8492 18656 8498
rect 18694 8463 18750 8472
rect 18604 8434 18656 8440
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18800 8362 18828 8910
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18144 8288 18196 8294
rect 18050 8256 18106 8265
rect 18432 8266 18644 8294
rect 18144 8230 18196 8236
rect 18050 8191 18106 8200
rect 18064 7750 18092 8191
rect 18257 8188 18565 8197
rect 18257 8186 18263 8188
rect 18319 8186 18343 8188
rect 18399 8186 18423 8188
rect 18479 8186 18503 8188
rect 18559 8186 18565 8188
rect 18319 8134 18321 8186
rect 18501 8134 18503 8186
rect 18257 8132 18263 8134
rect 18319 8132 18343 8134
rect 18399 8132 18423 8134
rect 18479 8132 18503 8134
rect 18559 8132 18565 8134
rect 18257 8123 18565 8132
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18052 7472 18104 7478
rect 18052 7414 18104 7420
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 17868 6248 17920 6254
rect 17868 6190 17920 6196
rect 17972 5710 18000 7346
rect 18064 7274 18092 7414
rect 18248 7410 18276 7822
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18052 7268 18104 7274
rect 18052 7210 18104 7216
rect 18257 7100 18565 7109
rect 18257 7098 18263 7100
rect 18319 7098 18343 7100
rect 18399 7098 18423 7100
rect 18479 7098 18503 7100
rect 18559 7098 18565 7100
rect 18319 7046 18321 7098
rect 18501 7046 18503 7098
rect 18257 7044 18263 7046
rect 18319 7044 18343 7046
rect 18399 7044 18423 7046
rect 18479 7044 18503 7046
rect 18559 7044 18565 7046
rect 18050 7032 18106 7041
rect 18257 7035 18565 7044
rect 18616 7002 18644 8266
rect 18892 8022 18920 9007
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18878 7712 18934 7721
rect 18050 6967 18106 6976
rect 18604 6996 18656 7002
rect 18064 6798 18092 6967
rect 18604 6938 18656 6944
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18420 6792 18472 6798
rect 18604 6792 18656 6798
rect 18420 6734 18472 6740
rect 18524 6752 18604 6780
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18156 6390 18184 6598
rect 18234 6488 18290 6497
rect 18234 6423 18290 6432
rect 18248 6390 18276 6423
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 18144 6384 18196 6390
rect 18144 6326 18196 6332
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 17960 5704 18012 5710
rect 17960 5646 18012 5652
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 17328 3998 17724 4026
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17328 3466 17356 3998
rect 17590 3904 17646 3913
rect 17590 3839 17646 3848
rect 17498 3768 17554 3777
rect 17498 3703 17554 3712
rect 17316 3460 17368 3466
rect 17316 3402 17368 3408
rect 17316 3188 17368 3194
rect 17316 3130 17368 3136
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17236 2514 17264 2790
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17132 1488 17184 1494
rect 17132 1430 17184 1436
rect 17132 1352 17184 1358
rect 17132 1294 17184 1300
rect 17144 160 17172 1294
rect 17236 1018 17264 2246
rect 17328 1737 17356 3130
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17314 1728 17370 1737
rect 17314 1663 17370 1672
rect 17420 1562 17448 2994
rect 17512 2514 17540 3703
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17500 1896 17552 1902
rect 17500 1838 17552 1844
rect 17408 1556 17460 1562
rect 17408 1498 17460 1504
rect 17316 1420 17368 1426
rect 17316 1362 17368 1368
rect 17224 1012 17276 1018
rect 17224 954 17276 960
rect 17328 160 17356 1362
rect 17512 160 17540 1838
rect 17604 649 17632 3839
rect 17788 3194 17816 4490
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 17880 2774 17908 5578
rect 17958 5400 18014 5409
rect 17958 5335 18014 5344
rect 17972 4078 18000 5335
rect 17960 4072 18012 4078
rect 17960 4014 18012 4020
rect 17960 3936 18012 3942
rect 17960 3878 18012 3884
rect 17972 3534 18000 3878
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17696 2746 17908 2774
rect 17590 640 17646 649
rect 17590 575 17646 584
rect 17696 160 17724 2746
rect 17972 2666 18000 3470
rect 17880 2638 18000 2666
rect 17774 2136 17830 2145
rect 17880 2122 17908 2638
rect 17958 2408 18014 2417
rect 17958 2343 18014 2352
rect 17830 2094 17908 2122
rect 17774 2071 17830 2080
rect 17972 1358 18000 2343
rect 18064 1562 18092 6326
rect 18144 6248 18196 6254
rect 18144 6190 18196 6196
rect 18156 5778 18184 6190
rect 18432 6186 18460 6734
rect 18524 6633 18552 6752
rect 18604 6734 18656 6740
rect 18604 6656 18656 6662
rect 18510 6624 18566 6633
rect 18604 6598 18656 6604
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18510 6559 18566 6568
rect 18510 6488 18566 6497
rect 18510 6423 18566 6432
rect 18524 6390 18552 6423
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18420 6180 18472 6186
rect 18420 6122 18472 6128
rect 18257 6012 18565 6021
rect 18257 6010 18263 6012
rect 18319 6010 18343 6012
rect 18399 6010 18423 6012
rect 18479 6010 18503 6012
rect 18559 6010 18565 6012
rect 18319 5958 18321 6010
rect 18501 5958 18503 6010
rect 18257 5956 18263 5958
rect 18319 5956 18343 5958
rect 18399 5956 18423 5958
rect 18479 5956 18503 5958
rect 18559 5956 18565 5958
rect 18257 5947 18565 5956
rect 18144 5772 18196 5778
rect 18144 5714 18196 5720
rect 18142 5536 18198 5545
rect 18142 5471 18198 5480
rect 18156 4690 18184 5471
rect 18616 5166 18644 6598
rect 18708 6322 18736 6598
rect 18696 6316 18748 6322
rect 18696 6258 18748 6264
rect 18604 5160 18656 5166
rect 18604 5102 18656 5108
rect 18708 5098 18736 6258
rect 18800 5914 18828 7686
rect 18878 7647 18934 7656
rect 18892 6798 18920 7647
rect 18984 7410 19012 11183
rect 19156 11154 19208 11160
rect 19062 11112 19118 11121
rect 19062 11047 19118 11056
rect 19076 9722 19104 11047
rect 19168 10130 19196 11154
rect 19260 10742 19288 12038
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19156 10124 19208 10130
rect 19156 10066 19208 10072
rect 19064 9716 19116 9722
rect 19064 9658 19116 9664
rect 19062 9580 19114 9586
rect 19062 9522 19114 9528
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18880 6656 18932 6662
rect 18880 6598 18932 6604
rect 18892 6497 18920 6598
rect 18878 6488 18934 6497
rect 18878 6423 18934 6432
rect 18880 6248 18932 6254
rect 19076 6236 19104 9522
rect 19168 9330 19196 10066
rect 19352 9353 19380 12135
rect 19444 11529 19472 12406
rect 19430 11520 19486 11529
rect 19430 11455 19486 11464
rect 19430 9752 19486 9761
rect 19430 9687 19486 9696
rect 19444 9432 19472 9687
rect 19536 9654 19564 12650
rect 19628 11082 19656 14214
rect 19720 13530 19748 14758
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19616 11076 19668 11082
rect 19616 11018 19668 11024
rect 19616 10600 19668 10606
rect 19616 10542 19668 10548
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19524 9444 19576 9450
rect 19444 9404 19524 9432
rect 19524 9386 19576 9392
rect 19338 9344 19394 9353
rect 19168 9302 19288 9330
rect 19154 9208 19210 9217
rect 19154 9143 19210 9152
rect 18880 6190 18932 6196
rect 18984 6208 19104 6236
rect 18788 5908 18840 5914
rect 18788 5850 18840 5856
rect 18788 5704 18840 5710
rect 18892 5658 18920 6190
rect 18840 5652 18920 5658
rect 18788 5646 18920 5652
rect 18800 5630 18920 5646
rect 18786 5536 18842 5545
rect 18786 5471 18842 5480
rect 18800 5234 18828 5471
rect 18892 5234 18920 5630
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18880 5228 18932 5234
rect 18880 5170 18932 5176
rect 18696 5092 18748 5098
rect 18696 5034 18748 5040
rect 18788 5024 18840 5030
rect 18788 4966 18840 4972
rect 18257 4924 18565 4933
rect 18257 4922 18263 4924
rect 18319 4922 18343 4924
rect 18399 4922 18423 4924
rect 18479 4922 18503 4924
rect 18559 4922 18565 4924
rect 18319 4870 18321 4922
rect 18501 4870 18503 4922
rect 18257 4868 18263 4870
rect 18319 4868 18343 4870
rect 18399 4868 18423 4870
rect 18479 4868 18503 4870
rect 18559 4868 18565 4870
rect 18257 4859 18565 4868
rect 18800 4826 18828 4966
rect 18788 4820 18840 4826
rect 18788 4762 18840 4768
rect 18234 4720 18290 4729
rect 18144 4684 18196 4690
rect 18234 4655 18290 4664
rect 18144 4626 18196 4632
rect 18248 4622 18276 4655
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18788 4480 18840 4486
rect 18788 4422 18840 4428
rect 18604 4140 18656 4146
rect 18604 4082 18656 4088
rect 18144 4072 18196 4078
rect 18144 4014 18196 4020
rect 18156 3670 18184 4014
rect 18257 3836 18565 3845
rect 18257 3834 18263 3836
rect 18319 3834 18343 3836
rect 18399 3834 18423 3836
rect 18479 3834 18503 3836
rect 18559 3834 18565 3836
rect 18319 3782 18321 3834
rect 18501 3782 18503 3834
rect 18257 3780 18263 3782
rect 18319 3780 18343 3782
rect 18399 3780 18423 3782
rect 18479 3780 18503 3782
rect 18559 3780 18565 3782
rect 18257 3771 18565 3780
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18234 3632 18290 3641
rect 18234 3567 18290 3576
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18052 1556 18104 1562
rect 18052 1498 18104 1504
rect 17960 1352 18012 1358
rect 17960 1294 18012 1300
rect 18050 1320 18106 1329
rect 18050 1255 18106 1264
rect 17776 1216 17828 1222
rect 17776 1158 17828 1164
rect 17788 950 17816 1158
rect 18064 1018 18092 1255
rect 18052 1012 18104 1018
rect 18052 954 18104 960
rect 17776 944 17828 950
rect 17776 886 17828 892
rect 17868 604 17920 610
rect 17868 546 17920 552
rect 17880 160 17908 546
rect 18156 513 18184 3470
rect 18248 3194 18276 3567
rect 18328 3528 18380 3534
rect 18616 3505 18644 4082
rect 18694 3904 18750 3913
rect 18694 3839 18750 3848
rect 18708 3738 18736 3839
rect 18696 3732 18748 3738
rect 18696 3674 18748 3680
rect 18328 3470 18380 3476
rect 18602 3496 18658 3505
rect 18236 3188 18288 3194
rect 18236 3130 18288 3136
rect 18340 3126 18368 3470
rect 18602 3431 18658 3440
rect 18602 3360 18658 3369
rect 18602 3295 18658 3304
rect 18616 3126 18644 3295
rect 18800 3194 18828 4422
rect 18892 4214 18920 5170
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 18892 3233 18920 4150
rect 18984 3466 19012 6208
rect 19064 4548 19116 4554
rect 19064 4490 19116 4496
rect 19076 4214 19104 4490
rect 19168 4282 19196 9143
rect 19260 9042 19288 9302
rect 19338 9279 19394 9288
rect 19522 9072 19578 9081
rect 19248 9036 19300 9042
rect 19300 8996 19380 9024
rect 19522 9007 19578 9016
rect 19248 8978 19300 8984
rect 19246 8800 19302 8809
rect 19246 8735 19302 8744
rect 19260 7834 19288 8735
rect 19352 8129 19380 8996
rect 19536 8974 19564 9007
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19628 8922 19656 10542
rect 19720 9994 19748 12174
rect 19812 11830 19840 14878
rect 19904 13138 19932 21014
rect 19996 20942 20024 22066
rect 20180 21978 20208 26846
rect 20260 26512 20312 26518
rect 20258 26480 20260 26489
rect 20312 26480 20314 26489
rect 20258 26415 20314 26424
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 20272 25498 20300 26318
rect 20260 25492 20312 25498
rect 20260 25434 20312 25440
rect 20260 24608 20312 24614
rect 20258 24576 20260 24585
rect 20312 24576 20314 24585
rect 20258 24511 20314 24520
rect 20364 24206 20392 29990
rect 20442 29951 20498 29960
rect 20444 29028 20496 29034
rect 20444 28970 20496 28976
rect 20456 28937 20484 28970
rect 20442 28928 20498 28937
rect 20442 28863 20498 28872
rect 20444 28416 20496 28422
rect 20442 28384 20444 28393
rect 20496 28384 20498 28393
rect 20442 28319 20498 28328
rect 20444 27872 20496 27878
rect 20442 27840 20444 27849
rect 20496 27840 20498 27849
rect 20442 27775 20498 27784
rect 20548 27554 20576 31436
rect 20628 31418 20680 31424
rect 20626 31240 20682 31249
rect 20626 31175 20682 31184
rect 20640 28082 20668 31175
rect 20729 30492 21037 30501
rect 20729 30490 20735 30492
rect 20791 30490 20815 30492
rect 20871 30490 20895 30492
rect 20951 30490 20975 30492
rect 21031 30490 21037 30492
rect 20791 30438 20793 30490
rect 20973 30438 20975 30490
rect 20729 30436 20735 30438
rect 20791 30436 20815 30438
rect 20871 30436 20895 30438
rect 20951 30436 20975 30438
rect 21031 30436 21037 30438
rect 20729 30427 21037 30436
rect 20729 29404 21037 29413
rect 20729 29402 20735 29404
rect 20791 29402 20815 29404
rect 20871 29402 20895 29404
rect 20951 29402 20975 29404
rect 21031 29402 21037 29404
rect 20791 29350 20793 29402
rect 20973 29350 20975 29402
rect 20729 29348 20735 29350
rect 20791 29348 20815 29350
rect 20871 29348 20895 29350
rect 20951 29348 20975 29350
rect 21031 29348 21037 29350
rect 20729 29339 21037 29348
rect 20729 28316 21037 28325
rect 20729 28314 20735 28316
rect 20791 28314 20815 28316
rect 20871 28314 20895 28316
rect 20951 28314 20975 28316
rect 21031 28314 21037 28316
rect 20791 28262 20793 28314
rect 20973 28262 20975 28314
rect 20729 28260 20735 28262
rect 20791 28260 20815 28262
rect 20871 28260 20895 28262
rect 20951 28260 20975 28262
rect 21031 28260 21037 28262
rect 20729 28251 21037 28260
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20456 27526 20576 27554
rect 20626 27568 20682 27577
rect 20456 26246 20484 27526
rect 20626 27503 20682 27512
rect 20536 27396 20588 27402
rect 20536 27338 20588 27344
rect 20548 26761 20576 27338
rect 20640 27010 20668 27503
rect 20729 27228 21037 27237
rect 20729 27226 20735 27228
rect 20791 27226 20815 27228
rect 20871 27226 20895 27228
rect 20951 27226 20975 27228
rect 21031 27226 21037 27228
rect 20791 27174 20793 27226
rect 20973 27174 20975 27226
rect 20729 27172 20735 27174
rect 20791 27172 20815 27174
rect 20871 27172 20895 27174
rect 20951 27172 20975 27174
rect 21031 27172 21037 27174
rect 20729 27163 21037 27172
rect 20640 26982 20760 27010
rect 20628 26784 20680 26790
rect 20534 26752 20590 26761
rect 20628 26726 20680 26732
rect 20534 26687 20590 26696
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20536 26240 20588 26246
rect 20536 26182 20588 26188
rect 20444 25696 20496 25702
rect 20444 25638 20496 25644
rect 20352 24200 20404 24206
rect 20456 24177 20484 25638
rect 20352 24142 20404 24148
rect 20442 24168 20498 24177
rect 20442 24103 20498 24112
rect 20260 24064 20312 24070
rect 20260 24006 20312 24012
rect 20272 23866 20300 24006
rect 20260 23860 20312 23866
rect 20260 23802 20312 23808
rect 20548 23712 20576 26182
rect 20640 25401 20668 26726
rect 20732 26246 20760 26982
rect 20720 26240 20772 26246
rect 20720 26182 20772 26188
rect 20729 26140 21037 26149
rect 20729 26138 20735 26140
rect 20791 26138 20815 26140
rect 20871 26138 20895 26140
rect 20951 26138 20975 26140
rect 21031 26138 21037 26140
rect 20791 26086 20793 26138
rect 20973 26086 20975 26138
rect 20729 26084 20735 26086
rect 20791 26084 20815 26086
rect 20871 26084 20895 26086
rect 20951 26084 20975 26086
rect 21031 26084 21037 26086
rect 20729 26075 21037 26084
rect 20626 25392 20682 25401
rect 20626 25327 20682 25336
rect 20729 25052 21037 25061
rect 20729 25050 20735 25052
rect 20791 25050 20815 25052
rect 20871 25050 20895 25052
rect 20951 25050 20975 25052
rect 21031 25050 21037 25052
rect 20791 24998 20793 25050
rect 20973 24998 20975 25050
rect 20729 24996 20735 24998
rect 20791 24996 20815 24998
rect 20871 24996 20895 24998
rect 20951 24996 20975 24998
rect 21031 24996 21037 24998
rect 20729 24987 21037 24996
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20456 23684 20576 23712
rect 20456 23610 20484 23684
rect 20456 23582 20576 23610
rect 20444 23520 20496 23526
rect 20442 23488 20444 23497
rect 20496 23488 20498 23497
rect 20442 23423 20498 23432
rect 20260 23248 20312 23254
rect 20312 23196 20392 23202
rect 20260 23190 20392 23196
rect 20272 23174 20392 23190
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20272 22234 20300 22986
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 20088 21950 20208 21978
rect 20088 21468 20116 21950
rect 20364 21842 20392 23174
rect 20444 22976 20496 22982
rect 20444 22918 20496 22924
rect 20456 22710 20484 22918
rect 20444 22704 20496 22710
rect 20444 22646 20496 22652
rect 20444 22432 20496 22438
rect 20442 22400 20444 22409
rect 20496 22400 20498 22409
rect 20442 22335 20498 22344
rect 20180 21814 20392 21842
rect 20180 21622 20208 21814
rect 20168 21616 20220 21622
rect 20168 21558 20220 21564
rect 20548 21554 20576 23582
rect 20536 21548 20588 21554
rect 20536 21490 20588 21496
rect 20444 21480 20496 21486
rect 20088 21440 20208 21468
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19996 20058 20024 20198
rect 20088 20058 20116 20402
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 20076 20052 20128 20058
rect 20076 19994 20128 20000
rect 19984 19440 20036 19446
rect 19984 19382 20036 19388
rect 19996 17202 20024 19382
rect 20076 19168 20128 19174
rect 20074 19136 20076 19145
rect 20128 19136 20130 19145
rect 20074 19071 20130 19080
rect 20180 18766 20208 21440
rect 20444 21422 20496 21428
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20260 20256 20312 20262
rect 20260 20198 20312 20204
rect 20272 19514 20300 20198
rect 20260 19508 20312 19514
rect 20260 19450 20312 19456
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 20168 18760 20220 18766
rect 20168 18702 20220 18708
rect 20272 17882 20300 19314
rect 20364 19310 20392 20946
rect 20352 19304 20404 19310
rect 20352 19246 20404 19252
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20364 18970 20392 19110
rect 20352 18964 20404 18970
rect 20352 18906 20404 18912
rect 20260 17876 20312 17882
rect 20260 17818 20312 17824
rect 20272 17542 20300 17818
rect 20260 17536 20312 17542
rect 20260 17478 20312 17484
rect 19984 17196 20036 17202
rect 19984 17138 20036 17144
rect 19982 17096 20038 17105
rect 19982 17031 20038 17040
rect 19996 15366 20024 17031
rect 20456 16776 20484 21422
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20548 17678 20576 19246
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20364 16748 20484 16776
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 20076 14884 20128 14890
rect 20076 14826 20128 14832
rect 19904 13110 20024 13138
rect 19996 12714 20024 13110
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 19892 12640 19944 12646
rect 19892 12582 19944 12588
rect 19904 12209 19932 12582
rect 19984 12368 20036 12374
rect 19984 12310 20036 12316
rect 19890 12200 19946 12209
rect 19890 12135 19946 12144
rect 19800 11824 19852 11830
rect 19800 11766 19852 11772
rect 19798 11656 19854 11665
rect 19798 11591 19854 11600
rect 19812 10538 19840 11591
rect 19800 10532 19852 10538
rect 19800 10474 19852 10480
rect 19708 9988 19760 9994
rect 19708 9930 19760 9936
rect 19706 9888 19762 9897
rect 19762 9846 19840 9874
rect 19706 9823 19762 9832
rect 19628 8894 19748 8922
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19430 8664 19486 8673
rect 19430 8599 19486 8608
rect 19444 8566 19472 8599
rect 19432 8560 19484 8566
rect 19432 8502 19484 8508
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19338 8120 19394 8129
rect 19338 8055 19394 8064
rect 19536 7954 19564 8230
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19628 7886 19656 8774
rect 19720 8566 19748 8894
rect 19708 8560 19760 8566
rect 19708 8502 19760 8508
rect 19616 7880 19668 7886
rect 19260 7806 19380 7834
rect 19616 7822 19668 7828
rect 19352 7750 19380 7806
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19616 7744 19668 7750
rect 19616 7686 19668 7692
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19248 6996 19300 7002
rect 19248 6938 19300 6944
rect 19260 4622 19288 6938
rect 19536 6882 19564 7482
rect 19628 6914 19656 7686
rect 19720 7410 19748 8502
rect 19812 7562 19840 9846
rect 19890 9480 19946 9489
rect 19890 9415 19946 9424
rect 19904 8022 19932 9415
rect 19892 8016 19944 8022
rect 19892 7958 19944 7964
rect 19892 7880 19944 7886
rect 19890 7848 19892 7857
rect 19944 7848 19946 7857
rect 19890 7783 19946 7792
rect 19812 7534 19932 7562
rect 19904 7478 19932 7534
rect 19892 7472 19944 7478
rect 19892 7414 19944 7420
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19628 6886 19840 6914
rect 19444 6854 19564 6882
rect 19444 6610 19472 6854
rect 19616 6792 19668 6798
rect 19668 6769 19748 6780
rect 19668 6760 19762 6769
rect 19668 6752 19706 6760
rect 19616 6734 19668 6740
rect 19706 6695 19762 6704
rect 19444 6582 19656 6610
rect 19522 6488 19578 6497
rect 19628 6458 19656 6582
rect 19522 6423 19578 6432
rect 19616 6452 19668 6458
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19444 5137 19472 5170
rect 19430 5128 19486 5137
rect 19430 5063 19486 5072
rect 19248 4616 19300 4622
rect 19248 4558 19300 4564
rect 19432 4548 19484 4554
rect 19432 4490 19484 4496
rect 19246 4312 19302 4321
rect 19156 4276 19208 4282
rect 19246 4247 19302 4256
rect 19156 4218 19208 4224
rect 19064 4208 19116 4214
rect 19064 4150 19116 4156
rect 19156 3936 19208 3942
rect 19156 3878 19208 3884
rect 19064 3528 19116 3534
rect 19064 3470 19116 3476
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18878 3224 18934 3233
rect 18788 3188 18840 3194
rect 18878 3159 18934 3168
rect 18788 3130 18840 3136
rect 18328 3120 18380 3126
rect 18328 3062 18380 3068
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18788 3052 18840 3058
rect 18892 3040 18920 3159
rect 18840 3012 18920 3040
rect 18788 2994 18840 3000
rect 18878 2816 18934 2825
rect 18257 2748 18565 2757
rect 18878 2751 18934 2760
rect 18257 2746 18263 2748
rect 18319 2746 18343 2748
rect 18399 2746 18423 2748
rect 18479 2746 18503 2748
rect 18559 2746 18565 2748
rect 18319 2694 18321 2746
rect 18501 2694 18503 2746
rect 18257 2692 18263 2694
rect 18319 2692 18343 2694
rect 18399 2692 18423 2694
rect 18479 2692 18503 2694
rect 18559 2692 18565 2694
rect 18257 2683 18565 2692
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18257 1660 18565 1669
rect 18257 1658 18263 1660
rect 18319 1658 18343 1660
rect 18399 1658 18423 1660
rect 18479 1658 18503 1660
rect 18559 1658 18565 1660
rect 18319 1606 18321 1658
rect 18501 1606 18503 1658
rect 18257 1604 18263 1606
rect 18319 1604 18343 1606
rect 18399 1604 18423 1606
rect 18479 1604 18503 1606
rect 18559 1604 18565 1606
rect 18257 1595 18565 1604
rect 18418 912 18474 921
rect 18418 847 18474 856
rect 18142 504 18198 513
rect 18142 439 18198 448
rect 18236 468 18288 474
rect 18236 410 18288 416
rect 17972 160 18092 184
rect 18248 160 18276 410
rect 18432 160 18460 847
rect 18708 610 18736 2450
rect 18892 1358 18920 2751
rect 18880 1352 18932 1358
rect 18880 1294 18932 1300
rect 18970 1048 19026 1057
rect 18970 983 19026 992
rect 18696 604 18748 610
rect 18696 546 18748 552
rect 18786 368 18842 377
rect 18786 303 18842 312
rect 18510 232 18566 241
rect 18510 167 18566 176
rect 16946 54 17080 82
rect 16578 -300 16634 54
rect 16762 -300 16818 54
rect 16946 -300 17002 54
rect 17130 -300 17186 160
rect 17314 -300 17370 160
rect 17498 -300 17554 160
rect 17682 -300 17738 160
rect 17866 -300 17922 160
rect 17972 156 18106 160
rect 17972 105 18000 156
rect 17956 96 18012 105
rect 17956 31 18012 40
rect 18050 -300 18106 156
rect 18234 -300 18290 160
rect 18418 -300 18474 160
rect 18524 82 18552 167
rect 18800 160 18828 303
rect 18984 160 19012 983
rect 19076 785 19104 3470
rect 19168 2378 19196 3878
rect 19260 2582 19288 4247
rect 19340 3732 19392 3738
rect 19340 3674 19392 3680
rect 19248 2576 19300 2582
rect 19248 2518 19300 2524
rect 19156 2372 19208 2378
rect 19156 2314 19208 2320
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19062 776 19118 785
rect 19062 711 19118 720
rect 19260 406 19288 2246
rect 19248 400 19300 406
rect 19248 342 19300 348
rect 19156 264 19208 270
rect 19156 206 19208 212
rect 19168 160 19196 206
rect 19352 160 19380 3674
rect 19444 338 19472 4490
rect 19536 3126 19564 6423
rect 19616 6394 19668 6400
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19616 5636 19668 5642
rect 19616 5578 19668 5584
rect 19628 4622 19656 5578
rect 19616 4616 19668 4622
rect 19616 4558 19668 4564
rect 19720 4146 19748 6258
rect 19812 5642 19840 6886
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 19904 6118 19932 6598
rect 19892 6112 19944 6118
rect 19892 6054 19944 6060
rect 19800 5636 19852 5642
rect 19800 5578 19852 5584
rect 19996 5370 20024 12310
rect 20088 11354 20116 14826
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20180 14074 20208 14214
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20180 12986 20208 13874
rect 20168 12980 20220 12986
rect 20168 12922 20220 12928
rect 20260 12232 20312 12238
rect 20260 12174 20312 12180
rect 20076 11348 20128 11354
rect 20076 11290 20128 11296
rect 20076 11076 20128 11082
rect 20076 11018 20128 11024
rect 20088 10452 20116 11018
rect 20272 10792 20300 12174
rect 20180 10764 20300 10792
rect 20180 10577 20208 10764
rect 20260 10668 20312 10674
rect 20260 10610 20312 10616
rect 20166 10568 20222 10577
rect 20166 10503 20222 10512
rect 20088 10424 20208 10452
rect 20076 9376 20128 9382
rect 20076 9318 20128 9324
rect 20088 9110 20116 9318
rect 20076 9104 20128 9110
rect 20076 9046 20128 9052
rect 20074 8392 20130 8401
rect 20074 8327 20130 8336
rect 20088 6934 20116 8327
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 19984 5364 20036 5370
rect 19984 5306 20036 5312
rect 20088 4758 20116 5850
rect 20180 5710 20208 10424
rect 20272 7546 20300 10610
rect 20364 9432 20392 16748
rect 20444 16652 20496 16658
rect 20444 16594 20496 16600
rect 20456 16561 20484 16594
rect 20442 16552 20498 16561
rect 20442 16487 20498 16496
rect 20444 15904 20496 15910
rect 20442 15872 20444 15881
rect 20496 15872 20498 15881
rect 20442 15807 20498 15816
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 20444 14816 20496 14822
rect 20442 14784 20444 14793
rect 20496 14784 20498 14793
rect 20442 14719 20498 14728
rect 20548 11898 20576 15098
rect 20536 11892 20588 11898
rect 20536 11834 20588 11840
rect 20534 10432 20590 10441
rect 20534 10367 20590 10376
rect 20364 9404 20484 9432
rect 20350 9344 20406 9353
rect 20350 9279 20406 9288
rect 20364 9178 20392 9279
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20260 7540 20312 7546
rect 20260 7482 20312 7488
rect 20456 6914 20484 9404
rect 20548 7546 20576 10367
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20640 7324 20668 24142
rect 20729 23964 21037 23973
rect 20729 23962 20735 23964
rect 20791 23962 20815 23964
rect 20871 23962 20895 23964
rect 20951 23962 20975 23964
rect 21031 23962 21037 23964
rect 20791 23910 20793 23962
rect 20973 23910 20975 23962
rect 20729 23908 20735 23910
rect 20791 23908 20815 23910
rect 20871 23908 20895 23910
rect 20951 23908 20975 23910
rect 21031 23908 21037 23910
rect 20729 23899 21037 23908
rect 20729 22876 21037 22885
rect 20729 22874 20735 22876
rect 20791 22874 20815 22876
rect 20871 22874 20895 22876
rect 20951 22874 20975 22876
rect 21031 22874 21037 22876
rect 20791 22822 20793 22874
rect 20973 22822 20975 22874
rect 20729 22820 20735 22822
rect 20791 22820 20815 22822
rect 20871 22820 20895 22822
rect 20951 22820 20975 22822
rect 21031 22820 21037 22822
rect 20729 22811 21037 22820
rect 20729 21788 21037 21797
rect 20729 21786 20735 21788
rect 20791 21786 20815 21788
rect 20871 21786 20895 21788
rect 20951 21786 20975 21788
rect 21031 21786 21037 21788
rect 20791 21734 20793 21786
rect 20973 21734 20975 21786
rect 20729 21732 20735 21734
rect 20791 21732 20815 21734
rect 20871 21732 20895 21734
rect 20951 21732 20975 21734
rect 21031 21732 21037 21734
rect 20729 21723 21037 21732
rect 20729 20700 21037 20709
rect 20729 20698 20735 20700
rect 20791 20698 20815 20700
rect 20871 20698 20895 20700
rect 20951 20698 20975 20700
rect 21031 20698 21037 20700
rect 20791 20646 20793 20698
rect 20973 20646 20975 20698
rect 20729 20644 20735 20646
rect 20791 20644 20815 20646
rect 20871 20644 20895 20646
rect 20951 20644 20975 20646
rect 21031 20644 21037 20646
rect 20729 20635 21037 20644
rect 21100 20482 21128 41074
rect 21272 40452 21324 40458
rect 21272 40394 21324 40400
rect 21284 40361 21312 40394
rect 21270 40352 21326 40361
rect 21270 40287 21326 40296
rect 21178 39400 21234 39409
rect 21178 39335 21234 39344
rect 21272 39364 21324 39370
rect 21192 33946 21220 39335
rect 21272 39306 21324 39312
rect 21284 39273 21312 39306
rect 21270 39264 21326 39273
rect 21270 39199 21326 39208
rect 21454 38312 21510 38321
rect 21272 38276 21324 38282
rect 21454 38247 21510 38256
rect 21272 38218 21324 38224
rect 21284 38185 21312 38218
rect 21270 38176 21326 38185
rect 21270 38111 21326 38120
rect 21272 36576 21324 36582
rect 21272 36518 21324 36524
rect 21284 36009 21312 36518
rect 21270 36000 21326 36009
rect 21270 35935 21326 35944
rect 21364 35488 21416 35494
rect 21364 35430 21416 35436
rect 21272 34944 21324 34950
rect 21270 34912 21272 34921
rect 21324 34912 21326 34921
rect 21270 34847 21326 34856
rect 21192 33918 21312 33946
rect 21180 33856 21232 33862
rect 21178 33824 21180 33833
rect 21232 33824 21234 33833
rect 21178 33759 21234 33768
rect 21284 33674 21312 33918
rect 21008 20454 21128 20482
rect 21192 33646 21312 33674
rect 21008 19718 21036 20454
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 20729 19612 21037 19621
rect 20729 19610 20735 19612
rect 20791 19610 20815 19612
rect 20871 19610 20895 19612
rect 20951 19610 20975 19612
rect 21031 19610 21037 19612
rect 20791 19558 20793 19610
rect 20973 19558 20975 19610
rect 20729 19556 20735 19558
rect 20791 19556 20815 19558
rect 20871 19556 20895 19558
rect 20951 19556 20975 19558
rect 21031 19556 21037 19558
rect 20729 19547 21037 19556
rect 20729 18524 21037 18533
rect 20729 18522 20735 18524
rect 20791 18522 20815 18524
rect 20871 18522 20895 18524
rect 20951 18522 20975 18524
rect 21031 18522 21037 18524
rect 20791 18470 20793 18522
rect 20973 18470 20975 18522
rect 20729 18468 20735 18470
rect 20791 18468 20815 18470
rect 20871 18468 20895 18470
rect 20951 18468 20975 18470
rect 21031 18468 21037 18470
rect 20729 18459 21037 18468
rect 20996 18080 21048 18086
rect 20994 18048 20996 18057
rect 21048 18048 21050 18057
rect 20994 17983 21050 17992
rect 20729 17436 21037 17445
rect 20729 17434 20735 17436
rect 20791 17434 20815 17436
rect 20871 17434 20895 17436
rect 20951 17434 20975 17436
rect 21031 17434 21037 17436
rect 20791 17382 20793 17434
rect 20973 17382 20975 17434
rect 20729 17380 20735 17382
rect 20791 17380 20815 17382
rect 20871 17380 20895 17382
rect 20951 17380 20975 17382
rect 21031 17380 21037 17382
rect 20729 17371 21037 17380
rect 20904 16992 20956 16998
rect 20902 16960 20904 16969
rect 20956 16960 20958 16969
rect 20902 16895 20958 16904
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 20729 16348 21037 16357
rect 20729 16346 20735 16348
rect 20791 16346 20815 16348
rect 20871 16346 20895 16348
rect 20951 16346 20975 16348
rect 21031 16346 21037 16348
rect 20791 16294 20793 16346
rect 20973 16294 20975 16346
rect 20729 16292 20735 16294
rect 20791 16292 20815 16294
rect 20871 16292 20895 16294
rect 20951 16292 20975 16294
rect 21031 16292 21037 16294
rect 20729 16283 21037 16292
rect 20729 15260 21037 15269
rect 20729 15258 20735 15260
rect 20791 15258 20815 15260
rect 20871 15258 20895 15260
rect 20951 15258 20975 15260
rect 21031 15258 21037 15260
rect 20791 15206 20793 15258
rect 20973 15206 20975 15258
rect 20729 15204 20735 15206
rect 20791 15204 20815 15206
rect 20871 15204 20895 15206
rect 20951 15204 20975 15206
rect 21031 15204 21037 15206
rect 20729 15195 21037 15204
rect 20729 14172 21037 14181
rect 20729 14170 20735 14172
rect 20791 14170 20815 14172
rect 20871 14170 20895 14172
rect 20951 14170 20975 14172
rect 21031 14170 21037 14172
rect 20791 14118 20793 14170
rect 20973 14118 20975 14170
rect 20729 14116 20735 14118
rect 20791 14116 20815 14118
rect 20871 14116 20895 14118
rect 20951 14116 20975 14118
rect 21031 14116 21037 14118
rect 20729 14107 21037 14116
rect 20729 13084 21037 13093
rect 20729 13082 20735 13084
rect 20791 13082 20815 13084
rect 20871 13082 20895 13084
rect 20951 13082 20975 13084
rect 21031 13082 21037 13084
rect 20791 13030 20793 13082
rect 20973 13030 20975 13082
rect 20729 13028 20735 13030
rect 20791 13028 20815 13030
rect 20871 13028 20895 13030
rect 20951 13028 20975 13030
rect 21031 13028 21037 13030
rect 20729 13019 21037 13028
rect 20729 11996 21037 12005
rect 20729 11994 20735 11996
rect 20791 11994 20815 11996
rect 20871 11994 20895 11996
rect 20951 11994 20975 11996
rect 21031 11994 21037 11996
rect 20791 11942 20793 11994
rect 20973 11942 20975 11994
rect 20729 11940 20735 11942
rect 20791 11940 20815 11942
rect 20871 11940 20895 11942
rect 20951 11940 20975 11942
rect 21031 11940 21037 11942
rect 20729 11931 21037 11940
rect 20729 10908 21037 10917
rect 20729 10906 20735 10908
rect 20791 10906 20815 10908
rect 20871 10906 20895 10908
rect 20951 10906 20975 10908
rect 21031 10906 21037 10908
rect 20791 10854 20793 10906
rect 20973 10854 20975 10906
rect 20729 10852 20735 10854
rect 20791 10852 20815 10854
rect 20871 10852 20895 10854
rect 20951 10852 20975 10854
rect 21031 10852 21037 10854
rect 20729 10843 21037 10852
rect 20729 9820 21037 9829
rect 20729 9818 20735 9820
rect 20791 9818 20815 9820
rect 20871 9818 20895 9820
rect 20951 9818 20975 9820
rect 21031 9818 21037 9820
rect 20791 9766 20793 9818
rect 20973 9766 20975 9818
rect 20729 9764 20735 9766
rect 20791 9764 20815 9766
rect 20871 9764 20895 9766
rect 20951 9764 20975 9766
rect 21031 9764 21037 9766
rect 20729 9755 21037 9764
rect 20729 8732 21037 8741
rect 20729 8730 20735 8732
rect 20791 8730 20815 8732
rect 20871 8730 20895 8732
rect 20951 8730 20975 8732
rect 21031 8730 21037 8732
rect 20791 8678 20793 8730
rect 20973 8678 20975 8730
rect 20729 8676 20735 8678
rect 20791 8676 20815 8678
rect 20871 8676 20895 8678
rect 20951 8676 20975 8678
rect 21031 8676 21037 8678
rect 20729 8667 21037 8676
rect 20729 7644 21037 7653
rect 20729 7642 20735 7644
rect 20791 7642 20815 7644
rect 20871 7642 20895 7644
rect 20951 7642 20975 7644
rect 21031 7642 21037 7644
rect 20791 7590 20793 7642
rect 20973 7590 20975 7642
rect 20729 7588 20735 7590
rect 20791 7588 20815 7590
rect 20871 7588 20895 7590
rect 20951 7588 20975 7590
rect 21031 7588 21037 7590
rect 20729 7579 21037 7588
rect 21100 7426 21128 16390
rect 21008 7398 21128 7426
rect 20640 7296 20760 7324
rect 20732 6914 20760 7296
rect 20272 6886 20484 6914
rect 20640 6886 20760 6914
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 19800 4752 19852 4758
rect 19800 4694 19852 4700
rect 20076 4752 20128 4758
rect 20076 4694 20128 4700
rect 19708 4140 19760 4146
rect 19708 4082 19760 4088
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19524 3120 19576 3126
rect 19524 3062 19576 3068
rect 19628 2961 19656 3470
rect 19614 2952 19670 2961
rect 19614 2887 19670 2896
rect 19614 2816 19670 2825
rect 19614 2751 19670 2760
rect 19628 1426 19656 2751
rect 19616 1420 19668 1426
rect 19616 1362 19668 1368
rect 19812 1358 19840 4694
rect 19890 4584 19946 4593
rect 19890 4519 19946 4528
rect 19904 4282 19932 4519
rect 19892 4276 19944 4282
rect 19892 4218 19944 4224
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20088 2650 20116 3470
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19800 1352 19852 1358
rect 19800 1294 19852 1300
rect 19996 746 20024 2246
rect 19984 740 20036 746
rect 19984 682 20036 688
rect 20180 678 20208 3538
rect 20272 2446 20300 6886
rect 20536 6656 20588 6662
rect 20536 6598 20588 6604
rect 20352 6316 20404 6322
rect 20352 6258 20404 6264
rect 20364 2774 20392 6258
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20456 5234 20484 6054
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20456 4282 20484 4626
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20364 2746 20484 2774
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 20364 814 20392 2246
rect 20352 808 20404 814
rect 20352 750 20404 756
rect 20168 672 20220 678
rect 20168 614 20220 620
rect 19432 332 19484 338
rect 19432 274 19484 280
rect 18602 82 18658 160
rect 18524 54 18658 82
rect 18602 -300 18658 54
rect 18786 -300 18842 160
rect 18970 -300 19026 160
rect 19154 -300 19210 160
rect 19338 -300 19394 160
rect 20456 134 20484 2746
rect 20548 1970 20576 6598
rect 20536 1964 20588 1970
rect 20536 1906 20588 1912
rect 20444 128 20496 134
rect 20444 70 20496 76
rect 20640 66 20668 6886
rect 21008 6662 21036 7398
rect 20996 6656 21048 6662
rect 20996 6598 21048 6604
rect 20729 6556 21037 6565
rect 20729 6554 20735 6556
rect 20791 6554 20815 6556
rect 20871 6554 20895 6556
rect 20951 6554 20975 6556
rect 21031 6554 21037 6556
rect 20791 6502 20793 6554
rect 20973 6502 20975 6554
rect 20729 6500 20735 6502
rect 20791 6500 20815 6502
rect 20871 6500 20895 6502
rect 20951 6500 20975 6502
rect 21031 6500 21037 6502
rect 20729 6491 21037 6500
rect 20729 5468 21037 5477
rect 20729 5466 20735 5468
rect 20791 5466 20815 5468
rect 20871 5466 20895 5468
rect 20951 5466 20975 5468
rect 21031 5466 21037 5468
rect 20791 5414 20793 5466
rect 20973 5414 20975 5466
rect 20729 5412 20735 5414
rect 20791 5412 20815 5414
rect 20871 5412 20895 5414
rect 20951 5412 20975 5414
rect 21031 5412 21037 5414
rect 20729 5403 21037 5412
rect 20729 4380 21037 4389
rect 20729 4378 20735 4380
rect 20791 4378 20815 4380
rect 20871 4378 20895 4380
rect 20951 4378 20975 4380
rect 21031 4378 21037 4380
rect 20791 4326 20793 4378
rect 20973 4326 20975 4378
rect 20729 4324 20735 4326
rect 20791 4324 20815 4326
rect 20871 4324 20895 4326
rect 20951 4324 20975 4326
rect 21031 4324 21037 4326
rect 20729 4315 21037 4324
rect 21192 4078 21220 33646
rect 21272 33040 21324 33046
rect 21272 32982 21324 32988
rect 21284 32745 21312 32982
rect 21270 32736 21326 32745
rect 21270 32671 21326 32680
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 21284 30569 21312 30602
rect 21270 30560 21326 30569
rect 21270 30495 21326 30504
rect 21272 29572 21324 29578
rect 21272 29514 21324 29520
rect 21284 29481 21312 29514
rect 21270 29472 21326 29481
rect 21270 29407 21326 29416
rect 21270 29200 21326 29209
rect 21270 29135 21326 29144
rect 21284 27674 21312 29135
rect 21272 27668 21324 27674
rect 21272 27610 21324 27616
rect 21272 27532 21324 27538
rect 21272 27474 21324 27480
rect 21284 27305 21312 27474
rect 21270 27296 21326 27305
rect 21270 27231 21326 27240
rect 21272 26376 21324 26382
rect 21272 26318 21324 26324
rect 21284 26217 21312 26318
rect 21270 26208 21326 26217
rect 21270 26143 21326 26152
rect 21272 23044 21324 23050
rect 21272 22986 21324 22992
rect 21284 22953 21312 22986
rect 21270 22944 21326 22953
rect 21270 22879 21326 22888
rect 21270 21856 21326 21865
rect 21270 21791 21326 21800
rect 21284 21690 21312 21791
rect 21272 21684 21324 21690
rect 21272 21626 21324 21632
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21284 20777 21312 20810
rect 21270 20768 21326 20777
rect 21270 20703 21326 20712
rect 21272 18828 21324 18834
rect 21272 18770 21324 18776
rect 21284 18601 21312 18770
rect 21270 18592 21326 18601
rect 21270 18527 21326 18536
rect 21270 17504 21326 17513
rect 21270 17439 21326 17448
rect 21284 17338 21312 17439
rect 21272 17332 21324 17338
rect 21272 17274 21324 17280
rect 21272 15428 21324 15434
rect 21272 15370 21324 15376
rect 21284 15337 21312 15370
rect 21270 15328 21326 15337
rect 21270 15263 21326 15272
rect 21270 14240 21326 14249
rect 21270 14175 21326 14184
rect 21284 14074 21312 14175
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21270 13152 21326 13161
rect 21270 13087 21326 13096
rect 21284 12986 21312 13087
rect 21272 12980 21324 12986
rect 21272 12922 21324 12928
rect 21376 12782 21404 35430
rect 21468 18737 21496 38247
rect 21548 37392 21600 37398
rect 21548 37334 21600 37340
rect 21560 27130 21588 37334
rect 21824 37324 21876 37330
rect 21824 37266 21876 37272
rect 21730 36680 21786 36689
rect 21730 36615 21786 36624
rect 21640 32768 21692 32774
rect 21640 32710 21692 32716
rect 21548 27124 21600 27130
rect 21548 27066 21600 27072
rect 21548 26920 21600 26926
rect 21548 26862 21600 26868
rect 21560 22030 21588 26862
rect 21652 23322 21680 32710
rect 21744 31362 21772 36615
rect 21836 31482 21864 37266
rect 21916 31748 21968 31754
rect 21916 31690 21968 31696
rect 21824 31476 21876 31482
rect 21824 31418 21876 31424
rect 21744 31334 21864 31362
rect 21732 31204 21784 31210
rect 21732 31146 21784 31152
rect 21640 23316 21692 23322
rect 21640 23258 21692 23264
rect 21744 23202 21772 31146
rect 21836 28121 21864 31334
rect 21822 28112 21878 28121
rect 21822 28047 21878 28056
rect 21824 27668 21876 27674
rect 21824 27610 21876 27616
rect 21652 23174 21772 23202
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21548 20800 21600 20806
rect 21548 20742 21600 20748
rect 21560 20233 21588 20742
rect 21546 20224 21602 20233
rect 21546 20159 21602 20168
rect 21546 19680 21602 19689
rect 21546 19615 21602 19624
rect 21560 18902 21588 19615
rect 21548 18896 21600 18902
rect 21548 18838 21600 18844
rect 21454 18728 21510 18737
rect 21652 18698 21680 23174
rect 21836 23066 21864 27610
rect 21928 26926 21956 31690
rect 21916 26920 21968 26926
rect 21916 26862 21968 26868
rect 21916 26240 21968 26246
rect 21916 26182 21968 26188
rect 21744 23038 21864 23066
rect 21744 21010 21772 23038
rect 21928 22094 21956 26182
rect 21836 22066 21956 22094
rect 21732 21004 21784 21010
rect 21732 20946 21784 20952
rect 21730 20904 21786 20913
rect 21730 20839 21786 20848
rect 21454 18663 21510 18672
rect 21640 18692 21692 18698
rect 21640 18634 21692 18640
rect 21744 18578 21772 20839
rect 21652 18550 21772 18578
rect 21364 12776 21416 12782
rect 21652 12753 21680 18550
rect 21836 18442 21864 22066
rect 21744 18414 21864 18442
rect 21744 16697 21772 18414
rect 21822 18320 21878 18329
rect 21822 18255 21878 18264
rect 21730 16688 21786 16697
rect 21730 16623 21786 16632
rect 21364 12718 21416 12724
rect 21638 12744 21694 12753
rect 21272 12708 21324 12714
rect 21638 12679 21694 12688
rect 21272 12650 21324 12656
rect 21284 11642 21312 12650
rect 21284 11614 21404 11642
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21284 10985 21312 11494
rect 21270 10976 21326 10985
rect 21270 10911 21326 10920
rect 21376 7682 21404 11614
rect 21364 7676 21416 7682
rect 21364 7618 21416 7624
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21468 4486 21496 7414
rect 21456 4480 21508 4486
rect 21456 4422 21508 4428
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21272 3392 21324 3398
rect 21270 3360 21272 3369
rect 21324 3360 21326 3369
rect 20729 3292 21037 3301
rect 21270 3295 21326 3304
rect 20729 3290 20735 3292
rect 20791 3290 20815 3292
rect 20871 3290 20895 3292
rect 20951 3290 20975 3292
rect 21031 3290 21037 3292
rect 20791 3238 20793 3290
rect 20973 3238 20975 3290
rect 20729 3236 20735 3238
rect 20791 3236 20815 3238
rect 20871 3236 20895 3238
rect 20951 3236 20975 3238
rect 21031 3236 21037 3238
rect 20729 3227 21037 3236
rect 21836 3194 21864 18255
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21928 9586 21956 14554
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21824 3188 21876 3194
rect 21824 3130 21876 3136
rect 20729 2204 21037 2213
rect 20729 2202 20735 2204
rect 20791 2202 20815 2204
rect 20871 2202 20895 2204
rect 20951 2202 20975 2204
rect 21031 2202 21037 2204
rect 20791 2150 20793 2202
rect 20973 2150 20975 2202
rect 20729 2148 20735 2150
rect 20791 2148 20815 2150
rect 20871 2148 20895 2150
rect 20951 2148 20975 2150
rect 21031 2148 21037 2150
rect 20729 2139 21037 2148
rect 21178 1184 21234 1193
rect 20729 1116 21037 1125
rect 21178 1119 21234 1128
rect 20729 1114 20735 1116
rect 20791 1114 20815 1116
rect 20871 1114 20895 1116
rect 20951 1114 20975 1116
rect 21031 1114 21037 1116
rect 20791 1062 20793 1114
rect 20973 1062 20975 1114
rect 20729 1060 20735 1062
rect 20791 1060 20815 1062
rect 20871 1060 20895 1062
rect 20951 1060 20975 1062
rect 21031 1060 21037 1062
rect 20729 1051 21037 1060
rect 21192 202 21220 1119
rect 21180 196 21232 202
rect 21180 138 21232 144
rect 20628 60 20680 66
rect 20628 2 20680 8
<< via2 >>
rect 202 41520 258 41576
rect 294 39752 350 39808
rect 294 27920 350 27976
rect 294 27376 350 27432
rect 478 32816 534 32872
rect 754 31864 810 31920
rect 570 29416 626 29472
rect 754 28872 810 28928
rect 1950 41384 2006 41440
rect 1398 39616 1454 39672
rect 1306 39208 1362 39264
rect 1214 38256 1270 38312
rect 1398 37848 1454 37904
rect 1306 37068 1308 37088
rect 1308 37068 1360 37088
rect 1360 37068 1362 37088
rect 1306 37032 1362 37068
rect 1214 36760 1270 36816
rect 1122 36624 1178 36680
rect 1306 36216 1362 36272
rect 1214 35944 1270 36000
rect 1490 37304 1546 37360
rect 1398 35808 1454 35864
rect 1214 35672 1270 35728
rect 1950 39344 2006 39400
rect 1674 36760 1730 36816
rect 1490 34720 1546 34776
rect 1306 33496 1362 33552
rect 1214 33088 1270 33144
rect 1398 32544 1454 32600
rect 1306 32136 1362 32192
rect 1030 30096 1086 30152
rect 1030 28736 1086 28792
rect 1398 31592 1454 31648
rect 1398 31048 1454 31104
rect 1214 29688 1270 29744
rect 1306 29008 1362 29064
rect 1950 37576 2006 37632
rect 2134 39752 2190 39808
rect 1950 34856 2006 34912
rect 1950 33224 2006 33280
rect 1766 31864 1822 31920
rect 2410 37168 2466 37224
rect 2318 36216 2374 36272
rect 2410 35264 2466 35320
rect 2686 40452 2742 40488
rect 2686 40432 2688 40452
rect 2688 40432 2740 40452
rect 2740 40432 2742 40452
rect 2778 38664 2834 38720
rect 3428 43002 3484 43004
rect 3508 43002 3564 43004
rect 3588 43002 3644 43004
rect 3668 43002 3724 43004
rect 3428 42950 3474 43002
rect 3474 42950 3484 43002
rect 3508 42950 3538 43002
rect 3538 42950 3550 43002
rect 3550 42950 3564 43002
rect 3588 42950 3602 43002
rect 3602 42950 3614 43002
rect 3614 42950 3644 43002
rect 3668 42950 3678 43002
rect 3678 42950 3724 43002
rect 3428 42948 3484 42950
rect 3508 42948 3564 42950
rect 3588 42948 3644 42950
rect 3668 42948 3724 42950
rect 3054 41556 3056 41576
rect 3056 41556 3108 41576
rect 3108 41556 3110 41576
rect 3054 41520 3110 41556
rect 3428 41914 3484 41916
rect 3508 41914 3564 41916
rect 3588 41914 3644 41916
rect 3668 41914 3724 41916
rect 3428 41862 3474 41914
rect 3474 41862 3484 41914
rect 3508 41862 3538 41914
rect 3538 41862 3550 41914
rect 3550 41862 3564 41914
rect 3588 41862 3602 41914
rect 3602 41862 3614 41914
rect 3614 41862 3644 41914
rect 3668 41862 3678 41914
rect 3678 41862 3724 41914
rect 3428 41860 3484 41862
rect 3508 41860 3564 41862
rect 3588 41860 3644 41862
rect 3668 41860 3724 41862
rect 4158 43832 4214 43888
rect 3606 40976 3662 41032
rect 3428 40826 3484 40828
rect 3508 40826 3564 40828
rect 3588 40826 3644 40828
rect 3668 40826 3724 40828
rect 3428 40774 3474 40826
rect 3474 40774 3484 40826
rect 3508 40774 3538 40826
rect 3538 40774 3550 40826
rect 3550 40774 3564 40826
rect 3588 40774 3602 40826
rect 3602 40774 3614 40826
rect 3614 40774 3644 40826
rect 3668 40774 3678 40826
rect 3678 40774 3724 40826
rect 3428 40772 3484 40774
rect 3508 40772 3564 40774
rect 3588 40772 3644 40774
rect 3668 40772 3724 40774
rect 3428 39738 3484 39740
rect 3508 39738 3564 39740
rect 3588 39738 3644 39740
rect 3668 39738 3724 39740
rect 3428 39686 3474 39738
rect 3474 39686 3484 39738
rect 3508 39686 3538 39738
rect 3538 39686 3550 39738
rect 3550 39686 3564 39738
rect 3588 39686 3602 39738
rect 3602 39686 3614 39738
rect 3614 39686 3644 39738
rect 3668 39686 3678 39738
rect 3678 39686 3724 39738
rect 3428 39684 3484 39686
rect 3508 39684 3564 39686
rect 3588 39684 3644 39686
rect 3668 39684 3724 39686
rect 3428 38650 3484 38652
rect 3508 38650 3564 38652
rect 3588 38650 3644 38652
rect 3668 38650 3724 38652
rect 3428 38598 3474 38650
rect 3474 38598 3484 38650
rect 3508 38598 3538 38650
rect 3538 38598 3550 38650
rect 3550 38598 3564 38650
rect 3588 38598 3602 38650
rect 3602 38598 3614 38650
rect 3614 38598 3644 38650
rect 3668 38598 3678 38650
rect 3678 38598 3724 38650
rect 3428 38596 3484 38598
rect 3508 38596 3564 38598
rect 3588 38596 3644 38598
rect 3668 38596 3724 38598
rect 3054 38392 3110 38448
rect 4618 42200 4674 42256
rect 4066 39380 4068 39400
rect 4068 39380 4120 39400
rect 4120 39380 4122 39400
rect 4066 39344 4122 39380
rect 2962 37868 3018 37904
rect 2962 37848 2964 37868
rect 2964 37848 3016 37868
rect 3016 37848 3018 37868
rect 3428 37562 3484 37564
rect 3508 37562 3564 37564
rect 3588 37562 3644 37564
rect 3668 37562 3724 37564
rect 3428 37510 3474 37562
rect 3474 37510 3484 37562
rect 3508 37510 3538 37562
rect 3538 37510 3550 37562
rect 3550 37510 3564 37562
rect 3588 37510 3602 37562
rect 3602 37510 3614 37562
rect 3614 37510 3644 37562
rect 3668 37510 3678 37562
rect 3678 37510 3724 37562
rect 3428 37508 3484 37510
rect 3508 37508 3564 37510
rect 3588 37508 3644 37510
rect 3668 37508 3724 37510
rect 4250 38972 4252 38992
rect 4252 38972 4304 38992
rect 4304 38972 4306 38992
rect 4250 38936 4306 38972
rect 4066 38392 4122 38448
rect 2226 31728 2282 31784
rect 1950 31456 2006 31512
rect 1858 30640 1914 30696
rect 1766 30096 1822 30152
rect 1674 29572 1730 29608
rect 1674 29552 1676 29572
rect 1676 29552 1728 29572
rect 1728 29552 1730 29572
rect 1582 29144 1638 29200
rect 1490 28600 1546 28656
rect 386 18944 442 19000
rect 294 15136 350 15192
rect 294 13776 350 13832
rect 754 24792 810 24848
rect 662 23976 718 24032
rect 478 14864 534 14920
rect 754 23432 810 23488
rect 754 22888 810 22944
rect 754 22344 810 22400
rect 846 21800 902 21856
rect 1122 26968 1178 27024
rect 1306 27784 1362 27840
rect 1306 27240 1362 27296
rect 1306 26696 1362 26752
rect 1214 26424 1270 26480
rect 1214 26288 1270 26344
rect 1122 25608 1178 25664
rect 1122 25472 1178 25528
rect 1214 25336 1270 25392
rect 1398 25744 1454 25800
rect 1674 28600 1730 28656
rect 1674 28484 1730 28520
rect 1674 28464 1676 28484
rect 1676 28464 1728 28484
rect 1728 28464 1730 28484
rect 1766 26424 1822 26480
rect 2042 27648 2098 27704
rect 2226 27920 2282 27976
rect 2778 33768 2834 33824
rect 2594 32544 2650 32600
rect 2502 31184 2558 31240
rect 3428 36474 3484 36476
rect 3508 36474 3564 36476
rect 3588 36474 3644 36476
rect 3668 36474 3724 36476
rect 3428 36422 3474 36474
rect 3474 36422 3484 36474
rect 3508 36422 3538 36474
rect 3538 36422 3550 36474
rect 3550 36422 3564 36474
rect 3588 36422 3602 36474
rect 3602 36422 3614 36474
rect 3614 36422 3644 36474
rect 3668 36422 3678 36474
rect 3678 36422 3724 36474
rect 3428 36420 3484 36422
rect 3508 36420 3564 36422
rect 3588 36420 3644 36422
rect 3668 36420 3724 36422
rect 3428 35386 3484 35388
rect 3508 35386 3564 35388
rect 3588 35386 3644 35388
rect 3668 35386 3724 35388
rect 3428 35334 3474 35386
rect 3474 35334 3484 35386
rect 3508 35334 3538 35386
rect 3538 35334 3550 35386
rect 3550 35334 3564 35386
rect 3588 35334 3602 35386
rect 3602 35334 3614 35386
rect 3614 35334 3644 35386
rect 3668 35334 3678 35386
rect 3678 35334 3724 35386
rect 3428 35332 3484 35334
rect 3508 35332 3564 35334
rect 3588 35332 3644 35334
rect 3668 35332 3724 35334
rect 3790 34448 3846 34504
rect 3428 34298 3484 34300
rect 3508 34298 3564 34300
rect 3588 34298 3644 34300
rect 3668 34298 3724 34300
rect 3428 34246 3474 34298
rect 3474 34246 3484 34298
rect 3508 34246 3538 34298
rect 3538 34246 3550 34298
rect 3550 34246 3564 34298
rect 3588 34246 3602 34298
rect 3602 34246 3614 34298
rect 3614 34246 3644 34298
rect 3668 34246 3678 34298
rect 3678 34246 3724 34298
rect 3428 34244 3484 34246
rect 3508 34244 3564 34246
rect 3588 34244 3644 34246
rect 3668 34244 3724 34246
rect 3330 34040 3386 34096
rect 2778 32680 2834 32736
rect 2778 32544 2834 32600
rect 2502 30368 2558 30424
rect 2410 29008 2466 29064
rect 3698 33532 3700 33552
rect 3700 33532 3752 33552
rect 3752 33532 3754 33552
rect 3698 33496 3754 33532
rect 4158 35980 4160 36000
rect 4160 35980 4212 36000
rect 4212 35980 4214 36000
rect 4158 35944 4214 35980
rect 4066 35536 4122 35592
rect 4066 34040 4122 34096
rect 4250 35128 4306 35184
rect 3428 33210 3484 33212
rect 3508 33210 3564 33212
rect 3588 33210 3644 33212
rect 3668 33210 3724 33212
rect 3428 33158 3474 33210
rect 3474 33158 3484 33210
rect 3508 33158 3538 33210
rect 3538 33158 3550 33210
rect 3550 33158 3564 33210
rect 3588 33158 3602 33210
rect 3602 33158 3614 33210
rect 3614 33158 3644 33210
rect 3668 33158 3678 33210
rect 3678 33158 3724 33210
rect 3428 33156 3484 33158
rect 3508 33156 3564 33158
rect 3588 33156 3644 33158
rect 3668 33156 3724 33158
rect 3882 32836 3938 32872
rect 3882 32816 3884 32836
rect 3884 32816 3936 32836
rect 3936 32816 3938 32836
rect 3514 32292 3570 32328
rect 3514 32272 3516 32292
rect 3516 32272 3568 32292
rect 3568 32272 3570 32292
rect 3428 32122 3484 32124
rect 3508 32122 3564 32124
rect 3588 32122 3644 32124
rect 3668 32122 3724 32124
rect 3428 32070 3474 32122
rect 3474 32070 3484 32122
rect 3508 32070 3538 32122
rect 3538 32070 3550 32122
rect 3550 32070 3564 32122
rect 3588 32070 3602 32122
rect 3602 32070 3614 32122
rect 3614 32070 3644 32122
rect 3668 32070 3678 32122
rect 3678 32070 3724 32122
rect 3428 32068 3484 32070
rect 3508 32068 3564 32070
rect 3588 32068 3644 32070
rect 3668 32068 3724 32070
rect 2962 31320 3018 31376
rect 2870 31048 2926 31104
rect 2778 30504 2834 30560
rect 2778 29824 2834 29880
rect 2778 29280 2834 29336
rect 3790 31592 3846 31648
rect 3428 31034 3484 31036
rect 3508 31034 3564 31036
rect 3588 31034 3644 31036
rect 3668 31034 3724 31036
rect 3428 30982 3474 31034
rect 3474 30982 3484 31034
rect 3508 30982 3538 31034
rect 3538 30982 3550 31034
rect 3550 30982 3564 31034
rect 3588 30982 3602 31034
rect 3602 30982 3614 31034
rect 3614 30982 3644 31034
rect 3668 30982 3678 31034
rect 3678 30982 3724 31034
rect 3428 30980 3484 30982
rect 3508 30980 3564 30982
rect 3588 30980 3644 30982
rect 3668 30980 3724 30982
rect 3606 30776 3662 30832
rect 3422 30232 3478 30288
rect 3428 29946 3484 29948
rect 3508 29946 3564 29948
rect 3588 29946 3644 29948
rect 3668 29946 3724 29948
rect 3428 29894 3474 29946
rect 3474 29894 3484 29946
rect 3508 29894 3538 29946
rect 3538 29894 3550 29946
rect 3550 29894 3564 29946
rect 3588 29894 3602 29946
rect 3602 29894 3614 29946
rect 3614 29894 3644 29946
rect 3668 29894 3678 29946
rect 3678 29894 3724 29946
rect 3428 29892 3484 29894
rect 3508 29892 3564 29894
rect 3588 29892 3644 29894
rect 3668 29892 3724 29894
rect 3330 29688 3386 29744
rect 2962 29416 3018 29472
rect 2594 28620 2650 28656
rect 2594 28600 2596 28620
rect 2596 28600 2648 28620
rect 2648 28600 2650 28620
rect 2410 28212 2466 28248
rect 2410 28192 2412 28212
rect 2412 28192 2464 28212
rect 2464 28192 2466 28212
rect 1950 26016 2006 26072
rect 1490 25472 1546 25528
rect 1306 25064 1362 25120
rect 1858 25200 1914 25256
rect 1306 24520 1362 24576
rect 1214 24248 1270 24304
rect 1306 23704 1362 23760
rect 1306 23568 1362 23624
rect 1490 23432 1546 23488
rect 1398 22616 1454 22672
rect 1214 21936 1270 21992
rect 938 21528 994 21584
rect 1122 21528 1178 21584
rect 754 20440 810 20496
rect 938 21120 994 21176
rect 754 18808 810 18864
rect 754 18536 810 18592
rect 754 18128 810 18184
rect 754 16496 810 16552
rect 662 16360 718 16416
rect 570 14456 626 14512
rect 846 16088 902 16144
rect 846 14728 902 14784
rect 1122 20984 1178 21040
rect 1214 19352 1270 19408
rect 1398 22072 1454 22128
rect 1214 18264 1270 18320
rect 1122 18128 1178 18184
rect 938 14320 994 14376
rect 846 10920 902 10976
rect 846 8336 902 8392
rect 846 8064 902 8120
rect 1030 10648 1086 10704
rect 570 7248 626 7304
rect 570 6568 626 6624
rect 478 2624 534 2680
rect 1030 7520 1086 7576
rect 1766 23976 1822 24032
rect 1674 23160 1730 23216
rect 1582 22616 1638 22672
rect 1674 20984 1730 21040
rect 1674 19216 1730 19272
rect 1490 18400 1546 18456
rect 1582 18264 1638 18320
rect 1490 17992 1546 18048
rect 2410 27104 2466 27160
rect 2134 24928 2190 24984
rect 2134 23740 2136 23760
rect 2136 23740 2188 23760
rect 2188 23740 2190 23760
rect 2134 23704 2190 23740
rect 3054 28192 3110 28248
rect 3054 27940 3110 27976
rect 3054 27920 3056 27940
rect 3056 27920 3108 27940
rect 3108 27920 3110 27940
rect 3054 27784 3110 27840
rect 3238 28872 3294 28928
rect 3238 27512 3294 27568
rect 3422 29280 3478 29336
rect 4158 33360 4214 33416
rect 3974 29960 4030 30016
rect 3974 29688 4030 29744
rect 3428 28858 3484 28860
rect 3508 28858 3564 28860
rect 3588 28858 3644 28860
rect 3668 28858 3724 28860
rect 3428 28806 3474 28858
rect 3474 28806 3484 28858
rect 3508 28806 3538 28858
rect 3538 28806 3550 28858
rect 3550 28806 3564 28858
rect 3588 28806 3602 28858
rect 3602 28806 3614 28858
rect 3614 28806 3644 28858
rect 3668 28806 3678 28858
rect 3678 28806 3724 28858
rect 3428 28804 3484 28806
rect 3508 28804 3564 28806
rect 3588 28804 3644 28806
rect 3668 28804 3724 28806
rect 3790 28056 3846 28112
rect 3428 27770 3484 27772
rect 3508 27770 3564 27772
rect 3588 27770 3644 27772
rect 3668 27770 3724 27772
rect 3428 27718 3474 27770
rect 3474 27718 3484 27770
rect 3508 27718 3538 27770
rect 3538 27718 3550 27770
rect 3550 27718 3564 27770
rect 3588 27718 3602 27770
rect 3602 27718 3614 27770
rect 3614 27718 3644 27770
rect 3668 27718 3678 27770
rect 3678 27718 3724 27770
rect 3428 27716 3484 27718
rect 3508 27716 3564 27718
rect 3588 27716 3644 27718
rect 3668 27716 3724 27718
rect 3698 27376 3754 27432
rect 2502 24676 2558 24712
rect 2502 24656 2504 24676
rect 2504 24656 2556 24676
rect 2556 24656 2558 24676
rect 2502 24248 2558 24304
rect 2134 22072 2190 22128
rect 1950 21292 1952 21312
rect 1952 21292 2004 21312
rect 2004 21292 2006 21312
rect 1950 21256 2006 21292
rect 1950 20576 2006 20632
rect 1858 19896 1914 19952
rect 1766 18944 1822 19000
rect 1582 17448 1638 17504
rect 2686 24928 2742 24984
rect 3146 27104 3202 27160
rect 3330 27240 3386 27296
rect 3054 26324 3056 26344
rect 3056 26324 3108 26344
rect 3108 26324 3110 26344
rect 3054 26288 3110 26324
rect 2870 25336 2926 25392
rect 2226 20032 2282 20088
rect 2134 19760 2190 19816
rect 2042 18692 2098 18728
rect 2042 18672 2044 18692
rect 2044 18672 2096 18692
rect 2096 18672 2098 18692
rect 1582 16904 1638 16960
rect 1766 16904 1822 16960
rect 1674 16768 1730 16824
rect 1766 16632 1822 16688
rect 1766 15952 1822 16008
rect 1674 15816 1730 15872
rect 1582 15272 1638 15328
rect 1398 14456 1454 14512
rect 1306 12960 1362 13016
rect 1490 13640 1546 13696
rect 2134 17176 2190 17232
rect 2318 17312 2374 17368
rect 2226 16360 2282 16416
rect 2042 15952 2098 16008
rect 2134 15544 2190 15600
rect 1950 15000 2006 15056
rect 2042 13912 2098 13968
rect 1766 13096 1822 13152
rect 1674 12280 1730 12336
rect 1582 12008 1638 12064
rect 1398 10920 1454 10976
rect 1306 9560 1362 9616
rect 1214 8472 1270 8528
rect 846 1944 902 2000
rect 1582 9288 1638 9344
rect 1398 7812 1454 7848
rect 1398 7792 1400 7812
rect 1400 7792 1452 7812
rect 1452 7792 1454 7812
rect 1398 7656 1454 7712
rect 1858 11736 1914 11792
rect 1766 9016 1822 9072
rect 1674 8336 1730 8392
rect 1398 5752 1454 5808
rect 1306 5208 1362 5264
rect 1950 11464 2006 11520
rect 2042 11056 2098 11112
rect 2778 22888 2834 22944
rect 2778 20848 2834 20904
rect 2962 23160 3018 23216
rect 2962 22208 3018 22264
rect 3146 25880 3202 25936
rect 3146 23160 3202 23216
rect 2686 19488 2742 19544
rect 2686 19352 2742 19408
rect 2594 18808 2650 18864
rect 2962 20440 3018 20496
rect 2870 18400 2926 18456
rect 3606 27004 3608 27024
rect 3608 27004 3660 27024
rect 3660 27004 3662 27024
rect 3606 26968 3662 27004
rect 3428 26682 3484 26684
rect 3508 26682 3564 26684
rect 3588 26682 3644 26684
rect 3668 26682 3724 26684
rect 3428 26630 3474 26682
rect 3474 26630 3484 26682
rect 3508 26630 3538 26682
rect 3538 26630 3550 26682
rect 3550 26630 3564 26682
rect 3588 26630 3602 26682
rect 3602 26630 3614 26682
rect 3614 26630 3644 26682
rect 3668 26630 3678 26682
rect 3678 26630 3724 26682
rect 3428 26628 3484 26630
rect 3508 26628 3564 26630
rect 3588 26628 3644 26630
rect 3668 26628 3724 26630
rect 3606 26188 3608 26208
rect 3608 26188 3660 26208
rect 3660 26188 3662 26208
rect 3606 26152 3662 26188
rect 3698 25744 3754 25800
rect 3974 27648 4030 27704
rect 3974 27512 4030 27568
rect 4250 33088 4306 33144
rect 4710 41792 4766 41848
rect 4894 40568 4950 40624
rect 4802 39072 4858 39128
rect 4986 38800 5042 38856
rect 4618 36760 4674 36816
rect 4526 36080 4582 36136
rect 4434 33360 4490 33416
rect 4158 29824 4214 29880
rect 4342 32428 4398 32464
rect 4342 32408 4344 32428
rect 4344 32408 4396 32428
rect 4396 32408 4398 32428
rect 4894 34584 4950 34640
rect 5446 41792 5502 41848
rect 5538 41656 5594 41712
rect 5446 41556 5448 41576
rect 5448 41556 5500 41576
rect 5500 41556 5502 41576
rect 5446 41520 5502 41556
rect 6274 43832 6330 43888
rect 5900 43546 5956 43548
rect 5980 43546 6036 43548
rect 6060 43546 6116 43548
rect 6140 43546 6196 43548
rect 5900 43494 5946 43546
rect 5946 43494 5956 43546
rect 5980 43494 6010 43546
rect 6010 43494 6022 43546
rect 6022 43494 6036 43546
rect 6060 43494 6074 43546
rect 6074 43494 6086 43546
rect 6086 43494 6116 43546
rect 6140 43494 6150 43546
rect 6150 43494 6196 43546
rect 5900 43492 5956 43494
rect 5980 43492 6036 43494
rect 6060 43492 6116 43494
rect 6140 43492 6196 43494
rect 5998 43052 6000 43072
rect 6000 43052 6052 43072
rect 6052 43052 6054 43072
rect 5998 43016 6054 43052
rect 5900 42458 5956 42460
rect 5980 42458 6036 42460
rect 6060 42458 6116 42460
rect 6140 42458 6196 42460
rect 5900 42406 5946 42458
rect 5946 42406 5956 42458
rect 5980 42406 6010 42458
rect 6010 42406 6022 42458
rect 6022 42406 6036 42458
rect 6060 42406 6074 42458
rect 6074 42406 6086 42458
rect 6086 42406 6116 42458
rect 6140 42406 6150 42458
rect 6150 42406 6196 42458
rect 5900 42404 5956 42406
rect 5980 42404 6036 42406
rect 6060 42404 6116 42406
rect 6140 42404 6196 42406
rect 5900 41370 5956 41372
rect 5980 41370 6036 41372
rect 6060 41370 6116 41372
rect 6140 41370 6196 41372
rect 5900 41318 5946 41370
rect 5946 41318 5956 41370
rect 5980 41318 6010 41370
rect 6010 41318 6022 41370
rect 6022 41318 6036 41370
rect 6060 41318 6074 41370
rect 6074 41318 6086 41370
rect 6086 41318 6116 41370
rect 6140 41318 6150 41370
rect 6150 41318 6196 41370
rect 5900 41316 5956 41318
rect 5980 41316 6036 41318
rect 6060 41316 6116 41318
rect 6140 41316 6196 41318
rect 6366 41520 6422 41576
rect 5900 40282 5956 40284
rect 5980 40282 6036 40284
rect 6060 40282 6116 40284
rect 6140 40282 6196 40284
rect 5900 40230 5946 40282
rect 5946 40230 5956 40282
rect 5980 40230 6010 40282
rect 6010 40230 6022 40282
rect 6022 40230 6036 40282
rect 6060 40230 6074 40282
rect 6074 40230 6086 40282
rect 6086 40230 6116 40282
rect 6140 40230 6150 40282
rect 6150 40230 6196 40282
rect 5900 40228 5956 40230
rect 5980 40228 6036 40230
rect 6060 40228 6116 40230
rect 6140 40228 6196 40230
rect 5262 38412 5318 38448
rect 5262 38392 5264 38412
rect 5264 38392 5316 38412
rect 5316 38392 5318 38412
rect 5262 37204 5264 37224
rect 5264 37204 5316 37224
rect 5316 37204 5318 37224
rect 5262 37168 5318 37204
rect 5538 37304 5594 37360
rect 5262 33940 5264 33960
rect 5264 33940 5316 33960
rect 5316 33940 5318 33960
rect 5262 33904 5318 33940
rect 4618 32000 4674 32056
rect 4434 30096 4490 30152
rect 4342 29416 4398 29472
rect 4250 26968 4306 27024
rect 3428 25594 3484 25596
rect 3508 25594 3564 25596
rect 3588 25594 3644 25596
rect 3668 25594 3724 25596
rect 3428 25542 3474 25594
rect 3474 25542 3484 25594
rect 3508 25542 3538 25594
rect 3538 25542 3550 25594
rect 3550 25542 3564 25594
rect 3588 25542 3602 25594
rect 3602 25542 3614 25594
rect 3614 25542 3644 25594
rect 3668 25542 3678 25594
rect 3678 25542 3724 25594
rect 3428 25540 3484 25542
rect 3508 25540 3564 25542
rect 3588 25540 3644 25542
rect 3668 25540 3724 25542
rect 3428 24506 3484 24508
rect 3508 24506 3564 24508
rect 3588 24506 3644 24508
rect 3668 24506 3724 24508
rect 3428 24454 3474 24506
rect 3474 24454 3484 24506
rect 3508 24454 3538 24506
rect 3538 24454 3550 24506
rect 3550 24454 3564 24506
rect 3588 24454 3602 24506
rect 3602 24454 3614 24506
rect 3614 24454 3644 24506
rect 3668 24454 3678 24506
rect 3678 24454 3724 24506
rect 3428 24452 3484 24454
rect 3508 24452 3564 24454
rect 3588 24452 3644 24454
rect 3668 24452 3724 24454
rect 4250 25744 4306 25800
rect 4250 25472 4306 25528
rect 4158 25336 4214 25392
rect 3428 23418 3484 23420
rect 3508 23418 3564 23420
rect 3588 23418 3644 23420
rect 3668 23418 3724 23420
rect 3428 23366 3474 23418
rect 3474 23366 3484 23418
rect 3508 23366 3538 23418
rect 3538 23366 3550 23418
rect 3550 23366 3564 23418
rect 3588 23366 3602 23418
rect 3602 23366 3614 23418
rect 3614 23366 3644 23418
rect 3668 23366 3678 23418
rect 3678 23366 3724 23418
rect 3428 23364 3484 23366
rect 3508 23364 3564 23366
rect 3588 23364 3644 23366
rect 3668 23364 3724 23366
rect 3330 23024 3386 23080
rect 4158 24384 4214 24440
rect 4066 23296 4122 23352
rect 3974 23160 4030 23216
rect 3606 22480 3662 22536
rect 3974 22772 4030 22808
rect 3974 22752 3976 22772
rect 3976 22752 4028 22772
rect 4028 22752 4030 22772
rect 3428 22330 3484 22332
rect 3508 22330 3564 22332
rect 3588 22330 3644 22332
rect 3668 22330 3724 22332
rect 3428 22278 3474 22330
rect 3474 22278 3484 22330
rect 3508 22278 3538 22330
rect 3538 22278 3550 22330
rect 3550 22278 3564 22330
rect 3588 22278 3602 22330
rect 3602 22278 3614 22330
rect 3614 22278 3644 22330
rect 3668 22278 3678 22330
rect 3678 22278 3724 22330
rect 3428 22276 3484 22278
rect 3508 22276 3564 22278
rect 3588 22276 3644 22278
rect 3668 22276 3724 22278
rect 3238 21664 3294 21720
rect 3422 21528 3478 21584
rect 3606 21936 3662 21992
rect 3974 22072 4030 22128
rect 4158 22344 4214 22400
rect 3428 21242 3484 21244
rect 3508 21242 3564 21244
rect 3588 21242 3644 21244
rect 3668 21242 3724 21244
rect 3428 21190 3474 21242
rect 3474 21190 3484 21242
rect 3508 21190 3538 21242
rect 3538 21190 3550 21242
rect 3550 21190 3564 21242
rect 3588 21190 3602 21242
rect 3602 21190 3614 21242
rect 3614 21190 3644 21242
rect 3668 21190 3678 21242
rect 3678 21190 3724 21242
rect 3428 21188 3484 21190
rect 3508 21188 3564 21190
rect 3588 21188 3644 21190
rect 3668 21188 3724 21190
rect 3330 20848 3386 20904
rect 3238 20168 3294 20224
rect 3238 20032 3294 20088
rect 3514 20304 3570 20360
rect 3698 20304 3754 20360
rect 3428 20154 3484 20156
rect 3508 20154 3564 20156
rect 3588 20154 3644 20156
rect 3668 20154 3724 20156
rect 3428 20102 3474 20154
rect 3474 20102 3484 20154
rect 3508 20102 3538 20154
rect 3538 20102 3550 20154
rect 3550 20102 3564 20154
rect 3588 20102 3602 20154
rect 3602 20102 3614 20154
rect 3614 20102 3644 20154
rect 3668 20102 3678 20154
rect 3678 20102 3724 20154
rect 3428 20100 3484 20102
rect 3508 20100 3564 20102
rect 3588 20100 3644 20102
rect 3668 20100 3724 20102
rect 3146 19624 3202 19680
rect 3054 18536 3110 18592
rect 3054 18400 3110 18456
rect 2686 17720 2742 17776
rect 3330 19352 3386 19408
rect 3428 19066 3484 19068
rect 3508 19066 3564 19068
rect 3588 19066 3644 19068
rect 3668 19066 3724 19068
rect 3428 19014 3474 19066
rect 3474 19014 3484 19066
rect 3508 19014 3538 19066
rect 3538 19014 3550 19066
rect 3550 19014 3564 19066
rect 3588 19014 3602 19066
rect 3602 19014 3614 19066
rect 3614 19014 3644 19066
rect 3668 19014 3678 19066
rect 3678 19014 3724 19066
rect 3428 19012 3484 19014
rect 3508 19012 3564 19014
rect 3588 19012 3644 19014
rect 3668 19012 3724 19014
rect 4066 21528 4122 21584
rect 3974 21120 4030 21176
rect 3606 18400 3662 18456
rect 4802 32136 4858 32192
rect 4802 30232 4858 30288
rect 4618 28328 4674 28384
rect 4802 29044 4804 29064
rect 4804 29044 4856 29064
rect 4856 29044 4858 29064
rect 4802 29008 4858 29044
rect 5170 32952 5226 33008
rect 5170 31456 5226 31512
rect 5900 39194 5956 39196
rect 5980 39194 6036 39196
rect 6060 39194 6116 39196
rect 6140 39194 6196 39196
rect 5900 39142 5946 39194
rect 5946 39142 5956 39194
rect 5980 39142 6010 39194
rect 6010 39142 6022 39194
rect 6022 39142 6036 39194
rect 6060 39142 6074 39194
rect 6074 39142 6086 39194
rect 6086 39142 6116 39194
rect 6140 39142 6150 39194
rect 6150 39142 6196 39194
rect 5900 39140 5956 39142
rect 5980 39140 6036 39142
rect 6060 39140 6116 39142
rect 6140 39140 6196 39142
rect 5722 36488 5778 36544
rect 5630 34448 5686 34504
rect 5446 32544 5502 32600
rect 5078 30232 5134 30288
rect 5354 30368 5410 30424
rect 5538 30232 5594 30288
rect 5078 28192 5134 28248
rect 4710 26832 4766 26888
rect 5446 30096 5502 30152
rect 5446 29280 5502 29336
rect 5538 29144 5594 29200
rect 4986 26288 5042 26344
rect 4618 24248 4674 24304
rect 4526 22888 4582 22944
rect 4710 22344 4766 22400
rect 5354 26852 5410 26888
rect 5354 26832 5356 26852
rect 5356 26832 5408 26852
rect 5408 26832 5410 26852
rect 5170 25900 5226 25936
rect 5170 25880 5172 25900
rect 5172 25880 5224 25900
rect 5224 25880 5226 25900
rect 5262 25200 5318 25256
rect 5900 38106 5956 38108
rect 5980 38106 6036 38108
rect 6060 38106 6116 38108
rect 6140 38106 6196 38108
rect 5900 38054 5946 38106
rect 5946 38054 5956 38106
rect 5980 38054 6010 38106
rect 6010 38054 6022 38106
rect 6022 38054 6036 38106
rect 6060 38054 6074 38106
rect 6074 38054 6086 38106
rect 6086 38054 6116 38106
rect 6140 38054 6150 38106
rect 6150 38054 6196 38106
rect 5900 38052 5956 38054
rect 5980 38052 6036 38054
rect 6060 38052 6116 38054
rect 6140 38052 6196 38054
rect 6458 37848 6514 37904
rect 6366 37712 6422 37768
rect 5900 37018 5956 37020
rect 5980 37018 6036 37020
rect 6060 37018 6116 37020
rect 6140 37018 6196 37020
rect 5900 36966 5946 37018
rect 5946 36966 5956 37018
rect 5980 36966 6010 37018
rect 6010 36966 6022 37018
rect 6022 36966 6036 37018
rect 6060 36966 6074 37018
rect 6074 36966 6086 37018
rect 6086 36966 6116 37018
rect 6140 36966 6150 37018
rect 6150 36966 6196 37018
rect 5900 36964 5956 36966
rect 5980 36964 6036 36966
rect 6060 36964 6116 36966
rect 6140 36964 6196 36966
rect 5900 35930 5956 35932
rect 5980 35930 6036 35932
rect 6060 35930 6116 35932
rect 6140 35930 6196 35932
rect 5900 35878 5946 35930
rect 5946 35878 5956 35930
rect 5980 35878 6010 35930
rect 6010 35878 6022 35930
rect 6022 35878 6036 35930
rect 6060 35878 6074 35930
rect 6074 35878 6086 35930
rect 6086 35878 6116 35930
rect 6140 35878 6150 35930
rect 6150 35878 6196 35930
rect 5900 35876 5956 35878
rect 5980 35876 6036 35878
rect 6060 35876 6116 35878
rect 6140 35876 6196 35878
rect 5906 35128 5962 35184
rect 5900 34842 5956 34844
rect 5980 34842 6036 34844
rect 6060 34842 6116 34844
rect 6140 34842 6196 34844
rect 5900 34790 5946 34842
rect 5946 34790 5956 34842
rect 5980 34790 6010 34842
rect 6010 34790 6022 34842
rect 6022 34790 6036 34842
rect 6060 34790 6074 34842
rect 6074 34790 6086 34842
rect 6086 34790 6116 34842
rect 6140 34790 6150 34842
rect 6150 34790 6196 34842
rect 5900 34788 5956 34790
rect 5980 34788 6036 34790
rect 6060 34788 6116 34790
rect 6140 34788 6196 34790
rect 6734 37304 6790 37360
rect 5900 33754 5956 33756
rect 5980 33754 6036 33756
rect 6060 33754 6116 33756
rect 6140 33754 6196 33756
rect 5900 33702 5946 33754
rect 5946 33702 5956 33754
rect 5980 33702 6010 33754
rect 6010 33702 6022 33754
rect 6022 33702 6036 33754
rect 6060 33702 6074 33754
rect 6074 33702 6086 33754
rect 6086 33702 6116 33754
rect 6140 33702 6150 33754
rect 6150 33702 6196 33754
rect 5900 33700 5956 33702
rect 5980 33700 6036 33702
rect 6060 33700 6116 33702
rect 6140 33700 6196 33702
rect 5900 32666 5956 32668
rect 5980 32666 6036 32668
rect 6060 32666 6116 32668
rect 6140 32666 6196 32668
rect 5900 32614 5946 32666
rect 5946 32614 5956 32666
rect 5980 32614 6010 32666
rect 6010 32614 6022 32666
rect 6022 32614 6036 32666
rect 6060 32614 6074 32666
rect 6074 32614 6086 32666
rect 6086 32614 6116 32666
rect 6140 32614 6150 32666
rect 6150 32614 6196 32666
rect 5900 32612 5956 32614
rect 5980 32612 6036 32614
rect 6060 32612 6116 32614
rect 6140 32612 6196 32614
rect 6550 34176 6606 34232
rect 6274 32000 6330 32056
rect 5900 31578 5956 31580
rect 5980 31578 6036 31580
rect 6060 31578 6116 31580
rect 6140 31578 6196 31580
rect 5900 31526 5946 31578
rect 5946 31526 5956 31578
rect 5980 31526 6010 31578
rect 6010 31526 6022 31578
rect 6022 31526 6036 31578
rect 6060 31526 6074 31578
rect 6074 31526 6086 31578
rect 6086 31526 6116 31578
rect 6140 31526 6150 31578
rect 6150 31526 6196 31578
rect 5900 31524 5956 31526
rect 5980 31524 6036 31526
rect 6060 31524 6116 31526
rect 6140 31524 6196 31526
rect 6274 31320 6330 31376
rect 5814 31048 5870 31104
rect 5900 30490 5956 30492
rect 5980 30490 6036 30492
rect 6060 30490 6116 30492
rect 6140 30490 6196 30492
rect 5900 30438 5946 30490
rect 5946 30438 5956 30490
rect 5980 30438 6010 30490
rect 6010 30438 6022 30490
rect 6022 30438 6036 30490
rect 6060 30438 6074 30490
rect 6074 30438 6086 30490
rect 6086 30438 6116 30490
rect 6140 30438 6150 30490
rect 6150 30438 6196 30490
rect 5900 30436 5956 30438
rect 5980 30436 6036 30438
rect 6060 30436 6116 30438
rect 6140 30436 6196 30438
rect 6734 33768 6790 33824
rect 6274 29416 6330 29472
rect 5900 29402 5956 29404
rect 5980 29402 6036 29404
rect 6060 29402 6116 29404
rect 6140 29402 6196 29404
rect 5900 29350 5946 29402
rect 5946 29350 5956 29402
rect 5980 29350 6010 29402
rect 6010 29350 6022 29402
rect 6022 29350 6036 29402
rect 6060 29350 6074 29402
rect 6074 29350 6086 29402
rect 6086 29350 6116 29402
rect 6140 29350 6150 29402
rect 6150 29350 6196 29402
rect 5900 29348 5956 29350
rect 5980 29348 6036 29350
rect 6060 29348 6116 29350
rect 6140 29348 6196 29350
rect 5900 28314 5956 28316
rect 5980 28314 6036 28316
rect 6060 28314 6116 28316
rect 6140 28314 6196 28316
rect 5900 28262 5946 28314
rect 5946 28262 5956 28314
rect 5980 28262 6010 28314
rect 6010 28262 6022 28314
rect 6022 28262 6036 28314
rect 6060 28262 6074 28314
rect 6074 28262 6086 28314
rect 6086 28262 6116 28314
rect 6140 28262 6150 28314
rect 6150 28262 6196 28314
rect 5900 28260 5956 28262
rect 5980 28260 6036 28262
rect 6060 28260 6116 28262
rect 6140 28260 6196 28262
rect 5906 28056 5962 28112
rect 5900 27226 5956 27228
rect 5980 27226 6036 27228
rect 6060 27226 6116 27228
rect 6140 27226 6196 27228
rect 5900 27174 5946 27226
rect 5946 27174 5956 27226
rect 5980 27174 6010 27226
rect 6010 27174 6022 27226
rect 6022 27174 6036 27226
rect 6060 27174 6074 27226
rect 6074 27174 6086 27226
rect 6086 27174 6116 27226
rect 6140 27174 6150 27226
rect 6150 27174 6196 27226
rect 5900 27172 5956 27174
rect 5980 27172 6036 27174
rect 6060 27172 6116 27174
rect 6140 27172 6196 27174
rect 6550 30232 6606 30288
rect 7194 40568 7250 40624
rect 8373 43002 8429 43004
rect 8453 43002 8509 43004
rect 8533 43002 8589 43004
rect 8613 43002 8669 43004
rect 8373 42950 8419 43002
rect 8419 42950 8429 43002
rect 8453 42950 8483 43002
rect 8483 42950 8495 43002
rect 8495 42950 8509 43002
rect 8533 42950 8547 43002
rect 8547 42950 8559 43002
rect 8559 42950 8589 43002
rect 8613 42950 8623 43002
rect 8623 42950 8669 43002
rect 8373 42948 8429 42950
rect 8453 42948 8509 42950
rect 8533 42948 8589 42950
rect 8613 42948 8669 42950
rect 8373 41914 8429 41916
rect 8453 41914 8509 41916
rect 8533 41914 8589 41916
rect 8613 41914 8669 41916
rect 8373 41862 8419 41914
rect 8419 41862 8429 41914
rect 8453 41862 8483 41914
rect 8483 41862 8495 41914
rect 8495 41862 8509 41914
rect 8533 41862 8547 41914
rect 8547 41862 8559 41914
rect 8559 41862 8589 41914
rect 8613 41862 8623 41914
rect 8623 41862 8669 41914
rect 8373 41860 8429 41862
rect 8453 41860 8509 41862
rect 8533 41860 8589 41862
rect 8613 41860 8669 41862
rect 8850 42472 8906 42528
rect 8850 42064 8906 42120
rect 7470 41520 7526 41576
rect 7378 37984 7434 38040
rect 7286 36624 7342 36680
rect 7286 34992 7342 35048
rect 7102 34176 7158 34232
rect 7010 31864 7066 31920
rect 7010 31592 7066 31648
rect 6918 31184 6974 31240
rect 7102 31204 7158 31240
rect 7102 31184 7104 31204
rect 7104 31184 7156 31204
rect 7156 31184 7158 31204
rect 8373 40826 8429 40828
rect 8453 40826 8509 40828
rect 8533 40826 8589 40828
rect 8613 40826 8669 40828
rect 8373 40774 8419 40826
rect 8419 40774 8429 40826
rect 8453 40774 8483 40826
rect 8483 40774 8495 40826
rect 8495 40774 8509 40826
rect 8533 40774 8547 40826
rect 8547 40774 8559 40826
rect 8559 40774 8589 40826
rect 8613 40774 8623 40826
rect 8623 40774 8669 40826
rect 8373 40772 8429 40774
rect 8453 40772 8509 40774
rect 8533 40772 8589 40774
rect 8613 40772 8669 40774
rect 7930 40024 7986 40080
rect 7838 38936 7894 38992
rect 8373 39738 8429 39740
rect 8453 39738 8509 39740
rect 8533 39738 8589 39740
rect 8613 39738 8669 39740
rect 8373 39686 8419 39738
rect 8419 39686 8429 39738
rect 8453 39686 8483 39738
rect 8483 39686 8495 39738
rect 8495 39686 8509 39738
rect 8533 39686 8547 39738
rect 8547 39686 8559 39738
rect 8559 39686 8589 39738
rect 8613 39686 8623 39738
rect 8623 39686 8669 39738
rect 8373 39684 8429 39686
rect 8453 39684 8509 39686
rect 8533 39684 8589 39686
rect 8613 39684 8669 39686
rect 7746 35808 7802 35864
rect 8373 38650 8429 38652
rect 8453 38650 8509 38652
rect 8533 38650 8589 38652
rect 8613 38650 8669 38652
rect 8373 38598 8419 38650
rect 8419 38598 8429 38650
rect 8453 38598 8483 38650
rect 8483 38598 8495 38650
rect 8495 38598 8509 38650
rect 8533 38598 8547 38650
rect 8547 38598 8559 38650
rect 8559 38598 8589 38650
rect 8613 38598 8623 38650
rect 8623 38598 8669 38650
rect 8373 38596 8429 38598
rect 8453 38596 8509 38598
rect 8533 38596 8589 38598
rect 8613 38596 8669 38598
rect 8758 37848 8814 37904
rect 8373 37562 8429 37564
rect 8453 37562 8509 37564
rect 8533 37562 8589 37564
rect 8613 37562 8669 37564
rect 8373 37510 8419 37562
rect 8419 37510 8429 37562
rect 8453 37510 8483 37562
rect 8483 37510 8495 37562
rect 8495 37510 8509 37562
rect 8533 37510 8547 37562
rect 8547 37510 8559 37562
rect 8559 37510 8589 37562
rect 8613 37510 8623 37562
rect 8623 37510 8669 37562
rect 8373 37508 8429 37510
rect 8453 37508 8509 37510
rect 8533 37508 8589 37510
rect 8613 37508 8669 37510
rect 8206 36488 8262 36544
rect 8373 36474 8429 36476
rect 8453 36474 8509 36476
rect 8533 36474 8589 36476
rect 8613 36474 8669 36476
rect 8373 36422 8419 36474
rect 8419 36422 8429 36474
rect 8453 36422 8483 36474
rect 8483 36422 8495 36474
rect 8495 36422 8509 36474
rect 8533 36422 8547 36474
rect 8547 36422 8559 36474
rect 8559 36422 8589 36474
rect 8613 36422 8623 36474
rect 8623 36422 8669 36474
rect 8373 36420 8429 36422
rect 8453 36420 8509 36422
rect 8533 36420 8589 36422
rect 8613 36420 8669 36422
rect 8373 35386 8429 35388
rect 8453 35386 8509 35388
rect 8533 35386 8589 35388
rect 8613 35386 8669 35388
rect 8373 35334 8419 35386
rect 8419 35334 8429 35386
rect 8453 35334 8483 35386
rect 8483 35334 8495 35386
rect 8495 35334 8509 35386
rect 8533 35334 8547 35386
rect 8547 35334 8559 35386
rect 8559 35334 8589 35386
rect 8613 35334 8623 35386
rect 8623 35334 8669 35386
rect 8373 35332 8429 35334
rect 8453 35332 8509 35334
rect 8533 35332 8589 35334
rect 8613 35332 8669 35334
rect 8022 34584 8078 34640
rect 7930 34176 7986 34232
rect 8206 34584 8262 34640
rect 8373 34298 8429 34300
rect 8453 34298 8509 34300
rect 8533 34298 8589 34300
rect 8613 34298 8669 34300
rect 8373 34246 8419 34298
rect 8419 34246 8429 34298
rect 8453 34246 8483 34298
rect 8483 34246 8495 34298
rect 8495 34246 8509 34298
rect 8533 34246 8547 34298
rect 8547 34246 8559 34298
rect 8559 34246 8589 34298
rect 8613 34246 8623 34298
rect 8623 34246 8669 34298
rect 8373 34244 8429 34246
rect 8453 34244 8509 34246
rect 8533 34244 8589 34246
rect 8613 34244 8669 34246
rect 7194 30660 7250 30696
rect 7194 30640 7196 30660
rect 7196 30640 7248 30660
rect 7248 30640 7250 30660
rect 6458 28736 6514 28792
rect 6366 27648 6422 27704
rect 6274 26152 6330 26208
rect 5900 26138 5956 26140
rect 5980 26138 6036 26140
rect 6060 26138 6116 26140
rect 6140 26138 6196 26140
rect 5900 26086 5946 26138
rect 5946 26086 5956 26138
rect 5980 26086 6010 26138
rect 6010 26086 6022 26138
rect 6022 26086 6036 26138
rect 6060 26086 6074 26138
rect 6074 26086 6086 26138
rect 6086 26086 6116 26138
rect 6140 26086 6150 26138
rect 6150 26086 6196 26138
rect 5900 26084 5956 26086
rect 5980 26084 6036 26086
rect 6060 26084 6116 26086
rect 6140 26084 6196 26086
rect 5170 23976 5226 24032
rect 5170 23840 5226 23896
rect 5538 24792 5594 24848
rect 5538 24248 5594 24304
rect 4526 21664 4582 21720
rect 4710 21256 4766 21312
rect 4158 19760 4214 19816
rect 3790 18128 3846 18184
rect 3428 17978 3484 17980
rect 3508 17978 3564 17980
rect 3588 17978 3644 17980
rect 3668 17978 3724 17980
rect 3428 17926 3474 17978
rect 3474 17926 3484 17978
rect 3508 17926 3538 17978
rect 3538 17926 3550 17978
rect 3550 17926 3564 17978
rect 3588 17926 3602 17978
rect 3602 17926 3614 17978
rect 3614 17926 3644 17978
rect 3668 17926 3678 17978
rect 3678 17926 3724 17978
rect 3428 17924 3484 17926
rect 3508 17924 3564 17926
rect 3588 17924 3644 17926
rect 3668 17924 3724 17926
rect 2594 16904 2650 16960
rect 2502 16496 2558 16552
rect 2686 16632 2742 16688
rect 3054 16768 3110 16824
rect 2870 16088 2926 16144
rect 2686 14592 2742 14648
rect 2594 14048 2650 14104
rect 2502 13232 2558 13288
rect 2594 12144 2650 12200
rect 2226 10784 2282 10840
rect 2502 11092 2504 11112
rect 2504 11092 2556 11112
rect 2556 11092 2558 11112
rect 2502 11056 2558 11092
rect 2226 10512 2282 10568
rect 2318 10376 2374 10432
rect 2042 8608 2098 8664
rect 1858 7812 1914 7848
rect 1858 7792 1860 7812
rect 1860 7792 1912 7812
rect 1912 7792 1914 7812
rect 1858 6296 1914 6352
rect 2042 7384 2098 7440
rect 2502 10920 2558 10976
rect 2594 10240 2650 10296
rect 2318 8744 2374 8800
rect 2226 8472 2282 8528
rect 2226 6976 2282 7032
rect 2226 6704 2282 6760
rect 1950 5616 2006 5672
rect 2410 8336 2466 8392
rect 2318 6160 2374 6216
rect 3514 17720 3570 17776
rect 3428 16890 3484 16892
rect 3508 16890 3564 16892
rect 3588 16890 3644 16892
rect 3668 16890 3724 16892
rect 3428 16838 3474 16890
rect 3474 16838 3484 16890
rect 3508 16838 3538 16890
rect 3538 16838 3550 16890
rect 3550 16838 3564 16890
rect 3588 16838 3602 16890
rect 3602 16838 3614 16890
rect 3614 16838 3644 16890
rect 3668 16838 3678 16890
rect 3678 16838 3724 16890
rect 3428 16836 3484 16838
rect 3508 16836 3564 16838
rect 3588 16836 3644 16838
rect 3668 16836 3724 16838
rect 3422 16496 3478 16552
rect 3790 16360 3846 16416
rect 3974 16532 3976 16552
rect 3976 16532 4028 16552
rect 4028 16532 4030 16552
rect 3974 16496 4030 16532
rect 3882 15852 3884 15872
rect 3884 15852 3936 15872
rect 3936 15852 3938 15872
rect 3428 15802 3484 15804
rect 3508 15802 3564 15804
rect 3588 15802 3644 15804
rect 3668 15802 3724 15804
rect 3428 15750 3474 15802
rect 3474 15750 3484 15802
rect 3508 15750 3538 15802
rect 3538 15750 3550 15802
rect 3550 15750 3564 15802
rect 3588 15750 3602 15802
rect 3602 15750 3614 15802
rect 3614 15750 3644 15802
rect 3668 15750 3678 15802
rect 3678 15750 3724 15802
rect 3428 15748 3484 15750
rect 3508 15748 3564 15750
rect 3588 15748 3644 15750
rect 3668 15748 3724 15750
rect 3882 15816 3938 15852
rect 3330 14864 3386 14920
rect 3428 14714 3484 14716
rect 3508 14714 3564 14716
rect 3588 14714 3644 14716
rect 3668 14714 3724 14716
rect 3428 14662 3474 14714
rect 3474 14662 3484 14714
rect 3508 14662 3538 14714
rect 3538 14662 3550 14714
rect 3550 14662 3564 14714
rect 3588 14662 3602 14714
rect 3602 14662 3614 14714
rect 3614 14662 3644 14714
rect 3668 14662 3678 14714
rect 3678 14662 3724 14714
rect 3428 14660 3484 14662
rect 3508 14660 3564 14662
rect 3588 14660 3644 14662
rect 3668 14660 3724 14662
rect 3428 13626 3484 13628
rect 3508 13626 3564 13628
rect 3588 13626 3644 13628
rect 3668 13626 3724 13628
rect 3428 13574 3474 13626
rect 3474 13574 3484 13626
rect 3508 13574 3538 13626
rect 3538 13574 3550 13626
rect 3550 13574 3564 13626
rect 3588 13574 3602 13626
rect 3602 13574 3614 13626
rect 3614 13574 3644 13626
rect 3668 13574 3678 13626
rect 3678 13574 3724 13626
rect 3428 13572 3484 13574
rect 3508 13572 3564 13574
rect 3588 13572 3644 13574
rect 3668 13572 3724 13574
rect 2870 12008 2926 12064
rect 3238 12960 3294 13016
rect 4250 18128 4306 18184
rect 4250 17856 4306 17912
rect 4158 16768 4214 16824
rect 4066 14048 4122 14104
rect 4342 17040 4398 17096
rect 4342 16224 4398 16280
rect 3882 13776 3938 13832
rect 3974 13368 4030 13424
rect 3974 13232 4030 13288
rect 4066 12824 4122 12880
rect 3882 12552 3938 12608
rect 3428 12538 3484 12540
rect 3508 12538 3564 12540
rect 3588 12538 3644 12540
rect 3668 12538 3724 12540
rect 3428 12486 3474 12538
rect 3474 12486 3484 12538
rect 3508 12486 3538 12538
rect 3538 12486 3550 12538
rect 3550 12486 3564 12538
rect 3588 12486 3602 12538
rect 3602 12486 3614 12538
rect 3614 12486 3644 12538
rect 3668 12486 3678 12538
rect 3678 12486 3724 12538
rect 3428 12484 3484 12486
rect 3508 12484 3564 12486
rect 3588 12484 3644 12486
rect 3668 12484 3724 12486
rect 3790 12382 3846 12438
rect 3428 11450 3484 11452
rect 3508 11450 3564 11452
rect 3588 11450 3644 11452
rect 3668 11450 3724 11452
rect 3428 11398 3474 11450
rect 3474 11398 3484 11450
rect 3508 11398 3538 11450
rect 3538 11398 3550 11450
rect 3550 11398 3564 11450
rect 3588 11398 3602 11450
rect 3602 11398 3614 11450
rect 3614 11398 3644 11450
rect 3668 11398 3678 11450
rect 3678 11398 3724 11450
rect 3428 11396 3484 11398
rect 3508 11396 3564 11398
rect 3588 11396 3644 11398
rect 3668 11396 3724 11398
rect 2778 9560 2834 9616
rect 2962 8336 3018 8392
rect 2686 7384 2742 7440
rect 2686 7248 2742 7304
rect 3428 10362 3484 10364
rect 3508 10362 3564 10364
rect 3588 10362 3644 10364
rect 3668 10362 3724 10364
rect 3428 10310 3474 10362
rect 3474 10310 3484 10362
rect 3508 10310 3538 10362
rect 3538 10310 3550 10362
rect 3550 10310 3564 10362
rect 3588 10310 3602 10362
rect 3602 10310 3614 10362
rect 3614 10310 3644 10362
rect 3668 10310 3678 10362
rect 3678 10310 3724 10362
rect 3428 10308 3484 10310
rect 3508 10308 3564 10310
rect 3588 10308 3644 10310
rect 3668 10308 3724 10310
rect 3330 9560 3386 9616
rect 3238 9288 3294 9344
rect 3146 8200 3202 8256
rect 3428 9274 3484 9276
rect 3508 9274 3564 9276
rect 3588 9274 3644 9276
rect 3668 9274 3724 9276
rect 3428 9222 3474 9274
rect 3474 9222 3484 9274
rect 3508 9222 3538 9274
rect 3538 9222 3550 9274
rect 3550 9222 3564 9274
rect 3588 9222 3602 9274
rect 3602 9222 3614 9274
rect 3614 9222 3644 9274
rect 3668 9222 3678 9274
rect 3678 9222 3724 9274
rect 3428 9220 3484 9222
rect 3508 9220 3564 9222
rect 3588 9220 3644 9222
rect 3668 9220 3724 9222
rect 3422 8492 3478 8528
rect 3422 8472 3424 8492
rect 3424 8472 3476 8492
rect 3476 8472 3478 8492
rect 3428 8186 3484 8188
rect 3508 8186 3564 8188
rect 3588 8186 3644 8188
rect 3668 8186 3724 8188
rect 3428 8134 3474 8186
rect 3474 8134 3484 8186
rect 3508 8134 3538 8186
rect 3538 8134 3550 8186
rect 3550 8134 3564 8186
rect 3588 8134 3602 8186
rect 3602 8134 3614 8186
rect 3614 8134 3644 8186
rect 3668 8134 3678 8186
rect 3678 8134 3724 8186
rect 3428 8132 3484 8134
rect 3508 8132 3564 8134
rect 3588 8132 3644 8134
rect 3668 8132 3724 8134
rect 2410 5344 2466 5400
rect 1858 2624 1914 2680
rect 386 720 442 776
rect 2962 7248 3018 7304
rect 2962 7112 3018 7168
rect 2870 5888 2926 5944
rect 2870 5208 2926 5264
rect 3698 7792 3754 7848
rect 3238 6976 3294 7032
rect 3146 6024 3202 6080
rect 3054 5752 3110 5808
rect 3054 5480 3110 5536
rect 2594 3576 2650 3632
rect 2410 3440 2466 3496
rect 2502 2624 2558 2680
rect 4066 11736 4122 11792
rect 4158 11464 4214 11520
rect 4066 11192 4122 11248
rect 3974 10648 4030 10704
rect 3974 10240 4030 10296
rect 4986 20576 5042 20632
rect 5078 20168 5134 20224
rect 4986 19896 5042 19952
rect 5262 20032 5318 20088
rect 5262 19624 5318 19680
rect 5078 17448 5134 17504
rect 4894 16360 4950 16416
rect 4618 14864 4674 14920
rect 4710 14476 4766 14512
rect 4710 14456 4712 14476
rect 4712 14456 4764 14476
rect 4764 14456 4766 14476
rect 4434 13932 4490 13968
rect 4434 13912 4436 13932
rect 4436 13912 4488 13932
rect 4488 13912 4490 13932
rect 4802 14320 4858 14376
rect 4434 12044 4436 12064
rect 4436 12044 4488 12064
rect 4488 12044 4490 12064
rect 4434 12008 4490 12044
rect 4986 13268 4988 13288
rect 4988 13268 5040 13288
rect 5040 13268 5042 13288
rect 4986 13232 5042 13268
rect 4986 12960 5042 13016
rect 4986 12552 5042 12608
rect 4894 12280 4950 12336
rect 4526 11464 4582 11520
rect 4526 11192 4582 11248
rect 4894 11464 4950 11520
rect 4894 11328 4950 11384
rect 4526 10920 4582 10976
rect 4802 11056 4858 11112
rect 4894 10920 4950 10976
rect 5900 25050 5956 25052
rect 5980 25050 6036 25052
rect 6060 25050 6116 25052
rect 6140 25050 6196 25052
rect 5900 24998 5946 25050
rect 5946 24998 5956 25050
rect 5980 24998 6010 25050
rect 6010 24998 6022 25050
rect 6022 24998 6036 25050
rect 6060 24998 6074 25050
rect 6074 24998 6086 25050
rect 6086 24998 6116 25050
rect 6140 24998 6150 25050
rect 6150 24998 6196 25050
rect 5900 24996 5956 24998
rect 5980 24996 6036 24998
rect 6060 24996 6116 24998
rect 6140 24996 6196 24998
rect 5900 23962 5956 23964
rect 5980 23962 6036 23964
rect 6060 23962 6116 23964
rect 6140 23962 6196 23964
rect 5900 23910 5946 23962
rect 5946 23910 5956 23962
rect 5980 23910 6010 23962
rect 6010 23910 6022 23962
rect 6022 23910 6036 23962
rect 6060 23910 6074 23962
rect 6074 23910 6086 23962
rect 6086 23910 6116 23962
rect 6140 23910 6150 23962
rect 6150 23910 6196 23962
rect 5900 23908 5956 23910
rect 5980 23908 6036 23910
rect 6060 23908 6116 23910
rect 6140 23908 6196 23910
rect 6458 24520 6514 24576
rect 5998 23432 6054 23488
rect 6274 22888 6330 22944
rect 5900 22874 5956 22876
rect 5980 22874 6036 22876
rect 6060 22874 6116 22876
rect 6140 22874 6196 22876
rect 5900 22822 5946 22874
rect 5946 22822 5956 22874
rect 5980 22822 6010 22874
rect 6010 22822 6022 22874
rect 6022 22822 6036 22874
rect 6060 22822 6074 22874
rect 6074 22822 6086 22874
rect 6086 22822 6116 22874
rect 6140 22822 6150 22874
rect 6150 22822 6196 22874
rect 5900 22820 5956 22822
rect 5980 22820 6036 22822
rect 6060 22820 6116 22822
rect 6140 22820 6196 22822
rect 5900 21786 5956 21788
rect 5980 21786 6036 21788
rect 6060 21786 6116 21788
rect 6140 21786 6196 21788
rect 5900 21734 5946 21786
rect 5946 21734 5956 21786
rect 5980 21734 6010 21786
rect 6010 21734 6022 21786
rect 6022 21734 6036 21786
rect 6060 21734 6074 21786
rect 6074 21734 6086 21786
rect 6086 21734 6116 21786
rect 6140 21734 6150 21786
rect 6150 21734 6196 21786
rect 5900 21732 5956 21734
rect 5980 21732 6036 21734
rect 6060 21732 6116 21734
rect 6140 21732 6196 21734
rect 5446 20440 5502 20496
rect 5906 21256 5962 21312
rect 5722 20712 5778 20768
rect 5900 20698 5956 20700
rect 5980 20698 6036 20700
rect 6060 20698 6116 20700
rect 6140 20698 6196 20700
rect 5900 20646 5946 20698
rect 5946 20646 5956 20698
rect 5980 20646 6010 20698
rect 6010 20646 6022 20698
rect 6022 20646 6036 20698
rect 6060 20646 6074 20698
rect 6074 20646 6086 20698
rect 6086 20646 6116 20698
rect 6140 20646 6150 20698
rect 6150 20646 6196 20698
rect 5900 20644 5956 20646
rect 5980 20644 6036 20646
rect 6060 20644 6116 20646
rect 6140 20644 6196 20646
rect 5538 19488 5594 19544
rect 5446 17720 5502 17776
rect 5446 16088 5502 16144
rect 5446 15544 5502 15600
rect 5538 15272 5594 15328
rect 5170 11056 5226 11112
rect 5354 12008 5410 12064
rect 4066 9696 4122 9752
rect 4158 9596 4160 9616
rect 4160 9596 4212 9616
rect 4212 9596 4214 9616
rect 4158 9560 4214 9596
rect 4066 9152 4122 9208
rect 3974 9016 4030 9072
rect 3790 7656 3846 7712
rect 4066 8064 4122 8120
rect 4066 7928 4122 7984
rect 4526 9968 4582 10024
rect 4434 8492 4490 8528
rect 4434 8472 4436 8492
rect 4436 8472 4488 8492
rect 4488 8472 4490 8492
rect 4710 9832 4766 9888
rect 4158 7792 4214 7848
rect 3882 7404 3938 7440
rect 3882 7384 3884 7404
rect 3884 7384 3936 7404
rect 3936 7384 3938 7404
rect 3974 7284 3976 7304
rect 3976 7284 4028 7304
rect 4028 7284 4030 7304
rect 3974 7248 4030 7284
rect 3428 7098 3484 7100
rect 3508 7098 3564 7100
rect 3588 7098 3644 7100
rect 3668 7098 3724 7100
rect 3428 7046 3474 7098
rect 3474 7046 3484 7098
rect 3508 7046 3538 7098
rect 3538 7046 3550 7098
rect 3550 7046 3564 7098
rect 3588 7046 3602 7098
rect 3602 7046 3614 7098
rect 3614 7046 3644 7098
rect 3668 7046 3678 7098
rect 3678 7046 3724 7098
rect 3428 7044 3484 7046
rect 3508 7044 3564 7046
rect 3588 7044 3644 7046
rect 3668 7044 3724 7046
rect 3974 6840 4030 6896
rect 3428 6010 3484 6012
rect 3508 6010 3564 6012
rect 3588 6010 3644 6012
rect 3668 6010 3724 6012
rect 3428 5958 3474 6010
rect 3474 5958 3484 6010
rect 3508 5958 3538 6010
rect 3538 5958 3550 6010
rect 3550 5958 3564 6010
rect 3588 5958 3602 6010
rect 3602 5958 3614 6010
rect 3614 5958 3644 6010
rect 3668 5958 3678 6010
rect 3678 5958 3724 6010
rect 3428 5956 3484 5958
rect 3508 5956 3564 5958
rect 3588 5956 3644 5958
rect 3668 5956 3724 5958
rect 3428 4922 3484 4924
rect 3508 4922 3564 4924
rect 3588 4922 3644 4924
rect 3668 4922 3724 4924
rect 3428 4870 3474 4922
rect 3474 4870 3484 4922
rect 3508 4870 3538 4922
rect 3538 4870 3550 4922
rect 3550 4870 3564 4922
rect 3588 4870 3602 4922
rect 3602 4870 3614 4922
rect 3614 4870 3644 4922
rect 3668 4870 3678 4922
rect 3678 4870 3724 4922
rect 3428 4868 3484 4870
rect 3508 4868 3564 4870
rect 3588 4868 3644 4870
rect 3668 4868 3724 4870
rect 3882 6024 3938 6080
rect 4158 7112 4214 7168
rect 4066 6568 4122 6624
rect 4066 6432 4122 6488
rect 4158 5616 4214 5672
rect 3606 4664 3662 4720
rect 3790 4664 3846 4720
rect 3974 4528 4030 4584
rect 3790 4392 3846 4448
rect 3428 3834 3484 3836
rect 3508 3834 3564 3836
rect 3588 3834 3644 3836
rect 3668 3834 3724 3836
rect 3428 3782 3474 3834
rect 3474 3782 3484 3834
rect 3508 3782 3538 3834
rect 3538 3782 3550 3834
rect 3550 3782 3564 3834
rect 3588 3782 3602 3834
rect 3602 3782 3614 3834
rect 3614 3782 3644 3834
rect 3668 3782 3678 3834
rect 3678 3782 3724 3834
rect 3428 3780 3484 3782
rect 3508 3780 3564 3782
rect 3588 3780 3644 3782
rect 3668 3780 3724 3782
rect 3428 2746 3484 2748
rect 3508 2746 3564 2748
rect 3588 2746 3644 2748
rect 3668 2746 3724 2748
rect 3428 2694 3474 2746
rect 3474 2694 3484 2746
rect 3508 2694 3538 2746
rect 3538 2694 3550 2746
rect 3550 2694 3564 2746
rect 3588 2694 3602 2746
rect 3602 2694 3614 2746
rect 3614 2694 3644 2746
rect 3668 2694 3678 2746
rect 3678 2694 3724 2746
rect 3428 2692 3484 2694
rect 3508 2692 3564 2694
rect 3588 2692 3644 2694
rect 3668 2692 3724 2694
rect 4158 4256 4214 4312
rect 4066 3984 4122 4040
rect 4158 3848 4214 3904
rect 4526 6296 4582 6352
rect 4434 5228 4490 5264
rect 4434 5208 4436 5228
rect 4436 5208 4488 5228
rect 4488 5208 4490 5228
rect 4526 4936 4582 4992
rect 4250 3712 4306 3768
rect 3790 2488 3846 2544
rect 4342 2624 4398 2680
rect 4710 9016 4766 9072
rect 4710 8880 4766 8936
rect 5078 9424 5134 9480
rect 4802 8608 4858 8664
rect 5538 13640 5594 13696
rect 5630 12552 5686 12608
rect 5900 19610 5956 19612
rect 5980 19610 6036 19612
rect 6060 19610 6116 19612
rect 6140 19610 6196 19612
rect 5900 19558 5946 19610
rect 5946 19558 5956 19610
rect 5980 19558 6010 19610
rect 6010 19558 6022 19610
rect 6022 19558 6036 19610
rect 6060 19558 6074 19610
rect 6074 19558 6086 19610
rect 6086 19558 6116 19610
rect 6140 19558 6150 19610
rect 6150 19558 6196 19610
rect 5900 19556 5956 19558
rect 5980 19556 6036 19558
rect 6060 19556 6116 19558
rect 6140 19556 6196 19558
rect 5900 18522 5956 18524
rect 5980 18522 6036 18524
rect 6060 18522 6116 18524
rect 6140 18522 6196 18524
rect 5900 18470 5946 18522
rect 5946 18470 5956 18522
rect 5980 18470 6010 18522
rect 6010 18470 6022 18522
rect 6022 18470 6036 18522
rect 6060 18470 6074 18522
rect 6074 18470 6086 18522
rect 6086 18470 6116 18522
rect 6140 18470 6150 18522
rect 6150 18470 6196 18522
rect 5900 18468 5956 18470
rect 5980 18468 6036 18470
rect 6060 18468 6116 18470
rect 6140 18468 6196 18470
rect 5906 18264 5962 18320
rect 5900 17434 5956 17436
rect 5980 17434 6036 17436
rect 6060 17434 6116 17436
rect 6140 17434 6196 17436
rect 5900 17382 5946 17434
rect 5946 17382 5956 17434
rect 5980 17382 6010 17434
rect 6010 17382 6022 17434
rect 6022 17382 6036 17434
rect 6060 17382 6074 17434
rect 6074 17382 6086 17434
rect 6086 17382 6116 17434
rect 6140 17382 6150 17434
rect 6150 17382 6196 17434
rect 5900 17380 5956 17382
rect 5980 17380 6036 17382
rect 6060 17380 6116 17382
rect 6140 17380 6196 17382
rect 6366 22072 6422 22128
rect 6366 20712 6422 20768
rect 6366 19352 6422 19408
rect 5906 16904 5962 16960
rect 6734 27124 6790 27160
rect 6734 27104 6736 27124
rect 6736 27104 6788 27124
rect 6788 27104 6790 27124
rect 7378 32428 7434 32464
rect 7378 32408 7380 32428
rect 7380 32408 7432 32428
rect 7432 32408 7434 32428
rect 7378 31592 7434 31648
rect 7378 29688 7434 29744
rect 7194 27648 7250 27704
rect 6918 26016 6974 26072
rect 6734 25472 6790 25528
rect 6734 24812 6790 24848
rect 6734 24792 6736 24812
rect 6736 24792 6788 24812
rect 6788 24792 6790 24812
rect 7286 26968 7342 27024
rect 7286 25880 7342 25936
rect 9632 42560 9688 42562
rect 9126 42508 9128 42528
rect 9128 42508 9180 42528
rect 9180 42508 9182 42528
rect 9126 42472 9182 42508
rect 9632 42508 9680 42560
rect 9680 42508 9688 42560
rect 9632 42506 9688 42508
rect 9126 41556 9128 41576
rect 9128 41556 9180 41576
rect 9180 41556 9182 41576
rect 9126 41520 9182 41556
rect 9770 41656 9826 41712
rect 9402 38800 9458 38856
rect 9034 34720 9090 34776
rect 8574 33904 8630 33960
rect 8850 33516 8906 33552
rect 9034 33768 9090 33824
rect 8850 33496 8852 33516
rect 8852 33496 8904 33516
rect 8904 33496 8906 33516
rect 8373 33210 8429 33212
rect 8453 33210 8509 33212
rect 8533 33210 8589 33212
rect 8613 33210 8669 33212
rect 8373 33158 8419 33210
rect 8419 33158 8429 33210
rect 8453 33158 8483 33210
rect 8483 33158 8495 33210
rect 8495 33158 8509 33210
rect 8533 33158 8547 33210
rect 8547 33158 8559 33210
rect 8559 33158 8589 33210
rect 8613 33158 8623 33210
rect 8623 33158 8669 33210
rect 8373 33156 8429 33158
rect 8453 33156 8509 33158
rect 8533 33156 8589 33158
rect 8613 33156 8669 33158
rect 8574 32988 8576 33008
rect 8576 32988 8628 33008
rect 8628 32988 8630 33008
rect 8574 32952 8630 32988
rect 7562 30368 7618 30424
rect 8022 31728 8078 31784
rect 8373 32122 8429 32124
rect 8453 32122 8509 32124
rect 8533 32122 8589 32124
rect 8613 32122 8669 32124
rect 8373 32070 8419 32122
rect 8419 32070 8429 32122
rect 8453 32070 8483 32122
rect 8483 32070 8495 32122
rect 8495 32070 8509 32122
rect 8533 32070 8547 32122
rect 8547 32070 8559 32122
rect 8559 32070 8589 32122
rect 8613 32070 8623 32122
rect 8623 32070 8669 32122
rect 8373 32068 8429 32070
rect 8453 32068 8509 32070
rect 8533 32068 8589 32070
rect 8613 32068 8669 32070
rect 8114 31456 8170 31512
rect 8206 31340 8262 31376
rect 8206 31320 8208 31340
rect 8208 31320 8260 31340
rect 8260 31320 8262 31340
rect 8114 30912 8170 30968
rect 8373 31034 8429 31036
rect 8453 31034 8509 31036
rect 8533 31034 8589 31036
rect 8613 31034 8669 31036
rect 8373 30982 8419 31034
rect 8419 30982 8429 31034
rect 8453 30982 8483 31034
rect 8483 30982 8495 31034
rect 8495 30982 8509 31034
rect 8533 30982 8547 31034
rect 8547 30982 8559 31034
rect 8559 30982 8589 31034
rect 8613 30982 8623 31034
rect 8623 30982 8669 31034
rect 8373 30980 8429 30982
rect 8453 30980 8509 30982
rect 8533 30980 8589 30982
rect 8613 30980 8669 30982
rect 7746 29144 7802 29200
rect 7562 25744 7618 25800
rect 7102 23840 7158 23896
rect 6642 20848 6698 20904
rect 6550 19488 6606 19544
rect 5900 16346 5956 16348
rect 5980 16346 6036 16348
rect 6060 16346 6116 16348
rect 6140 16346 6196 16348
rect 5900 16294 5946 16346
rect 5946 16294 5956 16346
rect 5980 16294 6010 16346
rect 6010 16294 6022 16346
rect 6022 16294 6036 16346
rect 6060 16294 6074 16346
rect 6074 16294 6086 16346
rect 6086 16294 6116 16346
rect 6140 16294 6150 16346
rect 6150 16294 6196 16346
rect 5900 16292 5956 16294
rect 5980 16292 6036 16294
rect 6060 16292 6116 16294
rect 6140 16292 6196 16294
rect 5906 15816 5962 15872
rect 5900 15258 5956 15260
rect 5980 15258 6036 15260
rect 6060 15258 6116 15260
rect 6140 15258 6196 15260
rect 5900 15206 5946 15258
rect 5946 15206 5956 15258
rect 5980 15206 6010 15258
rect 6010 15206 6022 15258
rect 6022 15206 6036 15258
rect 6060 15206 6074 15258
rect 6074 15206 6086 15258
rect 6086 15206 6116 15258
rect 6140 15206 6150 15258
rect 6150 15206 6196 15258
rect 5900 15204 5956 15206
rect 5980 15204 6036 15206
rect 6060 15204 6116 15206
rect 6140 15204 6196 15206
rect 6182 14728 6238 14784
rect 6274 14592 6330 14648
rect 5900 14170 5956 14172
rect 5980 14170 6036 14172
rect 6060 14170 6116 14172
rect 6140 14170 6196 14172
rect 5900 14118 5946 14170
rect 5946 14118 5956 14170
rect 5980 14118 6010 14170
rect 6010 14118 6022 14170
rect 6022 14118 6036 14170
rect 6060 14118 6074 14170
rect 6074 14118 6086 14170
rect 6086 14118 6116 14170
rect 6140 14118 6150 14170
rect 6150 14118 6196 14170
rect 5900 14116 5956 14118
rect 5980 14116 6036 14118
rect 6060 14116 6116 14118
rect 6140 14116 6196 14118
rect 5998 13504 6054 13560
rect 5814 13368 5870 13424
rect 5900 13082 5956 13084
rect 5980 13082 6036 13084
rect 6060 13082 6116 13084
rect 6140 13082 6196 13084
rect 5900 13030 5946 13082
rect 5946 13030 5956 13082
rect 5980 13030 6010 13082
rect 6010 13030 6022 13082
rect 6022 13030 6036 13082
rect 6060 13030 6074 13082
rect 6074 13030 6086 13082
rect 6086 13030 6116 13082
rect 6140 13030 6150 13082
rect 6150 13030 6196 13082
rect 5900 13028 5956 13030
rect 5980 13028 6036 13030
rect 6060 13028 6116 13030
rect 6140 13028 6196 13030
rect 5538 12008 5594 12064
rect 5538 11892 5594 11928
rect 5722 12008 5778 12064
rect 5538 11872 5540 11892
rect 5540 11872 5592 11892
rect 5592 11872 5594 11892
rect 5900 11994 5956 11996
rect 5980 11994 6036 11996
rect 6060 11994 6116 11996
rect 6140 11994 6196 11996
rect 5900 11942 5946 11994
rect 5946 11942 5956 11994
rect 5980 11942 6010 11994
rect 6010 11942 6022 11994
rect 6022 11942 6036 11994
rect 6060 11942 6074 11994
rect 6074 11942 6086 11994
rect 6086 11942 6116 11994
rect 6140 11942 6150 11994
rect 6150 11942 6196 11994
rect 5900 11940 5956 11942
rect 5980 11940 6036 11942
rect 6060 11940 6116 11942
rect 6140 11940 6196 11942
rect 5446 11328 5502 11384
rect 6182 11756 6238 11792
rect 6182 11736 6184 11756
rect 6184 11736 6236 11756
rect 6236 11736 6238 11756
rect 6734 15680 6790 15736
rect 6642 15544 6698 15600
rect 6550 15136 6606 15192
rect 6550 15000 6606 15056
rect 6366 14048 6422 14104
rect 6458 13096 6514 13152
rect 6366 12960 6422 13016
rect 6366 12708 6422 12744
rect 6366 12688 6368 12708
rect 6368 12688 6420 12708
rect 6420 12688 6422 12708
rect 6090 11328 6146 11384
rect 5446 11056 5502 11112
rect 5538 10376 5594 10432
rect 5354 9560 5410 9616
rect 5354 9288 5410 9344
rect 4802 7792 4858 7848
rect 4710 6568 4766 6624
rect 4710 4664 4766 4720
rect 4158 2352 4214 2408
rect 3428 1658 3484 1660
rect 3508 1658 3564 1660
rect 3588 1658 3644 1660
rect 3668 1658 3724 1660
rect 3428 1606 3474 1658
rect 3474 1606 3484 1658
rect 3508 1606 3538 1658
rect 3538 1606 3550 1658
rect 3550 1606 3564 1658
rect 3588 1606 3602 1658
rect 3602 1606 3614 1658
rect 3614 1606 3644 1658
rect 3668 1606 3678 1658
rect 3678 1606 3724 1658
rect 3428 1604 3484 1606
rect 3508 1604 3564 1606
rect 3588 1604 3644 1606
rect 3668 1604 3724 1606
rect 3882 584 3938 640
rect 4986 6296 5042 6352
rect 4894 6024 4950 6080
rect 5262 7928 5318 7984
rect 5170 7656 5226 7712
rect 5262 6840 5318 6896
rect 4986 4820 5042 4856
rect 4986 4800 4988 4820
rect 4988 4800 5040 4820
rect 5040 4800 5042 4820
rect 4986 3032 5042 3088
rect 5170 2352 5226 2408
rect 5900 10906 5956 10908
rect 5980 10906 6036 10908
rect 6060 10906 6116 10908
rect 6140 10906 6196 10908
rect 5900 10854 5946 10906
rect 5946 10854 5956 10906
rect 5980 10854 6010 10906
rect 6010 10854 6022 10906
rect 6022 10854 6036 10906
rect 6060 10854 6074 10906
rect 6074 10854 6086 10906
rect 6086 10854 6116 10906
rect 6140 10854 6150 10906
rect 6150 10854 6196 10906
rect 5900 10852 5956 10854
rect 5980 10852 6036 10854
rect 6060 10852 6116 10854
rect 6140 10852 6196 10854
rect 5900 9818 5956 9820
rect 5980 9818 6036 9820
rect 6060 9818 6116 9820
rect 6140 9818 6196 9820
rect 5900 9766 5946 9818
rect 5946 9766 5956 9818
rect 5980 9766 6010 9818
rect 6010 9766 6022 9818
rect 6022 9766 6036 9818
rect 6060 9766 6074 9818
rect 6074 9766 6086 9818
rect 6086 9766 6116 9818
rect 6140 9766 6150 9818
rect 6150 9766 6196 9818
rect 5900 9764 5956 9766
rect 5980 9764 6036 9766
rect 6060 9764 6116 9766
rect 6140 9764 6196 9766
rect 5998 9424 6054 9480
rect 6182 9560 6238 9616
rect 6366 11056 6422 11112
rect 6182 9152 6238 9208
rect 5722 8200 5778 8256
rect 5900 8730 5956 8732
rect 5980 8730 6036 8732
rect 6060 8730 6116 8732
rect 6140 8730 6196 8732
rect 5900 8678 5946 8730
rect 5946 8678 5956 8730
rect 5980 8678 6010 8730
rect 6010 8678 6022 8730
rect 6022 8678 6036 8730
rect 6060 8678 6074 8730
rect 6074 8678 6086 8730
rect 6086 8678 6116 8730
rect 6140 8678 6150 8730
rect 6150 8678 6196 8730
rect 5900 8676 5956 8678
rect 5980 8676 6036 8678
rect 6060 8676 6116 8678
rect 6140 8676 6196 8678
rect 6090 8508 6092 8528
rect 6092 8508 6144 8528
rect 6144 8508 6146 8528
rect 6090 8472 6146 8508
rect 5814 8064 5870 8120
rect 5998 8200 6054 8256
rect 6182 8084 6238 8120
rect 6182 8064 6184 8084
rect 6184 8064 6236 8084
rect 6236 8064 6238 8084
rect 5900 7642 5956 7644
rect 5980 7642 6036 7644
rect 6060 7642 6116 7644
rect 6140 7642 6196 7644
rect 5900 7590 5946 7642
rect 5946 7590 5956 7642
rect 5980 7590 6010 7642
rect 6010 7590 6022 7642
rect 6022 7590 6036 7642
rect 6060 7590 6074 7642
rect 6074 7590 6086 7642
rect 6086 7590 6116 7642
rect 6140 7590 6150 7642
rect 6150 7590 6196 7642
rect 5900 7588 5956 7590
rect 5980 7588 6036 7590
rect 6060 7588 6116 7590
rect 6140 7588 6196 7590
rect 5630 6452 5686 6488
rect 5630 6432 5632 6452
rect 5632 6432 5684 6452
rect 5684 6432 5686 6452
rect 5538 5652 5540 5672
rect 5540 5652 5592 5672
rect 5592 5652 5594 5672
rect 5538 5616 5594 5652
rect 5354 5344 5410 5400
rect 5446 4664 5502 4720
rect 6090 6840 6146 6896
rect 5900 6554 5956 6556
rect 5980 6554 6036 6556
rect 6060 6554 6116 6556
rect 6140 6554 6196 6556
rect 5900 6502 5946 6554
rect 5946 6502 5956 6554
rect 5980 6502 6010 6554
rect 6010 6502 6022 6554
rect 6022 6502 6036 6554
rect 6060 6502 6074 6554
rect 6074 6502 6086 6554
rect 6086 6502 6116 6554
rect 6140 6502 6150 6554
rect 6150 6502 6196 6554
rect 5900 6500 5956 6502
rect 5980 6500 6036 6502
rect 6060 6500 6116 6502
rect 6140 6500 6196 6502
rect 6826 15408 6882 15464
rect 6826 15000 6882 15056
rect 6734 13096 6790 13152
rect 6550 11056 6606 11112
rect 8850 33088 8906 33144
rect 9034 32952 9090 33008
rect 9034 32816 9090 32872
rect 8942 31728 8998 31784
rect 8206 30640 8262 30696
rect 8373 29946 8429 29948
rect 8453 29946 8509 29948
rect 8533 29946 8589 29948
rect 8613 29946 8669 29948
rect 8373 29894 8419 29946
rect 8419 29894 8429 29946
rect 8453 29894 8483 29946
rect 8483 29894 8495 29946
rect 8495 29894 8509 29946
rect 8533 29894 8547 29946
rect 8547 29894 8559 29946
rect 8559 29894 8589 29946
rect 8613 29894 8623 29946
rect 8623 29894 8669 29946
rect 8373 29892 8429 29894
rect 8453 29892 8509 29894
rect 8533 29892 8589 29894
rect 8613 29892 8669 29894
rect 8114 28464 8170 28520
rect 8298 29008 8354 29064
rect 8373 28858 8429 28860
rect 8453 28858 8509 28860
rect 8533 28858 8589 28860
rect 8613 28858 8669 28860
rect 8373 28806 8419 28858
rect 8419 28806 8429 28858
rect 8453 28806 8483 28858
rect 8483 28806 8495 28858
rect 8495 28806 8509 28858
rect 8533 28806 8547 28858
rect 8547 28806 8559 28858
rect 8559 28806 8589 28858
rect 8613 28806 8623 28858
rect 8623 28806 8669 28858
rect 8373 28804 8429 28806
rect 8453 28804 8509 28806
rect 8533 28804 8589 28806
rect 8613 28804 8669 28806
rect 8298 28600 8354 28656
rect 8373 27770 8429 27772
rect 8453 27770 8509 27772
rect 8533 27770 8589 27772
rect 8613 27770 8669 27772
rect 8373 27718 8419 27770
rect 8419 27718 8429 27770
rect 8453 27718 8483 27770
rect 8483 27718 8495 27770
rect 8495 27718 8509 27770
rect 8533 27718 8547 27770
rect 8547 27718 8559 27770
rect 8559 27718 8589 27770
rect 8613 27718 8623 27770
rect 8623 27718 8669 27770
rect 8373 27716 8429 27718
rect 8453 27716 8509 27718
rect 8533 27716 8589 27718
rect 8613 27716 8669 27718
rect 8206 26968 8262 27024
rect 8373 26682 8429 26684
rect 8453 26682 8509 26684
rect 8533 26682 8589 26684
rect 8613 26682 8669 26684
rect 8373 26630 8419 26682
rect 8419 26630 8429 26682
rect 8453 26630 8483 26682
rect 8483 26630 8495 26682
rect 8495 26630 8509 26682
rect 8533 26630 8547 26682
rect 8547 26630 8559 26682
rect 8559 26630 8589 26682
rect 8613 26630 8623 26682
rect 8623 26630 8669 26682
rect 8373 26628 8429 26630
rect 8453 26628 8509 26630
rect 8533 26628 8589 26630
rect 8613 26628 8669 26630
rect 8114 26308 8170 26344
rect 8114 26288 8116 26308
rect 8116 26288 8168 26308
rect 8168 26288 8170 26308
rect 7838 26152 7894 26208
rect 7838 25064 7894 25120
rect 7746 24928 7802 24984
rect 7654 24384 7710 24440
rect 8574 26288 8630 26344
rect 7470 23704 7526 23760
rect 7470 22208 7526 22264
rect 7470 20712 7526 20768
rect 7286 20576 7342 20632
rect 7378 20304 7434 20360
rect 7378 19896 7434 19952
rect 7378 19760 7434 19816
rect 7286 18808 7342 18864
rect 7654 22480 7710 22536
rect 8373 25594 8429 25596
rect 8453 25594 8509 25596
rect 8533 25594 8589 25596
rect 8613 25594 8669 25596
rect 8373 25542 8419 25594
rect 8419 25542 8429 25594
rect 8453 25542 8483 25594
rect 8483 25542 8495 25594
rect 8495 25542 8509 25594
rect 8533 25542 8547 25594
rect 8547 25542 8559 25594
rect 8559 25542 8589 25594
rect 8613 25542 8623 25594
rect 8623 25542 8669 25594
rect 8373 25540 8429 25542
rect 8453 25540 8509 25542
rect 8533 25540 8589 25542
rect 8613 25540 8669 25542
rect 8758 24928 8814 24984
rect 8373 24506 8429 24508
rect 8453 24506 8509 24508
rect 8533 24506 8589 24508
rect 8613 24506 8669 24508
rect 8373 24454 8419 24506
rect 8419 24454 8429 24506
rect 8453 24454 8483 24506
rect 8483 24454 8495 24506
rect 8495 24454 8509 24506
rect 8533 24454 8547 24506
rect 8547 24454 8559 24506
rect 8559 24454 8589 24506
rect 8613 24454 8623 24506
rect 8623 24454 8669 24506
rect 8373 24452 8429 24454
rect 8453 24452 8509 24454
rect 8533 24452 8589 24454
rect 8613 24452 8669 24454
rect 8206 23976 8262 24032
rect 7930 23568 7986 23624
rect 7102 16768 7158 16824
rect 7010 15680 7066 15736
rect 6918 13368 6974 13424
rect 6826 11736 6882 11792
rect 7010 12960 7066 13016
rect 7470 18284 7526 18320
rect 7470 18264 7472 18284
rect 7472 18264 7524 18284
rect 7524 18264 7526 18284
rect 8022 22072 8078 22128
rect 8373 23418 8429 23420
rect 8453 23418 8509 23420
rect 8533 23418 8589 23420
rect 8613 23418 8669 23420
rect 8373 23366 8419 23418
rect 8419 23366 8429 23418
rect 8453 23366 8483 23418
rect 8483 23366 8495 23418
rect 8495 23366 8509 23418
rect 8533 23366 8547 23418
rect 8547 23366 8559 23418
rect 8559 23366 8589 23418
rect 8613 23366 8623 23418
rect 8623 23366 8669 23418
rect 8373 23364 8429 23366
rect 8453 23364 8509 23366
rect 8533 23364 8589 23366
rect 8613 23364 8669 23366
rect 8114 21936 8170 21992
rect 8373 22330 8429 22332
rect 8453 22330 8509 22332
rect 8533 22330 8589 22332
rect 8613 22330 8669 22332
rect 8373 22278 8419 22330
rect 8419 22278 8429 22330
rect 8453 22278 8483 22330
rect 8483 22278 8495 22330
rect 8495 22278 8509 22330
rect 8533 22278 8547 22330
rect 8547 22278 8559 22330
rect 8559 22278 8589 22330
rect 8613 22278 8623 22330
rect 8623 22278 8669 22330
rect 8373 22276 8429 22278
rect 8453 22276 8509 22278
rect 8533 22276 8589 22278
rect 8613 22276 8669 22278
rect 7838 18808 7894 18864
rect 7838 17448 7894 17504
rect 7470 15544 7526 15600
rect 7838 16360 7894 16416
rect 7286 14456 7342 14512
rect 7286 14048 7342 14104
rect 7194 13776 7250 13832
rect 7010 11328 7066 11384
rect 7102 10920 7158 10976
rect 7286 13640 7342 13696
rect 6550 8608 6606 8664
rect 6458 7792 6514 7848
rect 6458 7520 6514 7576
rect 6458 6432 6514 6488
rect 6366 6160 6422 6216
rect 6550 6160 6606 6216
rect 6458 5888 6514 5944
rect 5900 5466 5956 5468
rect 5980 5466 6036 5468
rect 6060 5466 6116 5468
rect 6140 5466 6196 5468
rect 5900 5414 5946 5466
rect 5946 5414 5956 5466
rect 5980 5414 6010 5466
rect 6010 5414 6022 5466
rect 6022 5414 6036 5466
rect 6060 5414 6074 5466
rect 6074 5414 6086 5466
rect 6086 5414 6116 5466
rect 6140 5414 6150 5466
rect 6150 5414 6196 5466
rect 5900 5412 5956 5414
rect 5980 5412 6036 5414
rect 6060 5412 6116 5414
rect 6140 5412 6196 5414
rect 5900 4378 5956 4380
rect 5980 4378 6036 4380
rect 6060 4378 6116 4380
rect 6140 4378 6196 4380
rect 5900 4326 5946 4378
rect 5946 4326 5956 4378
rect 5980 4326 6010 4378
rect 6010 4326 6022 4378
rect 6022 4326 6036 4378
rect 6060 4326 6074 4378
rect 6074 4326 6086 4378
rect 6086 4326 6116 4378
rect 6140 4326 6150 4378
rect 6150 4326 6196 4378
rect 5900 4324 5956 4326
rect 5980 4324 6036 4326
rect 6060 4324 6116 4326
rect 6140 4324 6196 4326
rect 5354 1128 5410 1184
rect 5538 1264 5594 1320
rect 5900 3290 5956 3292
rect 5980 3290 6036 3292
rect 6060 3290 6116 3292
rect 6140 3290 6196 3292
rect 5900 3238 5946 3290
rect 5946 3238 5956 3290
rect 5980 3238 6010 3290
rect 6010 3238 6022 3290
rect 6022 3238 6036 3290
rect 6060 3238 6074 3290
rect 6074 3238 6086 3290
rect 6086 3238 6116 3290
rect 6140 3238 6150 3290
rect 6150 3238 6196 3290
rect 5900 3236 5956 3238
rect 5980 3236 6036 3238
rect 6060 3236 6116 3238
rect 6140 3236 6196 3238
rect 6274 3168 6330 3224
rect 6182 3032 6238 3088
rect 6550 3576 6606 3632
rect 6826 10376 6882 10432
rect 6918 9560 6974 9616
rect 6918 9052 6920 9072
rect 6920 9052 6972 9072
rect 6972 9052 6974 9072
rect 6918 9016 6974 9052
rect 7194 10376 7250 10432
rect 7378 13504 7434 13560
rect 7746 15000 7802 15056
rect 7654 14864 7710 14920
rect 7562 12280 7618 12336
rect 7194 9696 7250 9752
rect 7286 9424 7342 9480
rect 7746 14184 7802 14240
rect 9126 30096 9182 30152
rect 10230 43424 10286 43480
rect 10138 42644 10140 42664
rect 10140 42644 10192 42664
rect 10192 42644 10194 42664
rect 10138 42608 10194 42644
rect 9954 42064 10010 42120
rect 9862 39616 9918 39672
rect 9678 38120 9734 38176
rect 9402 37188 9458 37224
rect 9402 37168 9404 37188
rect 9404 37168 9456 37188
rect 9456 37168 9458 37188
rect 9402 36216 9458 36272
rect 9494 35672 9550 35728
rect 9770 35808 9826 35864
rect 10046 37868 10102 37904
rect 10046 37848 10048 37868
rect 10048 37848 10100 37868
rect 10100 37848 10102 37868
rect 9310 33904 9366 33960
rect 9954 35264 10010 35320
rect 9954 34992 10010 35048
rect 9586 32952 9642 33008
rect 9402 31864 9458 31920
rect 9402 31592 9458 31648
rect 9126 26968 9182 27024
rect 9034 25492 9090 25528
rect 9034 25472 9036 25492
rect 9036 25472 9088 25492
rect 9088 25472 9090 25492
rect 8373 21242 8429 21244
rect 8453 21242 8509 21244
rect 8533 21242 8589 21244
rect 8613 21242 8669 21244
rect 8373 21190 8419 21242
rect 8419 21190 8429 21242
rect 8453 21190 8483 21242
rect 8483 21190 8495 21242
rect 8495 21190 8509 21242
rect 8533 21190 8547 21242
rect 8547 21190 8559 21242
rect 8559 21190 8589 21242
rect 8613 21190 8623 21242
rect 8623 21190 8669 21242
rect 8373 21188 8429 21190
rect 8453 21188 8509 21190
rect 8533 21188 8589 21190
rect 8613 21188 8669 21190
rect 8666 20884 8668 20904
rect 8668 20884 8720 20904
rect 8720 20884 8722 20904
rect 8666 20848 8722 20884
rect 8373 20154 8429 20156
rect 8453 20154 8509 20156
rect 8533 20154 8589 20156
rect 8613 20154 8669 20156
rect 8373 20102 8419 20154
rect 8419 20102 8429 20154
rect 8453 20102 8483 20154
rect 8483 20102 8495 20154
rect 8495 20102 8509 20154
rect 8533 20102 8547 20154
rect 8547 20102 8559 20154
rect 8559 20102 8589 20154
rect 8613 20102 8623 20154
rect 8623 20102 8669 20154
rect 8373 20100 8429 20102
rect 8453 20100 8509 20102
rect 8533 20100 8589 20102
rect 8613 20100 8669 20102
rect 9034 23044 9090 23080
rect 9034 23024 9036 23044
rect 9036 23024 9088 23044
rect 9088 23024 9090 23044
rect 9034 22616 9090 22672
rect 9034 22480 9090 22536
rect 9034 21664 9090 21720
rect 8373 19066 8429 19068
rect 8453 19066 8509 19068
rect 8533 19066 8589 19068
rect 8613 19066 8669 19068
rect 8373 19014 8419 19066
rect 8419 19014 8429 19066
rect 8453 19014 8483 19066
rect 8483 19014 8495 19066
rect 8495 19014 8509 19066
rect 8533 19014 8547 19066
rect 8547 19014 8559 19066
rect 8559 19014 8589 19066
rect 8613 19014 8623 19066
rect 8623 19014 8669 19066
rect 8373 19012 8429 19014
rect 8453 19012 8509 19014
rect 8533 19012 8589 19014
rect 8613 19012 8669 19014
rect 8114 16088 8170 16144
rect 8022 14864 8078 14920
rect 7930 14456 7986 14512
rect 7930 13776 7986 13832
rect 7654 10920 7710 10976
rect 7654 10784 7710 10840
rect 7654 9968 7710 10024
rect 7654 9696 7710 9752
rect 7470 9424 7526 9480
rect 7194 8744 7250 8800
rect 6918 7248 6974 7304
rect 7102 6568 7158 6624
rect 7010 6160 7066 6216
rect 6734 5480 6790 5536
rect 6918 5752 6974 5808
rect 7562 8744 7618 8800
rect 7562 8472 7618 8528
rect 7470 8064 7526 8120
rect 7470 7792 7526 7848
rect 7838 9016 7894 9072
rect 7746 8064 7802 8120
rect 8373 17978 8429 17980
rect 8453 17978 8509 17980
rect 8533 17978 8589 17980
rect 8613 17978 8669 17980
rect 8373 17926 8419 17978
rect 8419 17926 8429 17978
rect 8453 17926 8483 17978
rect 8483 17926 8495 17978
rect 8495 17926 8509 17978
rect 8533 17926 8547 17978
rect 8547 17926 8559 17978
rect 8559 17926 8589 17978
rect 8613 17926 8623 17978
rect 8623 17926 8669 17978
rect 8373 17924 8429 17926
rect 8453 17924 8509 17926
rect 8533 17924 8589 17926
rect 8613 17924 8669 17926
rect 8942 19352 8998 19408
rect 8373 16890 8429 16892
rect 8453 16890 8509 16892
rect 8533 16890 8589 16892
rect 8613 16890 8669 16892
rect 8373 16838 8419 16890
rect 8419 16838 8429 16890
rect 8453 16838 8483 16890
rect 8483 16838 8495 16890
rect 8495 16838 8509 16890
rect 8533 16838 8547 16890
rect 8547 16838 8559 16890
rect 8559 16838 8589 16890
rect 8613 16838 8623 16890
rect 8623 16838 8669 16890
rect 8373 16836 8429 16838
rect 8453 16836 8509 16838
rect 8533 16836 8589 16838
rect 8613 16836 8669 16838
rect 8758 16088 8814 16144
rect 8373 15802 8429 15804
rect 8453 15802 8509 15804
rect 8533 15802 8589 15804
rect 8613 15802 8669 15804
rect 8373 15750 8419 15802
rect 8419 15750 8429 15802
rect 8453 15750 8483 15802
rect 8483 15750 8495 15802
rect 8495 15750 8509 15802
rect 8533 15750 8547 15802
rect 8547 15750 8559 15802
rect 8559 15750 8589 15802
rect 8613 15750 8623 15802
rect 8623 15750 8669 15802
rect 8373 15748 8429 15750
rect 8453 15748 8509 15750
rect 8533 15748 8589 15750
rect 8613 15748 8669 15750
rect 8666 15272 8722 15328
rect 8574 14884 8630 14920
rect 8574 14864 8576 14884
rect 8576 14864 8628 14884
rect 8628 14864 8630 14884
rect 8373 14714 8429 14716
rect 8453 14714 8509 14716
rect 8533 14714 8589 14716
rect 8613 14714 8669 14716
rect 8373 14662 8419 14714
rect 8419 14662 8429 14714
rect 8453 14662 8483 14714
rect 8483 14662 8495 14714
rect 8495 14662 8509 14714
rect 8533 14662 8547 14714
rect 8547 14662 8559 14714
rect 8559 14662 8589 14714
rect 8613 14662 8623 14714
rect 8623 14662 8669 14714
rect 8373 14660 8429 14662
rect 8453 14660 8509 14662
rect 8533 14660 8589 14662
rect 8613 14660 8669 14662
rect 8206 13776 8262 13832
rect 8758 14184 8814 14240
rect 8373 13626 8429 13628
rect 8453 13626 8509 13628
rect 8533 13626 8589 13628
rect 8613 13626 8669 13628
rect 8373 13574 8419 13626
rect 8419 13574 8429 13626
rect 8453 13574 8483 13626
rect 8483 13574 8495 13626
rect 8495 13574 8509 13626
rect 8533 13574 8547 13626
rect 8547 13574 8559 13626
rect 8559 13574 8589 13626
rect 8613 13574 8623 13626
rect 8623 13574 8669 13626
rect 8373 13572 8429 13574
rect 8453 13572 8509 13574
rect 8533 13572 8589 13574
rect 8613 13572 8669 13574
rect 8022 11600 8078 11656
rect 8298 13096 8354 13152
rect 8666 13368 8722 13424
rect 8666 12724 8668 12744
rect 8668 12724 8720 12744
rect 8720 12724 8722 12744
rect 8666 12688 8722 12724
rect 8373 12538 8429 12540
rect 8453 12538 8509 12540
rect 8533 12538 8589 12540
rect 8613 12538 8669 12540
rect 8373 12486 8419 12538
rect 8419 12486 8429 12538
rect 8453 12486 8483 12538
rect 8483 12486 8495 12538
rect 8495 12486 8509 12538
rect 8533 12486 8547 12538
rect 8547 12486 8559 12538
rect 8559 12486 8589 12538
rect 8613 12486 8623 12538
rect 8623 12486 8669 12538
rect 8373 12484 8429 12486
rect 8453 12484 8509 12486
rect 8533 12484 8589 12486
rect 8613 12484 8669 12486
rect 8022 10648 8078 10704
rect 8022 10376 8078 10432
rect 7562 7112 7618 7168
rect 7286 6568 7342 6624
rect 7286 6432 7342 6488
rect 7930 6704 7986 6760
rect 7286 6024 7342 6080
rect 6734 4548 6790 4584
rect 6734 4528 6736 4548
rect 6736 4528 6788 4548
rect 6788 4528 6790 4548
rect 6734 4392 6790 4448
rect 6826 3440 6882 3496
rect 6734 2896 6790 2952
rect 5900 2202 5956 2204
rect 5980 2202 6036 2204
rect 6060 2202 6116 2204
rect 6140 2202 6196 2204
rect 5900 2150 5946 2202
rect 5946 2150 5956 2202
rect 5980 2150 6010 2202
rect 6010 2150 6022 2202
rect 6022 2150 6036 2202
rect 6060 2150 6074 2202
rect 6074 2150 6086 2202
rect 6086 2150 6116 2202
rect 6140 2150 6150 2202
rect 6150 2150 6196 2202
rect 5900 2148 5956 2150
rect 5980 2148 6036 2150
rect 6060 2148 6116 2150
rect 6140 2148 6196 2150
rect 6090 1944 6146 2000
rect 6642 1944 6698 2000
rect 5900 1114 5956 1116
rect 5980 1114 6036 1116
rect 6060 1114 6116 1116
rect 6140 1114 6196 1116
rect 5900 1062 5946 1114
rect 5946 1062 5956 1114
rect 5980 1062 6010 1114
rect 6010 1062 6022 1114
rect 6022 1062 6036 1114
rect 6060 1062 6074 1114
rect 6074 1062 6086 1114
rect 6086 1062 6116 1114
rect 6140 1062 6150 1114
rect 6150 1062 6196 1114
rect 5900 1060 5956 1062
rect 5980 1060 6036 1062
rect 6060 1060 6116 1062
rect 6140 1060 6196 1062
rect 7010 4800 7066 4856
rect 7286 4392 7342 4448
rect 7286 3984 7342 4040
rect 7010 3304 7066 3360
rect 6918 3032 6974 3088
rect 7010 2352 7066 2408
rect 6826 1808 6882 1864
rect 7194 3168 7250 3224
rect 7654 5344 7710 5400
rect 7654 4936 7710 4992
rect 7930 6160 7986 6216
rect 7838 5208 7894 5264
rect 7838 3848 7894 3904
rect 8574 12008 8630 12064
rect 8373 11450 8429 11452
rect 8453 11450 8509 11452
rect 8533 11450 8589 11452
rect 8613 11450 8669 11452
rect 8373 11398 8419 11450
rect 8419 11398 8429 11450
rect 8453 11398 8483 11450
rect 8483 11398 8495 11450
rect 8495 11398 8509 11450
rect 8533 11398 8547 11450
rect 8547 11398 8559 11450
rect 8559 11398 8589 11450
rect 8613 11398 8623 11450
rect 8623 11398 8669 11450
rect 8373 11396 8429 11398
rect 8453 11396 8509 11398
rect 8533 11396 8589 11398
rect 8613 11396 8669 11398
rect 8373 10362 8429 10364
rect 8453 10362 8509 10364
rect 8533 10362 8589 10364
rect 8613 10362 8669 10364
rect 8373 10310 8419 10362
rect 8419 10310 8429 10362
rect 8453 10310 8483 10362
rect 8483 10310 8495 10362
rect 8495 10310 8509 10362
rect 8533 10310 8547 10362
rect 8547 10310 8559 10362
rect 8559 10310 8589 10362
rect 8613 10310 8623 10362
rect 8623 10310 8669 10362
rect 8373 10308 8429 10310
rect 8453 10308 8509 10310
rect 8533 10308 8589 10310
rect 8613 10308 8669 10310
rect 8206 9832 8262 9888
rect 8114 9696 8170 9752
rect 8298 9696 8354 9752
rect 8758 10124 8814 10160
rect 8758 10104 8760 10124
rect 8760 10104 8812 10124
rect 8812 10104 8814 10124
rect 8666 9696 8722 9752
rect 8206 9152 8262 9208
rect 8373 9274 8429 9276
rect 8453 9274 8509 9276
rect 8533 9274 8589 9276
rect 8613 9274 8669 9276
rect 8373 9222 8419 9274
rect 8419 9222 8429 9274
rect 8453 9222 8483 9274
rect 8483 9222 8495 9274
rect 8495 9222 8509 9274
rect 8533 9222 8547 9274
rect 8547 9222 8559 9274
rect 8559 9222 8589 9274
rect 8613 9222 8623 9274
rect 8623 9222 8669 9274
rect 8373 9220 8429 9222
rect 8453 9220 8509 9222
rect 8533 9220 8589 9222
rect 8613 9220 8669 9222
rect 8206 9036 8262 9072
rect 8206 9016 8208 9036
rect 8208 9016 8260 9036
rect 8260 9016 8262 9036
rect 8574 9016 8630 9072
rect 7286 2624 7342 2680
rect 7470 2216 7526 2272
rect 7930 3168 7986 3224
rect 8482 8608 8538 8664
rect 8390 8336 8446 8392
rect 8373 8186 8429 8188
rect 8453 8186 8509 8188
rect 8533 8186 8589 8188
rect 8613 8186 8669 8188
rect 8373 8134 8419 8186
rect 8419 8134 8429 8186
rect 8453 8134 8483 8186
rect 8483 8134 8495 8186
rect 8495 8134 8509 8186
rect 8533 8134 8547 8186
rect 8547 8134 8559 8186
rect 8559 8134 8589 8186
rect 8613 8134 8623 8186
rect 8623 8134 8669 8186
rect 8373 8132 8429 8134
rect 8453 8132 8509 8134
rect 8533 8132 8589 8134
rect 8613 8132 8669 8134
rect 8666 7792 8722 7848
rect 8666 7656 8722 7712
rect 8373 7098 8429 7100
rect 8453 7098 8509 7100
rect 8533 7098 8589 7100
rect 8613 7098 8669 7100
rect 8373 7046 8419 7098
rect 8419 7046 8429 7098
rect 8453 7046 8483 7098
rect 8483 7046 8495 7098
rect 8495 7046 8509 7098
rect 8533 7046 8547 7098
rect 8547 7046 8559 7098
rect 8559 7046 8589 7098
rect 8613 7046 8623 7098
rect 8623 7046 8669 7098
rect 8373 7044 8429 7046
rect 8453 7044 8509 7046
rect 8533 7044 8589 7046
rect 8613 7044 8669 7046
rect 8390 6568 8446 6624
rect 8574 6160 8630 6216
rect 8373 6010 8429 6012
rect 8453 6010 8509 6012
rect 8533 6010 8589 6012
rect 8613 6010 8669 6012
rect 8373 5958 8419 6010
rect 8419 5958 8429 6010
rect 8453 5958 8483 6010
rect 8483 5958 8495 6010
rect 8495 5958 8509 6010
rect 8533 5958 8547 6010
rect 8547 5958 8559 6010
rect 8559 5958 8589 6010
rect 8613 5958 8623 6010
rect 8623 5958 8669 6010
rect 8373 5956 8429 5958
rect 8453 5956 8509 5958
rect 8533 5956 8589 5958
rect 8613 5956 8669 5958
rect 8666 5752 8722 5808
rect 8206 4800 8262 4856
rect 8373 4922 8429 4924
rect 8453 4922 8509 4924
rect 8533 4922 8589 4924
rect 8613 4922 8669 4924
rect 8373 4870 8419 4922
rect 8419 4870 8429 4922
rect 8453 4870 8483 4922
rect 8483 4870 8495 4922
rect 8495 4870 8509 4922
rect 8533 4870 8547 4922
rect 8547 4870 8559 4922
rect 8559 4870 8589 4922
rect 8613 4870 8623 4922
rect 8623 4870 8669 4922
rect 8373 4868 8429 4870
rect 8453 4868 8509 4870
rect 8533 4868 8589 4870
rect 8613 4868 8669 4870
rect 8373 3834 8429 3836
rect 8453 3834 8509 3836
rect 8533 3834 8589 3836
rect 8613 3834 8669 3836
rect 8373 3782 8419 3834
rect 8419 3782 8429 3834
rect 8453 3782 8483 3834
rect 8483 3782 8495 3834
rect 8495 3782 8509 3834
rect 8533 3782 8547 3834
rect 8547 3782 8559 3834
rect 8559 3782 8589 3834
rect 8613 3782 8623 3834
rect 8623 3782 8669 3834
rect 8373 3780 8429 3782
rect 8453 3780 8509 3782
rect 8533 3780 8589 3782
rect 8613 3780 8669 3782
rect 8390 3576 8446 3632
rect 7562 720 7618 776
rect 8373 2746 8429 2748
rect 8453 2746 8509 2748
rect 8533 2746 8589 2748
rect 8613 2746 8669 2748
rect 8373 2694 8419 2746
rect 8419 2694 8429 2746
rect 8453 2694 8483 2746
rect 8483 2694 8495 2746
rect 8495 2694 8509 2746
rect 8533 2694 8547 2746
rect 8547 2694 8559 2746
rect 8559 2694 8589 2746
rect 8613 2694 8623 2746
rect 8623 2694 8669 2746
rect 8373 2692 8429 2694
rect 8453 2692 8509 2694
rect 8533 2692 8589 2694
rect 8613 2692 8669 2694
rect 8482 1980 8484 2000
rect 8484 1980 8536 2000
rect 8536 1980 8538 2000
rect 8482 1944 8538 1980
rect 8206 1708 8208 1728
rect 8208 1708 8260 1728
rect 8260 1708 8262 1728
rect 8206 1672 8262 1708
rect 8373 1658 8429 1660
rect 8453 1658 8509 1660
rect 8533 1658 8589 1660
rect 8613 1658 8669 1660
rect 8373 1606 8419 1658
rect 8419 1606 8429 1658
rect 8453 1606 8483 1658
rect 8483 1606 8495 1658
rect 8495 1606 8509 1658
rect 8533 1606 8547 1658
rect 8547 1606 8559 1658
rect 8559 1606 8589 1658
rect 8613 1606 8623 1658
rect 8623 1606 8669 1658
rect 8373 1604 8429 1606
rect 8453 1604 8509 1606
rect 8533 1604 8589 1606
rect 8613 1604 8669 1606
rect 8114 1536 8170 1592
rect 9402 29008 9458 29064
rect 9310 25064 9366 25120
rect 9678 32136 9734 32192
rect 9954 33768 10010 33824
rect 9954 32000 10010 32056
rect 10598 43288 10654 43344
rect 10845 43546 10901 43548
rect 10925 43546 10981 43548
rect 11005 43546 11061 43548
rect 11085 43546 11141 43548
rect 10845 43494 10891 43546
rect 10891 43494 10901 43546
rect 10925 43494 10955 43546
rect 10955 43494 10967 43546
rect 10967 43494 10981 43546
rect 11005 43494 11019 43546
rect 11019 43494 11031 43546
rect 11031 43494 11061 43546
rect 11085 43494 11095 43546
rect 11095 43494 11141 43546
rect 10845 43492 10901 43494
rect 10925 43492 10981 43494
rect 11005 43492 11061 43494
rect 11085 43492 11141 43494
rect 10782 42880 10838 42936
rect 10598 38256 10654 38312
rect 10506 38156 10508 38176
rect 10508 38156 10560 38176
rect 10560 38156 10562 38176
rect 10506 38120 10562 38156
rect 10414 36352 10470 36408
rect 10322 35808 10378 35864
rect 10138 34584 10194 34640
rect 10506 35808 10562 35864
rect 10506 35128 10562 35184
rect 10230 32000 10286 32056
rect 9770 30776 9826 30832
rect 9586 28600 9642 28656
rect 9862 28872 9918 28928
rect 10046 28328 10102 28384
rect 9954 26288 10010 26344
rect 9862 26016 9918 26072
rect 9770 25064 9826 25120
rect 9218 23568 9274 23624
rect 9310 23432 9366 23488
rect 9218 22772 9274 22808
rect 9218 22752 9220 22772
rect 9220 22752 9272 22772
rect 9272 22752 9274 22772
rect 9770 24792 9826 24848
rect 9310 21412 9366 21448
rect 9310 21392 9312 21412
rect 9312 21392 9364 21412
rect 9364 21392 9366 21412
rect 9402 18944 9458 19000
rect 9310 18128 9366 18184
rect 10138 26016 10194 26072
rect 10046 25744 10102 25800
rect 10138 25336 10194 25392
rect 10046 24792 10102 24848
rect 9954 24520 10010 24576
rect 9954 23840 10010 23896
rect 10414 31476 10470 31512
rect 10414 31456 10416 31476
rect 10416 31456 10468 31476
rect 10468 31456 10470 31476
rect 10322 29008 10378 29064
rect 10322 28600 10378 28656
rect 10322 26152 10378 26208
rect 10845 42458 10901 42460
rect 10925 42458 10981 42460
rect 11005 42458 11061 42460
rect 11085 42458 11141 42460
rect 10845 42406 10891 42458
rect 10891 42406 10901 42458
rect 10925 42406 10955 42458
rect 10955 42406 10967 42458
rect 10967 42406 10981 42458
rect 11005 42406 11019 42458
rect 11019 42406 11031 42458
rect 11031 42406 11061 42458
rect 11085 42406 11095 42458
rect 11095 42406 11141 42458
rect 10845 42404 10901 42406
rect 10925 42404 10981 42406
rect 11005 42404 11061 42406
rect 11085 42404 11141 42406
rect 10845 41370 10901 41372
rect 10925 41370 10981 41372
rect 11005 41370 11061 41372
rect 11085 41370 11141 41372
rect 10845 41318 10891 41370
rect 10891 41318 10901 41370
rect 10925 41318 10955 41370
rect 10955 41318 10967 41370
rect 10967 41318 10981 41370
rect 11005 41318 11019 41370
rect 11019 41318 11031 41370
rect 11031 41318 11061 41370
rect 11085 41318 11095 41370
rect 11095 41318 11141 41370
rect 10845 41316 10901 41318
rect 10925 41316 10981 41318
rect 11005 41316 11061 41318
rect 11085 41316 11141 41318
rect 10845 40282 10901 40284
rect 10925 40282 10981 40284
rect 11005 40282 11061 40284
rect 11085 40282 11141 40284
rect 10845 40230 10891 40282
rect 10891 40230 10901 40282
rect 10925 40230 10955 40282
rect 10955 40230 10967 40282
rect 10967 40230 10981 40282
rect 11005 40230 11019 40282
rect 11019 40230 11031 40282
rect 11031 40230 11061 40282
rect 11085 40230 11095 40282
rect 11095 40230 11141 40282
rect 10845 40228 10901 40230
rect 10925 40228 10981 40230
rect 11005 40228 11061 40230
rect 11085 40228 11141 40230
rect 10845 39194 10901 39196
rect 10925 39194 10981 39196
rect 11005 39194 11061 39196
rect 11085 39194 11141 39196
rect 10845 39142 10891 39194
rect 10891 39142 10901 39194
rect 10925 39142 10955 39194
rect 10955 39142 10967 39194
rect 10967 39142 10981 39194
rect 11005 39142 11019 39194
rect 11019 39142 11031 39194
rect 11031 39142 11061 39194
rect 11085 39142 11095 39194
rect 11095 39142 11141 39194
rect 10845 39140 10901 39142
rect 10925 39140 10981 39142
rect 11005 39140 11061 39142
rect 11085 39140 11141 39142
rect 10845 38106 10901 38108
rect 10925 38106 10981 38108
rect 11005 38106 11061 38108
rect 11085 38106 11141 38108
rect 10845 38054 10891 38106
rect 10891 38054 10901 38106
rect 10925 38054 10955 38106
rect 10955 38054 10967 38106
rect 10967 38054 10981 38106
rect 11005 38054 11019 38106
rect 11019 38054 11031 38106
rect 11031 38054 11061 38106
rect 11085 38054 11095 38106
rect 11095 38054 11141 38106
rect 10845 38052 10901 38054
rect 10925 38052 10981 38054
rect 11005 38052 11061 38054
rect 11085 38052 11141 38054
rect 10845 37018 10901 37020
rect 10925 37018 10981 37020
rect 11005 37018 11061 37020
rect 11085 37018 11141 37020
rect 10845 36966 10891 37018
rect 10891 36966 10901 37018
rect 10925 36966 10955 37018
rect 10955 36966 10967 37018
rect 10967 36966 10981 37018
rect 11005 36966 11019 37018
rect 11019 36966 11031 37018
rect 11031 36966 11061 37018
rect 11085 36966 11095 37018
rect 11095 36966 11141 37018
rect 10845 36964 10901 36966
rect 10925 36964 10981 36966
rect 11005 36964 11061 36966
rect 11085 36964 11141 36966
rect 11702 42608 11758 42664
rect 11518 37848 11574 37904
rect 10845 35930 10901 35932
rect 10925 35930 10981 35932
rect 11005 35930 11061 35932
rect 11085 35930 11141 35932
rect 10845 35878 10891 35930
rect 10891 35878 10901 35930
rect 10925 35878 10955 35930
rect 10955 35878 10967 35930
rect 10967 35878 10981 35930
rect 11005 35878 11019 35930
rect 11019 35878 11031 35930
rect 11031 35878 11061 35930
rect 11085 35878 11095 35930
rect 11095 35878 11141 35930
rect 10845 35876 10901 35878
rect 10925 35876 10981 35878
rect 11005 35876 11061 35878
rect 11085 35876 11141 35878
rect 10845 34842 10901 34844
rect 10925 34842 10981 34844
rect 11005 34842 11061 34844
rect 11085 34842 11141 34844
rect 10845 34790 10891 34842
rect 10891 34790 10901 34842
rect 10925 34790 10955 34842
rect 10955 34790 10967 34842
rect 10967 34790 10981 34842
rect 11005 34790 11019 34842
rect 11019 34790 11031 34842
rect 11031 34790 11061 34842
rect 11085 34790 11095 34842
rect 11095 34790 11141 34842
rect 10845 34788 10901 34790
rect 10925 34788 10981 34790
rect 11005 34788 11061 34790
rect 11085 34788 11141 34790
rect 11058 33904 11114 33960
rect 10845 33754 10901 33756
rect 10925 33754 10981 33756
rect 11005 33754 11061 33756
rect 11085 33754 11141 33756
rect 10845 33702 10891 33754
rect 10891 33702 10901 33754
rect 10925 33702 10955 33754
rect 10955 33702 10967 33754
rect 10967 33702 10981 33754
rect 11005 33702 11019 33754
rect 11019 33702 11031 33754
rect 11031 33702 11061 33754
rect 11085 33702 11095 33754
rect 11095 33702 11141 33754
rect 10845 33700 10901 33702
rect 10925 33700 10981 33702
rect 11005 33700 11061 33702
rect 11085 33700 11141 33702
rect 11242 33088 11298 33144
rect 10845 32666 10901 32668
rect 10925 32666 10981 32668
rect 11005 32666 11061 32668
rect 11085 32666 11141 32668
rect 10845 32614 10891 32666
rect 10891 32614 10901 32666
rect 10925 32614 10955 32666
rect 10955 32614 10967 32666
rect 10967 32614 10981 32666
rect 11005 32614 11019 32666
rect 11019 32614 11031 32666
rect 11031 32614 11061 32666
rect 11085 32614 11095 32666
rect 11095 32614 11141 32666
rect 10845 32612 10901 32614
rect 10925 32612 10981 32614
rect 11005 32612 11061 32614
rect 11085 32612 11141 32614
rect 11058 32172 11060 32192
rect 11060 32172 11112 32192
rect 11112 32172 11114 32192
rect 11058 32136 11114 32172
rect 10845 31578 10901 31580
rect 10925 31578 10981 31580
rect 11005 31578 11061 31580
rect 11085 31578 11141 31580
rect 10845 31526 10891 31578
rect 10891 31526 10901 31578
rect 10925 31526 10955 31578
rect 10955 31526 10967 31578
rect 10967 31526 10981 31578
rect 11005 31526 11019 31578
rect 11019 31526 11031 31578
rect 11031 31526 11061 31578
rect 11085 31526 11095 31578
rect 11095 31526 11141 31578
rect 10845 31524 10901 31526
rect 10925 31524 10981 31526
rect 11005 31524 11061 31526
rect 11085 31524 11141 31526
rect 10782 31320 10838 31376
rect 11058 31184 11114 31240
rect 10782 30640 10838 30696
rect 11610 34584 11666 34640
rect 11794 34584 11850 34640
rect 10845 30490 10901 30492
rect 10925 30490 10981 30492
rect 11005 30490 11061 30492
rect 11085 30490 11141 30492
rect 10845 30438 10891 30490
rect 10891 30438 10901 30490
rect 10925 30438 10955 30490
rect 10955 30438 10967 30490
rect 10967 30438 10981 30490
rect 11005 30438 11019 30490
rect 11019 30438 11031 30490
rect 11031 30438 11061 30490
rect 11085 30438 11095 30490
rect 11095 30438 11141 30490
rect 10845 30436 10901 30438
rect 10925 30436 10981 30438
rect 11005 30436 11061 30438
rect 11085 30436 11141 30438
rect 10845 29402 10901 29404
rect 10925 29402 10981 29404
rect 11005 29402 11061 29404
rect 11085 29402 11141 29404
rect 10845 29350 10891 29402
rect 10891 29350 10901 29402
rect 10925 29350 10955 29402
rect 10955 29350 10967 29402
rect 10967 29350 10981 29402
rect 11005 29350 11019 29402
rect 11019 29350 11031 29402
rect 11031 29350 11061 29402
rect 11085 29350 11095 29402
rect 11095 29350 11141 29402
rect 10845 29348 10901 29350
rect 10925 29348 10981 29350
rect 11005 29348 11061 29350
rect 11085 29348 11141 29350
rect 11242 29008 11298 29064
rect 10690 28464 10746 28520
rect 10845 28314 10901 28316
rect 10925 28314 10981 28316
rect 11005 28314 11061 28316
rect 11085 28314 11141 28316
rect 10845 28262 10891 28314
rect 10891 28262 10901 28314
rect 10925 28262 10955 28314
rect 10955 28262 10967 28314
rect 10967 28262 10981 28314
rect 11005 28262 11019 28314
rect 11019 28262 11031 28314
rect 11031 28262 11061 28314
rect 11085 28262 11095 28314
rect 11095 28262 11141 28314
rect 10845 28260 10901 28262
rect 10925 28260 10981 28262
rect 11005 28260 11061 28262
rect 11085 28260 11141 28262
rect 10845 27226 10901 27228
rect 10925 27226 10981 27228
rect 11005 27226 11061 27228
rect 11085 27226 11141 27228
rect 10845 27174 10891 27226
rect 10891 27174 10901 27226
rect 10925 27174 10955 27226
rect 10955 27174 10967 27226
rect 10967 27174 10981 27226
rect 11005 27174 11019 27226
rect 11019 27174 11031 27226
rect 11031 27174 11061 27226
rect 11085 27174 11095 27226
rect 11095 27174 11141 27226
rect 10845 27172 10901 27174
rect 10925 27172 10981 27174
rect 11005 27172 11061 27174
rect 11085 27172 11141 27174
rect 10966 26968 11022 27024
rect 10845 26138 10901 26140
rect 10925 26138 10981 26140
rect 11005 26138 11061 26140
rect 11085 26138 11141 26140
rect 10845 26086 10891 26138
rect 10891 26086 10901 26138
rect 10925 26086 10955 26138
rect 10955 26086 10967 26138
rect 10967 26086 10981 26138
rect 11005 26086 11019 26138
rect 11019 26086 11031 26138
rect 11031 26086 11061 26138
rect 11085 26086 11095 26138
rect 11095 26086 11141 26138
rect 10845 26084 10901 26086
rect 10925 26084 10981 26086
rect 11005 26084 11061 26086
rect 11085 26084 11141 26086
rect 12162 42200 12218 42256
rect 12346 41928 12402 41984
rect 12438 40976 12494 41032
rect 12438 38276 12494 38312
rect 12438 38256 12440 38276
rect 12440 38256 12492 38276
rect 12492 38256 12494 38276
rect 12438 37848 12494 37904
rect 12806 42064 12862 42120
rect 12714 37848 12770 37904
rect 12438 36760 12494 36816
rect 12438 36216 12494 36272
rect 12162 35808 12218 35864
rect 12162 35672 12218 35728
rect 12254 34856 12310 34912
rect 12530 34856 12586 34912
rect 13818 43832 13874 43888
rect 13542 43152 13598 43208
rect 13318 43002 13374 43004
rect 13398 43002 13454 43004
rect 13478 43002 13534 43004
rect 13558 43002 13614 43004
rect 13318 42950 13364 43002
rect 13364 42950 13374 43002
rect 13398 42950 13428 43002
rect 13428 42950 13440 43002
rect 13440 42950 13454 43002
rect 13478 42950 13492 43002
rect 13492 42950 13504 43002
rect 13504 42950 13534 43002
rect 13558 42950 13568 43002
rect 13568 42950 13614 43002
rect 13318 42948 13374 42950
rect 13398 42948 13454 42950
rect 13478 42948 13534 42950
rect 13558 42948 13614 42950
rect 13910 43288 13966 43344
rect 14186 43968 14242 44024
rect 14002 42744 14058 42800
rect 13318 41914 13374 41916
rect 13398 41914 13454 41916
rect 13478 41914 13534 41916
rect 13558 41914 13614 41916
rect 13318 41862 13364 41914
rect 13364 41862 13374 41914
rect 13398 41862 13428 41914
rect 13428 41862 13440 41914
rect 13440 41862 13454 41914
rect 13478 41862 13492 41914
rect 13492 41862 13504 41914
rect 13504 41862 13534 41914
rect 13558 41862 13568 41914
rect 13568 41862 13614 41914
rect 13318 41860 13374 41862
rect 13398 41860 13454 41862
rect 13478 41860 13534 41862
rect 13558 41860 13614 41862
rect 13174 41656 13230 41712
rect 13082 39072 13138 39128
rect 12990 38120 13046 38176
rect 12806 34720 12862 34776
rect 11794 31184 11850 31240
rect 11978 32952 12034 33008
rect 12070 31864 12126 31920
rect 11702 30096 11758 30152
rect 11702 29708 11758 29744
rect 11702 29688 11704 29708
rect 11704 29688 11756 29708
rect 11756 29688 11758 29708
rect 11794 28600 11850 28656
rect 11794 28056 11850 28112
rect 11426 26152 11482 26208
rect 11794 26696 11850 26752
rect 12438 30504 12494 30560
rect 12162 29008 12218 29064
rect 12438 28328 12494 28384
rect 12346 27648 12402 27704
rect 12346 26968 12402 27024
rect 12162 26560 12218 26616
rect 11978 26288 12034 26344
rect 10506 25336 10562 25392
rect 10414 24792 10470 24848
rect 9770 23432 9826 23488
rect 10322 23296 10378 23352
rect 9862 22616 9918 22672
rect 9770 21800 9826 21856
rect 9770 19080 9826 19136
rect 9494 17856 9550 17912
rect 9310 17040 9366 17096
rect 9218 16768 9274 16824
rect 9126 15680 9182 15736
rect 9126 15000 9182 15056
rect 9034 13812 9036 13832
rect 9036 13812 9088 13832
rect 9088 13812 9090 13832
rect 9034 13776 9090 13812
rect 9310 15816 9366 15872
rect 9310 15680 9366 15736
rect 9586 17584 9642 17640
rect 10230 21956 10286 21992
rect 10230 21936 10232 21956
rect 10232 21936 10284 21956
rect 10284 21936 10286 21956
rect 9954 20576 10010 20632
rect 10138 21392 10194 21448
rect 10230 20984 10286 21040
rect 10138 20712 10194 20768
rect 9954 19080 10010 19136
rect 10046 18808 10102 18864
rect 9862 17176 9918 17232
rect 9770 16904 9826 16960
rect 9954 17040 10010 17096
rect 9862 16768 9918 16824
rect 10230 19760 10286 19816
rect 10138 17312 10194 17368
rect 9678 16224 9734 16280
rect 9586 15272 9642 15328
rect 9218 11192 9274 11248
rect 9126 10376 9182 10432
rect 9034 5480 9090 5536
rect 9678 13776 9734 13832
rect 9586 13368 9642 13424
rect 9954 15272 10010 15328
rect 9862 14492 9864 14512
rect 9864 14492 9916 14512
rect 9916 14492 9918 14512
rect 9862 14456 9918 14492
rect 9954 14048 10010 14104
rect 9770 11736 9826 11792
rect 9770 10104 9826 10160
rect 10598 22752 10654 22808
rect 10506 22208 10562 22264
rect 10414 21800 10470 21856
rect 10506 19488 10562 19544
rect 10414 19216 10470 19272
rect 10506 18808 10562 18864
rect 11334 25744 11390 25800
rect 10845 25050 10901 25052
rect 10925 25050 10981 25052
rect 11005 25050 11061 25052
rect 11085 25050 11141 25052
rect 10845 24998 10891 25050
rect 10891 24998 10901 25050
rect 10925 24998 10955 25050
rect 10955 24998 10967 25050
rect 10967 24998 10981 25050
rect 11005 24998 11019 25050
rect 11019 24998 11031 25050
rect 11031 24998 11061 25050
rect 11085 24998 11095 25050
rect 11095 24998 11141 25050
rect 10845 24996 10901 24998
rect 10925 24996 10981 24998
rect 11005 24996 11061 24998
rect 11085 24996 11141 24998
rect 11058 24792 11114 24848
rect 11058 24248 11114 24304
rect 10845 23962 10901 23964
rect 10925 23962 10981 23964
rect 11005 23962 11061 23964
rect 11085 23962 11141 23964
rect 10845 23910 10891 23962
rect 10891 23910 10901 23962
rect 10925 23910 10955 23962
rect 10955 23910 10967 23962
rect 10967 23910 10981 23962
rect 11005 23910 11019 23962
rect 11019 23910 11031 23962
rect 11031 23910 11061 23962
rect 11085 23910 11095 23962
rect 11095 23910 11141 23962
rect 10845 23908 10901 23910
rect 10925 23908 10981 23910
rect 11005 23908 11061 23910
rect 11085 23908 11141 23910
rect 10782 23024 10838 23080
rect 11242 23432 11298 23488
rect 10845 22874 10901 22876
rect 10925 22874 10981 22876
rect 11005 22874 11061 22876
rect 11085 22874 11141 22876
rect 10845 22822 10891 22874
rect 10891 22822 10901 22874
rect 10925 22822 10955 22874
rect 10955 22822 10967 22874
rect 10967 22822 10981 22874
rect 11005 22822 11019 22874
rect 11019 22822 11031 22874
rect 11031 22822 11061 22874
rect 11085 22822 11095 22874
rect 11095 22822 11141 22874
rect 10845 22820 10901 22822
rect 10925 22820 10981 22822
rect 11005 22820 11061 22822
rect 11085 22820 11141 22822
rect 10845 21786 10901 21788
rect 10925 21786 10981 21788
rect 11005 21786 11061 21788
rect 11085 21786 11141 21788
rect 10845 21734 10891 21786
rect 10891 21734 10901 21786
rect 10925 21734 10955 21786
rect 10955 21734 10967 21786
rect 10967 21734 10981 21786
rect 11005 21734 11019 21786
rect 11019 21734 11031 21786
rect 11031 21734 11061 21786
rect 11085 21734 11095 21786
rect 11095 21734 11141 21786
rect 10845 21732 10901 21734
rect 10925 21732 10981 21734
rect 11005 21732 11061 21734
rect 11085 21732 11141 21734
rect 10845 20698 10901 20700
rect 10925 20698 10981 20700
rect 11005 20698 11061 20700
rect 11085 20698 11141 20700
rect 10845 20646 10891 20698
rect 10891 20646 10901 20698
rect 10925 20646 10955 20698
rect 10955 20646 10967 20698
rect 10967 20646 10981 20698
rect 11005 20646 11019 20698
rect 11019 20646 11031 20698
rect 11031 20646 11061 20698
rect 11085 20646 11095 20698
rect 11095 20646 11141 20698
rect 10845 20644 10901 20646
rect 10925 20644 10981 20646
rect 11005 20644 11061 20646
rect 11085 20644 11141 20646
rect 10874 19760 10930 19816
rect 10845 19610 10901 19612
rect 10925 19610 10981 19612
rect 11005 19610 11061 19612
rect 11085 19610 11141 19612
rect 10845 19558 10891 19610
rect 10891 19558 10901 19610
rect 10925 19558 10955 19610
rect 10955 19558 10967 19610
rect 10967 19558 10981 19610
rect 11005 19558 11019 19610
rect 11019 19558 11031 19610
rect 11031 19558 11061 19610
rect 11085 19558 11095 19610
rect 11095 19558 11141 19610
rect 10845 19556 10901 19558
rect 10925 19556 10981 19558
rect 11005 19556 11061 19558
rect 11085 19556 11141 19558
rect 11518 25472 11574 25528
rect 11426 24268 11482 24304
rect 11426 24248 11428 24268
rect 11428 24248 11480 24268
rect 11480 24248 11482 24268
rect 11886 24928 11942 24984
rect 11886 24384 11942 24440
rect 11886 23588 11942 23624
rect 11886 23568 11888 23588
rect 11888 23568 11940 23588
rect 11940 23568 11942 23588
rect 11702 21528 11758 21584
rect 10690 19216 10746 19272
rect 10845 18522 10901 18524
rect 10925 18522 10981 18524
rect 11005 18522 11061 18524
rect 11085 18522 11141 18524
rect 10845 18470 10891 18522
rect 10891 18470 10901 18522
rect 10925 18470 10955 18522
rect 10955 18470 10967 18522
rect 10967 18470 10981 18522
rect 11005 18470 11019 18522
rect 11019 18470 11031 18522
rect 11031 18470 11061 18522
rect 11085 18470 11095 18522
rect 11095 18470 11141 18522
rect 10845 18468 10901 18470
rect 10925 18468 10981 18470
rect 11005 18468 11061 18470
rect 11085 18468 11141 18470
rect 10690 18128 10746 18184
rect 10414 17040 10470 17096
rect 10598 14864 10654 14920
rect 10138 13096 10194 13152
rect 10414 13096 10470 13152
rect 10845 17434 10901 17436
rect 10925 17434 10981 17436
rect 11005 17434 11061 17436
rect 11085 17434 11141 17436
rect 10845 17382 10891 17434
rect 10891 17382 10901 17434
rect 10925 17382 10955 17434
rect 10955 17382 10967 17434
rect 10967 17382 10981 17434
rect 11005 17382 11019 17434
rect 11019 17382 11031 17434
rect 11031 17382 11061 17434
rect 11085 17382 11095 17434
rect 11095 17382 11141 17434
rect 10845 17380 10901 17382
rect 10925 17380 10981 17382
rect 11005 17380 11061 17382
rect 11085 17380 11141 17382
rect 10845 16346 10901 16348
rect 10925 16346 10981 16348
rect 11005 16346 11061 16348
rect 11085 16346 11141 16348
rect 10845 16294 10891 16346
rect 10891 16294 10901 16346
rect 10925 16294 10955 16346
rect 10955 16294 10967 16346
rect 10967 16294 10981 16346
rect 11005 16294 11019 16346
rect 11019 16294 11031 16346
rect 11031 16294 11061 16346
rect 11085 16294 11095 16346
rect 11095 16294 11141 16346
rect 10845 16292 10901 16294
rect 10925 16292 10981 16294
rect 11005 16292 11061 16294
rect 11085 16292 11141 16294
rect 11058 16088 11114 16144
rect 10845 15258 10901 15260
rect 10925 15258 10981 15260
rect 11005 15258 11061 15260
rect 11085 15258 11141 15260
rect 10845 15206 10891 15258
rect 10891 15206 10901 15258
rect 10925 15206 10955 15258
rect 10955 15206 10967 15258
rect 10967 15206 10981 15258
rect 11005 15206 11019 15258
rect 11019 15206 11031 15258
rect 11031 15206 11061 15258
rect 11085 15206 11095 15258
rect 11095 15206 11141 15258
rect 10845 15204 10901 15206
rect 10925 15204 10981 15206
rect 11005 15204 11061 15206
rect 11085 15204 11141 15206
rect 11058 14728 11114 14784
rect 10845 14170 10901 14172
rect 10925 14170 10981 14172
rect 11005 14170 11061 14172
rect 11085 14170 11141 14172
rect 10845 14118 10891 14170
rect 10891 14118 10901 14170
rect 10925 14118 10955 14170
rect 10955 14118 10967 14170
rect 10967 14118 10981 14170
rect 11005 14118 11019 14170
rect 11019 14118 11031 14170
rect 11031 14118 11061 14170
rect 11085 14118 11095 14170
rect 11095 14118 11141 14170
rect 10845 14116 10901 14118
rect 10925 14116 10981 14118
rect 11005 14116 11061 14118
rect 11085 14116 11141 14118
rect 10690 14048 10746 14104
rect 10598 13776 10654 13832
rect 10598 12416 10654 12472
rect 10230 11600 10286 11656
rect 10414 11056 10470 11112
rect 10046 10648 10102 10704
rect 9954 9288 10010 9344
rect 9218 7792 9274 7848
rect 9310 6160 9366 6216
rect 9218 5752 9274 5808
rect 9218 5652 9220 5672
rect 9220 5652 9272 5672
rect 9272 5652 9274 5672
rect 9218 5616 9274 5652
rect 9402 5208 9458 5264
rect 9310 5072 9366 5128
rect 9034 3304 9090 3360
rect 9310 3440 9366 3496
rect 9218 3168 9274 3224
rect 9310 2896 9366 2952
rect 9034 2352 9090 2408
rect 9126 2216 9182 2272
rect 9310 1808 9366 1864
rect 8114 1264 8170 1320
rect 8206 1128 8262 1184
rect 9310 1400 9366 1456
rect 10138 9832 10194 9888
rect 9678 7656 9734 7712
rect 10046 8608 10102 8664
rect 9862 7520 9918 7576
rect 9678 7112 9734 7168
rect 9678 6704 9734 6760
rect 9770 6296 9826 6352
rect 9770 5480 9826 5536
rect 12070 25608 12126 25664
rect 12346 26732 12348 26752
rect 12348 26732 12400 26752
rect 12400 26732 12402 26752
rect 12346 26696 12402 26732
rect 12714 29280 12770 29336
rect 12714 28872 12770 28928
rect 12070 23024 12126 23080
rect 12070 21548 12126 21584
rect 12070 21528 12072 21548
rect 12072 21528 12124 21548
rect 12124 21528 12126 21548
rect 11978 20848 12034 20904
rect 12346 23976 12402 24032
rect 12070 20460 12126 20496
rect 12070 20440 12072 20460
rect 12072 20440 12124 20460
rect 12124 20440 12126 20460
rect 11886 19508 11942 19544
rect 11886 19488 11888 19508
rect 11888 19488 11940 19508
rect 11940 19488 11942 19508
rect 11794 17040 11850 17096
rect 11794 16768 11850 16824
rect 11610 15680 11666 15736
rect 11518 14456 11574 14512
rect 11242 13096 11298 13152
rect 10845 13082 10901 13084
rect 10925 13082 10981 13084
rect 11005 13082 11061 13084
rect 11085 13082 11141 13084
rect 10845 13030 10891 13082
rect 10891 13030 10901 13082
rect 10925 13030 10955 13082
rect 10955 13030 10967 13082
rect 10967 13030 10981 13082
rect 11005 13030 11019 13082
rect 11019 13030 11031 13082
rect 11031 13030 11061 13082
rect 11085 13030 11095 13082
rect 11095 13030 11141 13082
rect 10845 13028 10901 13030
rect 10925 13028 10981 13030
rect 11005 13028 11061 13030
rect 11085 13028 11141 13030
rect 11058 12144 11114 12200
rect 11242 12144 11298 12200
rect 10845 11994 10901 11996
rect 10925 11994 10981 11996
rect 11005 11994 11061 11996
rect 11085 11994 11141 11996
rect 10845 11942 10891 11994
rect 10891 11942 10901 11994
rect 10925 11942 10955 11994
rect 10955 11942 10967 11994
rect 10967 11942 10981 11994
rect 11005 11942 11019 11994
rect 11019 11942 11031 11994
rect 11031 11942 11061 11994
rect 11085 11942 11095 11994
rect 11095 11942 11141 11994
rect 10845 11940 10901 11942
rect 10925 11940 10981 11942
rect 11005 11940 11061 11942
rect 11085 11940 11141 11942
rect 10845 10906 10901 10908
rect 10925 10906 10981 10908
rect 11005 10906 11061 10908
rect 11085 10906 11141 10908
rect 10845 10854 10891 10906
rect 10891 10854 10901 10906
rect 10925 10854 10955 10906
rect 10955 10854 10967 10906
rect 10967 10854 10981 10906
rect 11005 10854 11019 10906
rect 11019 10854 11031 10906
rect 11031 10854 11061 10906
rect 11085 10854 11095 10906
rect 11095 10854 11141 10906
rect 10845 10852 10901 10854
rect 10925 10852 10981 10854
rect 11005 10852 11061 10854
rect 11085 10852 11141 10854
rect 10690 10784 10746 10840
rect 11426 12688 11482 12744
rect 11610 12960 11666 13016
rect 11242 10512 11298 10568
rect 11242 10376 11298 10432
rect 10322 9696 10378 9752
rect 10506 9560 10562 9616
rect 10506 9288 10562 9344
rect 9770 4936 9826 4992
rect 9770 4800 9826 4856
rect 9862 3576 9918 3632
rect 10046 4528 10102 4584
rect 10414 7792 10470 7848
rect 11242 9832 11298 9888
rect 10845 9818 10901 9820
rect 10925 9818 10981 9820
rect 11005 9818 11061 9820
rect 11085 9818 11141 9820
rect 10845 9766 10891 9818
rect 10891 9766 10901 9818
rect 10925 9766 10955 9818
rect 10955 9766 10967 9818
rect 10967 9766 10981 9818
rect 11005 9766 11019 9818
rect 11019 9766 11031 9818
rect 11031 9766 11061 9818
rect 11085 9766 11095 9818
rect 11095 9766 11141 9818
rect 10845 9764 10901 9766
rect 10925 9764 10981 9766
rect 11005 9764 11061 9766
rect 11085 9764 11141 9766
rect 10966 9560 11022 9616
rect 10845 8730 10901 8732
rect 10925 8730 10981 8732
rect 11005 8730 11061 8732
rect 11085 8730 11141 8732
rect 10845 8678 10891 8730
rect 10891 8678 10901 8730
rect 10925 8678 10955 8730
rect 10955 8678 10967 8730
rect 10967 8678 10981 8730
rect 11005 8678 11019 8730
rect 11019 8678 11031 8730
rect 11031 8678 11061 8730
rect 11085 8678 11095 8730
rect 11095 8678 11141 8730
rect 10845 8676 10901 8678
rect 10925 8676 10981 8678
rect 11005 8676 11061 8678
rect 11085 8676 11141 8678
rect 10874 8200 10930 8256
rect 10874 7792 10930 7848
rect 11242 7792 11298 7848
rect 10845 7642 10901 7644
rect 10925 7642 10981 7644
rect 11005 7642 11061 7644
rect 11085 7642 11141 7644
rect 10845 7590 10891 7642
rect 10891 7590 10901 7642
rect 10925 7590 10955 7642
rect 10955 7590 10967 7642
rect 10967 7590 10981 7642
rect 11005 7590 11019 7642
rect 11019 7590 11031 7642
rect 11031 7590 11061 7642
rect 11085 7590 11095 7642
rect 11095 7590 11141 7642
rect 10845 7588 10901 7590
rect 10925 7588 10981 7590
rect 11005 7588 11061 7590
rect 11085 7588 11141 7590
rect 10506 6976 10562 7032
rect 10506 6296 10562 6352
rect 10874 7112 10930 7168
rect 10414 5888 10470 5944
rect 10414 5752 10470 5808
rect 10322 4936 10378 4992
rect 10046 3712 10102 3768
rect 10230 3848 10286 3904
rect 10506 4664 10562 4720
rect 11058 7112 11114 7168
rect 10966 6840 11022 6896
rect 10845 6554 10901 6556
rect 10925 6554 10981 6556
rect 11005 6554 11061 6556
rect 11085 6554 11141 6556
rect 10845 6502 10891 6554
rect 10891 6502 10901 6554
rect 10925 6502 10955 6554
rect 10955 6502 10967 6554
rect 10967 6502 10981 6554
rect 11005 6502 11019 6554
rect 11019 6502 11031 6554
rect 11031 6502 11061 6554
rect 11085 6502 11095 6554
rect 11095 6502 11141 6554
rect 10845 6500 10901 6502
rect 10925 6500 10981 6502
rect 11005 6500 11061 6502
rect 11085 6500 11141 6502
rect 10782 5888 10838 5944
rect 11150 6316 11206 6352
rect 11150 6296 11152 6316
rect 11152 6296 11204 6316
rect 11204 6296 11206 6316
rect 11058 6160 11114 6216
rect 11058 6024 11114 6080
rect 11610 10784 11666 10840
rect 11518 8744 11574 8800
rect 11334 7248 11390 7304
rect 12070 17040 12126 17096
rect 12714 25880 12770 25936
rect 12714 25608 12770 25664
rect 13318 40826 13374 40828
rect 13398 40826 13454 40828
rect 13478 40826 13534 40828
rect 13558 40826 13614 40828
rect 13318 40774 13364 40826
rect 13364 40774 13374 40826
rect 13398 40774 13428 40826
rect 13428 40774 13440 40826
rect 13440 40774 13454 40826
rect 13478 40774 13492 40826
rect 13492 40774 13504 40826
rect 13504 40774 13534 40826
rect 13558 40774 13568 40826
rect 13568 40774 13614 40826
rect 13318 40772 13374 40774
rect 13398 40772 13454 40774
rect 13478 40772 13534 40774
rect 13558 40772 13614 40774
rect 13542 40024 13598 40080
rect 13318 39738 13374 39740
rect 13398 39738 13454 39740
rect 13478 39738 13534 39740
rect 13558 39738 13614 39740
rect 13318 39686 13364 39738
rect 13364 39686 13374 39738
rect 13398 39686 13428 39738
rect 13428 39686 13440 39738
rect 13440 39686 13454 39738
rect 13478 39686 13492 39738
rect 13492 39686 13504 39738
rect 13504 39686 13534 39738
rect 13558 39686 13568 39738
rect 13568 39686 13614 39738
rect 13318 39684 13374 39686
rect 13398 39684 13454 39686
rect 13478 39684 13534 39686
rect 13558 39684 13614 39686
rect 13318 38650 13374 38652
rect 13398 38650 13454 38652
rect 13478 38650 13534 38652
rect 13558 38650 13614 38652
rect 13318 38598 13364 38650
rect 13364 38598 13374 38650
rect 13398 38598 13428 38650
rect 13428 38598 13440 38650
rect 13440 38598 13454 38650
rect 13478 38598 13492 38650
rect 13492 38598 13504 38650
rect 13504 38598 13534 38650
rect 13558 38598 13568 38650
rect 13568 38598 13614 38650
rect 13318 38596 13374 38598
rect 13398 38596 13454 38598
rect 13478 38596 13534 38598
rect 13558 38596 13614 38598
rect 13318 37562 13374 37564
rect 13398 37562 13454 37564
rect 13478 37562 13534 37564
rect 13558 37562 13614 37564
rect 13318 37510 13364 37562
rect 13364 37510 13374 37562
rect 13398 37510 13428 37562
rect 13428 37510 13440 37562
rect 13440 37510 13454 37562
rect 13478 37510 13492 37562
rect 13492 37510 13504 37562
rect 13504 37510 13534 37562
rect 13558 37510 13568 37562
rect 13568 37510 13614 37562
rect 13318 37508 13374 37510
rect 13398 37508 13454 37510
rect 13478 37508 13534 37510
rect 13558 37508 13614 37510
rect 14186 42880 14242 42936
rect 14370 42336 14426 42392
rect 14186 41692 14188 41712
rect 14188 41692 14240 41712
rect 14240 41692 14242 41712
rect 14186 41656 14242 41692
rect 14462 41928 14518 41984
rect 13318 36474 13374 36476
rect 13398 36474 13454 36476
rect 13478 36474 13534 36476
rect 13558 36474 13614 36476
rect 13318 36422 13364 36474
rect 13364 36422 13374 36474
rect 13398 36422 13428 36474
rect 13428 36422 13440 36474
rect 13440 36422 13454 36474
rect 13478 36422 13492 36474
rect 13492 36422 13504 36474
rect 13504 36422 13534 36474
rect 13558 36422 13568 36474
rect 13568 36422 13614 36474
rect 13318 36420 13374 36422
rect 13398 36420 13454 36422
rect 13478 36420 13534 36422
rect 13558 36420 13614 36422
rect 13542 36216 13598 36272
rect 13318 35386 13374 35388
rect 13398 35386 13454 35388
rect 13478 35386 13534 35388
rect 13558 35386 13614 35388
rect 13318 35334 13364 35386
rect 13364 35334 13374 35386
rect 13398 35334 13428 35386
rect 13428 35334 13440 35386
rect 13440 35334 13454 35386
rect 13478 35334 13492 35386
rect 13492 35334 13504 35386
rect 13504 35334 13534 35386
rect 13558 35334 13568 35386
rect 13568 35334 13614 35386
rect 13318 35332 13374 35334
rect 13398 35332 13454 35334
rect 13478 35332 13534 35334
rect 13558 35332 13614 35334
rect 13318 34298 13374 34300
rect 13398 34298 13454 34300
rect 13478 34298 13534 34300
rect 13558 34298 13614 34300
rect 13318 34246 13364 34298
rect 13364 34246 13374 34298
rect 13398 34246 13428 34298
rect 13428 34246 13440 34298
rect 13440 34246 13454 34298
rect 13478 34246 13492 34298
rect 13492 34246 13504 34298
rect 13504 34246 13534 34298
rect 13558 34246 13568 34298
rect 13568 34246 13614 34298
rect 13318 34244 13374 34246
rect 13398 34244 13454 34246
rect 13478 34244 13534 34246
rect 13558 34244 13614 34246
rect 13318 33210 13374 33212
rect 13398 33210 13454 33212
rect 13478 33210 13534 33212
rect 13558 33210 13614 33212
rect 13318 33158 13364 33210
rect 13364 33158 13374 33210
rect 13398 33158 13428 33210
rect 13428 33158 13440 33210
rect 13440 33158 13454 33210
rect 13478 33158 13492 33210
rect 13492 33158 13504 33210
rect 13504 33158 13534 33210
rect 13558 33158 13568 33210
rect 13568 33158 13614 33210
rect 13318 33156 13374 33158
rect 13398 33156 13454 33158
rect 13478 33156 13534 33158
rect 13558 33156 13614 33158
rect 13174 32952 13230 33008
rect 13082 32544 13138 32600
rect 13318 32122 13374 32124
rect 13398 32122 13454 32124
rect 13478 32122 13534 32124
rect 13558 32122 13614 32124
rect 13318 32070 13364 32122
rect 13364 32070 13374 32122
rect 13398 32070 13428 32122
rect 13428 32070 13440 32122
rect 13440 32070 13454 32122
rect 13478 32070 13492 32122
rect 13492 32070 13504 32122
rect 13504 32070 13534 32122
rect 13558 32070 13568 32122
rect 13568 32070 13614 32122
rect 13318 32068 13374 32070
rect 13398 32068 13454 32070
rect 13478 32068 13534 32070
rect 13558 32068 13614 32070
rect 13174 31592 13230 31648
rect 13318 31034 13374 31036
rect 13398 31034 13454 31036
rect 13478 31034 13534 31036
rect 13558 31034 13614 31036
rect 13318 30982 13364 31034
rect 13364 30982 13374 31034
rect 13398 30982 13428 31034
rect 13428 30982 13440 31034
rect 13440 30982 13454 31034
rect 13478 30982 13492 31034
rect 13492 30982 13504 31034
rect 13504 30982 13534 31034
rect 13558 30982 13568 31034
rect 13568 30982 13614 31034
rect 13318 30980 13374 30982
rect 13398 30980 13454 30982
rect 13478 30980 13534 30982
rect 13558 30980 13614 30982
rect 14002 37032 14058 37088
rect 13726 36216 13782 36272
rect 14646 43016 14702 43072
rect 15382 44512 15438 44568
rect 15474 43832 15530 43888
rect 15658 43696 15714 43752
rect 15790 43546 15846 43548
rect 15870 43546 15926 43548
rect 15950 43546 16006 43548
rect 16030 43546 16086 43548
rect 15790 43494 15836 43546
rect 15836 43494 15846 43546
rect 15870 43494 15900 43546
rect 15900 43494 15912 43546
rect 15912 43494 15926 43546
rect 15950 43494 15964 43546
rect 15964 43494 15976 43546
rect 15976 43494 16006 43546
rect 16030 43494 16040 43546
rect 16040 43494 16086 43546
rect 15790 43492 15846 43494
rect 15870 43492 15926 43494
rect 15950 43492 16006 43494
rect 16030 43492 16086 43494
rect 14830 42336 14886 42392
rect 14830 41520 14886 41576
rect 15566 42336 15622 42392
rect 15474 41792 15530 41848
rect 16118 43152 16174 43208
rect 16210 42644 16212 42664
rect 16212 42644 16264 42664
rect 16264 42644 16266 42664
rect 16210 42608 16266 42644
rect 15790 42458 15846 42460
rect 15870 42458 15926 42460
rect 15950 42458 16006 42460
rect 16030 42458 16086 42460
rect 15790 42406 15836 42458
rect 15836 42406 15846 42458
rect 15870 42406 15900 42458
rect 15900 42406 15912 42458
rect 15912 42406 15926 42458
rect 15950 42406 15964 42458
rect 15964 42406 15976 42458
rect 15976 42406 16006 42458
rect 16030 42406 16040 42458
rect 16040 42406 16086 42458
rect 15790 42404 15846 42406
rect 15870 42404 15926 42406
rect 15950 42404 16006 42406
rect 16030 42404 16086 42406
rect 16578 42744 16634 42800
rect 16394 42200 16450 42256
rect 16302 42064 16358 42120
rect 15750 41792 15806 41848
rect 15198 41384 15254 41440
rect 14554 41132 14610 41168
rect 14554 41112 14556 41132
rect 14556 41112 14608 41132
rect 14608 41112 14610 41132
rect 14830 41112 14886 41168
rect 15198 41112 15254 41168
rect 16026 41520 16082 41576
rect 14922 40876 14924 40896
rect 14924 40876 14976 40896
rect 14976 40876 14978 40896
rect 14922 40840 14978 40876
rect 14462 39752 14518 39808
rect 14278 37712 14334 37768
rect 13726 34176 13782 34232
rect 13818 33768 13874 33824
rect 13818 33632 13874 33688
rect 13818 30776 13874 30832
rect 13318 29946 13374 29948
rect 13398 29946 13454 29948
rect 13478 29946 13534 29948
rect 13558 29946 13614 29948
rect 13318 29894 13364 29946
rect 13364 29894 13374 29946
rect 13398 29894 13428 29946
rect 13428 29894 13440 29946
rect 13440 29894 13454 29946
rect 13478 29894 13492 29946
rect 13492 29894 13504 29946
rect 13504 29894 13534 29946
rect 13558 29894 13568 29946
rect 13568 29894 13614 29946
rect 13318 29892 13374 29894
rect 13398 29892 13454 29894
rect 13478 29892 13534 29894
rect 13558 29892 13614 29894
rect 13174 28872 13230 28928
rect 12898 27956 12900 27976
rect 12900 27956 12952 27976
rect 12952 27956 12954 27976
rect 12898 27920 12954 27956
rect 12898 26560 12954 26616
rect 13318 28858 13374 28860
rect 13398 28858 13454 28860
rect 13478 28858 13534 28860
rect 13558 28858 13614 28860
rect 13318 28806 13364 28858
rect 13364 28806 13374 28858
rect 13398 28806 13428 28858
rect 13428 28806 13440 28858
rect 13440 28806 13454 28858
rect 13478 28806 13492 28858
rect 13492 28806 13504 28858
rect 13504 28806 13534 28858
rect 13558 28806 13568 28858
rect 13568 28806 13614 28858
rect 13318 28804 13374 28806
rect 13398 28804 13454 28806
rect 13478 28804 13534 28806
rect 13558 28804 13614 28806
rect 13542 28328 13598 28384
rect 13318 27770 13374 27772
rect 13398 27770 13454 27772
rect 13478 27770 13534 27772
rect 13558 27770 13614 27772
rect 13318 27718 13364 27770
rect 13364 27718 13374 27770
rect 13398 27718 13428 27770
rect 13428 27718 13440 27770
rect 13440 27718 13454 27770
rect 13478 27718 13492 27770
rect 13492 27718 13504 27770
rect 13504 27718 13534 27770
rect 13558 27718 13568 27770
rect 13568 27718 13614 27770
rect 13318 27716 13374 27718
rect 13398 27716 13454 27718
rect 13478 27716 13534 27718
rect 13558 27716 13614 27718
rect 13082 27648 13138 27704
rect 13318 26682 13374 26684
rect 13398 26682 13454 26684
rect 13478 26682 13534 26684
rect 13558 26682 13614 26684
rect 13318 26630 13364 26682
rect 13364 26630 13374 26682
rect 13398 26630 13428 26682
rect 13428 26630 13440 26682
rect 13440 26630 13454 26682
rect 13478 26630 13492 26682
rect 13492 26630 13504 26682
rect 13504 26630 13534 26682
rect 13558 26630 13568 26682
rect 13568 26630 13614 26682
rect 13318 26628 13374 26630
rect 13398 26628 13454 26630
rect 13478 26628 13534 26630
rect 13558 26628 13614 26630
rect 15106 40296 15162 40352
rect 15790 41370 15846 41372
rect 15870 41370 15926 41372
rect 15950 41370 16006 41372
rect 16030 41370 16086 41372
rect 15790 41318 15836 41370
rect 15836 41318 15846 41370
rect 15870 41318 15900 41370
rect 15900 41318 15912 41370
rect 15912 41318 15926 41370
rect 15950 41318 15964 41370
rect 15964 41318 15976 41370
rect 15976 41318 16006 41370
rect 16030 41318 16040 41370
rect 16040 41318 16086 41370
rect 15790 41316 15846 41318
rect 15870 41316 15926 41318
rect 15950 41316 16006 41318
rect 16030 41316 16086 41318
rect 16578 41248 16634 41304
rect 16210 40724 16266 40760
rect 16210 40704 16212 40724
rect 16212 40704 16264 40724
rect 16264 40704 16266 40724
rect 15790 40282 15846 40284
rect 15870 40282 15926 40284
rect 15950 40282 16006 40284
rect 16030 40282 16086 40284
rect 15790 40230 15836 40282
rect 15836 40230 15846 40282
rect 15870 40230 15900 40282
rect 15900 40230 15912 40282
rect 15912 40230 15926 40282
rect 15950 40230 15964 40282
rect 15964 40230 15976 40282
rect 15976 40230 16006 40282
rect 16030 40230 16040 40282
rect 16040 40230 16086 40282
rect 15790 40228 15846 40230
rect 15870 40228 15926 40230
rect 15950 40228 16006 40230
rect 16030 40228 16086 40230
rect 14554 35128 14610 35184
rect 14278 34720 14334 34776
rect 14370 34448 14426 34504
rect 14462 34176 14518 34232
rect 14278 31728 14334 31784
rect 14094 30776 14150 30832
rect 14094 30640 14150 30696
rect 13818 29416 13874 29472
rect 13818 28600 13874 28656
rect 13818 28056 13874 28112
rect 14094 28464 14150 28520
rect 13910 27512 13966 27568
rect 13542 25880 13598 25936
rect 13542 25744 13598 25800
rect 13318 25594 13374 25596
rect 13398 25594 13454 25596
rect 13478 25594 13534 25596
rect 13558 25594 13614 25596
rect 13318 25542 13364 25594
rect 13364 25542 13374 25594
rect 13398 25542 13428 25594
rect 13428 25542 13440 25594
rect 13440 25542 13454 25594
rect 13478 25542 13492 25594
rect 13492 25542 13504 25594
rect 13504 25542 13534 25594
rect 13558 25542 13568 25594
rect 13568 25542 13614 25594
rect 13318 25540 13374 25542
rect 13398 25540 13454 25542
rect 13478 25540 13534 25542
rect 13558 25540 13614 25542
rect 12438 23704 12494 23760
rect 12806 23704 12862 23760
rect 12530 23604 12532 23624
rect 12532 23604 12584 23624
rect 12584 23604 12586 23624
rect 12530 23568 12586 23604
rect 12990 24656 13046 24712
rect 12346 18944 12402 19000
rect 12346 18672 12402 18728
rect 12714 20168 12770 20224
rect 12346 17992 12402 18048
rect 12162 16360 12218 16416
rect 12162 15136 12218 15192
rect 12346 15544 12402 15600
rect 12162 15020 12218 15056
rect 12162 15000 12164 15020
rect 12164 15000 12216 15020
rect 12216 15000 12218 15020
rect 12070 14592 12126 14648
rect 12070 14048 12126 14104
rect 11886 11872 11942 11928
rect 11886 11600 11942 11656
rect 11794 10648 11850 10704
rect 11886 9152 11942 9208
rect 12070 11056 12126 11112
rect 11978 8744 12034 8800
rect 12622 17040 12678 17096
rect 12622 14592 12678 14648
rect 12714 13504 12770 13560
rect 12346 9288 12402 9344
rect 12346 9152 12402 9208
rect 12254 8472 12310 8528
rect 11518 7248 11574 7304
rect 11518 6976 11574 7032
rect 11702 6840 11758 6896
rect 11610 6160 11666 6216
rect 11426 6024 11482 6080
rect 11058 5616 11114 5672
rect 10845 5466 10901 5468
rect 10925 5466 10981 5468
rect 11005 5466 11061 5468
rect 11085 5466 11141 5468
rect 10845 5414 10891 5466
rect 10891 5414 10901 5466
rect 10925 5414 10955 5466
rect 10955 5414 10967 5466
rect 10967 5414 10981 5466
rect 11005 5414 11019 5466
rect 11019 5414 11031 5466
rect 11031 5414 11061 5466
rect 11085 5414 11095 5466
rect 11095 5414 11141 5466
rect 10845 5412 10901 5414
rect 10925 5412 10981 5414
rect 11005 5412 11061 5414
rect 11085 5412 11141 5414
rect 10782 5208 10838 5264
rect 10874 4936 10930 4992
rect 10874 4664 10930 4720
rect 11058 5072 11114 5128
rect 11058 4528 11114 4584
rect 10845 4378 10901 4380
rect 10925 4378 10981 4380
rect 11005 4378 11061 4380
rect 11085 4378 11141 4380
rect 10845 4326 10891 4378
rect 10891 4326 10901 4378
rect 10925 4326 10955 4378
rect 10955 4326 10967 4378
rect 10967 4326 10981 4378
rect 11005 4326 11019 4378
rect 11019 4326 11031 4378
rect 11031 4326 11061 4378
rect 11085 4326 11095 4378
rect 11095 4326 11141 4378
rect 10845 4324 10901 4326
rect 10925 4324 10981 4326
rect 11005 4324 11061 4326
rect 11085 4324 11141 4326
rect 10506 3576 10562 3632
rect 10138 2488 10194 2544
rect 10414 2932 10416 2952
rect 10416 2932 10468 2952
rect 10468 2932 10470 2952
rect 10414 2896 10470 2932
rect 10414 2796 10416 2816
rect 10416 2796 10468 2816
rect 10468 2796 10470 2816
rect 10414 2760 10470 2796
rect 11150 3984 11206 4040
rect 11334 5072 11390 5128
rect 11518 5480 11574 5536
rect 11794 6160 11850 6216
rect 11702 5364 11758 5400
rect 11702 5344 11704 5364
rect 11704 5344 11756 5364
rect 11756 5344 11758 5364
rect 12162 7520 12218 7576
rect 12346 8200 12402 8256
rect 13910 25880 13966 25936
rect 13818 24928 13874 24984
rect 13318 24506 13374 24508
rect 13398 24506 13454 24508
rect 13478 24506 13534 24508
rect 13558 24506 13614 24508
rect 13318 24454 13364 24506
rect 13364 24454 13374 24506
rect 13398 24454 13428 24506
rect 13428 24454 13440 24506
rect 13440 24454 13454 24506
rect 13478 24454 13492 24506
rect 13492 24454 13504 24506
rect 13504 24454 13534 24506
rect 13558 24454 13568 24506
rect 13568 24454 13614 24506
rect 13318 24452 13374 24454
rect 13398 24452 13454 24454
rect 13478 24452 13534 24454
rect 13558 24452 13614 24454
rect 13174 23704 13230 23760
rect 13318 23418 13374 23420
rect 13398 23418 13454 23420
rect 13478 23418 13534 23420
rect 13558 23418 13614 23420
rect 13318 23366 13364 23418
rect 13364 23366 13374 23418
rect 13398 23366 13428 23418
rect 13428 23366 13440 23418
rect 13440 23366 13454 23418
rect 13478 23366 13492 23418
rect 13492 23366 13504 23418
rect 13504 23366 13534 23418
rect 13558 23366 13568 23418
rect 13568 23366 13614 23418
rect 13318 23364 13374 23366
rect 13398 23364 13454 23366
rect 13478 23364 13534 23366
rect 13558 23364 13614 23366
rect 12990 22480 13046 22536
rect 13318 22330 13374 22332
rect 13398 22330 13454 22332
rect 13478 22330 13534 22332
rect 13558 22330 13614 22332
rect 13318 22278 13364 22330
rect 13364 22278 13374 22330
rect 13398 22278 13428 22330
rect 13428 22278 13440 22330
rect 13440 22278 13454 22330
rect 13478 22278 13492 22330
rect 13492 22278 13504 22330
rect 13504 22278 13534 22330
rect 13558 22278 13568 22330
rect 13568 22278 13614 22330
rect 13318 22276 13374 22278
rect 13398 22276 13454 22278
rect 13478 22276 13534 22278
rect 13558 22276 13614 22278
rect 13174 22072 13230 22128
rect 12990 20984 13046 21040
rect 13634 21936 13690 21992
rect 13318 21242 13374 21244
rect 13398 21242 13454 21244
rect 13478 21242 13534 21244
rect 13558 21242 13614 21244
rect 13318 21190 13364 21242
rect 13364 21190 13374 21242
rect 13398 21190 13428 21242
rect 13428 21190 13440 21242
rect 13440 21190 13454 21242
rect 13478 21190 13492 21242
rect 13492 21190 13504 21242
rect 13504 21190 13534 21242
rect 13558 21190 13568 21242
rect 13568 21190 13614 21242
rect 13318 21188 13374 21190
rect 13398 21188 13454 21190
rect 13478 21188 13534 21190
rect 13558 21188 13614 21190
rect 13542 21020 13544 21040
rect 13544 21020 13596 21040
rect 13596 21020 13598 21040
rect 13542 20984 13598 21020
rect 13542 20712 13598 20768
rect 13318 20154 13374 20156
rect 13398 20154 13454 20156
rect 13478 20154 13534 20156
rect 13558 20154 13614 20156
rect 13318 20102 13364 20154
rect 13364 20102 13374 20154
rect 13398 20102 13428 20154
rect 13428 20102 13440 20154
rect 13440 20102 13454 20154
rect 13478 20102 13492 20154
rect 13492 20102 13504 20154
rect 13504 20102 13534 20154
rect 13558 20102 13568 20154
rect 13568 20102 13614 20154
rect 13318 20100 13374 20102
rect 13398 20100 13454 20102
rect 13478 20100 13534 20102
rect 13558 20100 13614 20102
rect 13358 19488 13414 19544
rect 13318 19066 13374 19068
rect 13398 19066 13454 19068
rect 13478 19066 13534 19068
rect 13558 19066 13614 19068
rect 13318 19014 13364 19066
rect 13364 19014 13374 19066
rect 13398 19014 13428 19066
rect 13428 19014 13440 19066
rect 13440 19014 13454 19066
rect 13478 19014 13492 19066
rect 13492 19014 13504 19066
rect 13504 19014 13534 19066
rect 13558 19014 13568 19066
rect 13568 19014 13614 19066
rect 13318 19012 13374 19014
rect 13398 19012 13454 19014
rect 13478 19012 13534 19014
rect 13558 19012 13614 19014
rect 13910 23180 13966 23216
rect 13910 23160 13912 23180
rect 13912 23160 13964 23180
rect 13964 23160 13966 23180
rect 13910 22344 13966 22400
rect 13818 21256 13874 21312
rect 13634 18264 13690 18320
rect 13318 17978 13374 17980
rect 13398 17978 13454 17980
rect 13478 17978 13534 17980
rect 13558 17978 13614 17980
rect 13318 17926 13364 17978
rect 13364 17926 13374 17978
rect 13398 17926 13428 17978
rect 13428 17926 13440 17978
rect 13440 17926 13454 17978
rect 13478 17926 13492 17978
rect 13492 17926 13504 17978
rect 13504 17926 13534 17978
rect 13558 17926 13568 17978
rect 13568 17926 13614 17978
rect 13318 17924 13374 17926
rect 13398 17924 13454 17926
rect 13478 17924 13534 17926
rect 13558 17924 13614 17926
rect 12898 14864 12954 14920
rect 13318 16890 13374 16892
rect 13398 16890 13454 16892
rect 13478 16890 13534 16892
rect 13558 16890 13614 16892
rect 13318 16838 13364 16890
rect 13364 16838 13374 16890
rect 13398 16838 13428 16890
rect 13428 16838 13440 16890
rect 13440 16838 13454 16890
rect 13478 16838 13492 16890
rect 13492 16838 13504 16890
rect 13504 16838 13534 16890
rect 13558 16838 13568 16890
rect 13568 16838 13614 16890
rect 13318 16836 13374 16838
rect 13398 16836 13454 16838
rect 13478 16836 13534 16838
rect 13558 16836 13614 16838
rect 13174 15816 13230 15872
rect 13318 15802 13374 15804
rect 13398 15802 13454 15804
rect 13478 15802 13534 15804
rect 13558 15802 13614 15804
rect 13318 15750 13364 15802
rect 13364 15750 13374 15802
rect 13398 15750 13428 15802
rect 13428 15750 13440 15802
rect 13440 15750 13454 15802
rect 13478 15750 13492 15802
rect 13492 15750 13504 15802
rect 13504 15750 13534 15802
rect 13558 15750 13568 15802
rect 13568 15750 13614 15802
rect 13318 15748 13374 15750
rect 13398 15748 13454 15750
rect 13478 15748 13534 15750
rect 13558 15748 13614 15750
rect 14186 25880 14242 25936
rect 14738 34176 14794 34232
rect 16210 39208 16266 39264
rect 15790 39194 15846 39196
rect 15870 39194 15926 39196
rect 15950 39194 16006 39196
rect 16030 39194 16086 39196
rect 15790 39142 15836 39194
rect 15836 39142 15846 39194
rect 15870 39142 15900 39194
rect 15900 39142 15912 39194
rect 15912 39142 15926 39194
rect 15950 39142 15964 39194
rect 15964 39142 15976 39194
rect 15976 39142 16006 39194
rect 16030 39142 16040 39194
rect 16040 39142 16086 39194
rect 15790 39140 15846 39142
rect 15870 39140 15926 39142
rect 15950 39140 16006 39142
rect 16030 39140 16086 39142
rect 15790 38106 15846 38108
rect 15870 38106 15926 38108
rect 15950 38106 16006 38108
rect 16030 38106 16086 38108
rect 15790 38054 15836 38106
rect 15836 38054 15846 38106
rect 15870 38054 15900 38106
rect 15900 38054 15912 38106
rect 15912 38054 15926 38106
rect 15950 38054 15964 38106
rect 15964 38054 15976 38106
rect 15976 38054 16006 38106
rect 16030 38054 16040 38106
rect 16040 38054 16086 38106
rect 15790 38052 15846 38054
rect 15870 38052 15926 38054
rect 15950 38052 16006 38054
rect 16030 38052 16086 38054
rect 15658 37984 15714 38040
rect 15290 37712 15346 37768
rect 15790 37018 15846 37020
rect 15870 37018 15926 37020
rect 15950 37018 16006 37020
rect 16030 37018 16086 37020
rect 15790 36966 15836 37018
rect 15836 36966 15846 37018
rect 15870 36966 15900 37018
rect 15900 36966 15912 37018
rect 15912 36966 15926 37018
rect 15950 36966 15964 37018
rect 15964 36966 15976 37018
rect 15976 36966 16006 37018
rect 16030 36966 16040 37018
rect 16040 36966 16086 37018
rect 15790 36964 15846 36966
rect 15870 36964 15926 36966
rect 15950 36964 16006 36966
rect 16030 36964 16086 36966
rect 15106 35808 15162 35864
rect 15566 35944 15622 36000
rect 15382 35672 15438 35728
rect 15790 35930 15846 35932
rect 15870 35930 15926 35932
rect 15950 35930 16006 35932
rect 16030 35930 16086 35932
rect 15790 35878 15836 35930
rect 15836 35878 15846 35930
rect 15870 35878 15900 35930
rect 15900 35878 15912 35930
rect 15912 35878 15926 35930
rect 15950 35878 15964 35930
rect 15964 35878 15976 35930
rect 15976 35878 16006 35930
rect 16030 35878 16040 35930
rect 16040 35878 16086 35930
rect 15790 35876 15846 35878
rect 15870 35876 15926 35878
rect 15950 35876 16006 35878
rect 16030 35876 16086 35878
rect 15198 34176 15254 34232
rect 15014 33768 15070 33824
rect 14830 32816 14886 32872
rect 14738 32000 14794 32056
rect 14738 31592 14794 31648
rect 15842 35672 15898 35728
rect 15474 34720 15530 34776
rect 15382 34584 15438 34640
rect 15658 35128 15714 35184
rect 15790 34842 15846 34844
rect 15870 34842 15926 34844
rect 15950 34842 16006 34844
rect 16030 34842 16086 34844
rect 15790 34790 15836 34842
rect 15836 34790 15846 34842
rect 15870 34790 15900 34842
rect 15900 34790 15912 34842
rect 15912 34790 15926 34842
rect 15950 34790 15964 34842
rect 15964 34790 15976 34842
rect 15976 34790 16006 34842
rect 16030 34790 16040 34842
rect 16040 34790 16086 34842
rect 15790 34788 15846 34790
rect 15870 34788 15926 34790
rect 15950 34788 16006 34790
rect 16030 34788 16086 34790
rect 15790 33754 15846 33756
rect 15870 33754 15926 33756
rect 15950 33754 16006 33756
rect 16030 33754 16086 33756
rect 15790 33702 15836 33754
rect 15836 33702 15846 33754
rect 15870 33702 15900 33754
rect 15900 33702 15912 33754
rect 15912 33702 15926 33754
rect 15950 33702 15964 33754
rect 15964 33702 15976 33754
rect 15976 33702 16006 33754
rect 16030 33702 16040 33754
rect 16040 33702 16086 33754
rect 15790 33700 15846 33702
rect 15870 33700 15926 33702
rect 15950 33700 16006 33702
rect 16030 33700 16086 33702
rect 15658 33632 15714 33688
rect 15106 31884 15162 31920
rect 15106 31864 15108 31884
rect 15108 31864 15160 31884
rect 15160 31864 15162 31884
rect 15014 31728 15070 31784
rect 14646 30912 14702 30968
rect 16210 32952 16266 33008
rect 14094 23568 14150 23624
rect 15106 29688 15162 29744
rect 14738 26696 14794 26752
rect 14462 25064 14518 25120
rect 14462 24248 14518 24304
rect 14002 20168 14058 20224
rect 14002 19216 14058 19272
rect 14278 18400 14334 18456
rect 13318 14714 13374 14716
rect 13398 14714 13454 14716
rect 13478 14714 13534 14716
rect 13558 14714 13614 14716
rect 13318 14662 13364 14714
rect 13364 14662 13374 14714
rect 13398 14662 13428 14714
rect 13428 14662 13440 14714
rect 13440 14662 13454 14714
rect 13478 14662 13492 14714
rect 13492 14662 13504 14714
rect 13504 14662 13534 14714
rect 13558 14662 13568 14714
rect 13568 14662 13614 14714
rect 13318 14660 13374 14662
rect 13398 14660 13454 14662
rect 13478 14660 13534 14662
rect 13558 14660 13614 14662
rect 13318 13626 13374 13628
rect 13398 13626 13454 13628
rect 13478 13626 13534 13628
rect 13558 13626 13614 13628
rect 13318 13574 13364 13626
rect 13364 13574 13374 13626
rect 13398 13574 13428 13626
rect 13428 13574 13440 13626
rect 13440 13574 13454 13626
rect 13478 13574 13492 13626
rect 13492 13574 13504 13626
rect 13504 13574 13534 13626
rect 13558 13574 13568 13626
rect 13568 13574 13614 13626
rect 13318 13572 13374 13574
rect 13398 13572 13454 13574
rect 13478 13572 13534 13574
rect 13558 13572 13614 13574
rect 13082 11328 13138 11384
rect 12806 10376 12862 10432
rect 13318 12538 13374 12540
rect 13398 12538 13454 12540
rect 13478 12538 13534 12540
rect 13558 12538 13614 12540
rect 13318 12486 13364 12538
rect 13364 12486 13374 12538
rect 13398 12486 13428 12538
rect 13428 12486 13440 12538
rect 13440 12486 13454 12538
rect 13478 12486 13492 12538
rect 13492 12486 13504 12538
rect 13504 12486 13534 12538
rect 13558 12486 13568 12538
rect 13568 12486 13614 12538
rect 13318 12484 13374 12486
rect 13398 12484 13454 12486
rect 13478 12484 13534 12486
rect 13558 12484 13614 12486
rect 14278 15136 14334 15192
rect 14738 23568 14794 23624
rect 14646 22616 14702 22672
rect 14738 22072 14794 22128
rect 14646 21936 14702 21992
rect 15198 29008 15254 29064
rect 15198 28600 15254 28656
rect 15014 24112 15070 24168
rect 15790 32666 15846 32668
rect 15870 32666 15926 32668
rect 15950 32666 16006 32668
rect 16030 32666 16086 32668
rect 15790 32614 15836 32666
rect 15836 32614 15846 32666
rect 15870 32614 15900 32666
rect 15900 32614 15912 32666
rect 15912 32614 15926 32666
rect 15950 32614 15964 32666
rect 15964 32614 15976 32666
rect 15976 32614 16006 32666
rect 16030 32614 16040 32666
rect 16040 32614 16086 32666
rect 15790 32612 15846 32614
rect 15870 32612 15926 32614
rect 15950 32612 16006 32614
rect 16030 32612 16086 32614
rect 17038 41112 17094 41168
rect 16486 39208 16542 39264
rect 16946 40060 16948 40080
rect 16948 40060 17000 40080
rect 17000 40060 17002 40080
rect 16946 40024 17002 40060
rect 16394 34584 16450 34640
rect 17774 42608 17830 42664
rect 17406 41656 17462 41712
rect 17682 42064 17738 42120
rect 17222 39072 17278 39128
rect 17130 38664 17186 38720
rect 17314 37440 17370 37496
rect 17038 36760 17094 36816
rect 16946 35264 17002 35320
rect 17314 35808 17370 35864
rect 15790 31578 15846 31580
rect 15870 31578 15926 31580
rect 15950 31578 16006 31580
rect 16030 31578 16086 31580
rect 15790 31526 15836 31578
rect 15836 31526 15846 31578
rect 15870 31526 15900 31578
rect 15900 31526 15912 31578
rect 15912 31526 15926 31578
rect 15950 31526 15964 31578
rect 15964 31526 15976 31578
rect 15976 31526 16006 31578
rect 16030 31526 16040 31578
rect 16040 31526 16086 31578
rect 15790 31524 15846 31526
rect 15870 31524 15926 31526
rect 15950 31524 16006 31526
rect 16030 31524 16086 31526
rect 15474 31320 15530 31376
rect 15658 31320 15714 31376
rect 16302 31048 16358 31104
rect 15474 30096 15530 30152
rect 15658 30640 15714 30696
rect 15790 30490 15846 30492
rect 15870 30490 15926 30492
rect 15950 30490 16006 30492
rect 16030 30490 16086 30492
rect 15790 30438 15836 30490
rect 15836 30438 15846 30490
rect 15870 30438 15900 30490
rect 15900 30438 15912 30490
rect 15912 30438 15926 30490
rect 15950 30438 15964 30490
rect 15964 30438 15976 30490
rect 15976 30438 16006 30490
rect 16030 30438 16040 30490
rect 16040 30438 16086 30490
rect 15790 30436 15846 30438
rect 15870 30436 15926 30438
rect 15950 30436 16006 30438
rect 16030 30436 16086 30438
rect 15790 29402 15846 29404
rect 15870 29402 15926 29404
rect 15950 29402 16006 29404
rect 16030 29402 16086 29404
rect 15790 29350 15836 29402
rect 15836 29350 15846 29402
rect 15870 29350 15900 29402
rect 15900 29350 15912 29402
rect 15912 29350 15926 29402
rect 15950 29350 15964 29402
rect 15964 29350 15976 29402
rect 15976 29350 16006 29402
rect 16030 29350 16040 29402
rect 16040 29350 16086 29402
rect 15790 29348 15846 29350
rect 15870 29348 15926 29350
rect 15950 29348 16006 29350
rect 16030 29348 16086 29350
rect 15790 28314 15846 28316
rect 15870 28314 15926 28316
rect 15950 28314 16006 28316
rect 16030 28314 16086 28316
rect 15790 28262 15836 28314
rect 15836 28262 15846 28314
rect 15870 28262 15900 28314
rect 15900 28262 15912 28314
rect 15912 28262 15926 28314
rect 15950 28262 15964 28314
rect 15964 28262 15976 28314
rect 15976 28262 16006 28314
rect 16030 28262 16040 28314
rect 16040 28262 16086 28314
rect 15790 28260 15846 28262
rect 15870 28260 15926 28262
rect 15950 28260 16006 28262
rect 16030 28260 16086 28262
rect 15658 27648 15714 27704
rect 15382 24112 15438 24168
rect 15198 23568 15254 23624
rect 15014 21664 15070 21720
rect 15790 27226 15846 27228
rect 15870 27226 15926 27228
rect 15950 27226 16006 27228
rect 16030 27226 16086 27228
rect 15790 27174 15836 27226
rect 15836 27174 15846 27226
rect 15870 27174 15900 27226
rect 15900 27174 15912 27226
rect 15912 27174 15926 27226
rect 15950 27174 15964 27226
rect 15964 27174 15976 27226
rect 15976 27174 16006 27226
rect 16030 27174 16040 27226
rect 16040 27174 16086 27226
rect 15790 27172 15846 27174
rect 15870 27172 15926 27174
rect 15950 27172 16006 27174
rect 16030 27172 16086 27174
rect 15566 25100 15568 25120
rect 15568 25100 15620 25120
rect 15620 25100 15622 25120
rect 15566 25064 15622 25100
rect 15790 26138 15846 26140
rect 15870 26138 15926 26140
rect 15950 26138 16006 26140
rect 16030 26138 16086 26140
rect 15790 26086 15836 26138
rect 15836 26086 15846 26138
rect 15870 26086 15900 26138
rect 15900 26086 15912 26138
rect 15912 26086 15926 26138
rect 15950 26086 15964 26138
rect 15964 26086 15976 26138
rect 15976 26086 16006 26138
rect 16030 26086 16040 26138
rect 16040 26086 16086 26138
rect 15790 26084 15846 26086
rect 15870 26084 15926 26086
rect 15950 26084 16006 26086
rect 16030 26084 16086 26086
rect 16210 30368 16266 30424
rect 17130 33360 17186 33416
rect 16210 26152 16266 26208
rect 16210 25200 16266 25256
rect 15790 25050 15846 25052
rect 15870 25050 15926 25052
rect 15950 25050 16006 25052
rect 16030 25050 16086 25052
rect 15790 24998 15836 25050
rect 15836 24998 15846 25050
rect 15870 24998 15900 25050
rect 15900 24998 15912 25050
rect 15912 24998 15926 25050
rect 15950 24998 15964 25050
rect 15964 24998 15976 25050
rect 15976 24998 16006 25050
rect 16030 24998 16040 25050
rect 16040 24998 16086 25050
rect 15790 24996 15846 24998
rect 15870 24996 15926 24998
rect 15950 24996 16006 24998
rect 16030 24996 16086 24998
rect 15790 23962 15846 23964
rect 15870 23962 15926 23964
rect 15950 23962 16006 23964
rect 16030 23962 16086 23964
rect 15790 23910 15836 23962
rect 15836 23910 15846 23962
rect 15870 23910 15900 23962
rect 15900 23910 15912 23962
rect 15912 23910 15926 23962
rect 15950 23910 15964 23962
rect 15964 23910 15976 23962
rect 15976 23910 16006 23962
rect 16030 23910 16040 23962
rect 16040 23910 16086 23962
rect 15790 23908 15846 23910
rect 15870 23908 15926 23910
rect 15950 23908 16006 23910
rect 16030 23908 16086 23910
rect 15750 23568 15806 23624
rect 14922 20848 14978 20904
rect 14922 19896 14978 19952
rect 15290 19760 15346 19816
rect 14922 18828 14978 18864
rect 14922 18808 14924 18828
rect 14924 18808 14976 18828
rect 14976 18808 14978 18828
rect 14462 16088 14518 16144
rect 14278 14320 14334 14376
rect 13818 12416 13874 12472
rect 13266 11872 13322 11928
rect 13318 11450 13374 11452
rect 13398 11450 13454 11452
rect 13478 11450 13534 11452
rect 13558 11450 13614 11452
rect 13318 11398 13364 11450
rect 13364 11398 13374 11450
rect 13398 11398 13428 11450
rect 13428 11398 13440 11450
rect 13440 11398 13454 11450
rect 13478 11398 13492 11450
rect 13492 11398 13504 11450
rect 13504 11398 13534 11450
rect 13558 11398 13568 11450
rect 13568 11398 13614 11450
rect 13318 11396 13374 11398
rect 13398 11396 13454 11398
rect 13478 11396 13534 11398
rect 13558 11396 13614 11398
rect 13318 10362 13374 10364
rect 13398 10362 13454 10364
rect 13478 10362 13534 10364
rect 13558 10362 13614 10364
rect 13318 10310 13364 10362
rect 13364 10310 13374 10362
rect 13398 10310 13428 10362
rect 13428 10310 13440 10362
rect 13440 10310 13454 10362
rect 13478 10310 13492 10362
rect 13492 10310 13504 10362
rect 13504 10310 13534 10362
rect 13558 10310 13568 10362
rect 13568 10310 13614 10362
rect 13318 10308 13374 10310
rect 13398 10308 13454 10310
rect 13478 10308 13534 10310
rect 13558 10308 13614 10310
rect 12530 9832 12586 9888
rect 12806 9832 12862 9888
rect 12530 8064 12586 8120
rect 13082 9832 13138 9888
rect 12898 8880 12954 8936
rect 12806 8472 12862 8528
rect 12530 7792 12586 7848
rect 12254 7248 12310 7304
rect 12714 7112 12770 7168
rect 12622 6976 12678 7032
rect 12714 6740 12716 6760
rect 12716 6740 12768 6760
rect 12768 6740 12770 6760
rect 12714 6704 12770 6740
rect 12346 6316 12402 6352
rect 12346 6296 12348 6316
rect 12348 6296 12400 6316
rect 12400 6296 12402 6316
rect 12346 6160 12402 6216
rect 12806 6432 12862 6488
rect 12346 5888 12402 5944
rect 11610 5072 11666 5128
rect 11702 4800 11758 4856
rect 11426 4528 11482 4584
rect 11610 4528 11666 4584
rect 11242 3576 11298 3632
rect 10690 3304 10746 3360
rect 10845 3290 10901 3292
rect 10925 3290 10981 3292
rect 11005 3290 11061 3292
rect 11085 3290 11141 3292
rect 10845 3238 10891 3290
rect 10891 3238 10901 3290
rect 10925 3238 10955 3290
rect 10955 3238 10967 3290
rect 10967 3238 10981 3290
rect 11005 3238 11019 3290
rect 11019 3238 11031 3290
rect 11031 3238 11061 3290
rect 11085 3238 11095 3290
rect 11095 3238 11141 3290
rect 10845 3236 10901 3238
rect 10925 3236 10981 3238
rect 11005 3236 11061 3238
rect 11085 3236 11141 3238
rect 10782 3052 10838 3088
rect 10782 3032 10784 3052
rect 10784 3032 10836 3052
rect 10836 3032 10838 3052
rect 10690 2796 10692 2816
rect 10692 2796 10744 2816
rect 10744 2796 10746 2816
rect 10690 2760 10746 2796
rect 10046 1128 10102 1184
rect 10230 1128 10286 1184
rect 10046 992 10102 1048
rect 10046 856 10102 912
rect 10230 992 10286 1048
rect 10230 740 10286 776
rect 10230 720 10232 740
rect 10232 720 10284 740
rect 10284 720 10286 740
rect 7470 40 7526 96
rect 8574 40 8630 96
rect 10874 2624 10930 2680
rect 11058 2896 11114 2952
rect 11150 2760 11206 2816
rect 11150 2388 11152 2408
rect 11152 2388 11204 2408
rect 11204 2388 11206 2408
rect 11150 2352 11206 2388
rect 10845 2202 10901 2204
rect 10925 2202 10981 2204
rect 11005 2202 11061 2204
rect 11085 2202 11141 2204
rect 10845 2150 10891 2202
rect 10891 2150 10901 2202
rect 10925 2150 10955 2202
rect 10955 2150 10967 2202
rect 10967 2150 10981 2202
rect 11005 2150 11019 2202
rect 11019 2150 11031 2202
rect 11031 2150 11061 2202
rect 11085 2150 11095 2202
rect 11095 2150 11141 2202
rect 10845 2148 10901 2150
rect 10925 2148 10981 2150
rect 11005 2148 11061 2150
rect 11085 2148 11141 2150
rect 10874 1536 10930 1592
rect 11886 5072 11942 5128
rect 12530 5616 12586 5672
rect 12714 5752 12770 5808
rect 12070 4800 12126 4856
rect 11978 4392 12034 4448
rect 11886 4256 11942 4312
rect 11610 3576 11666 3632
rect 11518 3304 11574 3360
rect 11794 3848 11850 3904
rect 11702 2896 11758 2952
rect 11426 2252 11428 2272
rect 11428 2252 11480 2272
rect 11480 2252 11482 2272
rect 11426 2216 11482 2252
rect 12990 8472 13046 8528
rect 12990 6704 13046 6760
rect 13318 9274 13374 9276
rect 13398 9274 13454 9276
rect 13478 9274 13534 9276
rect 13558 9274 13614 9276
rect 13318 9222 13364 9274
rect 13364 9222 13374 9274
rect 13398 9222 13428 9274
rect 13428 9222 13440 9274
rect 13440 9222 13454 9274
rect 13478 9222 13492 9274
rect 13492 9222 13504 9274
rect 13504 9222 13534 9274
rect 13558 9222 13568 9274
rect 13568 9222 13614 9274
rect 13318 9220 13374 9222
rect 13398 9220 13454 9222
rect 13478 9220 13534 9222
rect 13558 9220 13614 9222
rect 13910 11872 13966 11928
rect 13726 11464 13782 11520
rect 13726 10376 13782 10432
rect 14094 12300 14150 12336
rect 14094 12280 14096 12300
rect 14096 12280 14148 12300
rect 14148 12280 14150 12300
rect 14094 11328 14150 11384
rect 14094 10920 14150 10976
rect 14094 10784 14150 10840
rect 14554 15272 14610 15328
rect 15474 19760 15530 19816
rect 15790 22874 15846 22876
rect 15870 22874 15926 22876
rect 15950 22874 16006 22876
rect 16030 22874 16086 22876
rect 15790 22822 15836 22874
rect 15836 22822 15846 22874
rect 15870 22822 15900 22874
rect 15900 22822 15912 22874
rect 15912 22822 15926 22874
rect 15950 22822 15964 22874
rect 15964 22822 15976 22874
rect 15976 22822 16006 22874
rect 16030 22822 16040 22874
rect 16040 22822 16086 22874
rect 15790 22820 15846 22822
rect 15870 22820 15926 22822
rect 15950 22820 16006 22822
rect 16030 22820 16086 22822
rect 15790 21786 15846 21788
rect 15870 21786 15926 21788
rect 15950 21786 16006 21788
rect 16030 21786 16086 21788
rect 15790 21734 15836 21786
rect 15836 21734 15846 21786
rect 15870 21734 15900 21786
rect 15900 21734 15912 21786
rect 15912 21734 15926 21786
rect 15950 21734 15964 21786
rect 15964 21734 15976 21786
rect 15976 21734 16006 21786
rect 16030 21734 16040 21786
rect 16040 21734 16086 21786
rect 15790 21732 15846 21734
rect 15870 21732 15926 21734
rect 15950 21732 16006 21734
rect 16030 21732 16086 21734
rect 16578 23296 16634 23352
rect 16946 31320 17002 31376
rect 17314 34992 17370 35048
rect 17130 32408 17186 32464
rect 17406 31864 17462 31920
rect 17130 30776 17186 30832
rect 17038 29144 17094 29200
rect 17406 29008 17462 29064
rect 16854 26560 16910 26616
rect 16762 25200 16818 25256
rect 16946 24792 17002 24848
rect 16854 22208 16910 22264
rect 16486 21392 16542 21448
rect 16302 20984 16358 21040
rect 15790 20698 15846 20700
rect 15870 20698 15926 20700
rect 15950 20698 16006 20700
rect 16030 20698 16086 20700
rect 15790 20646 15836 20698
rect 15836 20646 15846 20698
rect 15870 20646 15900 20698
rect 15900 20646 15912 20698
rect 15912 20646 15926 20698
rect 15950 20646 15964 20698
rect 15964 20646 15976 20698
rect 15976 20646 16006 20698
rect 16030 20646 16040 20698
rect 16040 20646 16086 20698
rect 15790 20644 15846 20646
rect 15870 20644 15926 20646
rect 15950 20644 16006 20646
rect 16030 20644 16086 20646
rect 15790 19610 15846 19612
rect 15870 19610 15926 19612
rect 15950 19610 16006 19612
rect 16030 19610 16086 19612
rect 15790 19558 15836 19610
rect 15836 19558 15846 19610
rect 15870 19558 15900 19610
rect 15900 19558 15912 19610
rect 15912 19558 15926 19610
rect 15950 19558 15964 19610
rect 15964 19558 15976 19610
rect 15976 19558 16006 19610
rect 16030 19558 16040 19610
rect 16040 19558 16086 19610
rect 15790 19556 15846 19558
rect 15870 19556 15926 19558
rect 15950 19556 16006 19558
rect 16030 19556 16086 19558
rect 14922 15272 14978 15328
rect 15014 14456 15070 14512
rect 14830 14320 14886 14376
rect 15198 16496 15254 16552
rect 15474 18128 15530 18184
rect 15790 18522 15846 18524
rect 15870 18522 15926 18524
rect 15950 18522 16006 18524
rect 16030 18522 16086 18524
rect 15790 18470 15836 18522
rect 15836 18470 15846 18522
rect 15870 18470 15900 18522
rect 15900 18470 15912 18522
rect 15912 18470 15926 18522
rect 15950 18470 15964 18522
rect 15964 18470 15976 18522
rect 15976 18470 16006 18522
rect 16030 18470 16040 18522
rect 16040 18470 16086 18522
rect 15790 18468 15846 18470
rect 15870 18468 15926 18470
rect 15950 18468 16006 18470
rect 16030 18468 16086 18470
rect 15382 17076 15384 17096
rect 15384 17076 15436 17096
rect 15436 17076 15438 17096
rect 15382 17040 15438 17076
rect 15198 15136 15254 15192
rect 14738 12552 14794 12608
rect 14646 11736 14702 11792
rect 14002 9288 14058 9344
rect 13910 9152 13966 9208
rect 13318 8186 13374 8188
rect 13398 8186 13454 8188
rect 13478 8186 13534 8188
rect 13558 8186 13614 8188
rect 13318 8134 13364 8186
rect 13364 8134 13374 8186
rect 13398 8134 13428 8186
rect 13428 8134 13440 8186
rect 13440 8134 13454 8186
rect 13478 8134 13492 8186
rect 13492 8134 13504 8186
rect 13504 8134 13534 8186
rect 13558 8134 13568 8186
rect 13568 8134 13614 8186
rect 13318 8132 13374 8134
rect 13398 8132 13454 8134
rect 13478 8132 13534 8134
rect 13558 8132 13614 8134
rect 14002 8200 14058 8256
rect 14002 8064 14058 8120
rect 13318 7098 13374 7100
rect 13398 7098 13454 7100
rect 13478 7098 13534 7100
rect 13558 7098 13614 7100
rect 13318 7046 13364 7098
rect 13364 7046 13374 7098
rect 13398 7046 13428 7098
rect 13428 7046 13440 7098
rect 13440 7046 13454 7098
rect 13478 7046 13492 7098
rect 13492 7046 13504 7098
rect 13504 7046 13534 7098
rect 13558 7046 13568 7098
rect 13568 7046 13614 7098
rect 13318 7044 13374 7046
rect 13398 7044 13454 7046
rect 13478 7044 13534 7046
rect 13558 7044 13614 7046
rect 13082 6296 13138 6352
rect 12898 6024 12954 6080
rect 13634 6296 13690 6352
rect 13318 6010 13374 6012
rect 13398 6010 13454 6012
rect 13478 6010 13534 6012
rect 13558 6010 13614 6012
rect 13318 5958 13364 6010
rect 13364 5958 13374 6010
rect 13398 5958 13428 6010
rect 13428 5958 13440 6010
rect 13440 5958 13454 6010
rect 13478 5958 13492 6010
rect 13492 5958 13504 6010
rect 13504 5958 13534 6010
rect 13558 5958 13568 6010
rect 13568 5958 13614 6010
rect 13318 5956 13374 5958
rect 13398 5956 13454 5958
rect 13478 5956 13534 5958
rect 13558 5956 13614 5958
rect 12898 5344 12954 5400
rect 12438 4800 12494 4856
rect 12162 4664 12218 4720
rect 12346 4664 12402 4720
rect 12254 4256 12310 4312
rect 12806 5072 12862 5128
rect 12714 4800 12770 4856
rect 13542 5344 13598 5400
rect 13910 7384 13966 7440
rect 13910 7112 13966 7168
rect 14186 9460 14188 9480
rect 14188 9460 14240 9480
rect 14240 9460 14242 9480
rect 14186 9424 14242 9460
rect 14278 9288 14334 9344
rect 14462 10104 14518 10160
rect 14646 10104 14702 10160
rect 14554 9152 14610 9208
rect 14278 7928 14334 7984
rect 14186 6976 14242 7032
rect 14094 6568 14150 6624
rect 13910 6024 13966 6080
rect 14002 5888 14058 5944
rect 14186 5888 14242 5944
rect 15106 14320 15162 14376
rect 15106 13096 15162 13152
rect 15106 11736 15162 11792
rect 15790 17434 15846 17436
rect 15870 17434 15926 17436
rect 15950 17434 16006 17436
rect 16030 17434 16086 17436
rect 15790 17382 15836 17434
rect 15836 17382 15846 17434
rect 15870 17382 15900 17434
rect 15900 17382 15912 17434
rect 15912 17382 15926 17434
rect 15950 17382 15964 17434
rect 15964 17382 15976 17434
rect 15976 17382 16006 17434
rect 16030 17382 16040 17434
rect 16040 17382 16086 17434
rect 15790 17380 15846 17382
rect 15870 17380 15926 17382
rect 15950 17380 16006 17382
rect 16030 17380 16086 17382
rect 16026 16652 16082 16688
rect 16026 16632 16028 16652
rect 16028 16632 16080 16652
rect 16080 16632 16082 16652
rect 15790 16346 15846 16348
rect 15870 16346 15926 16348
rect 15950 16346 16006 16348
rect 16030 16346 16086 16348
rect 15790 16294 15836 16346
rect 15836 16294 15846 16346
rect 15870 16294 15900 16346
rect 15900 16294 15912 16346
rect 15912 16294 15926 16346
rect 15950 16294 15964 16346
rect 15964 16294 15976 16346
rect 15976 16294 16006 16346
rect 16030 16294 16040 16346
rect 16040 16294 16086 16346
rect 15790 16292 15846 16294
rect 15870 16292 15926 16294
rect 15950 16292 16006 16294
rect 16030 16292 16086 16294
rect 15566 15408 15622 15464
rect 15474 14048 15530 14104
rect 15790 15258 15846 15260
rect 15870 15258 15926 15260
rect 15950 15258 16006 15260
rect 16030 15258 16086 15260
rect 15790 15206 15836 15258
rect 15836 15206 15846 15258
rect 15870 15206 15900 15258
rect 15900 15206 15912 15258
rect 15912 15206 15926 15258
rect 15950 15206 15964 15258
rect 15964 15206 15976 15258
rect 15976 15206 16006 15258
rect 16030 15206 16040 15258
rect 16040 15206 16086 15258
rect 15790 15204 15846 15206
rect 15870 15204 15926 15206
rect 15950 15204 16006 15206
rect 16030 15204 16086 15206
rect 15790 14170 15846 14172
rect 15870 14170 15926 14172
rect 15950 14170 16006 14172
rect 16030 14170 16086 14172
rect 15790 14118 15836 14170
rect 15836 14118 15846 14170
rect 15870 14118 15900 14170
rect 15900 14118 15912 14170
rect 15912 14118 15926 14170
rect 15950 14118 15964 14170
rect 15964 14118 15976 14170
rect 15976 14118 16006 14170
rect 16030 14118 16040 14170
rect 16040 14118 16086 14170
rect 15790 14116 15846 14118
rect 15870 14116 15926 14118
rect 15950 14116 16006 14118
rect 16030 14116 16086 14118
rect 15290 12416 15346 12472
rect 15290 12008 15346 12064
rect 15382 11736 15438 11792
rect 15934 13252 15990 13288
rect 15934 13232 15936 13252
rect 15936 13232 15988 13252
rect 15988 13232 15990 13252
rect 15790 13082 15846 13084
rect 15870 13082 15926 13084
rect 15950 13082 16006 13084
rect 16030 13082 16086 13084
rect 15790 13030 15836 13082
rect 15836 13030 15846 13082
rect 15870 13030 15900 13082
rect 15900 13030 15912 13082
rect 15912 13030 15926 13082
rect 15950 13030 15964 13082
rect 15964 13030 15976 13082
rect 15976 13030 16006 13082
rect 16030 13030 16040 13082
rect 16040 13030 16086 13082
rect 15790 13028 15846 13030
rect 15870 13028 15926 13030
rect 15950 13028 16006 13030
rect 16030 13028 16086 13030
rect 16210 14592 16266 14648
rect 16486 20712 16542 20768
rect 16486 20576 16542 20632
rect 16302 14320 16358 14376
rect 17314 26732 17316 26752
rect 17316 26732 17368 26752
rect 17368 26732 17370 26752
rect 17314 26696 17370 26732
rect 17130 22480 17186 22536
rect 17130 21936 17186 21992
rect 16578 18128 16634 18184
rect 16486 16768 16542 16824
rect 16486 16496 16542 16552
rect 16670 15680 16726 15736
rect 15658 12416 15714 12472
rect 16118 12708 16174 12744
rect 16118 12688 16120 12708
rect 16120 12688 16172 12708
rect 16172 12688 16174 12708
rect 15790 11994 15846 11996
rect 15870 11994 15926 11996
rect 15950 11994 16006 11996
rect 16030 11994 16086 11996
rect 15790 11942 15836 11994
rect 15836 11942 15846 11994
rect 15870 11942 15900 11994
rect 15900 11942 15912 11994
rect 15912 11942 15926 11994
rect 15950 11942 15964 11994
rect 15964 11942 15976 11994
rect 15976 11942 16006 11994
rect 16030 11942 16040 11994
rect 16040 11942 16086 11994
rect 15790 11940 15846 11942
rect 15870 11940 15926 11942
rect 15950 11940 16006 11942
rect 16030 11940 16086 11942
rect 15290 10784 15346 10840
rect 14922 9152 14978 9208
rect 14646 7520 14702 7576
rect 14830 7384 14886 7440
rect 15290 9560 15346 9616
rect 16302 12552 16358 12608
rect 16302 12416 16358 12472
rect 16302 12008 16358 12064
rect 15658 10920 15714 10976
rect 15790 10906 15846 10908
rect 15870 10906 15926 10908
rect 15950 10906 16006 10908
rect 16030 10906 16086 10908
rect 15790 10854 15836 10906
rect 15836 10854 15846 10906
rect 15870 10854 15900 10906
rect 15900 10854 15912 10906
rect 15912 10854 15926 10906
rect 15950 10854 15964 10906
rect 15964 10854 15976 10906
rect 15976 10854 16006 10906
rect 16030 10854 16040 10906
rect 16040 10854 16086 10906
rect 15790 10852 15846 10854
rect 15870 10852 15926 10854
rect 15950 10852 16006 10854
rect 16030 10852 16086 10854
rect 16210 10784 16266 10840
rect 16946 18264 17002 18320
rect 16946 16124 16948 16144
rect 16948 16124 17000 16144
rect 17000 16124 17002 16144
rect 16946 16088 17002 16124
rect 16946 15408 17002 15464
rect 16670 13268 16672 13288
rect 16672 13268 16724 13288
rect 16724 13268 16726 13288
rect 16670 13232 16726 13268
rect 16670 12688 16726 12744
rect 16946 13640 17002 13696
rect 16946 12552 17002 12608
rect 15014 7656 15070 7712
rect 15658 9832 15714 9888
rect 15790 9818 15846 9820
rect 15870 9818 15926 9820
rect 15950 9818 16006 9820
rect 16030 9818 16086 9820
rect 15790 9766 15836 9818
rect 15836 9766 15846 9818
rect 15870 9766 15900 9818
rect 15900 9766 15912 9818
rect 15912 9766 15926 9818
rect 15950 9766 15964 9818
rect 15964 9766 15976 9818
rect 15976 9766 16006 9818
rect 16030 9766 16040 9818
rect 16040 9766 16086 9818
rect 15790 9764 15846 9766
rect 15870 9764 15926 9766
rect 15950 9764 16006 9766
rect 16030 9764 16086 9766
rect 16302 10512 16358 10568
rect 16302 9832 16358 9888
rect 15658 9424 15714 9480
rect 15750 9152 15806 9208
rect 15290 8608 15346 8664
rect 14830 6704 14886 6760
rect 15474 8880 15530 8936
rect 16394 8916 16396 8936
rect 16396 8916 16448 8936
rect 16448 8916 16450 8936
rect 16394 8880 16450 8916
rect 15790 8730 15846 8732
rect 15870 8730 15926 8732
rect 15950 8730 16006 8732
rect 16030 8730 16086 8732
rect 15790 8678 15836 8730
rect 15836 8678 15846 8730
rect 15870 8678 15900 8730
rect 15900 8678 15912 8730
rect 15912 8678 15926 8730
rect 15950 8678 15964 8730
rect 15964 8678 15976 8730
rect 15976 8678 16006 8730
rect 16030 8678 16040 8730
rect 16040 8678 16086 8730
rect 15790 8676 15846 8678
rect 15870 8676 15926 8678
rect 15950 8676 16006 8678
rect 16030 8676 16086 8678
rect 16210 8628 16266 8664
rect 16210 8608 16212 8628
rect 16212 8608 16264 8628
rect 16264 8608 16266 8628
rect 16210 8064 16266 8120
rect 15790 7642 15846 7644
rect 15870 7642 15926 7644
rect 15950 7642 16006 7644
rect 16030 7642 16086 7644
rect 15790 7590 15836 7642
rect 15836 7590 15846 7642
rect 15870 7590 15900 7642
rect 15900 7590 15912 7642
rect 15912 7590 15926 7642
rect 15950 7590 15964 7642
rect 15964 7590 15976 7642
rect 15976 7590 16006 7642
rect 16030 7590 16040 7642
rect 16040 7590 16086 7642
rect 15790 7588 15846 7590
rect 15870 7588 15926 7590
rect 15950 7588 16006 7590
rect 16030 7588 16086 7590
rect 16394 7928 16450 7984
rect 16670 8084 16726 8120
rect 16670 8064 16672 8084
rect 16672 8064 16724 8084
rect 16724 8064 16726 8084
rect 16210 7656 16266 7712
rect 16394 7656 16450 7712
rect 15290 6704 15346 6760
rect 13318 4922 13374 4924
rect 13398 4922 13454 4924
rect 13478 4922 13534 4924
rect 13558 4922 13614 4924
rect 13318 4870 13364 4922
rect 13364 4870 13374 4922
rect 13398 4870 13428 4922
rect 13428 4870 13440 4922
rect 13440 4870 13454 4922
rect 13478 4870 13492 4922
rect 13492 4870 13504 4922
rect 13504 4870 13534 4922
rect 13558 4870 13568 4922
rect 13568 4870 13614 4922
rect 13318 4868 13374 4870
rect 13398 4868 13454 4870
rect 13478 4868 13534 4870
rect 13558 4868 13614 4870
rect 13174 4800 13230 4856
rect 12438 4392 12494 4448
rect 12898 4392 12954 4448
rect 13174 4684 13230 4720
rect 13174 4664 13176 4684
rect 13176 4664 13228 4684
rect 13228 4664 13230 4684
rect 13174 4120 13230 4176
rect 12438 3984 12494 4040
rect 13358 4120 13414 4176
rect 13266 3984 13322 4040
rect 14554 5888 14610 5944
rect 14186 5208 14242 5264
rect 14186 4936 14242 4992
rect 14554 5072 14610 5128
rect 14094 4664 14150 4720
rect 14370 4800 14426 4856
rect 14554 4936 14610 4992
rect 14830 5752 14886 5808
rect 15014 6160 15070 6216
rect 15014 5752 15070 5808
rect 15290 6432 15346 6488
rect 15290 6024 15346 6080
rect 14738 5072 14794 5128
rect 15198 5108 15200 5128
rect 15200 5108 15252 5128
rect 15252 5108 15254 5128
rect 15198 5072 15254 5108
rect 15566 6432 15622 6488
rect 15790 6554 15846 6556
rect 15870 6554 15926 6556
rect 15950 6554 16006 6556
rect 16030 6554 16086 6556
rect 15790 6502 15836 6554
rect 15836 6502 15846 6554
rect 15870 6502 15900 6554
rect 15900 6502 15912 6554
rect 15912 6502 15926 6554
rect 15950 6502 15964 6554
rect 15964 6502 15976 6554
rect 15976 6502 16006 6554
rect 16030 6502 16040 6554
rect 16040 6502 16086 6554
rect 15790 6500 15846 6502
rect 15870 6500 15926 6502
rect 15950 6500 16006 6502
rect 16030 6500 16086 6502
rect 16210 6432 16266 6488
rect 17222 20304 17278 20360
rect 17958 41792 18014 41848
rect 18694 43308 18750 43344
rect 18694 43288 18696 43308
rect 18696 43288 18748 43308
rect 18748 43288 18750 43308
rect 18263 43002 18319 43004
rect 18343 43002 18399 43004
rect 18423 43002 18479 43004
rect 18503 43002 18559 43004
rect 18263 42950 18309 43002
rect 18309 42950 18319 43002
rect 18343 42950 18373 43002
rect 18373 42950 18385 43002
rect 18385 42950 18399 43002
rect 18423 42950 18437 43002
rect 18437 42950 18449 43002
rect 18449 42950 18479 43002
rect 18503 42950 18513 43002
rect 18513 42950 18559 43002
rect 18263 42948 18319 42950
rect 18343 42948 18399 42950
rect 18423 42948 18479 42950
rect 18503 42948 18559 42950
rect 18326 42608 18382 42664
rect 18234 42064 18290 42120
rect 18263 41914 18319 41916
rect 18343 41914 18399 41916
rect 18423 41914 18479 41916
rect 18503 41914 18559 41916
rect 18263 41862 18309 41914
rect 18309 41862 18319 41914
rect 18343 41862 18373 41914
rect 18373 41862 18385 41914
rect 18385 41862 18399 41914
rect 18423 41862 18437 41914
rect 18437 41862 18449 41914
rect 18449 41862 18479 41914
rect 18503 41862 18513 41914
rect 18513 41862 18559 41914
rect 18263 41860 18319 41862
rect 18343 41860 18399 41862
rect 18423 41860 18479 41862
rect 18503 41860 18559 41862
rect 18878 43152 18934 43208
rect 19062 42764 19118 42800
rect 19062 42744 19064 42764
rect 19064 42744 19116 42764
rect 19116 42744 19118 42764
rect 18694 41112 18750 41168
rect 17682 39752 17738 39808
rect 18263 40826 18319 40828
rect 18343 40826 18399 40828
rect 18423 40826 18479 40828
rect 18503 40826 18559 40828
rect 18263 40774 18309 40826
rect 18309 40774 18319 40826
rect 18343 40774 18373 40826
rect 18373 40774 18385 40826
rect 18385 40774 18399 40826
rect 18423 40774 18437 40826
rect 18437 40774 18449 40826
rect 18449 40774 18479 40826
rect 18503 40774 18513 40826
rect 18513 40774 18559 40826
rect 18263 40772 18319 40774
rect 18343 40772 18399 40774
rect 18423 40772 18479 40774
rect 18503 40772 18559 40774
rect 18326 40568 18382 40624
rect 18234 40432 18290 40488
rect 18142 40024 18198 40080
rect 18418 40160 18474 40216
rect 18602 40024 18658 40080
rect 18263 39738 18319 39740
rect 18343 39738 18399 39740
rect 18423 39738 18479 39740
rect 18503 39738 18559 39740
rect 18263 39686 18309 39738
rect 18309 39686 18319 39738
rect 18343 39686 18373 39738
rect 18373 39686 18385 39738
rect 18385 39686 18399 39738
rect 18423 39686 18437 39738
rect 18437 39686 18449 39738
rect 18449 39686 18479 39738
rect 18503 39686 18513 39738
rect 18513 39686 18559 39738
rect 18263 39684 18319 39686
rect 18343 39684 18399 39686
rect 18423 39684 18479 39686
rect 18503 39684 18559 39686
rect 17958 39208 18014 39264
rect 18326 39364 18382 39400
rect 18326 39344 18328 39364
rect 18328 39344 18380 39364
rect 18380 39344 18382 39364
rect 18326 39092 18382 39128
rect 18326 39072 18328 39092
rect 18328 39072 18380 39092
rect 18380 39072 18382 39092
rect 18050 38956 18106 38992
rect 18694 39616 18750 39672
rect 19982 43968 20038 44024
rect 19338 41964 19340 41984
rect 19340 41964 19392 41984
rect 19392 41964 19394 41984
rect 19338 41928 19394 41964
rect 18878 40976 18934 41032
rect 18602 39208 18658 39264
rect 18050 38936 18052 38956
rect 18052 38936 18104 38956
rect 18104 38936 18106 38956
rect 18263 38650 18319 38652
rect 18343 38650 18399 38652
rect 18423 38650 18479 38652
rect 18503 38650 18559 38652
rect 18263 38598 18309 38650
rect 18309 38598 18319 38650
rect 18343 38598 18373 38650
rect 18373 38598 18385 38650
rect 18385 38598 18399 38650
rect 18423 38598 18437 38650
rect 18437 38598 18449 38650
rect 18449 38598 18479 38650
rect 18503 38598 18513 38650
rect 18513 38598 18559 38650
rect 18263 38596 18319 38598
rect 18343 38596 18399 38598
rect 18423 38596 18479 38598
rect 18503 38596 18559 38598
rect 18263 37562 18319 37564
rect 18343 37562 18399 37564
rect 18423 37562 18479 37564
rect 18503 37562 18559 37564
rect 18263 37510 18309 37562
rect 18309 37510 18319 37562
rect 18343 37510 18373 37562
rect 18373 37510 18385 37562
rect 18385 37510 18399 37562
rect 18423 37510 18437 37562
rect 18437 37510 18449 37562
rect 18449 37510 18479 37562
rect 18503 37510 18513 37562
rect 18513 37510 18559 37562
rect 18263 37508 18319 37510
rect 18343 37508 18399 37510
rect 18423 37508 18479 37510
rect 18503 37508 18559 37510
rect 18142 36624 18198 36680
rect 18418 36896 18474 36952
rect 18326 36624 18382 36680
rect 18263 36474 18319 36476
rect 18343 36474 18399 36476
rect 18423 36474 18479 36476
rect 18503 36474 18559 36476
rect 18263 36422 18309 36474
rect 18309 36422 18319 36474
rect 18343 36422 18373 36474
rect 18373 36422 18385 36474
rect 18385 36422 18399 36474
rect 18423 36422 18437 36474
rect 18437 36422 18449 36474
rect 18449 36422 18479 36474
rect 18503 36422 18513 36474
rect 18513 36422 18559 36474
rect 18263 36420 18319 36422
rect 18343 36420 18399 36422
rect 18423 36420 18479 36422
rect 18503 36420 18559 36422
rect 19062 39616 19118 39672
rect 18878 38936 18934 38992
rect 18786 37204 18788 37224
rect 18788 37204 18840 37224
rect 18840 37204 18842 37224
rect 18786 37168 18842 37204
rect 18694 36352 18750 36408
rect 18418 36116 18420 36136
rect 18420 36116 18472 36136
rect 18472 36116 18474 36136
rect 18418 36080 18474 36116
rect 18970 37984 19026 38040
rect 19246 39380 19248 39400
rect 19248 39380 19300 39400
rect 19300 39380 19302 39400
rect 19246 39344 19302 39380
rect 21178 43560 21234 43616
rect 20735 43546 20791 43548
rect 20815 43546 20871 43548
rect 20895 43546 20951 43548
rect 20975 43546 21031 43548
rect 20735 43494 20781 43546
rect 20781 43494 20791 43546
rect 20815 43494 20845 43546
rect 20845 43494 20857 43546
rect 20857 43494 20871 43546
rect 20895 43494 20909 43546
rect 20909 43494 20921 43546
rect 20921 43494 20951 43546
rect 20975 43494 20985 43546
rect 20985 43494 21031 43546
rect 20735 43492 20791 43494
rect 20815 43492 20871 43494
rect 20895 43492 20951 43494
rect 20975 43492 21031 43494
rect 19982 43016 20038 43072
rect 19798 41384 19854 41440
rect 19706 41112 19762 41168
rect 19706 39888 19762 39944
rect 19706 39480 19762 39536
rect 18970 36760 19026 36816
rect 18786 35672 18842 35728
rect 18263 35386 18319 35388
rect 18343 35386 18399 35388
rect 18423 35386 18479 35388
rect 18503 35386 18559 35388
rect 18263 35334 18309 35386
rect 18309 35334 18319 35386
rect 18343 35334 18373 35386
rect 18373 35334 18385 35386
rect 18385 35334 18399 35386
rect 18423 35334 18437 35386
rect 18437 35334 18449 35386
rect 18449 35334 18479 35386
rect 18503 35334 18513 35386
rect 18513 35334 18559 35386
rect 18263 35332 18319 35334
rect 18343 35332 18399 35334
rect 18423 35332 18479 35334
rect 18503 35332 18559 35334
rect 18263 34298 18319 34300
rect 18343 34298 18399 34300
rect 18423 34298 18479 34300
rect 18503 34298 18559 34300
rect 18263 34246 18309 34298
rect 18309 34246 18319 34298
rect 18343 34246 18373 34298
rect 18373 34246 18385 34298
rect 18385 34246 18399 34298
rect 18423 34246 18437 34298
rect 18437 34246 18449 34298
rect 18449 34246 18479 34298
rect 18503 34246 18513 34298
rect 18513 34246 18559 34298
rect 18263 34244 18319 34246
rect 18343 34244 18399 34246
rect 18423 34244 18479 34246
rect 18503 34244 18559 34246
rect 18970 34448 19026 34504
rect 18510 33904 18566 33960
rect 18142 33496 18198 33552
rect 18050 32408 18106 32464
rect 18263 33210 18319 33212
rect 18343 33210 18399 33212
rect 18423 33210 18479 33212
rect 18503 33210 18559 33212
rect 18263 33158 18309 33210
rect 18309 33158 18319 33210
rect 18343 33158 18373 33210
rect 18373 33158 18385 33210
rect 18385 33158 18399 33210
rect 18423 33158 18437 33210
rect 18437 33158 18449 33210
rect 18449 33158 18479 33210
rect 18503 33158 18513 33210
rect 18513 33158 18559 33210
rect 18263 33156 18319 33158
rect 18343 33156 18399 33158
rect 18423 33156 18479 33158
rect 18503 33156 18559 33158
rect 18786 34040 18842 34096
rect 18694 33496 18750 33552
rect 18694 32952 18750 33008
rect 18694 32816 18750 32872
rect 19154 37712 19210 37768
rect 19246 35264 19302 35320
rect 20735 42458 20791 42460
rect 20815 42458 20871 42460
rect 20895 42458 20951 42460
rect 20975 42458 21031 42460
rect 20735 42406 20781 42458
rect 20781 42406 20791 42458
rect 20815 42406 20845 42458
rect 20845 42406 20857 42458
rect 20857 42406 20871 42458
rect 20895 42406 20909 42458
rect 20909 42406 20921 42458
rect 20921 42406 20951 42458
rect 20975 42406 20985 42458
rect 20985 42406 21031 42458
rect 20735 42404 20791 42406
rect 20815 42404 20871 42406
rect 20895 42404 20951 42406
rect 20975 42404 21031 42406
rect 21270 42472 21326 42528
rect 19798 36488 19854 36544
rect 18234 32272 18290 32328
rect 18263 32122 18319 32124
rect 18343 32122 18399 32124
rect 18423 32122 18479 32124
rect 18503 32122 18559 32124
rect 18263 32070 18309 32122
rect 18309 32070 18319 32122
rect 18343 32070 18373 32122
rect 18373 32070 18385 32122
rect 18385 32070 18399 32122
rect 18423 32070 18437 32122
rect 18437 32070 18449 32122
rect 18449 32070 18479 32122
rect 18503 32070 18513 32122
rect 18513 32070 18559 32122
rect 18263 32068 18319 32070
rect 18343 32068 18399 32070
rect 18423 32068 18479 32070
rect 18503 32068 18559 32070
rect 17590 29008 17646 29064
rect 18234 31728 18290 31784
rect 18418 31320 18474 31376
rect 18142 31184 18198 31240
rect 18326 31184 18382 31240
rect 18263 31034 18319 31036
rect 18343 31034 18399 31036
rect 18423 31034 18479 31036
rect 18503 31034 18559 31036
rect 18263 30982 18309 31034
rect 18309 30982 18319 31034
rect 18343 30982 18373 31034
rect 18373 30982 18385 31034
rect 18385 30982 18399 31034
rect 18423 30982 18437 31034
rect 18437 30982 18449 31034
rect 18449 30982 18479 31034
rect 18503 30982 18513 31034
rect 18513 30982 18559 31034
rect 18263 30980 18319 30982
rect 18343 30980 18399 30982
rect 18423 30980 18479 30982
rect 18503 30980 18559 30982
rect 18234 30096 18290 30152
rect 18263 29946 18319 29948
rect 18343 29946 18399 29948
rect 18423 29946 18479 29948
rect 18503 29946 18559 29948
rect 18263 29894 18309 29946
rect 18309 29894 18319 29946
rect 18343 29894 18373 29946
rect 18373 29894 18385 29946
rect 18385 29894 18399 29946
rect 18423 29894 18437 29946
rect 18437 29894 18449 29946
rect 18449 29894 18479 29946
rect 18503 29894 18513 29946
rect 18513 29894 18559 29946
rect 18263 29892 18319 29894
rect 18343 29892 18399 29894
rect 18423 29892 18479 29894
rect 18503 29892 18559 29894
rect 18694 31084 18696 31104
rect 18696 31084 18748 31104
rect 18748 31084 18750 31104
rect 18694 31048 18750 31084
rect 18786 30912 18842 30968
rect 19062 33496 19118 33552
rect 20534 40840 20590 40896
rect 21270 41384 21326 41440
rect 20735 41370 20791 41372
rect 20815 41370 20871 41372
rect 20895 41370 20951 41372
rect 20975 41370 21031 41372
rect 20735 41318 20781 41370
rect 20781 41318 20791 41370
rect 20815 41318 20845 41370
rect 20845 41318 20857 41370
rect 20857 41318 20871 41370
rect 20895 41318 20909 41370
rect 20909 41318 20921 41370
rect 20921 41318 20951 41370
rect 20975 41318 20985 41370
rect 20985 41318 21031 41370
rect 20735 41316 20791 41318
rect 20815 41316 20871 41318
rect 20895 41316 20951 41318
rect 20975 41316 21031 41318
rect 20735 40282 20791 40284
rect 20815 40282 20871 40284
rect 20895 40282 20951 40284
rect 20975 40282 21031 40284
rect 20735 40230 20781 40282
rect 20781 40230 20791 40282
rect 20815 40230 20845 40282
rect 20845 40230 20857 40282
rect 20857 40230 20871 40282
rect 20895 40230 20909 40282
rect 20909 40230 20921 40282
rect 20921 40230 20951 40282
rect 20975 40230 20985 40282
rect 20985 40230 21031 40282
rect 20735 40228 20791 40230
rect 20815 40228 20871 40230
rect 20895 40228 20951 40230
rect 20975 40228 21031 40230
rect 20994 39788 20996 39808
rect 20996 39788 21048 39808
rect 21048 39788 21050 39808
rect 20994 39752 21050 39788
rect 20735 39194 20791 39196
rect 20815 39194 20871 39196
rect 20895 39194 20951 39196
rect 20975 39194 21031 39196
rect 20735 39142 20781 39194
rect 20781 39142 20791 39194
rect 20815 39142 20845 39194
rect 20845 39142 20857 39194
rect 20857 39142 20871 39194
rect 20895 39142 20909 39194
rect 20909 39142 20921 39194
rect 20921 39142 20951 39194
rect 20975 39142 20985 39194
rect 20985 39142 21031 39194
rect 20735 39140 20791 39142
rect 20815 39140 20871 39142
rect 20895 39140 20951 39142
rect 20975 39140 21031 39142
rect 20442 38700 20444 38720
rect 20444 38700 20496 38720
rect 20496 38700 20498 38720
rect 20442 38664 20498 38700
rect 20442 37612 20444 37632
rect 20444 37612 20496 37632
rect 20496 37612 20498 37632
rect 20442 37576 20498 37612
rect 20258 37168 20314 37224
rect 20735 38106 20791 38108
rect 20815 38106 20871 38108
rect 20895 38106 20951 38108
rect 20975 38106 21031 38108
rect 20735 38054 20781 38106
rect 20781 38054 20791 38106
rect 20815 38054 20845 38106
rect 20845 38054 20857 38106
rect 20857 38054 20871 38106
rect 20895 38054 20909 38106
rect 20909 38054 20921 38106
rect 20921 38054 20951 38106
rect 20975 38054 20985 38106
rect 20985 38054 21031 38106
rect 20735 38052 20791 38054
rect 20815 38052 20871 38054
rect 20895 38052 20951 38054
rect 20975 38052 21031 38054
rect 20735 37018 20791 37020
rect 20815 37018 20871 37020
rect 20895 37018 20951 37020
rect 20975 37018 21031 37020
rect 20735 36966 20781 37018
rect 20781 36966 20791 37018
rect 20815 36966 20845 37018
rect 20845 36966 20857 37018
rect 20857 36966 20871 37018
rect 20895 36966 20909 37018
rect 20909 36966 20921 37018
rect 20921 36966 20951 37018
rect 20975 36966 20985 37018
rect 20985 36966 21031 37018
rect 20735 36964 20791 36966
rect 20815 36964 20871 36966
rect 20895 36964 20951 36966
rect 20975 36964 21031 36966
rect 20735 35930 20791 35932
rect 20815 35930 20871 35932
rect 20895 35930 20951 35932
rect 20975 35930 21031 35932
rect 20735 35878 20781 35930
rect 20781 35878 20791 35930
rect 20815 35878 20845 35930
rect 20845 35878 20857 35930
rect 20857 35878 20871 35930
rect 20895 35878 20909 35930
rect 20909 35878 20921 35930
rect 20921 35878 20951 35930
rect 20975 35878 20985 35930
rect 20985 35878 21031 35930
rect 20735 35876 20791 35878
rect 20815 35876 20871 35878
rect 20895 35876 20951 35878
rect 20975 35876 21031 35878
rect 19430 34040 19486 34096
rect 19338 33260 19340 33280
rect 19340 33260 19392 33280
rect 19392 33260 19394 33280
rect 19338 33224 19394 33260
rect 19522 33768 19578 33824
rect 19706 33904 19762 33960
rect 19062 31884 19118 31920
rect 19062 31864 19064 31884
rect 19064 31864 19116 31884
rect 19116 31864 19118 31884
rect 19062 31048 19118 31104
rect 19430 32716 19432 32736
rect 19432 32716 19484 32736
rect 19484 32716 19486 32736
rect 19430 32680 19486 32716
rect 19706 33224 19762 33280
rect 19430 32408 19486 32464
rect 19246 31048 19302 31104
rect 20350 35400 20406 35456
rect 20442 34348 20444 34368
rect 20444 34348 20496 34368
rect 20496 34348 20498 34368
rect 20074 32680 20130 32736
rect 19890 31728 19946 31784
rect 19154 30776 19210 30832
rect 18263 28858 18319 28860
rect 18343 28858 18399 28860
rect 18423 28858 18479 28860
rect 18503 28858 18559 28860
rect 18263 28806 18309 28858
rect 18309 28806 18319 28858
rect 18343 28806 18373 28858
rect 18373 28806 18385 28858
rect 18385 28806 18399 28858
rect 18423 28806 18437 28858
rect 18437 28806 18449 28858
rect 18449 28806 18479 28858
rect 18503 28806 18513 28858
rect 18513 28806 18559 28858
rect 18263 28804 18319 28806
rect 18343 28804 18399 28806
rect 18423 28804 18479 28806
rect 18503 28804 18559 28806
rect 17774 28056 17830 28112
rect 17866 25200 17922 25256
rect 17774 23296 17830 23352
rect 18263 27770 18319 27772
rect 18343 27770 18399 27772
rect 18423 27770 18479 27772
rect 18503 27770 18559 27772
rect 18263 27718 18309 27770
rect 18309 27718 18319 27770
rect 18343 27718 18373 27770
rect 18373 27718 18385 27770
rect 18385 27718 18399 27770
rect 18423 27718 18437 27770
rect 18437 27718 18449 27770
rect 18449 27718 18479 27770
rect 18503 27718 18513 27770
rect 18513 27718 18559 27770
rect 18263 27716 18319 27718
rect 18343 27716 18399 27718
rect 18423 27716 18479 27718
rect 18503 27716 18559 27718
rect 18602 26968 18658 27024
rect 18263 26682 18319 26684
rect 18343 26682 18399 26684
rect 18423 26682 18479 26684
rect 18503 26682 18559 26684
rect 18263 26630 18309 26682
rect 18309 26630 18319 26682
rect 18343 26630 18373 26682
rect 18373 26630 18385 26682
rect 18385 26630 18399 26682
rect 18423 26630 18437 26682
rect 18437 26630 18449 26682
rect 18449 26630 18479 26682
rect 18503 26630 18513 26682
rect 18513 26630 18559 26682
rect 18263 26628 18319 26630
rect 18343 26628 18399 26630
rect 18423 26628 18479 26630
rect 18503 26628 18559 26630
rect 19062 29144 19118 29200
rect 19246 30096 19302 30152
rect 19246 29144 19302 29200
rect 19246 28192 19302 28248
rect 19246 28056 19302 28112
rect 18878 26832 18934 26888
rect 18510 25880 18566 25936
rect 18263 25594 18319 25596
rect 18343 25594 18399 25596
rect 18423 25594 18479 25596
rect 18503 25594 18559 25596
rect 18263 25542 18309 25594
rect 18309 25542 18319 25594
rect 18343 25542 18373 25594
rect 18373 25542 18385 25594
rect 18385 25542 18399 25594
rect 18423 25542 18437 25594
rect 18437 25542 18449 25594
rect 18449 25542 18479 25594
rect 18503 25542 18513 25594
rect 18513 25542 18559 25594
rect 18263 25540 18319 25542
rect 18343 25540 18399 25542
rect 18423 25540 18479 25542
rect 18503 25540 18559 25542
rect 19062 26152 19118 26208
rect 17774 21392 17830 21448
rect 17774 19896 17830 19952
rect 17590 17584 17646 17640
rect 18263 24506 18319 24508
rect 18343 24506 18399 24508
rect 18423 24506 18479 24508
rect 18503 24506 18559 24508
rect 18263 24454 18309 24506
rect 18309 24454 18319 24506
rect 18343 24454 18373 24506
rect 18373 24454 18385 24506
rect 18385 24454 18399 24506
rect 18423 24454 18437 24506
rect 18437 24454 18449 24506
rect 18449 24454 18479 24506
rect 18503 24454 18513 24506
rect 18513 24454 18559 24506
rect 18263 24452 18319 24454
rect 18343 24452 18399 24454
rect 18423 24452 18479 24454
rect 18503 24452 18559 24454
rect 18263 23418 18319 23420
rect 18343 23418 18399 23420
rect 18423 23418 18479 23420
rect 18503 23418 18559 23420
rect 18263 23366 18309 23418
rect 18309 23366 18319 23418
rect 18343 23366 18373 23418
rect 18373 23366 18385 23418
rect 18385 23366 18399 23418
rect 18423 23366 18437 23418
rect 18437 23366 18449 23418
rect 18449 23366 18479 23418
rect 18503 23366 18513 23418
rect 18513 23366 18559 23418
rect 18263 23364 18319 23366
rect 18343 23364 18399 23366
rect 18423 23364 18479 23366
rect 18503 23364 18559 23366
rect 18263 22330 18319 22332
rect 18343 22330 18399 22332
rect 18423 22330 18479 22332
rect 18503 22330 18559 22332
rect 18263 22278 18309 22330
rect 18309 22278 18319 22330
rect 18343 22278 18373 22330
rect 18373 22278 18385 22330
rect 18385 22278 18399 22330
rect 18423 22278 18437 22330
rect 18437 22278 18449 22330
rect 18449 22278 18479 22330
rect 18503 22278 18513 22330
rect 18513 22278 18559 22330
rect 18263 22276 18319 22278
rect 18343 22276 18399 22278
rect 18423 22276 18479 22278
rect 18503 22276 18559 22278
rect 18263 21242 18319 21244
rect 18343 21242 18399 21244
rect 18423 21242 18479 21244
rect 18503 21242 18559 21244
rect 18263 21190 18309 21242
rect 18309 21190 18319 21242
rect 18343 21190 18373 21242
rect 18373 21190 18385 21242
rect 18385 21190 18399 21242
rect 18423 21190 18437 21242
rect 18437 21190 18449 21242
rect 18449 21190 18479 21242
rect 18503 21190 18513 21242
rect 18513 21190 18559 21242
rect 18263 21188 18319 21190
rect 18343 21188 18399 21190
rect 18423 21188 18479 21190
rect 18503 21188 18559 21190
rect 18263 20154 18319 20156
rect 18343 20154 18399 20156
rect 18423 20154 18479 20156
rect 18503 20154 18559 20156
rect 18263 20102 18309 20154
rect 18309 20102 18319 20154
rect 18343 20102 18373 20154
rect 18373 20102 18385 20154
rect 18385 20102 18399 20154
rect 18423 20102 18437 20154
rect 18437 20102 18449 20154
rect 18449 20102 18479 20154
rect 18503 20102 18513 20154
rect 18513 20102 18559 20154
rect 18263 20100 18319 20102
rect 18343 20100 18399 20102
rect 18423 20100 18479 20102
rect 18503 20100 18559 20102
rect 18263 19066 18319 19068
rect 18343 19066 18399 19068
rect 18423 19066 18479 19068
rect 18503 19066 18559 19068
rect 18263 19014 18309 19066
rect 18309 19014 18319 19066
rect 18343 19014 18373 19066
rect 18373 19014 18385 19066
rect 18385 19014 18399 19066
rect 18423 19014 18437 19066
rect 18437 19014 18449 19066
rect 18449 19014 18479 19066
rect 18503 19014 18513 19066
rect 18513 19014 18559 19066
rect 18263 19012 18319 19014
rect 18343 19012 18399 19014
rect 18423 19012 18479 19014
rect 18503 19012 18559 19014
rect 18263 17978 18319 17980
rect 18343 17978 18399 17980
rect 18423 17978 18479 17980
rect 18503 17978 18559 17980
rect 18263 17926 18309 17978
rect 18309 17926 18319 17978
rect 18343 17926 18373 17978
rect 18373 17926 18385 17978
rect 18385 17926 18399 17978
rect 18423 17926 18437 17978
rect 18437 17926 18449 17978
rect 18449 17926 18479 17978
rect 18503 17926 18513 17978
rect 18513 17926 18559 17978
rect 18263 17924 18319 17926
rect 18343 17924 18399 17926
rect 18423 17924 18479 17926
rect 18503 17924 18559 17926
rect 18050 17040 18106 17096
rect 17774 15952 17830 16008
rect 17406 14864 17462 14920
rect 17314 13776 17370 13832
rect 17314 12144 17370 12200
rect 17222 11464 17278 11520
rect 17682 14320 17738 14376
rect 17590 13504 17646 13560
rect 17038 10668 17094 10704
rect 17038 10648 17040 10668
rect 17040 10648 17092 10668
rect 17092 10648 17094 10668
rect 17038 10240 17094 10296
rect 17038 9288 17094 9344
rect 16578 7248 16634 7304
rect 16394 6976 16450 7032
rect 17682 12824 17738 12880
rect 17682 12280 17738 12336
rect 17866 11872 17922 11928
rect 18263 16890 18319 16892
rect 18343 16890 18399 16892
rect 18423 16890 18479 16892
rect 18503 16890 18559 16892
rect 18263 16838 18309 16890
rect 18309 16838 18319 16890
rect 18343 16838 18373 16890
rect 18373 16838 18385 16890
rect 18385 16838 18399 16890
rect 18423 16838 18437 16890
rect 18437 16838 18449 16890
rect 18449 16838 18479 16890
rect 18503 16838 18513 16890
rect 18513 16838 18559 16890
rect 18263 16836 18319 16838
rect 18343 16836 18399 16838
rect 18423 16836 18479 16838
rect 18503 16836 18559 16838
rect 18050 16496 18106 16552
rect 18263 15802 18319 15804
rect 18343 15802 18399 15804
rect 18423 15802 18479 15804
rect 18503 15802 18559 15804
rect 18263 15750 18309 15802
rect 18309 15750 18319 15802
rect 18343 15750 18373 15802
rect 18373 15750 18385 15802
rect 18385 15750 18399 15802
rect 18423 15750 18437 15802
rect 18437 15750 18449 15802
rect 18449 15750 18479 15802
rect 18503 15750 18513 15802
rect 18513 15750 18559 15802
rect 18263 15748 18319 15750
rect 18343 15748 18399 15750
rect 18423 15748 18479 15750
rect 18503 15748 18559 15750
rect 18418 15544 18474 15600
rect 19798 30912 19854 30968
rect 19522 29552 19578 29608
rect 19338 26460 19340 26480
rect 19340 26460 19392 26480
rect 19392 26460 19394 26480
rect 19338 26424 19394 26460
rect 19246 25064 19302 25120
rect 19338 23296 19394 23352
rect 19062 21392 19118 21448
rect 18970 20984 19026 21040
rect 19706 27648 19762 27704
rect 20258 33360 20314 33416
rect 20442 34312 20498 34348
rect 20442 33260 20444 33280
rect 20444 33260 20496 33280
rect 20496 33260 20498 33280
rect 20442 33224 20498 33260
rect 20350 32816 20406 32872
rect 20534 32136 20590 32192
rect 20735 34842 20791 34844
rect 20815 34842 20871 34844
rect 20895 34842 20951 34844
rect 20975 34842 21031 34844
rect 20735 34790 20781 34842
rect 20781 34790 20791 34842
rect 20815 34790 20845 34842
rect 20845 34790 20857 34842
rect 20857 34790 20871 34842
rect 20895 34790 20909 34842
rect 20909 34790 20921 34842
rect 20921 34790 20951 34842
rect 20975 34790 20985 34842
rect 20985 34790 21031 34842
rect 20735 34788 20791 34790
rect 20815 34788 20871 34790
rect 20895 34788 20951 34790
rect 20975 34788 21031 34790
rect 20735 33754 20791 33756
rect 20815 33754 20871 33756
rect 20895 33754 20951 33756
rect 20975 33754 21031 33756
rect 20735 33702 20781 33754
rect 20781 33702 20791 33754
rect 20815 33702 20845 33754
rect 20845 33702 20857 33754
rect 20857 33702 20871 33754
rect 20895 33702 20909 33754
rect 20909 33702 20921 33754
rect 20921 33702 20951 33754
rect 20975 33702 20985 33754
rect 20985 33702 21031 33754
rect 20735 33700 20791 33702
rect 20815 33700 20871 33702
rect 20895 33700 20951 33702
rect 20975 33700 21031 33702
rect 20735 32666 20791 32668
rect 20815 32666 20871 32668
rect 20895 32666 20951 32668
rect 20975 32666 21031 32668
rect 20735 32614 20781 32666
rect 20781 32614 20791 32666
rect 20815 32614 20845 32666
rect 20845 32614 20857 32666
rect 20857 32614 20871 32666
rect 20895 32614 20909 32666
rect 20909 32614 20921 32666
rect 20921 32614 20951 32666
rect 20975 32614 20985 32666
rect 20985 32614 21031 32666
rect 20735 32612 20791 32614
rect 20815 32612 20871 32614
rect 20895 32612 20951 32614
rect 20975 32612 21031 32614
rect 20735 31578 20791 31580
rect 20815 31578 20871 31580
rect 20895 31578 20951 31580
rect 20975 31578 21031 31580
rect 20735 31526 20781 31578
rect 20781 31526 20791 31578
rect 20815 31526 20845 31578
rect 20845 31526 20857 31578
rect 20857 31526 20871 31578
rect 20895 31526 20909 31578
rect 20909 31526 20921 31578
rect 20921 31526 20951 31578
rect 20975 31526 20985 31578
rect 20985 31526 21031 31578
rect 20735 31524 20791 31526
rect 20815 31524 20871 31526
rect 20895 31524 20951 31526
rect 20975 31524 21031 31526
rect 20442 31084 20444 31104
rect 20444 31084 20496 31104
rect 20496 31084 20498 31104
rect 20442 31048 20498 31084
rect 19614 24792 19670 24848
rect 19890 25608 19946 25664
rect 19522 22480 19578 22536
rect 19522 22344 19578 22400
rect 19706 22480 19762 22536
rect 18694 16088 18750 16144
rect 18694 15136 18750 15192
rect 18263 14714 18319 14716
rect 18343 14714 18399 14716
rect 18423 14714 18479 14716
rect 18503 14714 18559 14716
rect 18263 14662 18309 14714
rect 18309 14662 18319 14714
rect 18343 14662 18373 14714
rect 18373 14662 18385 14714
rect 18385 14662 18399 14714
rect 18423 14662 18437 14714
rect 18437 14662 18449 14714
rect 18449 14662 18479 14714
rect 18503 14662 18513 14714
rect 18513 14662 18559 14714
rect 18263 14660 18319 14662
rect 18343 14660 18399 14662
rect 18423 14660 18479 14662
rect 18503 14660 18559 14662
rect 18234 14320 18290 14376
rect 18263 13626 18319 13628
rect 18343 13626 18399 13628
rect 18423 13626 18479 13628
rect 18503 13626 18559 13628
rect 18263 13574 18309 13626
rect 18309 13574 18319 13626
rect 18343 13574 18373 13626
rect 18373 13574 18385 13626
rect 18385 13574 18399 13626
rect 18423 13574 18437 13626
rect 18437 13574 18449 13626
rect 18449 13574 18479 13626
rect 18503 13574 18513 13626
rect 18513 13574 18559 13626
rect 18263 13572 18319 13574
rect 18343 13572 18399 13574
rect 18423 13572 18479 13574
rect 18503 13572 18559 13574
rect 18263 12538 18319 12540
rect 18343 12538 18399 12540
rect 18423 12538 18479 12540
rect 18503 12538 18559 12540
rect 18263 12486 18309 12538
rect 18309 12486 18319 12538
rect 18343 12486 18373 12538
rect 18373 12486 18385 12538
rect 18385 12486 18399 12538
rect 18423 12486 18437 12538
rect 18437 12486 18449 12538
rect 18449 12486 18479 12538
rect 18503 12486 18513 12538
rect 18513 12486 18559 12538
rect 18263 12484 18319 12486
rect 18343 12484 18399 12486
rect 18423 12484 18479 12486
rect 18503 12484 18559 12486
rect 17774 11600 17830 11656
rect 17774 10412 17776 10432
rect 17776 10412 17828 10432
rect 17828 10412 17830 10432
rect 17774 10376 17830 10412
rect 17682 10004 17684 10024
rect 17684 10004 17736 10024
rect 17736 10004 17738 10024
rect 17682 9968 17738 10004
rect 17958 11328 18014 11384
rect 17866 9968 17922 10024
rect 17314 8064 17370 8120
rect 17130 7248 17186 7304
rect 16854 6704 16910 6760
rect 15382 5208 15438 5264
rect 15790 5466 15846 5468
rect 15870 5466 15926 5468
rect 15950 5466 16006 5468
rect 16030 5466 16086 5468
rect 15790 5414 15836 5466
rect 15836 5414 15846 5466
rect 15870 5414 15900 5466
rect 15900 5414 15912 5466
rect 15912 5414 15926 5466
rect 15950 5414 15964 5466
rect 15964 5414 15976 5466
rect 15976 5414 16006 5466
rect 16030 5414 16040 5466
rect 16040 5414 16086 5466
rect 15790 5412 15846 5414
rect 15870 5412 15926 5414
rect 15950 5412 16006 5414
rect 16030 5412 16086 5414
rect 15750 5208 15806 5264
rect 16210 5480 16266 5536
rect 16762 6296 16818 6352
rect 14186 4428 14188 4448
rect 14188 4428 14240 4448
rect 14240 4428 14242 4448
rect 14186 4392 14242 4428
rect 14646 4528 14702 4584
rect 15658 4392 15714 4448
rect 15790 4378 15846 4380
rect 15870 4378 15926 4380
rect 15950 4378 16006 4380
rect 16030 4378 16086 4380
rect 15790 4326 15836 4378
rect 15836 4326 15846 4378
rect 15870 4326 15900 4378
rect 15900 4326 15912 4378
rect 15912 4326 15926 4378
rect 15950 4326 15964 4378
rect 15964 4326 15976 4378
rect 15976 4326 16006 4378
rect 16030 4326 16040 4378
rect 16040 4326 16086 4378
rect 15790 4324 15846 4326
rect 15870 4324 15926 4326
rect 15950 4324 16006 4326
rect 16030 4324 16086 4326
rect 15290 4256 15346 4312
rect 12806 3848 12862 3904
rect 13015 3848 13071 3904
rect 12438 3612 12440 3632
rect 12440 3612 12492 3632
rect 12492 3612 12494 3632
rect 11886 3168 11942 3224
rect 11886 3052 11942 3088
rect 11886 3032 11888 3052
rect 11888 3032 11940 3052
rect 11940 3032 11942 3052
rect 11794 2488 11850 2544
rect 12438 3576 12494 3612
rect 12898 3712 12954 3768
rect 13450 3984 13506 4040
rect 13910 3848 13966 3904
rect 13318 3834 13374 3836
rect 13398 3834 13454 3836
rect 13478 3834 13534 3836
rect 13558 3834 13614 3836
rect 13318 3782 13364 3834
rect 13364 3782 13374 3834
rect 13398 3782 13428 3834
rect 13428 3782 13440 3834
rect 13440 3782 13454 3834
rect 13478 3782 13492 3834
rect 13492 3782 13504 3834
rect 13504 3782 13534 3834
rect 13558 3782 13568 3834
rect 13568 3782 13614 3834
rect 13318 3780 13374 3782
rect 13398 3780 13454 3782
rect 13478 3780 13534 3782
rect 13558 3780 13614 3782
rect 12070 3052 12126 3088
rect 12070 3032 12072 3052
rect 12072 3032 12124 3052
rect 12124 3032 12126 3052
rect 12254 2760 12310 2816
rect 12438 3304 12494 3360
rect 12438 2760 12494 2816
rect 12714 3304 12770 3360
rect 12806 2896 12862 2952
rect 12990 3168 13046 3224
rect 12714 2488 12770 2544
rect 11794 1808 11850 1864
rect 11978 1808 12034 1864
rect 11794 1368 11796 1408
rect 11796 1368 11848 1408
rect 11848 1368 11850 1408
rect 11794 1352 11850 1368
rect 10845 1114 10901 1116
rect 10925 1114 10981 1116
rect 11005 1114 11061 1116
rect 11085 1114 11141 1116
rect 10845 1062 10891 1114
rect 10891 1062 10901 1114
rect 10925 1062 10955 1114
rect 10955 1062 10967 1114
rect 10967 1062 10981 1114
rect 11005 1062 11019 1114
rect 11019 1062 11031 1114
rect 11031 1062 11061 1114
rect 11085 1062 11095 1114
rect 11095 1062 11141 1114
rect 10845 1060 10901 1062
rect 10925 1060 10981 1062
rect 11005 1060 11061 1062
rect 11085 1060 11141 1062
rect 11150 856 11206 912
rect 11518 720 11574 776
rect 12438 2352 12494 2408
rect 14094 3712 14150 3768
rect 14738 3712 14794 3768
rect 14186 3168 14242 3224
rect 14370 3188 14426 3224
rect 14370 3168 14372 3188
rect 14372 3168 14424 3188
rect 14424 3168 14426 3188
rect 14830 3168 14886 3224
rect 13726 2760 13782 2816
rect 13318 2746 13374 2748
rect 13398 2746 13454 2748
rect 13478 2746 13534 2748
rect 13558 2746 13614 2748
rect 13318 2694 13364 2746
rect 13364 2694 13374 2746
rect 13398 2694 13428 2746
rect 13428 2694 13440 2746
rect 13440 2694 13454 2746
rect 13478 2694 13492 2746
rect 13492 2694 13504 2746
rect 13504 2694 13534 2746
rect 13558 2694 13568 2746
rect 13568 2694 13614 2746
rect 13318 2692 13374 2694
rect 13398 2692 13454 2694
rect 13478 2692 13534 2694
rect 13558 2692 13614 2694
rect 13818 2624 13874 2680
rect 14002 2624 14058 2680
rect 13726 2488 13782 2544
rect 12806 2216 12862 2272
rect 12990 2352 13046 2408
rect 13358 2216 13414 2272
rect 12622 2080 12678 2136
rect 12898 2080 12954 2136
rect 14002 2488 14058 2544
rect 14370 2760 14426 2816
rect 12622 1672 12678 1728
rect 12070 992 12126 1048
rect 12806 1672 12862 1728
rect 12530 1128 12586 1184
rect 12898 584 12954 640
rect 13318 1658 13374 1660
rect 13398 1658 13454 1660
rect 13478 1658 13534 1660
rect 13558 1658 13614 1660
rect 13318 1606 13364 1658
rect 13364 1606 13374 1658
rect 13398 1606 13428 1658
rect 13428 1606 13440 1658
rect 13440 1606 13454 1658
rect 13478 1606 13492 1658
rect 13492 1606 13504 1658
rect 13504 1606 13534 1658
rect 13558 1606 13568 1658
rect 13568 1606 13614 1658
rect 13318 1604 13374 1606
rect 13398 1604 13454 1606
rect 13478 1604 13534 1606
rect 13558 1604 13614 1606
rect 13358 1264 13414 1320
rect 13542 1300 13544 1320
rect 13544 1300 13596 1320
rect 13596 1300 13598 1320
rect 13542 1264 13598 1300
rect 13358 720 13414 776
rect 13542 756 13544 776
rect 13544 756 13596 776
rect 13596 756 13598 776
rect 13542 720 13598 756
rect 13266 620 13268 640
rect 13268 620 13320 640
rect 13320 620 13322 640
rect 13266 584 13322 620
rect 14186 1536 14242 1592
rect 14554 1944 14610 2000
rect 15106 3576 15162 3632
rect 15106 3304 15162 3360
rect 15106 3168 15162 3224
rect 15750 3848 15806 3904
rect 15474 3304 15530 3360
rect 15474 3168 15530 3224
rect 16302 4392 16358 4448
rect 16486 5228 16542 5264
rect 16486 5208 16488 5228
rect 16488 5208 16540 5228
rect 16540 5208 16542 5228
rect 16670 5752 16726 5808
rect 16854 5752 16910 5808
rect 16854 5208 16910 5264
rect 16854 4664 16910 4720
rect 17038 5344 17094 5400
rect 17038 4936 17094 4992
rect 16486 4120 16542 4176
rect 15842 3476 15844 3496
rect 15844 3476 15896 3496
rect 15896 3476 15898 3496
rect 15842 3440 15898 3476
rect 16026 3440 16082 3496
rect 16486 3848 16542 3904
rect 15790 3290 15846 3292
rect 15870 3290 15926 3292
rect 15950 3290 16006 3292
rect 16030 3290 16086 3292
rect 15790 3238 15836 3290
rect 15836 3238 15846 3290
rect 15870 3238 15900 3290
rect 15900 3238 15912 3290
rect 15912 3238 15926 3290
rect 15950 3238 15964 3290
rect 15964 3238 15976 3290
rect 15976 3238 16006 3290
rect 16030 3238 16040 3290
rect 16040 3238 16086 3290
rect 15790 3236 15846 3238
rect 15870 3236 15926 3238
rect 15950 3236 16006 3238
rect 16030 3236 16086 3238
rect 15658 3168 15714 3224
rect 16394 3304 16450 3360
rect 16302 3068 16304 3088
rect 16304 3068 16356 3088
rect 16356 3068 16358 3088
rect 14922 1980 14924 2000
rect 14924 1980 14976 2000
rect 14976 1980 14978 2000
rect 14922 1944 14978 1980
rect 14738 1264 14794 1320
rect 15382 2760 15438 2816
rect 16302 3032 16358 3068
rect 14646 312 14702 368
rect 15290 312 15346 368
rect 15790 2202 15846 2204
rect 15870 2202 15926 2204
rect 15950 2202 16006 2204
rect 16030 2202 16086 2204
rect 15790 2150 15836 2202
rect 15836 2150 15846 2202
rect 15870 2150 15900 2202
rect 15900 2150 15912 2202
rect 15912 2150 15926 2202
rect 15950 2150 15964 2202
rect 15964 2150 15976 2202
rect 15976 2150 16006 2202
rect 16030 2150 16040 2202
rect 16040 2150 16086 2202
rect 15790 2148 15846 2150
rect 15870 2148 15926 2150
rect 15950 2148 16006 2150
rect 16030 2148 16086 2150
rect 16946 3984 17002 4040
rect 16762 3712 16818 3768
rect 16762 3304 16818 3360
rect 16486 3168 16542 3224
rect 16670 3168 16726 3224
rect 16578 2896 16634 2952
rect 16486 2524 16488 2544
rect 16488 2524 16540 2544
rect 16540 2524 16542 2544
rect 16486 2488 16542 2524
rect 16486 2388 16488 2408
rect 16488 2388 16540 2408
rect 16540 2388 16542 2408
rect 16486 2352 16542 2388
rect 16210 2216 16266 2272
rect 15934 1400 15990 1456
rect 15790 1114 15846 1116
rect 15870 1114 15926 1116
rect 15950 1114 16006 1116
rect 16030 1114 16086 1116
rect 15790 1062 15836 1114
rect 15836 1062 15846 1114
rect 15870 1062 15900 1114
rect 15900 1062 15912 1114
rect 15912 1062 15926 1114
rect 15950 1062 15964 1114
rect 15964 1062 15976 1114
rect 15976 1062 16006 1114
rect 16030 1062 16040 1114
rect 16040 1062 16086 1114
rect 15790 1060 15846 1062
rect 15870 1060 15926 1062
rect 15950 1060 16006 1062
rect 16030 1060 16086 1062
rect 15750 312 15806 368
rect 16302 1300 16304 1320
rect 16304 1300 16356 1320
rect 16356 1300 16358 1320
rect 16302 1264 16358 1300
rect 16302 1164 16304 1184
rect 16304 1164 16356 1184
rect 16356 1164 16358 1184
rect 16302 1128 16358 1164
rect 16210 992 16266 1048
rect 16762 2352 16818 2408
rect 16946 2216 17002 2272
rect 16946 1536 17002 1592
rect 16762 740 16818 776
rect 16762 720 16764 740
rect 16764 720 16816 740
rect 16816 720 16818 740
rect 18263 11450 18319 11452
rect 18343 11450 18399 11452
rect 18423 11450 18479 11452
rect 18503 11450 18559 11452
rect 18263 11398 18309 11450
rect 18309 11398 18319 11450
rect 18343 11398 18373 11450
rect 18373 11398 18385 11450
rect 18385 11398 18399 11450
rect 18423 11398 18437 11450
rect 18437 11398 18449 11450
rect 18449 11398 18479 11450
rect 18503 11398 18513 11450
rect 18513 11398 18559 11450
rect 18263 11396 18319 11398
rect 18343 11396 18399 11398
rect 18423 11396 18479 11398
rect 18503 11396 18559 11398
rect 19062 12552 19118 12608
rect 20442 29996 20444 30016
rect 20444 29996 20496 30016
rect 20496 29996 20498 30016
rect 19890 21292 19892 21312
rect 19892 21292 19944 21312
rect 19944 21292 19946 21312
rect 19890 21256 19946 21292
rect 19798 17040 19854 17096
rect 19522 15952 19578 16008
rect 19522 13640 19578 13696
rect 19338 12144 19394 12200
rect 18970 11192 19026 11248
rect 18263 10362 18319 10364
rect 18343 10362 18399 10364
rect 18423 10362 18479 10364
rect 18503 10362 18559 10364
rect 18263 10310 18309 10362
rect 18309 10310 18319 10362
rect 18343 10310 18373 10362
rect 18373 10310 18385 10362
rect 18385 10310 18399 10362
rect 18423 10310 18437 10362
rect 18437 10310 18449 10362
rect 18449 10310 18479 10362
rect 18503 10310 18513 10362
rect 18513 10310 18559 10362
rect 18263 10308 18319 10310
rect 18343 10308 18399 10310
rect 18423 10308 18479 10310
rect 18503 10308 18559 10310
rect 18510 9968 18566 10024
rect 18786 10920 18842 10976
rect 18694 9968 18750 10024
rect 18050 9152 18106 9208
rect 17682 7384 17738 7440
rect 17590 7248 17646 7304
rect 17682 6024 17738 6080
rect 17682 5752 17738 5808
rect 17498 4800 17554 4856
rect 18263 9274 18319 9276
rect 18343 9274 18399 9276
rect 18423 9274 18479 9276
rect 18503 9274 18559 9276
rect 18263 9222 18309 9274
rect 18309 9222 18319 9274
rect 18343 9222 18373 9274
rect 18373 9222 18385 9274
rect 18385 9222 18399 9274
rect 18423 9222 18437 9274
rect 18437 9222 18449 9274
rect 18449 9222 18479 9274
rect 18503 9222 18513 9274
rect 18513 9222 18559 9274
rect 18263 9220 18319 9222
rect 18343 9220 18399 9222
rect 18423 9220 18479 9222
rect 18503 9220 18559 9222
rect 18694 9152 18750 9208
rect 18326 8900 18382 8936
rect 18326 8880 18328 8900
rect 18328 8880 18380 8900
rect 18380 8880 18382 8900
rect 18878 9016 18934 9072
rect 18694 8472 18750 8528
rect 18050 8200 18106 8256
rect 18263 8186 18319 8188
rect 18343 8186 18399 8188
rect 18423 8186 18479 8188
rect 18503 8186 18559 8188
rect 18263 8134 18309 8186
rect 18309 8134 18319 8186
rect 18343 8134 18373 8186
rect 18373 8134 18385 8186
rect 18385 8134 18399 8186
rect 18423 8134 18437 8186
rect 18437 8134 18449 8186
rect 18449 8134 18479 8186
rect 18503 8134 18513 8186
rect 18513 8134 18559 8186
rect 18263 8132 18319 8134
rect 18343 8132 18399 8134
rect 18423 8132 18479 8134
rect 18503 8132 18559 8134
rect 18263 7098 18319 7100
rect 18343 7098 18399 7100
rect 18423 7098 18479 7100
rect 18503 7098 18559 7100
rect 18263 7046 18309 7098
rect 18309 7046 18319 7098
rect 18343 7046 18373 7098
rect 18373 7046 18385 7098
rect 18385 7046 18399 7098
rect 18423 7046 18437 7098
rect 18437 7046 18449 7098
rect 18449 7046 18479 7098
rect 18503 7046 18513 7098
rect 18513 7046 18559 7098
rect 18263 7044 18319 7046
rect 18343 7044 18399 7046
rect 18423 7044 18479 7046
rect 18503 7044 18559 7046
rect 18050 6976 18106 7032
rect 18234 6432 18290 6488
rect 17590 3848 17646 3904
rect 17498 3712 17554 3768
rect 17314 1672 17370 1728
rect 17958 5344 18014 5400
rect 17590 584 17646 640
rect 17774 2080 17830 2136
rect 17958 2352 18014 2408
rect 18510 6568 18566 6624
rect 18510 6432 18566 6488
rect 18263 6010 18319 6012
rect 18343 6010 18399 6012
rect 18423 6010 18479 6012
rect 18503 6010 18559 6012
rect 18263 5958 18309 6010
rect 18309 5958 18319 6010
rect 18343 5958 18373 6010
rect 18373 5958 18385 6010
rect 18385 5958 18399 6010
rect 18423 5958 18437 6010
rect 18437 5958 18449 6010
rect 18449 5958 18479 6010
rect 18503 5958 18513 6010
rect 18513 5958 18559 6010
rect 18263 5956 18319 5958
rect 18343 5956 18399 5958
rect 18423 5956 18479 5958
rect 18503 5956 18559 5958
rect 18142 5480 18198 5536
rect 18878 7656 18934 7712
rect 19062 11056 19118 11112
rect 18878 6432 18934 6488
rect 19430 11464 19486 11520
rect 19430 9696 19486 9752
rect 19154 9152 19210 9208
rect 18786 5480 18842 5536
rect 18263 4922 18319 4924
rect 18343 4922 18399 4924
rect 18423 4922 18479 4924
rect 18503 4922 18559 4924
rect 18263 4870 18309 4922
rect 18309 4870 18319 4922
rect 18343 4870 18373 4922
rect 18373 4870 18385 4922
rect 18385 4870 18399 4922
rect 18423 4870 18437 4922
rect 18437 4870 18449 4922
rect 18449 4870 18479 4922
rect 18503 4870 18513 4922
rect 18513 4870 18559 4922
rect 18263 4868 18319 4870
rect 18343 4868 18399 4870
rect 18423 4868 18479 4870
rect 18503 4868 18559 4870
rect 18234 4664 18290 4720
rect 18263 3834 18319 3836
rect 18343 3834 18399 3836
rect 18423 3834 18479 3836
rect 18503 3834 18559 3836
rect 18263 3782 18309 3834
rect 18309 3782 18319 3834
rect 18343 3782 18373 3834
rect 18373 3782 18385 3834
rect 18385 3782 18399 3834
rect 18423 3782 18437 3834
rect 18437 3782 18449 3834
rect 18449 3782 18479 3834
rect 18503 3782 18513 3834
rect 18513 3782 18559 3834
rect 18263 3780 18319 3782
rect 18343 3780 18399 3782
rect 18423 3780 18479 3782
rect 18503 3780 18559 3782
rect 18234 3576 18290 3632
rect 18050 1264 18106 1320
rect 18694 3848 18750 3904
rect 18602 3440 18658 3496
rect 18602 3304 18658 3360
rect 19338 9288 19394 9344
rect 19522 9016 19578 9072
rect 19246 8744 19302 8800
rect 20258 26460 20260 26480
rect 20260 26460 20312 26480
rect 20312 26460 20314 26480
rect 20258 26424 20314 26460
rect 20258 24556 20260 24576
rect 20260 24556 20312 24576
rect 20312 24556 20314 24576
rect 20258 24520 20314 24556
rect 20442 29960 20498 29996
rect 20442 28872 20498 28928
rect 20442 28364 20444 28384
rect 20444 28364 20496 28384
rect 20496 28364 20498 28384
rect 20442 28328 20498 28364
rect 20442 27820 20444 27840
rect 20444 27820 20496 27840
rect 20496 27820 20498 27840
rect 20442 27784 20498 27820
rect 20626 31184 20682 31240
rect 20735 30490 20791 30492
rect 20815 30490 20871 30492
rect 20895 30490 20951 30492
rect 20975 30490 21031 30492
rect 20735 30438 20781 30490
rect 20781 30438 20791 30490
rect 20815 30438 20845 30490
rect 20845 30438 20857 30490
rect 20857 30438 20871 30490
rect 20895 30438 20909 30490
rect 20909 30438 20921 30490
rect 20921 30438 20951 30490
rect 20975 30438 20985 30490
rect 20985 30438 21031 30490
rect 20735 30436 20791 30438
rect 20815 30436 20871 30438
rect 20895 30436 20951 30438
rect 20975 30436 21031 30438
rect 20735 29402 20791 29404
rect 20815 29402 20871 29404
rect 20895 29402 20951 29404
rect 20975 29402 21031 29404
rect 20735 29350 20781 29402
rect 20781 29350 20791 29402
rect 20815 29350 20845 29402
rect 20845 29350 20857 29402
rect 20857 29350 20871 29402
rect 20895 29350 20909 29402
rect 20909 29350 20921 29402
rect 20921 29350 20951 29402
rect 20975 29350 20985 29402
rect 20985 29350 21031 29402
rect 20735 29348 20791 29350
rect 20815 29348 20871 29350
rect 20895 29348 20951 29350
rect 20975 29348 21031 29350
rect 20735 28314 20791 28316
rect 20815 28314 20871 28316
rect 20895 28314 20951 28316
rect 20975 28314 21031 28316
rect 20735 28262 20781 28314
rect 20781 28262 20791 28314
rect 20815 28262 20845 28314
rect 20845 28262 20857 28314
rect 20857 28262 20871 28314
rect 20895 28262 20909 28314
rect 20909 28262 20921 28314
rect 20921 28262 20951 28314
rect 20975 28262 20985 28314
rect 20985 28262 21031 28314
rect 20735 28260 20791 28262
rect 20815 28260 20871 28262
rect 20895 28260 20951 28262
rect 20975 28260 21031 28262
rect 20626 27512 20682 27568
rect 20735 27226 20791 27228
rect 20815 27226 20871 27228
rect 20895 27226 20951 27228
rect 20975 27226 21031 27228
rect 20735 27174 20781 27226
rect 20781 27174 20791 27226
rect 20815 27174 20845 27226
rect 20845 27174 20857 27226
rect 20857 27174 20871 27226
rect 20895 27174 20909 27226
rect 20909 27174 20921 27226
rect 20921 27174 20951 27226
rect 20975 27174 20985 27226
rect 20985 27174 21031 27226
rect 20735 27172 20791 27174
rect 20815 27172 20871 27174
rect 20895 27172 20951 27174
rect 20975 27172 21031 27174
rect 20534 26696 20590 26752
rect 20442 24112 20498 24168
rect 20735 26138 20791 26140
rect 20815 26138 20871 26140
rect 20895 26138 20951 26140
rect 20975 26138 21031 26140
rect 20735 26086 20781 26138
rect 20781 26086 20791 26138
rect 20815 26086 20845 26138
rect 20845 26086 20857 26138
rect 20857 26086 20871 26138
rect 20895 26086 20909 26138
rect 20909 26086 20921 26138
rect 20921 26086 20951 26138
rect 20975 26086 20985 26138
rect 20985 26086 21031 26138
rect 20735 26084 20791 26086
rect 20815 26084 20871 26086
rect 20895 26084 20951 26086
rect 20975 26084 21031 26086
rect 20626 25336 20682 25392
rect 20735 25050 20791 25052
rect 20815 25050 20871 25052
rect 20895 25050 20951 25052
rect 20975 25050 21031 25052
rect 20735 24998 20781 25050
rect 20781 24998 20791 25050
rect 20815 24998 20845 25050
rect 20845 24998 20857 25050
rect 20857 24998 20871 25050
rect 20895 24998 20909 25050
rect 20909 24998 20921 25050
rect 20921 24998 20951 25050
rect 20975 24998 20985 25050
rect 20985 24998 21031 25050
rect 20735 24996 20791 24998
rect 20815 24996 20871 24998
rect 20895 24996 20951 24998
rect 20975 24996 21031 24998
rect 20442 23468 20444 23488
rect 20444 23468 20496 23488
rect 20496 23468 20498 23488
rect 20442 23432 20498 23468
rect 20442 22380 20444 22400
rect 20444 22380 20496 22400
rect 20496 22380 20498 22400
rect 20442 22344 20498 22380
rect 20074 19116 20076 19136
rect 20076 19116 20128 19136
rect 20128 19116 20130 19136
rect 20074 19080 20130 19116
rect 19982 17040 20038 17096
rect 19890 12144 19946 12200
rect 19798 11600 19854 11656
rect 19706 9832 19762 9888
rect 19430 8608 19486 8664
rect 19338 8064 19394 8120
rect 19890 9424 19946 9480
rect 19890 7828 19892 7848
rect 19892 7828 19944 7848
rect 19944 7828 19946 7848
rect 19890 7792 19946 7828
rect 19706 6704 19762 6760
rect 19522 6432 19578 6488
rect 19430 5072 19486 5128
rect 19246 4256 19302 4312
rect 18878 3168 18934 3224
rect 18878 2760 18934 2816
rect 18263 2746 18319 2748
rect 18343 2746 18399 2748
rect 18423 2746 18479 2748
rect 18503 2746 18559 2748
rect 18263 2694 18309 2746
rect 18309 2694 18319 2746
rect 18343 2694 18373 2746
rect 18373 2694 18385 2746
rect 18385 2694 18399 2746
rect 18423 2694 18437 2746
rect 18437 2694 18449 2746
rect 18449 2694 18479 2746
rect 18503 2694 18513 2746
rect 18513 2694 18559 2746
rect 18263 2692 18319 2694
rect 18343 2692 18399 2694
rect 18423 2692 18479 2694
rect 18503 2692 18559 2694
rect 18263 1658 18319 1660
rect 18343 1658 18399 1660
rect 18423 1658 18479 1660
rect 18503 1658 18559 1660
rect 18263 1606 18309 1658
rect 18309 1606 18319 1658
rect 18343 1606 18373 1658
rect 18373 1606 18385 1658
rect 18385 1606 18399 1658
rect 18423 1606 18437 1658
rect 18437 1606 18449 1658
rect 18449 1606 18479 1658
rect 18503 1606 18513 1658
rect 18513 1606 18559 1658
rect 18263 1604 18319 1606
rect 18343 1604 18399 1606
rect 18423 1604 18479 1606
rect 18503 1604 18559 1606
rect 18418 856 18474 912
rect 18142 448 18198 504
rect 18970 992 19026 1048
rect 18786 312 18842 368
rect 18510 176 18566 232
rect 17956 40 18012 96
rect 19062 720 19118 776
rect 20166 10512 20222 10568
rect 20074 8336 20130 8392
rect 20442 16496 20498 16552
rect 20442 15852 20444 15872
rect 20444 15852 20496 15872
rect 20496 15852 20498 15872
rect 20442 15816 20498 15852
rect 20442 14764 20444 14784
rect 20444 14764 20496 14784
rect 20496 14764 20498 14784
rect 20442 14728 20498 14764
rect 20534 10376 20590 10432
rect 20350 9288 20406 9344
rect 20735 23962 20791 23964
rect 20815 23962 20871 23964
rect 20895 23962 20951 23964
rect 20975 23962 21031 23964
rect 20735 23910 20781 23962
rect 20781 23910 20791 23962
rect 20815 23910 20845 23962
rect 20845 23910 20857 23962
rect 20857 23910 20871 23962
rect 20895 23910 20909 23962
rect 20909 23910 20921 23962
rect 20921 23910 20951 23962
rect 20975 23910 20985 23962
rect 20985 23910 21031 23962
rect 20735 23908 20791 23910
rect 20815 23908 20871 23910
rect 20895 23908 20951 23910
rect 20975 23908 21031 23910
rect 20735 22874 20791 22876
rect 20815 22874 20871 22876
rect 20895 22874 20951 22876
rect 20975 22874 21031 22876
rect 20735 22822 20781 22874
rect 20781 22822 20791 22874
rect 20815 22822 20845 22874
rect 20845 22822 20857 22874
rect 20857 22822 20871 22874
rect 20895 22822 20909 22874
rect 20909 22822 20921 22874
rect 20921 22822 20951 22874
rect 20975 22822 20985 22874
rect 20985 22822 21031 22874
rect 20735 22820 20791 22822
rect 20815 22820 20871 22822
rect 20895 22820 20951 22822
rect 20975 22820 21031 22822
rect 20735 21786 20791 21788
rect 20815 21786 20871 21788
rect 20895 21786 20951 21788
rect 20975 21786 21031 21788
rect 20735 21734 20781 21786
rect 20781 21734 20791 21786
rect 20815 21734 20845 21786
rect 20845 21734 20857 21786
rect 20857 21734 20871 21786
rect 20895 21734 20909 21786
rect 20909 21734 20921 21786
rect 20921 21734 20951 21786
rect 20975 21734 20985 21786
rect 20985 21734 21031 21786
rect 20735 21732 20791 21734
rect 20815 21732 20871 21734
rect 20895 21732 20951 21734
rect 20975 21732 21031 21734
rect 20735 20698 20791 20700
rect 20815 20698 20871 20700
rect 20895 20698 20951 20700
rect 20975 20698 21031 20700
rect 20735 20646 20781 20698
rect 20781 20646 20791 20698
rect 20815 20646 20845 20698
rect 20845 20646 20857 20698
rect 20857 20646 20871 20698
rect 20895 20646 20909 20698
rect 20909 20646 20921 20698
rect 20921 20646 20951 20698
rect 20975 20646 20985 20698
rect 20985 20646 21031 20698
rect 20735 20644 20791 20646
rect 20815 20644 20871 20646
rect 20895 20644 20951 20646
rect 20975 20644 21031 20646
rect 21270 40296 21326 40352
rect 21178 39344 21234 39400
rect 21270 39208 21326 39264
rect 21454 38256 21510 38312
rect 21270 38120 21326 38176
rect 21270 35944 21326 36000
rect 21270 34892 21272 34912
rect 21272 34892 21324 34912
rect 21324 34892 21326 34912
rect 21270 34856 21326 34892
rect 21178 33804 21180 33824
rect 21180 33804 21232 33824
rect 21232 33804 21234 33824
rect 21178 33768 21234 33804
rect 20735 19610 20791 19612
rect 20815 19610 20871 19612
rect 20895 19610 20951 19612
rect 20975 19610 21031 19612
rect 20735 19558 20781 19610
rect 20781 19558 20791 19610
rect 20815 19558 20845 19610
rect 20845 19558 20857 19610
rect 20857 19558 20871 19610
rect 20895 19558 20909 19610
rect 20909 19558 20921 19610
rect 20921 19558 20951 19610
rect 20975 19558 20985 19610
rect 20985 19558 21031 19610
rect 20735 19556 20791 19558
rect 20815 19556 20871 19558
rect 20895 19556 20951 19558
rect 20975 19556 21031 19558
rect 20735 18522 20791 18524
rect 20815 18522 20871 18524
rect 20895 18522 20951 18524
rect 20975 18522 21031 18524
rect 20735 18470 20781 18522
rect 20781 18470 20791 18522
rect 20815 18470 20845 18522
rect 20845 18470 20857 18522
rect 20857 18470 20871 18522
rect 20895 18470 20909 18522
rect 20909 18470 20921 18522
rect 20921 18470 20951 18522
rect 20975 18470 20985 18522
rect 20985 18470 21031 18522
rect 20735 18468 20791 18470
rect 20815 18468 20871 18470
rect 20895 18468 20951 18470
rect 20975 18468 21031 18470
rect 20994 18028 20996 18048
rect 20996 18028 21048 18048
rect 21048 18028 21050 18048
rect 20994 17992 21050 18028
rect 20735 17434 20791 17436
rect 20815 17434 20871 17436
rect 20895 17434 20951 17436
rect 20975 17434 21031 17436
rect 20735 17382 20781 17434
rect 20781 17382 20791 17434
rect 20815 17382 20845 17434
rect 20845 17382 20857 17434
rect 20857 17382 20871 17434
rect 20895 17382 20909 17434
rect 20909 17382 20921 17434
rect 20921 17382 20951 17434
rect 20975 17382 20985 17434
rect 20985 17382 21031 17434
rect 20735 17380 20791 17382
rect 20815 17380 20871 17382
rect 20895 17380 20951 17382
rect 20975 17380 21031 17382
rect 20902 16940 20904 16960
rect 20904 16940 20956 16960
rect 20956 16940 20958 16960
rect 20902 16904 20958 16940
rect 20735 16346 20791 16348
rect 20815 16346 20871 16348
rect 20895 16346 20951 16348
rect 20975 16346 21031 16348
rect 20735 16294 20781 16346
rect 20781 16294 20791 16346
rect 20815 16294 20845 16346
rect 20845 16294 20857 16346
rect 20857 16294 20871 16346
rect 20895 16294 20909 16346
rect 20909 16294 20921 16346
rect 20921 16294 20951 16346
rect 20975 16294 20985 16346
rect 20985 16294 21031 16346
rect 20735 16292 20791 16294
rect 20815 16292 20871 16294
rect 20895 16292 20951 16294
rect 20975 16292 21031 16294
rect 20735 15258 20791 15260
rect 20815 15258 20871 15260
rect 20895 15258 20951 15260
rect 20975 15258 21031 15260
rect 20735 15206 20781 15258
rect 20781 15206 20791 15258
rect 20815 15206 20845 15258
rect 20845 15206 20857 15258
rect 20857 15206 20871 15258
rect 20895 15206 20909 15258
rect 20909 15206 20921 15258
rect 20921 15206 20951 15258
rect 20975 15206 20985 15258
rect 20985 15206 21031 15258
rect 20735 15204 20791 15206
rect 20815 15204 20871 15206
rect 20895 15204 20951 15206
rect 20975 15204 21031 15206
rect 20735 14170 20791 14172
rect 20815 14170 20871 14172
rect 20895 14170 20951 14172
rect 20975 14170 21031 14172
rect 20735 14118 20781 14170
rect 20781 14118 20791 14170
rect 20815 14118 20845 14170
rect 20845 14118 20857 14170
rect 20857 14118 20871 14170
rect 20895 14118 20909 14170
rect 20909 14118 20921 14170
rect 20921 14118 20951 14170
rect 20975 14118 20985 14170
rect 20985 14118 21031 14170
rect 20735 14116 20791 14118
rect 20815 14116 20871 14118
rect 20895 14116 20951 14118
rect 20975 14116 21031 14118
rect 20735 13082 20791 13084
rect 20815 13082 20871 13084
rect 20895 13082 20951 13084
rect 20975 13082 21031 13084
rect 20735 13030 20781 13082
rect 20781 13030 20791 13082
rect 20815 13030 20845 13082
rect 20845 13030 20857 13082
rect 20857 13030 20871 13082
rect 20895 13030 20909 13082
rect 20909 13030 20921 13082
rect 20921 13030 20951 13082
rect 20975 13030 20985 13082
rect 20985 13030 21031 13082
rect 20735 13028 20791 13030
rect 20815 13028 20871 13030
rect 20895 13028 20951 13030
rect 20975 13028 21031 13030
rect 20735 11994 20791 11996
rect 20815 11994 20871 11996
rect 20895 11994 20951 11996
rect 20975 11994 21031 11996
rect 20735 11942 20781 11994
rect 20781 11942 20791 11994
rect 20815 11942 20845 11994
rect 20845 11942 20857 11994
rect 20857 11942 20871 11994
rect 20895 11942 20909 11994
rect 20909 11942 20921 11994
rect 20921 11942 20951 11994
rect 20975 11942 20985 11994
rect 20985 11942 21031 11994
rect 20735 11940 20791 11942
rect 20815 11940 20871 11942
rect 20895 11940 20951 11942
rect 20975 11940 21031 11942
rect 20735 10906 20791 10908
rect 20815 10906 20871 10908
rect 20895 10906 20951 10908
rect 20975 10906 21031 10908
rect 20735 10854 20781 10906
rect 20781 10854 20791 10906
rect 20815 10854 20845 10906
rect 20845 10854 20857 10906
rect 20857 10854 20871 10906
rect 20895 10854 20909 10906
rect 20909 10854 20921 10906
rect 20921 10854 20951 10906
rect 20975 10854 20985 10906
rect 20985 10854 21031 10906
rect 20735 10852 20791 10854
rect 20815 10852 20871 10854
rect 20895 10852 20951 10854
rect 20975 10852 21031 10854
rect 20735 9818 20791 9820
rect 20815 9818 20871 9820
rect 20895 9818 20951 9820
rect 20975 9818 21031 9820
rect 20735 9766 20781 9818
rect 20781 9766 20791 9818
rect 20815 9766 20845 9818
rect 20845 9766 20857 9818
rect 20857 9766 20871 9818
rect 20895 9766 20909 9818
rect 20909 9766 20921 9818
rect 20921 9766 20951 9818
rect 20975 9766 20985 9818
rect 20985 9766 21031 9818
rect 20735 9764 20791 9766
rect 20815 9764 20871 9766
rect 20895 9764 20951 9766
rect 20975 9764 21031 9766
rect 20735 8730 20791 8732
rect 20815 8730 20871 8732
rect 20895 8730 20951 8732
rect 20975 8730 21031 8732
rect 20735 8678 20781 8730
rect 20781 8678 20791 8730
rect 20815 8678 20845 8730
rect 20845 8678 20857 8730
rect 20857 8678 20871 8730
rect 20895 8678 20909 8730
rect 20909 8678 20921 8730
rect 20921 8678 20951 8730
rect 20975 8678 20985 8730
rect 20985 8678 21031 8730
rect 20735 8676 20791 8678
rect 20815 8676 20871 8678
rect 20895 8676 20951 8678
rect 20975 8676 21031 8678
rect 20735 7642 20791 7644
rect 20815 7642 20871 7644
rect 20895 7642 20951 7644
rect 20975 7642 21031 7644
rect 20735 7590 20781 7642
rect 20781 7590 20791 7642
rect 20815 7590 20845 7642
rect 20845 7590 20857 7642
rect 20857 7590 20871 7642
rect 20895 7590 20909 7642
rect 20909 7590 20921 7642
rect 20921 7590 20951 7642
rect 20975 7590 20985 7642
rect 20985 7590 21031 7642
rect 20735 7588 20791 7590
rect 20815 7588 20871 7590
rect 20895 7588 20951 7590
rect 20975 7588 21031 7590
rect 19614 2896 19670 2952
rect 19614 2760 19670 2816
rect 19890 4528 19946 4584
rect 20735 6554 20791 6556
rect 20815 6554 20871 6556
rect 20895 6554 20951 6556
rect 20975 6554 21031 6556
rect 20735 6502 20781 6554
rect 20781 6502 20791 6554
rect 20815 6502 20845 6554
rect 20845 6502 20857 6554
rect 20857 6502 20871 6554
rect 20895 6502 20909 6554
rect 20909 6502 20921 6554
rect 20921 6502 20951 6554
rect 20975 6502 20985 6554
rect 20985 6502 21031 6554
rect 20735 6500 20791 6502
rect 20815 6500 20871 6502
rect 20895 6500 20951 6502
rect 20975 6500 21031 6502
rect 20735 5466 20791 5468
rect 20815 5466 20871 5468
rect 20895 5466 20951 5468
rect 20975 5466 21031 5468
rect 20735 5414 20781 5466
rect 20781 5414 20791 5466
rect 20815 5414 20845 5466
rect 20845 5414 20857 5466
rect 20857 5414 20871 5466
rect 20895 5414 20909 5466
rect 20909 5414 20921 5466
rect 20921 5414 20951 5466
rect 20975 5414 20985 5466
rect 20985 5414 21031 5466
rect 20735 5412 20791 5414
rect 20815 5412 20871 5414
rect 20895 5412 20951 5414
rect 20975 5412 21031 5414
rect 20735 4378 20791 4380
rect 20815 4378 20871 4380
rect 20895 4378 20951 4380
rect 20975 4378 21031 4380
rect 20735 4326 20781 4378
rect 20781 4326 20791 4378
rect 20815 4326 20845 4378
rect 20845 4326 20857 4378
rect 20857 4326 20871 4378
rect 20895 4326 20909 4378
rect 20909 4326 20921 4378
rect 20921 4326 20951 4378
rect 20975 4326 20985 4378
rect 20985 4326 21031 4378
rect 20735 4324 20791 4326
rect 20815 4324 20871 4326
rect 20895 4324 20951 4326
rect 20975 4324 21031 4326
rect 21270 32680 21326 32736
rect 21270 30504 21326 30560
rect 21270 29416 21326 29472
rect 21270 29144 21326 29200
rect 21270 27240 21326 27296
rect 21270 26152 21326 26208
rect 21270 22888 21326 22944
rect 21270 21800 21326 21856
rect 21270 20712 21326 20768
rect 21270 18536 21326 18592
rect 21270 17448 21326 17504
rect 21270 15272 21326 15328
rect 21270 14184 21326 14240
rect 21270 13096 21326 13152
rect 21730 36624 21786 36680
rect 21822 28056 21878 28112
rect 21546 20168 21602 20224
rect 21546 19624 21602 19680
rect 21454 18672 21510 18728
rect 21730 20848 21786 20904
rect 21822 18264 21878 18320
rect 21730 16632 21786 16688
rect 21638 12688 21694 12744
rect 21270 10920 21326 10976
rect 21270 3340 21272 3360
rect 21272 3340 21324 3360
rect 21324 3340 21326 3360
rect 21270 3304 21326 3340
rect 20735 3290 20791 3292
rect 20815 3290 20871 3292
rect 20895 3290 20951 3292
rect 20975 3290 21031 3292
rect 20735 3238 20781 3290
rect 20781 3238 20791 3290
rect 20815 3238 20845 3290
rect 20845 3238 20857 3290
rect 20857 3238 20871 3290
rect 20895 3238 20909 3290
rect 20909 3238 20921 3290
rect 20921 3238 20951 3290
rect 20975 3238 20985 3290
rect 20985 3238 21031 3290
rect 20735 3236 20791 3238
rect 20815 3236 20871 3238
rect 20895 3236 20951 3238
rect 20975 3236 21031 3238
rect 20735 2202 20791 2204
rect 20815 2202 20871 2204
rect 20895 2202 20951 2204
rect 20975 2202 21031 2204
rect 20735 2150 20781 2202
rect 20781 2150 20791 2202
rect 20815 2150 20845 2202
rect 20845 2150 20857 2202
rect 20857 2150 20871 2202
rect 20895 2150 20909 2202
rect 20909 2150 20921 2202
rect 20921 2150 20951 2202
rect 20975 2150 20985 2202
rect 20985 2150 21031 2202
rect 20735 2148 20791 2150
rect 20815 2148 20871 2150
rect 20895 2148 20951 2150
rect 20975 2148 21031 2150
rect 21178 1128 21234 1184
rect 20735 1114 20791 1116
rect 20815 1114 20871 1116
rect 20895 1114 20951 1116
rect 20975 1114 21031 1116
rect 20735 1062 20781 1114
rect 20781 1062 20791 1114
rect 20815 1062 20845 1114
rect 20845 1062 20857 1114
rect 20857 1062 20871 1114
rect 20895 1062 20909 1114
rect 20909 1062 20921 1114
rect 20921 1062 20951 1114
rect 20975 1062 20985 1114
rect 20985 1062 21031 1114
rect 20735 1060 20791 1062
rect 20815 1060 20871 1062
rect 20895 1060 20951 1062
rect 20975 1060 21031 1062
<< metal3 >>
rect 14590 44508 14596 44572
rect 14660 44570 14666 44572
rect 15377 44570 15443 44573
rect 14660 44568 15443 44570
rect 14660 44512 15382 44568
rect 15438 44512 15443 44568
rect 14660 44510 15443 44512
rect 14660 44508 14666 44510
rect 15377 44507 15443 44510
rect 14181 44026 14247 44029
rect 19977 44026 20043 44029
rect 14181 44024 20043 44026
rect 14181 43968 14186 44024
rect 14242 43968 19982 44024
rect 20038 43968 20043 44024
rect 14181 43966 20043 43968
rect 14181 43963 14247 43966
rect 19977 43963 20043 43966
rect 4153 43890 4219 43893
rect 6269 43890 6335 43893
rect 4153 43888 6335 43890
rect 4153 43832 4158 43888
rect 4214 43832 6274 43888
rect 6330 43832 6335 43888
rect 4153 43830 6335 43832
rect 4153 43827 4219 43830
rect 6269 43827 6335 43830
rect 13813 43890 13879 43893
rect 15469 43890 15535 43893
rect 13813 43888 15535 43890
rect 13813 43832 13818 43888
rect 13874 43832 15474 43888
rect 15530 43832 15535 43888
rect 13813 43830 15535 43832
rect 13813 43827 13879 43830
rect 15469 43827 15535 43830
rect 15653 43754 15719 43757
rect 16614 43754 16620 43756
rect 15653 43752 16620 43754
rect 15653 43696 15658 43752
rect 15714 43696 16620 43752
rect 15653 43694 16620 43696
rect 15653 43691 15719 43694
rect 16614 43692 16620 43694
rect 16684 43692 16690 43756
rect 21173 43618 21239 43621
rect 21840 43618 22300 43648
rect 21173 43616 22300 43618
rect 21173 43560 21178 43616
rect 21234 43560 22300 43616
rect 21173 43558 22300 43560
rect 21173 43555 21239 43558
rect 5890 43552 6206 43553
rect 5890 43488 5896 43552
rect 5960 43488 5976 43552
rect 6040 43488 6056 43552
rect 6120 43488 6136 43552
rect 6200 43488 6206 43552
rect 5890 43487 6206 43488
rect 10835 43552 11151 43553
rect 10835 43488 10841 43552
rect 10905 43488 10921 43552
rect 10985 43488 11001 43552
rect 11065 43488 11081 43552
rect 11145 43488 11151 43552
rect 10835 43487 11151 43488
rect 15780 43552 16096 43553
rect 15780 43488 15786 43552
rect 15850 43488 15866 43552
rect 15930 43488 15946 43552
rect 16010 43488 16026 43552
rect 16090 43488 16096 43552
rect 15780 43487 16096 43488
rect 20725 43552 21041 43553
rect 20725 43488 20731 43552
rect 20795 43488 20811 43552
rect 20875 43488 20891 43552
rect 20955 43488 20971 43552
rect 21035 43488 21041 43552
rect 21840 43528 22300 43558
rect 20725 43487 21041 43488
rect 10225 43482 10291 43485
rect 10225 43480 10426 43482
rect 10225 43424 10230 43480
rect 10286 43424 10426 43480
rect 10225 43422 10426 43424
rect 10225 43419 10291 43422
rect 10366 43346 10426 43422
rect 10593 43346 10659 43349
rect 10366 43344 10659 43346
rect 10366 43288 10598 43344
rect 10654 43288 10659 43344
rect 10366 43286 10659 43288
rect 10593 43283 10659 43286
rect 13905 43346 13971 43349
rect 18689 43346 18755 43349
rect 13905 43344 18755 43346
rect 13905 43288 13910 43344
rect 13966 43288 18694 43344
rect 18750 43288 18755 43344
rect 13905 43286 18755 43288
rect 13905 43283 13971 43286
rect 18689 43283 18755 43286
rect 5022 43148 5028 43212
rect 5092 43210 5098 43212
rect 13537 43210 13603 43213
rect 5092 43208 13603 43210
rect 5092 43152 13542 43208
rect 13598 43152 13603 43208
rect 5092 43150 13603 43152
rect 5092 43148 5098 43150
rect 13537 43147 13603 43150
rect 16113 43210 16179 43213
rect 16246 43210 16252 43212
rect 16113 43208 16252 43210
rect 16113 43152 16118 43208
rect 16174 43152 16252 43208
rect 16113 43150 16252 43152
rect 16113 43147 16179 43150
rect 16246 43148 16252 43150
rect 16316 43148 16322 43212
rect 18873 43210 18939 43213
rect 16392 43208 18939 43210
rect 16392 43152 18878 43208
rect 18934 43152 18939 43208
rect 16392 43150 18939 43152
rect 5574 43012 5580 43076
rect 5644 43074 5650 43076
rect 5993 43074 6059 43077
rect 5644 43072 6059 43074
rect 5644 43016 5998 43072
rect 6054 43016 6059 43072
rect 5644 43014 6059 43016
rect 5644 43012 5650 43014
rect 5993 43011 6059 43014
rect 14641 43074 14707 43077
rect 16392 43074 16452 43150
rect 18873 43147 18939 43150
rect 14641 43072 16452 43074
rect 14641 43016 14646 43072
rect 14702 43016 16452 43072
rect 14641 43014 16452 43016
rect 19977 43074 20043 43077
rect 21840 43074 22300 43104
rect 19977 43072 22300 43074
rect 19977 43016 19982 43072
rect 20038 43016 22300 43072
rect 19977 43014 22300 43016
rect 14641 43011 14707 43014
rect 19977 43011 20043 43014
rect 3418 43008 3734 43009
rect 3418 42944 3424 43008
rect 3488 42944 3504 43008
rect 3568 42944 3584 43008
rect 3648 42944 3664 43008
rect 3728 42944 3734 43008
rect 3418 42943 3734 42944
rect 8363 43008 8679 43009
rect 8363 42944 8369 43008
rect 8433 42944 8449 43008
rect 8513 42944 8529 43008
rect 8593 42944 8609 43008
rect 8673 42944 8679 43008
rect 8363 42943 8679 42944
rect 13308 43008 13624 43009
rect 13308 42944 13314 43008
rect 13378 42944 13394 43008
rect 13458 42944 13474 43008
rect 13538 42944 13554 43008
rect 13618 42944 13624 43008
rect 13308 42943 13624 42944
rect 18253 43008 18569 43009
rect 18253 42944 18259 43008
rect 18323 42944 18339 43008
rect 18403 42944 18419 43008
rect 18483 42944 18499 43008
rect 18563 42944 18569 43008
rect 21840 42984 22300 43014
rect 18253 42943 18569 42944
rect 10542 42876 10548 42940
rect 10612 42938 10618 42940
rect 10777 42938 10843 42941
rect 10612 42936 10843 42938
rect 10612 42880 10782 42936
rect 10838 42880 10843 42936
rect 10612 42878 10843 42880
rect 10612 42876 10618 42878
rect 10777 42875 10843 42878
rect 14181 42938 14247 42941
rect 14181 42936 16866 42938
rect 14181 42880 14186 42936
rect 14242 42880 16866 42936
rect 14181 42878 16866 42880
rect 14181 42875 14247 42878
rect 13997 42802 14063 42805
rect 16573 42802 16639 42805
rect 13997 42800 16639 42802
rect 13997 42744 14002 42800
rect 14058 42744 16578 42800
rect 16634 42744 16639 42800
rect 13997 42742 16639 42744
rect 16806 42802 16866 42878
rect 19057 42802 19123 42805
rect 16806 42800 19123 42802
rect 16806 42744 19062 42800
rect 19118 42744 19123 42800
rect 16806 42742 19123 42744
rect 13997 42739 14063 42742
rect 16573 42739 16639 42742
rect 19057 42739 19123 42742
rect 10133 42666 10199 42669
rect 11697 42666 11763 42669
rect 10133 42664 11763 42666
rect 10133 42608 10138 42664
rect 10194 42608 11702 42664
rect 11758 42608 11763 42664
rect 10133 42606 11763 42608
rect 10133 42603 10199 42606
rect 11697 42603 11763 42606
rect 15510 42604 15516 42668
rect 15580 42666 15586 42668
rect 16205 42666 16271 42669
rect 15580 42664 16271 42666
rect 15580 42608 16210 42664
rect 16266 42608 16271 42664
rect 15580 42606 16271 42608
rect 15580 42604 15586 42606
rect 16205 42603 16271 42606
rect 17769 42666 17835 42669
rect 18321 42666 18387 42669
rect 17769 42664 18387 42666
rect 17769 42608 17774 42664
rect 17830 42608 18326 42664
rect 18382 42608 18387 42664
rect 17769 42606 18387 42608
rect 17769 42603 17835 42606
rect 18321 42603 18387 42606
rect 9627 42562 9693 42567
rect 8845 42530 8911 42533
rect 9121 42530 9187 42533
rect 8845 42528 9187 42530
rect 8845 42472 8850 42528
rect 8906 42472 9126 42528
rect 9182 42472 9187 42528
rect 9627 42506 9632 42562
rect 9688 42506 9693 42562
rect 9627 42501 9693 42506
rect 21265 42530 21331 42533
rect 21840 42530 22300 42560
rect 21265 42528 22300 42530
rect 8845 42470 9187 42472
rect 8845 42467 8911 42470
rect 9121 42467 9187 42470
rect 5890 42464 6206 42465
rect 5890 42400 5896 42464
rect 5960 42400 5976 42464
rect 6040 42400 6056 42464
rect 6120 42400 6136 42464
rect 6200 42400 6206 42464
rect 5890 42399 6206 42400
rect 9630 42394 9690 42501
rect 21265 42472 21270 42528
rect 21326 42472 22300 42528
rect 21265 42470 22300 42472
rect 21265 42467 21331 42470
rect 10835 42464 11151 42465
rect 10835 42400 10841 42464
rect 10905 42400 10921 42464
rect 10985 42400 11001 42464
rect 11065 42400 11081 42464
rect 11145 42400 11151 42464
rect 10835 42399 11151 42400
rect 15780 42464 16096 42465
rect 15780 42400 15786 42464
rect 15850 42400 15866 42464
rect 15930 42400 15946 42464
rect 16010 42400 16026 42464
rect 16090 42400 16096 42464
rect 15780 42399 16096 42400
rect 20725 42464 21041 42465
rect 20725 42400 20731 42464
rect 20795 42400 20811 42464
rect 20875 42400 20891 42464
rect 20955 42400 20971 42464
rect 21035 42400 21041 42464
rect 21840 42440 22300 42470
rect 20725 42399 21041 42400
rect 14365 42394 14431 42397
rect 6272 42334 9690 42394
rect 11286 42392 14431 42394
rect 11286 42336 14370 42392
rect 14426 42336 14431 42392
rect 11286 42334 14431 42336
rect 4613 42258 4679 42261
rect 6272 42258 6332 42334
rect 4613 42256 6332 42258
rect 4613 42200 4618 42256
rect 4674 42200 6332 42256
rect 4613 42198 6332 42200
rect 4613 42195 4679 42198
rect 7414 42196 7420 42260
rect 7484 42258 7490 42260
rect 11286 42258 11346 42334
rect 14365 42331 14431 42334
rect 14825 42394 14891 42397
rect 15561 42394 15627 42397
rect 14825 42392 15627 42394
rect 14825 42336 14830 42392
rect 14886 42336 15566 42392
rect 15622 42336 15627 42392
rect 14825 42334 15627 42336
rect 14825 42331 14891 42334
rect 15561 42331 15627 42334
rect 7484 42198 11346 42258
rect 12157 42258 12223 42261
rect 16389 42258 16455 42261
rect 12157 42256 16455 42258
rect 12157 42200 12162 42256
rect 12218 42200 16394 42256
rect 16450 42200 16455 42256
rect 12157 42198 16455 42200
rect 7484 42196 7490 42198
rect 12157 42195 12223 42198
rect 16389 42195 16455 42198
rect 5390 42060 5396 42124
rect 5460 42122 5466 42124
rect 8845 42122 8911 42125
rect 5460 42120 8911 42122
rect 5460 42064 8850 42120
rect 8906 42064 8911 42120
rect 5460 42062 8911 42064
rect 5460 42060 5466 42062
rect 8845 42059 8911 42062
rect 9438 42060 9444 42124
rect 9508 42122 9514 42124
rect 9949 42122 10015 42125
rect 9508 42120 10015 42122
rect 9508 42064 9954 42120
rect 10010 42064 10015 42120
rect 9508 42062 10015 42064
rect 9508 42060 9514 42062
rect 9949 42059 10015 42062
rect 12801 42122 12867 42125
rect 12934 42122 12940 42124
rect 12801 42120 12940 42122
rect 12801 42064 12806 42120
rect 12862 42064 12940 42120
rect 12801 42062 12940 42064
rect 12801 42059 12867 42062
rect 12934 42060 12940 42062
rect 13004 42060 13010 42124
rect 16297 42122 16363 42125
rect 17677 42122 17743 42125
rect 13172 42120 16363 42122
rect 13172 42064 16302 42120
rect 16358 42064 16363 42120
rect 13172 42062 16363 42064
rect 12341 41986 12407 41989
rect 13172 41986 13232 42062
rect 16297 42059 16363 42062
rect 16438 42120 17743 42122
rect 16438 42064 17682 42120
rect 17738 42064 17743 42120
rect 16438 42062 17743 42064
rect 12341 41984 13232 41986
rect 12341 41928 12346 41984
rect 12402 41928 13232 41984
rect 12341 41926 13232 41928
rect 14457 41986 14523 41989
rect 16438 41986 16498 42062
rect 17677 42059 17743 42062
rect 18086 42060 18092 42124
rect 18156 42122 18162 42124
rect 18229 42122 18295 42125
rect 18156 42120 18295 42122
rect 18156 42064 18234 42120
rect 18290 42064 18295 42120
rect 18156 42062 18295 42064
rect 18156 42060 18162 42062
rect 18229 42059 18295 42062
rect 14457 41984 16498 41986
rect 14457 41928 14462 41984
rect 14518 41928 16498 41984
rect 14457 41926 16498 41928
rect 19333 41986 19399 41989
rect 21840 41986 22300 42016
rect 19333 41984 22300 41986
rect 19333 41928 19338 41984
rect 19394 41928 22300 41984
rect 19333 41926 22300 41928
rect 12341 41923 12407 41926
rect 14457 41923 14523 41926
rect 19333 41923 19399 41926
rect 3418 41920 3734 41921
rect 3418 41856 3424 41920
rect 3488 41856 3504 41920
rect 3568 41856 3584 41920
rect 3648 41856 3664 41920
rect 3728 41856 3734 41920
rect 3418 41855 3734 41856
rect 8363 41920 8679 41921
rect 8363 41856 8369 41920
rect 8433 41856 8449 41920
rect 8513 41856 8529 41920
rect 8593 41856 8609 41920
rect 8673 41856 8679 41920
rect 8363 41855 8679 41856
rect 13308 41920 13624 41921
rect 13308 41856 13314 41920
rect 13378 41856 13394 41920
rect 13458 41856 13474 41920
rect 13538 41856 13554 41920
rect 13618 41856 13624 41920
rect 13308 41855 13624 41856
rect 18253 41920 18569 41921
rect 18253 41856 18259 41920
rect 18323 41856 18339 41920
rect 18403 41856 18419 41920
rect 18483 41856 18499 41920
rect 18563 41856 18569 41920
rect 21840 41896 22300 41926
rect 18253 41855 18569 41856
rect 4705 41850 4771 41853
rect 5441 41850 5507 41853
rect 4705 41848 5507 41850
rect 4705 41792 4710 41848
rect 4766 41792 5446 41848
rect 5502 41792 5507 41848
rect 4705 41790 5507 41792
rect 4705 41787 4771 41790
rect 5441 41787 5507 41790
rect 15326 41788 15332 41852
rect 15396 41850 15402 41852
rect 15469 41850 15535 41853
rect 15396 41848 15535 41850
rect 15396 41792 15474 41848
rect 15530 41792 15535 41848
rect 15396 41790 15535 41792
rect 15396 41788 15402 41790
rect 15469 41787 15535 41790
rect 15745 41850 15811 41853
rect 17953 41850 18019 41853
rect 15745 41848 18019 41850
rect 15745 41792 15750 41848
rect 15806 41792 17958 41848
rect 18014 41792 18019 41848
rect 15745 41790 18019 41792
rect 15745 41787 15811 41790
rect 17953 41787 18019 41790
rect 1158 41652 1164 41716
rect 1228 41714 1234 41716
rect 5533 41714 5599 41717
rect 1228 41712 5599 41714
rect 1228 41656 5538 41712
rect 5594 41656 5599 41712
rect 1228 41654 5599 41656
rect 1228 41652 1234 41654
rect 5533 41651 5599 41654
rect 6494 41652 6500 41716
rect 6564 41714 6570 41716
rect 9765 41714 9831 41717
rect 13169 41716 13235 41717
rect 13118 41714 13124 41716
rect 6564 41712 9831 41714
rect 6564 41656 9770 41712
rect 9826 41656 9831 41712
rect 6564 41654 9831 41656
rect 13078 41654 13124 41714
rect 13188 41712 13235 41716
rect 13230 41656 13235 41712
rect 6564 41652 6570 41654
rect 9765 41651 9831 41654
rect 13118 41652 13124 41654
rect 13188 41652 13235 41656
rect 13169 41651 13235 41652
rect 14181 41714 14247 41717
rect 17401 41714 17467 41717
rect 14181 41712 17467 41714
rect 14181 41656 14186 41712
rect 14242 41656 17406 41712
rect 17462 41656 17467 41712
rect 14181 41654 17467 41656
rect 14181 41651 14247 41654
rect 17401 41651 17467 41654
rect 197 41578 263 41581
rect 3049 41578 3115 41581
rect 3918 41578 3924 41580
rect 197 41576 2790 41578
rect 197 41520 202 41576
rect 258 41520 2790 41576
rect 197 41518 2790 41520
rect 197 41515 263 41518
rect 1945 41442 2011 41445
rect 2078 41442 2084 41444
rect 1945 41440 2084 41442
rect 1945 41384 1950 41440
rect 2006 41384 2084 41440
rect 1945 41382 2084 41384
rect 1945 41379 2011 41382
rect 2078 41380 2084 41382
rect 2148 41380 2154 41444
rect 2730 41442 2790 41518
rect 3049 41576 3924 41578
rect 3049 41520 3054 41576
rect 3110 41520 3924 41576
rect 3049 41518 3924 41520
rect 3049 41515 3115 41518
rect 3918 41516 3924 41518
rect 3988 41516 3994 41580
rect 5441 41578 5507 41581
rect 4110 41576 5507 41578
rect 4110 41520 5446 41576
rect 5502 41520 5507 41576
rect 4110 41518 5507 41520
rect 4110 41442 4170 41518
rect 5441 41515 5507 41518
rect 6361 41578 6427 41581
rect 7465 41578 7531 41581
rect 6361 41576 7531 41578
rect 6361 41520 6366 41576
rect 6422 41520 7470 41576
rect 7526 41520 7531 41576
rect 6361 41518 7531 41520
rect 6361 41515 6427 41518
rect 7465 41515 7531 41518
rect 9121 41578 9187 41581
rect 9254 41578 9260 41580
rect 9121 41576 9260 41578
rect 9121 41520 9126 41576
rect 9182 41520 9260 41576
rect 9121 41518 9260 41520
rect 9121 41515 9187 41518
rect 9254 41516 9260 41518
rect 9324 41516 9330 41580
rect 11646 41516 11652 41580
rect 11716 41578 11722 41580
rect 14825 41578 14891 41581
rect 11716 41576 14891 41578
rect 11716 41520 14830 41576
rect 14886 41520 14891 41576
rect 11716 41518 14891 41520
rect 11716 41516 11722 41518
rect 14825 41515 14891 41518
rect 16021 41578 16087 41581
rect 16021 41576 16268 41578
rect 16021 41520 16026 41576
rect 16082 41520 16268 41576
rect 16021 41518 16268 41520
rect 16021 41515 16087 41518
rect 2730 41382 4170 41442
rect 15193 41442 15259 41445
rect 15510 41442 15516 41444
rect 15193 41440 15516 41442
rect 15193 41384 15198 41440
rect 15254 41384 15516 41440
rect 15193 41382 15516 41384
rect 15193 41379 15259 41382
rect 15510 41380 15516 41382
rect 15580 41380 15586 41444
rect 16208 41442 16268 41518
rect 19793 41442 19859 41445
rect 16208 41440 19859 41442
rect 16208 41384 19798 41440
rect 19854 41384 19859 41440
rect 16208 41382 19859 41384
rect 19793 41379 19859 41382
rect 21265 41442 21331 41445
rect 21840 41442 22300 41472
rect 21265 41440 22300 41442
rect 21265 41384 21270 41440
rect 21326 41384 22300 41440
rect 21265 41382 22300 41384
rect 21265 41379 21331 41382
rect 5890 41376 6206 41377
rect 5890 41312 5896 41376
rect 5960 41312 5976 41376
rect 6040 41312 6056 41376
rect 6120 41312 6136 41376
rect 6200 41312 6206 41376
rect 5890 41311 6206 41312
rect 10835 41376 11151 41377
rect 10835 41312 10841 41376
rect 10905 41312 10921 41376
rect 10985 41312 11001 41376
rect 11065 41312 11081 41376
rect 11145 41312 11151 41376
rect 10835 41311 11151 41312
rect 15780 41376 16096 41377
rect 15780 41312 15786 41376
rect 15850 41312 15866 41376
rect 15930 41312 15946 41376
rect 16010 41312 16026 41376
rect 16090 41312 16096 41376
rect 15780 41311 16096 41312
rect 20725 41376 21041 41377
rect 20725 41312 20731 41376
rect 20795 41312 20811 41376
rect 20875 41312 20891 41376
rect 20955 41312 20971 41376
rect 21035 41312 21041 41376
rect 21840 41352 22300 41382
rect 20725 41311 21041 41312
rect 16430 41244 16436 41308
rect 16500 41306 16506 41308
rect 16573 41306 16639 41309
rect 16500 41304 16639 41306
rect 16500 41248 16578 41304
rect 16634 41248 16639 41304
rect 16500 41246 16639 41248
rect 16500 41244 16506 41246
rect 16573 41243 16639 41246
rect 14549 41172 14615 41173
rect 14549 41168 14596 41172
rect 14660 41170 14666 41172
rect 14825 41170 14891 41173
rect 14958 41170 14964 41172
rect 14549 41112 14554 41168
rect 14549 41108 14596 41112
rect 14660 41110 14706 41170
rect 14825 41168 14964 41170
rect 14825 41112 14830 41168
rect 14886 41112 14964 41168
rect 14825 41110 14964 41112
rect 14660 41108 14666 41110
rect 14549 41107 14615 41108
rect 14825 41107 14891 41110
rect 14958 41108 14964 41110
rect 15028 41108 15034 41172
rect 15193 41170 15259 41173
rect 17033 41170 17099 41173
rect 15193 41168 17099 41170
rect 15193 41112 15198 41168
rect 15254 41112 17038 41168
rect 17094 41112 17099 41168
rect 15193 41110 17099 41112
rect 15193 41107 15259 41110
rect 17033 41107 17099 41110
rect 18689 41170 18755 41173
rect 19701 41170 19767 41173
rect 18689 41168 19767 41170
rect 18689 41112 18694 41168
rect 18750 41112 19706 41168
rect 19762 41112 19767 41168
rect 18689 41110 19767 41112
rect 18689 41107 18755 41110
rect 19701 41107 19767 41110
rect 3182 40972 3188 41036
rect 3252 41034 3258 41036
rect 3601 41034 3667 41037
rect 3252 41032 3667 41034
rect 3252 40976 3606 41032
rect 3662 40976 3667 41032
rect 3252 40974 3667 40976
rect 3252 40972 3258 40974
rect 3601 40971 3667 40974
rect 12433 41034 12499 41037
rect 18873 41034 18939 41037
rect 12433 41032 18939 41034
rect 12433 40976 12438 41032
rect 12494 40976 18878 41032
rect 18934 40976 18939 41032
rect 12433 40974 18939 40976
rect 12433 40971 12499 40974
rect 18873 40971 18939 40974
rect 14917 40898 14983 40901
rect 18086 40898 18092 40900
rect 14917 40896 18092 40898
rect 14917 40840 14922 40896
rect 14978 40840 18092 40896
rect 14917 40838 18092 40840
rect 14917 40835 14983 40838
rect 18086 40836 18092 40838
rect 18156 40836 18162 40900
rect 20529 40898 20595 40901
rect 21840 40898 22300 40928
rect 20529 40896 22300 40898
rect 20529 40840 20534 40896
rect 20590 40840 22300 40896
rect 20529 40838 22300 40840
rect 20529 40835 20595 40838
rect 3418 40832 3734 40833
rect 3418 40768 3424 40832
rect 3488 40768 3504 40832
rect 3568 40768 3584 40832
rect 3648 40768 3664 40832
rect 3728 40768 3734 40832
rect 3418 40767 3734 40768
rect 8363 40832 8679 40833
rect 8363 40768 8369 40832
rect 8433 40768 8449 40832
rect 8513 40768 8529 40832
rect 8593 40768 8609 40832
rect 8673 40768 8679 40832
rect 8363 40767 8679 40768
rect 13308 40832 13624 40833
rect 13308 40768 13314 40832
rect 13378 40768 13394 40832
rect 13458 40768 13474 40832
rect 13538 40768 13554 40832
rect 13618 40768 13624 40832
rect 13308 40767 13624 40768
rect 18253 40832 18569 40833
rect 18253 40768 18259 40832
rect 18323 40768 18339 40832
rect 18403 40768 18419 40832
rect 18483 40768 18499 40832
rect 18563 40768 18569 40832
rect 21840 40808 22300 40838
rect 18253 40767 18569 40768
rect 16205 40762 16271 40765
rect 16614 40762 16620 40764
rect 16205 40760 16620 40762
rect 16205 40704 16210 40760
rect 16266 40704 16620 40760
rect 16205 40702 16620 40704
rect 16205 40699 16271 40702
rect 16614 40700 16620 40702
rect 16684 40700 16690 40764
rect 4889 40626 4955 40629
rect 7189 40626 7255 40629
rect 12198 40626 12204 40628
rect 4889 40624 12204 40626
rect 4889 40568 4894 40624
rect 4950 40568 7194 40624
rect 7250 40568 12204 40624
rect 4889 40566 12204 40568
rect 4889 40563 4955 40566
rect 7189 40563 7255 40566
rect 12198 40564 12204 40566
rect 12268 40626 12274 40628
rect 18321 40626 18387 40629
rect 12268 40624 18387 40626
rect 12268 40568 18326 40624
rect 18382 40568 18387 40624
rect 12268 40566 18387 40568
rect 12268 40564 12274 40566
rect 18321 40563 18387 40566
rect 1710 40428 1716 40492
rect 1780 40490 1786 40492
rect 2681 40490 2747 40493
rect 18229 40490 18295 40493
rect 1780 40488 18295 40490
rect 1780 40432 2686 40488
rect 2742 40432 18234 40488
rect 18290 40432 18295 40488
rect 1780 40430 18295 40432
rect 1780 40428 1786 40430
rect 2681 40427 2747 40430
rect 18229 40427 18295 40430
rect 15101 40354 15167 40357
rect 15326 40354 15332 40356
rect 15101 40352 15332 40354
rect 15101 40296 15106 40352
rect 15162 40296 15332 40352
rect 15101 40294 15332 40296
rect 15101 40291 15167 40294
rect 15326 40292 15332 40294
rect 15396 40292 15402 40356
rect 21265 40354 21331 40357
rect 21840 40354 22300 40384
rect 21265 40352 22300 40354
rect 21265 40296 21270 40352
rect 21326 40296 22300 40352
rect 21265 40294 22300 40296
rect 21265 40291 21331 40294
rect 5890 40288 6206 40289
rect 5890 40224 5896 40288
rect 5960 40224 5976 40288
rect 6040 40224 6056 40288
rect 6120 40224 6136 40288
rect 6200 40224 6206 40288
rect 5890 40223 6206 40224
rect 10835 40288 11151 40289
rect 10835 40224 10841 40288
rect 10905 40224 10921 40288
rect 10985 40224 11001 40288
rect 11065 40224 11081 40288
rect 11145 40224 11151 40288
rect 10835 40223 11151 40224
rect 15780 40288 16096 40289
rect 15780 40224 15786 40288
rect 15850 40224 15866 40288
rect 15930 40224 15946 40288
rect 16010 40224 16026 40288
rect 16090 40224 16096 40288
rect 15780 40223 16096 40224
rect 20725 40288 21041 40289
rect 20725 40224 20731 40288
rect 20795 40224 20811 40288
rect 20875 40224 20891 40288
rect 20955 40224 20971 40288
rect 21035 40224 21041 40288
rect 21840 40264 22300 40294
rect 20725 40223 21041 40224
rect 18413 40218 18479 40221
rect 16806 40216 18479 40218
rect 16806 40160 18418 40216
rect 18474 40160 18479 40216
rect 16806 40158 18479 40160
rect 7925 40084 7991 40085
rect 7925 40080 7972 40084
rect 8036 40082 8042 40084
rect 7925 40024 7930 40080
rect 7925 40020 7972 40024
rect 8036 40022 8082 40082
rect 8036 40020 8042 40022
rect 12750 40020 12756 40084
rect 12820 40082 12826 40084
rect 13537 40082 13603 40085
rect 16806 40082 16866 40158
rect 18413 40155 18479 40158
rect 12820 40080 16866 40082
rect 12820 40024 13542 40080
rect 13598 40024 16866 40080
rect 12820 40022 16866 40024
rect 16941 40084 17007 40085
rect 16941 40080 16988 40084
rect 17052 40082 17058 40084
rect 16941 40024 16946 40080
rect 12820 40020 12826 40022
rect 7925 40019 7991 40020
rect 13537 40019 13603 40022
rect 16941 40020 16988 40024
rect 17052 40022 17098 40082
rect 17052 40020 17058 40022
rect 17902 40020 17908 40084
rect 17972 40082 17978 40084
rect 18137 40082 18203 40085
rect 17972 40080 18203 40082
rect 17972 40024 18142 40080
rect 18198 40024 18203 40080
rect 17972 40022 18203 40024
rect 17972 40020 17978 40022
rect 16941 40019 17007 40020
rect 18137 40019 18203 40022
rect 18597 40084 18663 40085
rect 18597 40080 18644 40084
rect 18708 40082 18714 40084
rect 18597 40024 18602 40080
rect 18597 40020 18644 40024
rect 18708 40022 18754 40082
rect 18708 40020 18714 40022
rect 18597 40019 18663 40020
rect 19701 39946 19767 39949
rect 18094 39944 19767 39946
rect 18094 39888 19706 39944
rect 19762 39888 19767 39944
rect 18094 39886 19767 39888
rect 289 39810 355 39813
rect 2129 39810 2195 39813
rect 14457 39810 14523 39813
rect 17534 39810 17540 39812
rect 289 39808 2790 39810
rect 289 39752 294 39808
rect 350 39752 2134 39808
rect 2190 39752 2790 39808
rect 289 39750 2790 39752
rect 289 39747 355 39750
rect 2129 39747 2195 39750
rect 1393 39674 1459 39677
rect 246 39672 1459 39674
rect 246 39616 1398 39672
rect 1454 39616 1459 39672
rect 246 39614 1459 39616
rect -300 39538 160 39568
rect 246 39538 306 39614
rect 1393 39611 1459 39614
rect -300 39478 306 39538
rect 2730 39538 2790 39750
rect 14457 39808 17540 39810
rect 14457 39752 14462 39808
rect 14518 39752 17540 39808
rect 14457 39750 17540 39752
rect 14457 39747 14523 39750
rect 17534 39748 17540 39750
rect 17604 39748 17610 39812
rect 17677 39810 17743 39813
rect 18094 39810 18154 39886
rect 19701 39883 19767 39886
rect 17677 39808 18154 39810
rect 17677 39752 17682 39808
rect 17738 39752 18154 39808
rect 17677 39750 18154 39752
rect 20989 39810 21055 39813
rect 21840 39810 22300 39840
rect 20989 39808 22300 39810
rect 20989 39752 20994 39808
rect 21050 39752 22300 39808
rect 20989 39750 22300 39752
rect 17677 39747 17743 39750
rect 20989 39747 21055 39750
rect 3418 39744 3734 39745
rect 3418 39680 3424 39744
rect 3488 39680 3504 39744
rect 3568 39680 3584 39744
rect 3648 39680 3664 39744
rect 3728 39680 3734 39744
rect 3418 39679 3734 39680
rect 8363 39744 8679 39745
rect 8363 39680 8369 39744
rect 8433 39680 8449 39744
rect 8513 39680 8529 39744
rect 8593 39680 8609 39744
rect 8673 39680 8679 39744
rect 8363 39679 8679 39680
rect 13308 39744 13624 39745
rect 13308 39680 13314 39744
rect 13378 39680 13394 39744
rect 13458 39680 13474 39744
rect 13538 39680 13554 39744
rect 13618 39680 13624 39744
rect 13308 39679 13624 39680
rect 18253 39744 18569 39745
rect 18253 39680 18259 39744
rect 18323 39680 18339 39744
rect 18403 39680 18419 39744
rect 18483 39680 18499 39744
rect 18563 39680 18569 39744
rect 21840 39720 22300 39750
rect 18253 39679 18569 39680
rect 9857 39674 9923 39677
rect 9990 39674 9996 39676
rect 9857 39672 9996 39674
rect 9857 39616 9862 39672
rect 9918 39616 9996 39672
rect 9857 39614 9996 39616
rect 9857 39611 9923 39614
rect 9990 39612 9996 39614
rect 10060 39612 10066 39676
rect 18689 39674 18755 39677
rect 19057 39674 19123 39677
rect 18689 39672 19123 39674
rect 18689 39616 18694 39672
rect 18750 39616 19062 39672
rect 19118 39616 19123 39672
rect 18689 39614 19123 39616
rect 18689 39611 18755 39614
rect 19057 39611 19123 39614
rect 19701 39538 19767 39541
rect 2730 39536 19767 39538
rect 2730 39480 19706 39536
rect 19762 39480 19767 39536
rect 2730 39478 19767 39480
rect -300 39448 160 39478
rect 19701 39475 19767 39478
rect 1945 39400 2011 39405
rect 1945 39344 1950 39400
rect 2006 39344 2011 39400
rect 1945 39339 2011 39344
rect 4061 39402 4127 39405
rect 18321 39402 18387 39405
rect 4061 39400 18387 39402
rect 4061 39344 4066 39400
rect 4122 39344 18326 39400
rect 18382 39344 18387 39400
rect 4061 39342 18387 39344
rect 4061 39339 4127 39342
rect 18321 39339 18387 39342
rect 19241 39402 19307 39405
rect 21173 39402 21239 39405
rect 19241 39400 21239 39402
rect 19241 39344 19246 39400
rect 19302 39344 21178 39400
rect 21234 39344 21239 39400
rect 19241 39342 21239 39344
rect 19241 39339 19307 39342
rect 21173 39339 21239 39342
rect -300 39266 160 39296
rect 1301 39266 1367 39269
rect -300 39264 1367 39266
rect -300 39208 1306 39264
rect 1362 39208 1367 39264
rect -300 39206 1367 39208
rect -300 39176 160 39206
rect 1301 39203 1367 39206
rect -300 38994 160 39024
rect 1948 38994 2008 39339
rect 16205 39268 16271 39269
rect 16205 39264 16252 39268
rect 16316 39266 16322 39268
rect 16481 39266 16547 39269
rect 17953 39266 18019 39269
rect 18597 39268 18663 39269
rect 18597 39266 18644 39268
rect 16205 39208 16210 39264
rect 16205 39204 16252 39208
rect 16316 39206 16362 39266
rect 16481 39264 18019 39266
rect 16481 39208 16486 39264
rect 16542 39208 17958 39264
rect 18014 39208 18019 39264
rect 16481 39206 18019 39208
rect 18552 39264 18644 39266
rect 18552 39208 18602 39264
rect 18552 39206 18644 39208
rect 16316 39204 16322 39206
rect 16205 39203 16271 39204
rect 16481 39203 16547 39206
rect 17953 39203 18019 39206
rect 18597 39204 18644 39206
rect 18708 39204 18714 39268
rect 21265 39266 21331 39269
rect 21840 39266 22300 39296
rect 21265 39264 22300 39266
rect 21265 39208 21270 39264
rect 21326 39208 22300 39264
rect 21265 39206 22300 39208
rect 18597 39203 18663 39204
rect 21265 39203 21331 39206
rect 5890 39200 6206 39201
rect 5890 39136 5896 39200
rect 5960 39136 5976 39200
rect 6040 39136 6056 39200
rect 6120 39136 6136 39200
rect 6200 39136 6206 39200
rect 5890 39135 6206 39136
rect 10835 39200 11151 39201
rect 10835 39136 10841 39200
rect 10905 39136 10921 39200
rect 10985 39136 11001 39200
rect 11065 39136 11081 39200
rect 11145 39136 11151 39200
rect 10835 39135 11151 39136
rect 15780 39200 16096 39201
rect 15780 39136 15786 39200
rect 15850 39136 15866 39200
rect 15930 39136 15946 39200
rect 16010 39136 16026 39200
rect 16090 39136 16096 39200
rect 15780 39135 16096 39136
rect 20725 39200 21041 39201
rect 20725 39136 20731 39200
rect 20795 39136 20811 39200
rect 20875 39136 20891 39200
rect 20955 39136 20971 39200
rect 21035 39136 21041 39200
rect 21840 39176 22300 39206
rect 20725 39135 21041 39136
rect 4797 39130 4863 39133
rect 5022 39130 5028 39132
rect 4797 39128 5028 39130
rect 4797 39072 4802 39128
rect 4858 39072 5028 39128
rect 4797 39070 5028 39072
rect 4797 39067 4863 39070
rect 5022 39068 5028 39070
rect 5092 39068 5098 39132
rect 13077 39130 13143 39133
rect 13854 39130 13860 39132
rect 13077 39128 13860 39130
rect 13077 39072 13082 39128
rect 13138 39072 13860 39128
rect 13077 39070 13860 39072
rect 13077 39067 13143 39070
rect 13854 39068 13860 39070
rect 13924 39068 13930 39132
rect 17217 39130 17283 39133
rect 18321 39130 18387 39133
rect 17217 39128 18387 39130
rect 17217 39072 17222 39128
rect 17278 39072 18326 39128
rect 18382 39072 18387 39128
rect 17217 39070 18387 39072
rect 17217 39067 17283 39070
rect 18321 39067 18387 39070
rect -300 38934 2008 38994
rect 4245 38994 4311 38997
rect 7833 38994 7899 38997
rect 4245 38992 7899 38994
rect 4245 38936 4250 38992
rect 4306 38936 7838 38992
rect 7894 38936 7899 38992
rect 4245 38934 7899 38936
rect -300 38904 160 38934
rect 4245 38931 4311 38934
rect 7833 38931 7899 38934
rect 18045 38994 18111 38997
rect 18873 38994 18939 38997
rect 18045 38992 18939 38994
rect 18045 38936 18050 38992
rect 18106 38936 18878 38992
rect 18934 38936 18939 38992
rect 18045 38934 18939 38936
rect 18045 38931 18111 38934
rect 18873 38931 18939 38934
rect 974 38796 980 38860
rect 1044 38858 1050 38860
rect 4981 38858 5047 38861
rect 1044 38856 5047 38858
rect 1044 38800 4986 38856
rect 5042 38800 5047 38856
rect 1044 38798 5047 38800
rect 1044 38796 1050 38798
rect 4981 38795 5047 38798
rect 9397 38858 9463 38861
rect 9397 38856 15578 38858
rect 9397 38800 9402 38856
rect 9458 38800 15578 38856
rect 9397 38798 15578 38800
rect 9397 38795 9463 38798
rect -300 38722 160 38752
rect 2773 38722 2839 38725
rect -300 38720 2839 38722
rect -300 38664 2778 38720
rect 2834 38664 2839 38720
rect -300 38662 2839 38664
rect -300 38632 160 38662
rect 2773 38659 2839 38662
rect 3418 38656 3734 38657
rect 3418 38592 3424 38656
rect 3488 38592 3504 38656
rect 3568 38592 3584 38656
rect 3648 38592 3664 38656
rect 3728 38592 3734 38656
rect 3418 38591 3734 38592
rect 8363 38656 8679 38657
rect 8363 38592 8369 38656
rect 8433 38592 8449 38656
rect 8513 38592 8529 38656
rect 8593 38592 8609 38656
rect 8673 38592 8679 38656
rect 8363 38591 8679 38592
rect 13308 38656 13624 38657
rect 13308 38592 13314 38656
rect 13378 38592 13394 38656
rect 13458 38592 13474 38656
rect 13538 38592 13554 38656
rect 13618 38592 13624 38656
rect 13308 38591 13624 38592
rect -300 38450 160 38480
rect 3049 38450 3115 38453
rect -300 38448 3115 38450
rect -300 38392 3054 38448
rect 3110 38392 3115 38448
rect -300 38390 3115 38392
rect -300 38360 160 38390
rect 3049 38387 3115 38390
rect 4061 38450 4127 38453
rect 5257 38450 5323 38453
rect 4061 38448 5323 38450
rect 4061 38392 4066 38448
rect 4122 38392 5262 38448
rect 5318 38392 5323 38448
rect 4061 38390 5323 38392
rect 4061 38387 4127 38390
rect 5257 38387 5323 38390
rect 1209 38314 1275 38317
rect 798 38312 1275 38314
rect 798 38256 1214 38312
rect 1270 38256 1275 38312
rect 798 38254 1275 38256
rect -300 38178 160 38208
rect 798 38178 858 38254
rect 1209 38251 1275 38254
rect 10593 38314 10659 38317
rect 12433 38314 12499 38317
rect 10593 38312 12499 38314
rect 10593 38256 10598 38312
rect 10654 38256 12438 38312
rect 12494 38256 12499 38312
rect 10593 38254 12499 38256
rect 15518 38314 15578 38798
rect 17125 38724 17191 38725
rect 17125 38720 17172 38724
rect 17236 38722 17242 38724
rect 20437 38722 20503 38725
rect 21840 38722 22300 38752
rect 17125 38664 17130 38720
rect 17125 38660 17172 38664
rect 17236 38662 17282 38722
rect 20437 38720 22300 38722
rect 20437 38664 20442 38720
rect 20498 38664 22300 38720
rect 20437 38662 22300 38664
rect 17236 38660 17242 38662
rect 17125 38659 17191 38660
rect 20437 38659 20503 38662
rect 18253 38656 18569 38657
rect 18253 38592 18259 38656
rect 18323 38592 18339 38656
rect 18403 38592 18419 38656
rect 18483 38592 18499 38656
rect 18563 38592 18569 38656
rect 21840 38632 22300 38662
rect 18253 38591 18569 38592
rect 21449 38314 21515 38317
rect 15518 38312 21515 38314
rect 15518 38256 21454 38312
rect 21510 38256 21515 38312
rect 15518 38254 21515 38256
rect 10593 38251 10659 38254
rect 12433 38251 12499 38254
rect 21449 38251 21515 38254
rect -300 38118 858 38178
rect 9673 38178 9739 38181
rect 10501 38178 10567 38181
rect 9673 38176 10567 38178
rect 9673 38120 9678 38176
rect 9734 38120 10506 38176
rect 10562 38120 10567 38176
rect 9673 38118 10567 38120
rect -300 38088 160 38118
rect 9673 38115 9739 38118
rect 10501 38115 10567 38118
rect 12566 38116 12572 38180
rect 12636 38178 12642 38180
rect 12985 38178 13051 38181
rect 12636 38176 13051 38178
rect 12636 38120 12990 38176
rect 13046 38120 13051 38176
rect 12636 38118 13051 38120
rect 12636 38116 12642 38118
rect 12985 38115 13051 38118
rect 21265 38178 21331 38181
rect 21840 38178 22300 38208
rect 21265 38176 22300 38178
rect 21265 38120 21270 38176
rect 21326 38120 22300 38176
rect 21265 38118 22300 38120
rect 21265 38115 21331 38118
rect 5890 38112 6206 38113
rect 5890 38048 5896 38112
rect 5960 38048 5976 38112
rect 6040 38048 6056 38112
rect 6120 38048 6136 38112
rect 6200 38048 6206 38112
rect 5890 38047 6206 38048
rect 10835 38112 11151 38113
rect 10835 38048 10841 38112
rect 10905 38048 10921 38112
rect 10985 38048 11001 38112
rect 11065 38048 11081 38112
rect 11145 38048 11151 38112
rect 10835 38047 11151 38048
rect 15780 38112 16096 38113
rect 15780 38048 15786 38112
rect 15850 38048 15866 38112
rect 15930 38048 15946 38112
rect 16010 38048 16026 38112
rect 16090 38048 16096 38112
rect 15780 38047 16096 38048
rect 20725 38112 21041 38113
rect 20725 38048 20731 38112
rect 20795 38048 20811 38112
rect 20875 38048 20891 38112
rect 20955 38048 20971 38112
rect 21035 38048 21041 38112
rect 21840 38088 22300 38118
rect 20725 38047 21041 38048
rect 7373 38042 7439 38045
rect 15653 38042 15719 38045
rect 6318 38040 7439 38042
rect 6318 37984 7378 38040
rect 7434 37984 7439 38040
rect 6318 37982 7439 37984
rect -300 37906 160 37936
rect 1393 37906 1459 37909
rect -300 37904 1459 37906
rect -300 37848 1398 37904
rect 1454 37848 1459 37904
rect -300 37846 1459 37848
rect -300 37816 160 37846
rect 1393 37843 1459 37846
rect 2957 37906 3023 37909
rect 6318 37906 6378 37982
rect 7373 37979 7439 37982
rect 11240 38040 15719 38042
rect 11240 37984 15658 38040
rect 15714 37984 15719 38040
rect 11240 37982 15719 37984
rect 2957 37904 6378 37906
rect 2957 37848 2962 37904
rect 3018 37848 6378 37904
rect 2957 37846 6378 37848
rect 6453 37906 6519 37909
rect 8753 37906 8819 37909
rect 6453 37904 8819 37906
rect 6453 37848 6458 37904
rect 6514 37848 8758 37904
rect 8814 37848 8819 37904
rect 6453 37846 8819 37848
rect 2957 37843 3023 37846
rect 6453 37843 6519 37846
rect 8753 37843 8819 37846
rect 10041 37906 10107 37909
rect 11240 37906 11300 37982
rect 15653 37979 15719 37982
rect 18965 38042 19031 38045
rect 18965 38040 19074 38042
rect 18965 37984 18970 38040
rect 19026 37984 19074 38040
rect 18965 37979 19074 37984
rect 10041 37904 11300 37906
rect 10041 37848 10046 37904
rect 10102 37848 11300 37904
rect 10041 37846 11300 37848
rect 11513 37906 11579 37909
rect 12433 37906 12499 37909
rect 11513 37904 12499 37906
rect 11513 37848 11518 37904
rect 11574 37848 12438 37904
rect 12494 37848 12499 37904
rect 11513 37846 12499 37848
rect 10041 37843 10107 37846
rect 11513 37843 11579 37846
rect 12433 37843 12499 37846
rect 12709 37906 12775 37909
rect 19014 37908 19074 37979
rect 16430 37906 16436 37908
rect 12709 37904 16436 37906
rect 12709 37848 12714 37904
rect 12770 37848 16436 37904
rect 12709 37846 16436 37848
rect 12709 37843 12775 37846
rect 16430 37844 16436 37846
rect 16500 37844 16506 37908
rect 19006 37844 19012 37908
rect 19076 37844 19082 37908
rect 6361 37770 6427 37773
rect 14273 37770 14339 37773
rect 6361 37768 14339 37770
rect 6361 37712 6366 37768
rect 6422 37712 14278 37768
rect 14334 37712 14339 37768
rect 6361 37710 14339 37712
rect 6361 37707 6427 37710
rect 14273 37707 14339 37710
rect 15285 37770 15351 37773
rect 19149 37770 19215 37773
rect 15285 37768 19215 37770
rect 15285 37712 15290 37768
rect 15346 37712 19154 37768
rect 19210 37712 19215 37768
rect 15285 37710 19215 37712
rect 15285 37707 15351 37710
rect 19149 37707 19215 37710
rect -300 37634 160 37664
rect 1945 37634 2011 37637
rect -300 37632 2011 37634
rect -300 37576 1950 37632
rect 2006 37576 2011 37632
rect -300 37574 2011 37576
rect -300 37544 160 37574
rect 1945 37571 2011 37574
rect 20437 37634 20503 37637
rect 21840 37634 22300 37664
rect 20437 37632 22300 37634
rect 20437 37576 20442 37632
rect 20498 37576 22300 37632
rect 20437 37574 22300 37576
rect 20437 37571 20503 37574
rect 3418 37568 3734 37569
rect 3418 37504 3424 37568
rect 3488 37504 3504 37568
rect 3568 37504 3584 37568
rect 3648 37504 3664 37568
rect 3728 37504 3734 37568
rect 3418 37503 3734 37504
rect 8363 37568 8679 37569
rect 8363 37504 8369 37568
rect 8433 37504 8449 37568
rect 8513 37504 8529 37568
rect 8593 37504 8609 37568
rect 8673 37504 8679 37568
rect 8363 37503 8679 37504
rect 13308 37568 13624 37569
rect 13308 37504 13314 37568
rect 13378 37504 13394 37568
rect 13458 37504 13474 37568
rect 13538 37504 13554 37568
rect 13618 37504 13624 37568
rect 13308 37503 13624 37504
rect 18253 37568 18569 37569
rect 18253 37504 18259 37568
rect 18323 37504 18339 37568
rect 18403 37504 18419 37568
rect 18483 37504 18499 37568
rect 18563 37504 18569 37568
rect 21840 37544 22300 37574
rect 18253 37503 18569 37504
rect 16798 37436 16804 37500
rect 16868 37498 16874 37500
rect 17309 37498 17375 37501
rect 16868 37496 17375 37498
rect 16868 37440 17314 37496
rect 17370 37440 17375 37496
rect 16868 37438 17375 37440
rect 16868 37436 16874 37438
rect 17309 37435 17375 37438
rect -300 37362 160 37392
rect 1485 37362 1551 37365
rect 5533 37362 5599 37365
rect -300 37360 1551 37362
rect -300 37304 1490 37360
rect 1546 37304 1551 37360
rect -300 37302 1551 37304
rect -300 37272 160 37302
rect 1485 37299 1551 37302
rect 2730 37360 5599 37362
rect 2730 37304 5538 37360
rect 5594 37304 5599 37360
rect 2730 37302 5599 37304
rect 2405 37226 2471 37229
rect 2730 37226 2790 37302
rect 5533 37299 5599 37302
rect 6729 37362 6795 37365
rect 6862 37362 6868 37364
rect 6729 37360 6868 37362
rect 6729 37304 6734 37360
rect 6790 37304 6868 37360
rect 6729 37302 6868 37304
rect 6729 37299 6795 37302
rect 6862 37300 6868 37302
rect 6932 37362 6938 37364
rect 6932 37302 9690 37362
rect 6932 37300 6938 37302
rect 2405 37224 2790 37226
rect 2405 37168 2410 37224
rect 2466 37168 2790 37224
rect 2405 37166 2790 37168
rect 5257 37226 5323 37229
rect 9397 37226 9463 37229
rect 5257 37224 9463 37226
rect 5257 37168 5262 37224
rect 5318 37168 9402 37224
rect 9458 37168 9463 37224
rect 5257 37166 9463 37168
rect 9630 37226 9690 37302
rect 13118 37300 13124 37364
rect 13188 37362 13194 37364
rect 19926 37362 19932 37364
rect 13188 37302 19932 37362
rect 13188 37300 13194 37302
rect 19926 37300 19932 37302
rect 19996 37300 20002 37364
rect 18781 37226 18847 37229
rect 9630 37224 18847 37226
rect 9630 37168 18786 37224
rect 18842 37168 18847 37224
rect 9630 37166 18847 37168
rect 2405 37163 2471 37166
rect 5257 37163 5323 37166
rect 9397 37163 9463 37166
rect 18781 37163 18847 37166
rect 20253 37226 20319 37229
rect 20253 37224 21282 37226
rect 20253 37168 20258 37224
rect 20314 37168 21282 37224
rect 20253 37166 21282 37168
rect 20253 37163 20319 37166
rect -300 37090 160 37120
rect 1301 37090 1367 37093
rect -300 37088 1367 37090
rect -300 37032 1306 37088
rect 1362 37032 1367 37088
rect -300 37030 1367 37032
rect -300 37000 160 37030
rect 1301 37027 1367 37030
rect 12198 37028 12204 37092
rect 12268 37090 12274 37092
rect 13997 37090 14063 37093
rect 12268 37088 14063 37090
rect 12268 37032 14002 37088
rect 14058 37032 14063 37088
rect 12268 37030 14063 37032
rect 21222 37090 21282 37166
rect 21840 37090 22300 37120
rect 21222 37030 22300 37090
rect 12268 37028 12274 37030
rect 13997 37027 14063 37030
rect 5890 37024 6206 37025
rect 5890 36960 5896 37024
rect 5960 36960 5976 37024
rect 6040 36960 6056 37024
rect 6120 36960 6136 37024
rect 6200 36960 6206 37024
rect 5890 36959 6206 36960
rect 10835 37024 11151 37025
rect 10835 36960 10841 37024
rect 10905 36960 10921 37024
rect 10985 36960 11001 37024
rect 11065 36960 11081 37024
rect 11145 36960 11151 37024
rect 10835 36959 11151 36960
rect 15780 37024 16096 37025
rect 15780 36960 15786 37024
rect 15850 36960 15866 37024
rect 15930 36960 15946 37024
rect 16010 36960 16026 37024
rect 16090 36960 16096 37024
rect 15780 36959 16096 36960
rect 20725 37024 21041 37025
rect 20725 36960 20731 37024
rect 20795 36960 20811 37024
rect 20875 36960 20891 37024
rect 20955 36960 20971 37024
rect 21035 36960 21041 37024
rect 21840 37000 22300 37030
rect 20725 36959 21041 36960
rect 18086 36892 18092 36956
rect 18156 36954 18162 36956
rect 18413 36954 18479 36957
rect 18156 36952 18479 36954
rect 18156 36896 18418 36952
rect 18474 36896 18479 36952
rect 18156 36894 18479 36896
rect 18156 36892 18162 36894
rect 18413 36891 18479 36894
rect -300 36818 160 36848
rect 1209 36818 1275 36821
rect -300 36816 1275 36818
rect -300 36760 1214 36816
rect 1270 36760 1275 36816
rect -300 36758 1275 36760
rect -300 36728 160 36758
rect 1209 36755 1275 36758
rect 1669 36818 1735 36821
rect 4613 36818 4679 36821
rect 1669 36816 9690 36818
rect 1669 36760 1674 36816
rect 1730 36760 4618 36816
rect 4674 36760 9690 36816
rect 1669 36758 9690 36760
rect 1669 36755 1735 36758
rect 4613 36755 4679 36758
rect 1117 36682 1183 36685
rect 798 36680 1183 36682
rect 798 36624 1122 36680
rect 1178 36624 1183 36680
rect 798 36622 1183 36624
rect -300 36546 160 36576
rect 798 36546 858 36622
rect 1117 36619 1183 36622
rect 5390 36620 5396 36684
rect 5460 36682 5466 36684
rect 7281 36682 7347 36685
rect 5460 36680 7347 36682
rect 5460 36624 7286 36680
rect 7342 36624 7347 36680
rect 5460 36622 7347 36624
rect 9630 36682 9690 36758
rect 10542 36756 10548 36820
rect 10612 36818 10618 36820
rect 12433 36818 12499 36821
rect 10612 36816 12499 36818
rect 10612 36760 12438 36816
rect 12494 36760 12499 36816
rect 10612 36758 12499 36760
rect 10612 36756 10618 36758
rect 12433 36755 12499 36758
rect 17033 36818 17099 36821
rect 18965 36818 19031 36821
rect 17033 36816 19031 36818
rect 17033 36760 17038 36816
rect 17094 36760 18970 36816
rect 19026 36760 19031 36816
rect 17033 36758 19031 36760
rect 17033 36755 17099 36758
rect 18965 36755 19031 36758
rect 18137 36682 18203 36685
rect 9630 36680 18203 36682
rect 9630 36624 18142 36680
rect 18198 36624 18203 36680
rect 9630 36622 18203 36624
rect 5460 36620 5466 36622
rect 7281 36619 7347 36622
rect 18137 36619 18203 36622
rect 18321 36682 18387 36685
rect 21725 36682 21791 36685
rect 18321 36680 21791 36682
rect 18321 36624 18326 36680
rect 18382 36624 21730 36680
rect 21786 36624 21791 36680
rect 18321 36622 21791 36624
rect 18321 36619 18387 36622
rect 21725 36619 21791 36622
rect -300 36486 858 36546
rect 5717 36546 5783 36549
rect 8201 36546 8267 36549
rect 5717 36544 8267 36546
rect 5717 36488 5722 36544
rect 5778 36488 8206 36544
rect 8262 36488 8267 36544
rect 5717 36486 8267 36488
rect -300 36456 160 36486
rect 5717 36483 5783 36486
rect 8201 36483 8267 36486
rect 19793 36546 19859 36549
rect 21840 36546 22300 36576
rect 19793 36544 22300 36546
rect 19793 36488 19798 36544
rect 19854 36488 22300 36544
rect 19793 36486 22300 36488
rect 19793 36483 19859 36486
rect 3418 36480 3734 36481
rect 3418 36416 3424 36480
rect 3488 36416 3504 36480
rect 3568 36416 3584 36480
rect 3648 36416 3664 36480
rect 3728 36416 3734 36480
rect 3418 36415 3734 36416
rect 8363 36480 8679 36481
rect 8363 36416 8369 36480
rect 8433 36416 8449 36480
rect 8513 36416 8529 36480
rect 8593 36416 8609 36480
rect 8673 36416 8679 36480
rect 8363 36415 8679 36416
rect 13308 36480 13624 36481
rect 13308 36416 13314 36480
rect 13378 36416 13394 36480
rect 13458 36416 13474 36480
rect 13538 36416 13554 36480
rect 13618 36416 13624 36480
rect 13308 36415 13624 36416
rect 18253 36480 18569 36481
rect 18253 36416 18259 36480
rect 18323 36416 18339 36480
rect 18403 36416 18419 36480
rect 18483 36416 18499 36480
rect 18563 36416 18569 36480
rect 21840 36456 22300 36486
rect 18253 36415 18569 36416
rect 10409 36410 10475 36413
rect 18689 36412 18755 36413
rect 10409 36408 12312 36410
rect 10409 36352 10414 36408
rect 10470 36352 12312 36408
rect 10409 36350 12312 36352
rect 10409 36347 10475 36350
rect -300 36274 160 36304
rect 1301 36274 1367 36277
rect -300 36272 1367 36274
rect -300 36216 1306 36272
rect 1362 36216 1367 36272
rect -300 36214 1367 36216
rect -300 36184 160 36214
rect 1301 36211 1367 36214
rect 2313 36274 2379 36277
rect 8150 36274 8156 36276
rect 2313 36272 8156 36274
rect 2313 36216 2318 36272
rect 2374 36216 8156 36272
rect 2313 36214 8156 36216
rect 2313 36211 2379 36214
rect 8150 36212 8156 36214
rect 8220 36274 8226 36276
rect 9397 36274 9463 36277
rect 8220 36272 12082 36274
rect 8220 36216 9402 36272
rect 9458 36216 12082 36272
rect 8220 36214 12082 36216
rect 8220 36212 8226 36214
rect 9397 36211 9463 36214
rect 4521 36138 4587 36141
rect 4478 36136 4587 36138
rect 4478 36080 4526 36136
rect 4582 36080 4587 36136
rect 4478 36075 4587 36080
rect -300 36002 160 36032
rect 1209 36002 1275 36005
rect -300 36000 1275 36002
rect -300 35944 1214 36000
rect 1270 35944 1275 36000
rect -300 35942 1275 35944
rect -300 35912 160 35942
rect 1209 35939 1275 35942
rect 4153 36002 4219 36005
rect 4478 36004 4538 36075
rect 4470 36002 4476 36004
rect 4153 36000 4476 36002
rect 4153 35944 4158 36000
rect 4214 35944 4476 36000
rect 4153 35942 4476 35944
rect 4153 35939 4219 35942
rect 4470 35940 4476 35942
rect 4540 35940 4546 36004
rect 12022 36002 12082 36214
rect 12252 36138 12312 36350
rect 18638 36348 18644 36412
rect 18708 36410 18755 36412
rect 18708 36408 18800 36410
rect 18750 36352 18800 36408
rect 18708 36350 18800 36352
rect 18708 36348 18755 36350
rect 18689 36347 18755 36348
rect 12433 36274 12499 36277
rect 13537 36274 13603 36277
rect 12433 36272 13603 36274
rect 12433 36216 12438 36272
rect 12494 36216 13542 36272
rect 13598 36216 13603 36272
rect 12433 36214 13603 36216
rect 12433 36211 12499 36214
rect 13537 36211 13603 36214
rect 13721 36274 13787 36277
rect 19006 36274 19012 36276
rect 13721 36272 19012 36274
rect 13721 36216 13726 36272
rect 13782 36216 19012 36272
rect 13721 36214 19012 36216
rect 13721 36211 13787 36214
rect 19006 36212 19012 36214
rect 19076 36212 19082 36276
rect 18413 36138 18479 36141
rect 18822 36138 18828 36140
rect 12252 36136 18828 36138
rect 12252 36080 18418 36136
rect 18474 36080 18828 36136
rect 12252 36078 18828 36080
rect 18413 36075 18479 36078
rect 18822 36076 18828 36078
rect 18892 36076 18898 36140
rect 15561 36002 15627 36005
rect 12022 36000 15627 36002
rect 12022 35944 15566 36000
rect 15622 35944 15627 36000
rect 12022 35942 15627 35944
rect 15561 35939 15627 35942
rect 21265 36002 21331 36005
rect 21840 36002 22300 36032
rect 21265 36000 22300 36002
rect 21265 35944 21270 36000
rect 21326 35944 22300 36000
rect 21265 35942 22300 35944
rect 21265 35939 21331 35942
rect 5890 35936 6206 35937
rect 5890 35872 5896 35936
rect 5960 35872 5976 35936
rect 6040 35872 6056 35936
rect 6120 35872 6136 35936
rect 6200 35872 6206 35936
rect 5890 35871 6206 35872
rect 10835 35936 11151 35937
rect 10835 35872 10841 35936
rect 10905 35872 10921 35936
rect 10985 35872 11001 35936
rect 11065 35872 11081 35936
rect 11145 35872 11151 35936
rect 10835 35871 11151 35872
rect 15780 35936 16096 35937
rect 15780 35872 15786 35936
rect 15850 35872 15866 35936
rect 15930 35872 15946 35936
rect 16010 35872 16026 35936
rect 16090 35872 16096 35936
rect 15780 35871 16096 35872
rect 20725 35936 21041 35937
rect 20725 35872 20731 35936
rect 20795 35872 20811 35936
rect 20875 35872 20891 35936
rect 20955 35872 20971 35936
rect 21035 35872 21041 35936
rect 21840 35912 22300 35942
rect 20725 35871 21041 35872
rect 1393 35864 1459 35869
rect 1393 35808 1398 35864
rect 1454 35808 1459 35864
rect 1393 35803 1459 35808
rect 7741 35866 7807 35869
rect 9070 35866 9076 35868
rect 7741 35864 9076 35866
rect 7741 35808 7746 35864
rect 7802 35808 9076 35864
rect 7741 35806 9076 35808
rect 7741 35803 7807 35806
rect 9070 35804 9076 35806
rect 9140 35804 9146 35868
rect 9765 35866 9831 35869
rect 10317 35866 10383 35869
rect 9765 35864 10383 35866
rect 9765 35808 9770 35864
rect 9826 35808 10322 35864
rect 10378 35808 10383 35864
rect 9765 35806 10383 35808
rect 9765 35803 9831 35806
rect 10317 35803 10383 35806
rect 10501 35866 10567 35869
rect 12157 35866 12223 35869
rect 10501 35864 10610 35866
rect 10501 35808 10506 35864
rect 10562 35808 10610 35864
rect 10501 35803 10610 35808
rect 12157 35864 12450 35866
rect 12157 35808 12162 35864
rect 12218 35808 12450 35864
rect 12157 35806 12450 35808
rect 12157 35803 12223 35806
rect -300 35730 160 35760
rect 1209 35730 1275 35733
rect -300 35728 1275 35730
rect -300 35672 1214 35728
rect 1270 35672 1275 35728
rect -300 35670 1275 35672
rect -300 35640 160 35670
rect 1209 35667 1275 35670
rect -300 35458 160 35488
rect 1396 35458 1456 35803
rect 8886 35668 8892 35732
rect 8956 35730 8962 35732
rect 9489 35730 9555 35733
rect 8956 35728 9555 35730
rect 8956 35672 9494 35728
rect 9550 35672 9555 35728
rect 8956 35670 9555 35672
rect 10550 35730 10610 35803
rect 12157 35730 12223 35733
rect 10550 35728 12223 35730
rect 10550 35672 12162 35728
rect 12218 35672 12223 35728
rect 10550 35670 12223 35672
rect 12390 35730 12450 35806
rect 14406 35804 14412 35868
rect 14476 35866 14482 35868
rect 15101 35866 15167 35869
rect 14476 35864 15167 35866
rect 14476 35808 15106 35864
rect 15162 35808 15167 35864
rect 14476 35806 15167 35808
rect 14476 35804 14482 35806
rect 15101 35803 15167 35806
rect 17309 35866 17375 35869
rect 19190 35866 19196 35868
rect 17309 35864 19196 35866
rect 17309 35808 17314 35864
rect 17370 35808 19196 35864
rect 17309 35806 19196 35808
rect 17309 35803 17375 35806
rect 19190 35804 19196 35806
rect 19260 35804 19266 35868
rect 15377 35730 15443 35733
rect 12390 35728 15443 35730
rect 12390 35672 15382 35728
rect 15438 35672 15443 35728
rect 12390 35670 15443 35672
rect 8956 35668 8962 35670
rect 9489 35667 9555 35670
rect 12157 35667 12223 35670
rect 15377 35667 15443 35670
rect 15837 35730 15903 35733
rect 18781 35730 18847 35733
rect 15837 35728 18847 35730
rect 15837 35672 15842 35728
rect 15898 35672 18786 35728
rect 18842 35672 18847 35728
rect 15837 35670 18847 35672
rect 15837 35667 15903 35670
rect 18781 35667 18847 35670
rect 4061 35594 4127 35597
rect 11462 35594 11468 35596
rect 4061 35592 11468 35594
rect 4061 35536 4066 35592
rect 4122 35536 11468 35592
rect 4061 35534 11468 35536
rect 4061 35531 4127 35534
rect 11462 35532 11468 35534
rect 11532 35532 11538 35596
rect -300 35398 1456 35458
rect 20345 35458 20411 35461
rect 21840 35458 22300 35488
rect 20345 35456 22300 35458
rect 20345 35400 20350 35456
rect 20406 35400 22300 35456
rect 20345 35398 22300 35400
rect -300 35368 160 35398
rect 20345 35395 20411 35398
rect 3418 35392 3734 35393
rect 3418 35328 3424 35392
rect 3488 35328 3504 35392
rect 3568 35328 3584 35392
rect 3648 35328 3664 35392
rect 3728 35328 3734 35392
rect 3418 35327 3734 35328
rect 8363 35392 8679 35393
rect 8363 35328 8369 35392
rect 8433 35328 8449 35392
rect 8513 35328 8529 35392
rect 8593 35328 8609 35392
rect 8673 35328 8679 35392
rect 8363 35327 8679 35328
rect 13308 35392 13624 35393
rect 13308 35328 13314 35392
rect 13378 35328 13394 35392
rect 13458 35328 13474 35392
rect 13538 35328 13554 35392
rect 13618 35328 13624 35392
rect 13308 35327 13624 35328
rect 18253 35392 18569 35393
rect 18253 35328 18259 35392
rect 18323 35328 18339 35392
rect 18403 35328 18419 35392
rect 18483 35328 18499 35392
rect 18563 35328 18569 35392
rect 21840 35368 22300 35398
rect 18253 35327 18569 35328
rect 790 35260 796 35324
rect 860 35322 866 35324
rect 2405 35322 2471 35325
rect 860 35320 2471 35322
rect 860 35264 2410 35320
rect 2466 35264 2471 35320
rect 860 35262 2471 35264
rect 860 35260 866 35262
rect 2405 35259 2471 35262
rect 9949 35322 10015 35325
rect 11278 35322 11284 35324
rect 9949 35320 11284 35322
rect 9949 35264 9954 35320
rect 10010 35264 11284 35320
rect 9949 35262 11284 35264
rect 9949 35259 10015 35262
rect 11278 35260 11284 35262
rect 11348 35260 11354 35324
rect 14038 35260 14044 35324
rect 14108 35322 14114 35324
rect 16941 35322 17007 35325
rect 14108 35320 17007 35322
rect 14108 35264 16946 35320
rect 17002 35264 17007 35320
rect 14108 35262 17007 35264
rect 14108 35260 14114 35262
rect 16941 35259 17007 35262
rect 19241 35320 19307 35325
rect 19241 35264 19246 35320
rect 19302 35264 19307 35320
rect 19241 35259 19307 35264
rect -300 35186 160 35216
rect 4245 35186 4311 35189
rect -300 35184 4311 35186
rect -300 35128 4250 35184
rect 4306 35128 4311 35184
rect -300 35126 4311 35128
rect -300 35096 160 35126
rect 4245 35123 4311 35126
rect 5901 35186 5967 35189
rect 7782 35186 7788 35188
rect 5901 35184 7788 35186
rect 5901 35128 5906 35184
rect 5962 35128 7788 35184
rect 5901 35126 7788 35128
rect 5901 35123 5967 35126
rect 7782 35124 7788 35126
rect 7852 35186 7858 35188
rect 10501 35186 10567 35189
rect 7852 35184 10567 35186
rect 7852 35128 10506 35184
rect 10562 35128 10567 35184
rect 7852 35126 10567 35128
rect 7852 35124 7858 35126
rect 10501 35123 10567 35126
rect 14549 35188 14615 35189
rect 14549 35184 14596 35188
rect 14660 35186 14666 35188
rect 15653 35186 15719 35189
rect 19244 35186 19304 35259
rect 14549 35128 14554 35184
rect 14549 35124 14596 35128
rect 14660 35126 14706 35186
rect 15653 35184 19304 35186
rect 15653 35128 15658 35184
rect 15714 35128 19304 35184
rect 15653 35126 19304 35128
rect 14660 35124 14666 35126
rect 14549 35123 14615 35124
rect 15653 35123 15719 35126
rect 7281 35050 7347 35053
rect 9949 35050 10015 35053
rect 17309 35050 17375 35053
rect 7281 35048 7850 35050
rect 7281 34992 7286 35048
rect 7342 34992 7850 35048
rect 7281 34990 7850 34992
rect 7281 34987 7347 34990
rect -300 34914 160 34944
rect 1945 34914 2011 34917
rect -300 34912 2011 34914
rect -300 34856 1950 34912
rect 2006 34856 2011 34912
rect -300 34854 2011 34856
rect 7790 34914 7850 34990
rect 9949 35048 17375 35050
rect 9949 34992 9954 35048
rect 10010 34992 17314 35048
rect 17370 34992 17375 35048
rect 9949 34990 17375 34992
rect 9949 34987 10015 34990
rect 17309 34987 17375 34990
rect 12249 34914 12315 34917
rect 12525 34914 12591 34917
rect 7790 34854 10610 34914
rect -300 34824 160 34854
rect 1945 34851 2011 34854
rect 5890 34848 6206 34849
rect 5890 34784 5896 34848
rect 5960 34784 5976 34848
rect 6040 34784 6056 34848
rect 6120 34784 6136 34848
rect 6200 34784 6206 34848
rect 5890 34783 6206 34784
rect 1485 34778 1551 34781
rect 9029 34778 9095 34781
rect 798 34776 1551 34778
rect 798 34720 1490 34776
rect 1546 34720 1551 34776
rect 798 34718 1551 34720
rect -300 34642 160 34672
rect 798 34642 858 34718
rect 1485 34715 1551 34718
rect 8020 34776 9095 34778
rect 8020 34720 9034 34776
rect 9090 34720 9095 34776
rect 8020 34718 9095 34720
rect 8020 34645 8080 34718
rect 9029 34715 9095 34718
rect -300 34582 858 34642
rect 4889 34642 4955 34645
rect 8017 34642 8083 34645
rect 8201 34642 8267 34645
rect 4889 34640 8083 34642
rect 4889 34584 4894 34640
rect 4950 34584 8022 34640
rect 8078 34584 8083 34640
rect 4889 34582 8083 34584
rect -300 34552 160 34582
rect 4889 34579 4955 34582
rect 8017 34579 8083 34582
rect 8158 34640 8267 34642
rect 8158 34584 8206 34640
rect 8262 34584 8267 34640
rect 8158 34579 8267 34584
rect 10133 34644 10199 34645
rect 10133 34640 10180 34644
rect 10244 34642 10250 34644
rect 10133 34584 10138 34640
rect 10133 34580 10180 34584
rect 10244 34582 10290 34642
rect 10244 34580 10250 34582
rect 10133 34579 10199 34580
rect 3785 34506 3851 34509
rect 2730 34504 3851 34506
rect 2730 34448 3790 34504
rect 3846 34448 3851 34504
rect 2730 34446 3851 34448
rect -300 34370 160 34400
rect 2730 34370 2790 34446
rect 3785 34443 3851 34446
rect 5625 34506 5691 34509
rect 6494 34506 6500 34508
rect 5625 34504 6500 34506
rect 5625 34448 5630 34504
rect 5686 34448 6500 34504
rect 5625 34446 6500 34448
rect 5625 34443 5691 34446
rect 6494 34444 6500 34446
rect 6564 34444 6570 34508
rect 8158 34506 8218 34579
rect 10358 34506 10364 34508
rect 8158 34446 10364 34506
rect 10358 34444 10364 34446
rect 10428 34444 10434 34508
rect 10550 34506 10610 34854
rect 12249 34912 12591 34914
rect 12249 34856 12254 34912
rect 12310 34856 12530 34912
rect 12586 34856 12591 34912
rect 12249 34854 12591 34856
rect 12249 34851 12315 34854
rect 12525 34851 12591 34854
rect 21265 34914 21331 34917
rect 21840 34914 22300 34944
rect 21265 34912 22300 34914
rect 21265 34856 21270 34912
rect 21326 34856 22300 34912
rect 21265 34854 22300 34856
rect 21265 34851 21331 34854
rect 10835 34848 11151 34849
rect 10835 34784 10841 34848
rect 10905 34784 10921 34848
rect 10985 34784 11001 34848
rect 11065 34784 11081 34848
rect 11145 34784 11151 34848
rect 10835 34783 11151 34784
rect 15780 34848 16096 34849
rect 15780 34784 15786 34848
rect 15850 34784 15866 34848
rect 15930 34784 15946 34848
rect 16010 34784 16026 34848
rect 16090 34784 16096 34848
rect 15780 34783 16096 34784
rect 20725 34848 21041 34849
rect 20725 34784 20731 34848
rect 20795 34784 20811 34848
rect 20875 34784 20891 34848
rect 20955 34784 20971 34848
rect 21035 34784 21041 34848
rect 21840 34824 22300 34854
rect 20725 34783 21041 34784
rect 11646 34716 11652 34780
rect 11716 34778 11722 34780
rect 12801 34778 12867 34781
rect 11716 34776 12867 34778
rect 11716 34720 12806 34776
rect 12862 34720 12867 34776
rect 11716 34718 12867 34720
rect 11716 34716 11722 34718
rect 12801 34715 12867 34718
rect 14273 34778 14339 34781
rect 15469 34780 15535 34781
rect 15142 34778 15148 34780
rect 14273 34776 15148 34778
rect 14273 34720 14278 34776
rect 14334 34720 15148 34776
rect 14273 34718 15148 34720
rect 14273 34715 14339 34718
rect 15142 34716 15148 34718
rect 15212 34716 15218 34780
rect 15469 34778 15516 34780
rect 15424 34776 15516 34778
rect 15424 34720 15474 34776
rect 15424 34718 15516 34720
rect 15469 34716 15516 34718
rect 15580 34716 15586 34780
rect 15469 34715 15535 34716
rect 11605 34644 11671 34645
rect 11605 34642 11652 34644
rect 11560 34640 11652 34642
rect 11560 34584 11610 34640
rect 11560 34582 11652 34584
rect 11605 34580 11652 34582
rect 11716 34580 11722 34644
rect 11789 34642 11855 34645
rect 12014 34642 12020 34644
rect 11789 34640 12020 34642
rect 11789 34584 11794 34640
rect 11850 34584 12020 34640
rect 11789 34582 12020 34584
rect 11605 34579 11671 34580
rect 11789 34579 11855 34582
rect 12014 34580 12020 34582
rect 12084 34580 12090 34644
rect 15377 34642 15443 34645
rect 16389 34642 16455 34645
rect 15377 34640 16455 34642
rect 15377 34584 15382 34640
rect 15438 34584 16394 34640
rect 16450 34584 16455 34640
rect 15377 34582 16455 34584
rect 15377 34579 15443 34582
rect 16389 34579 16455 34582
rect 12198 34506 12204 34508
rect 10550 34446 12204 34506
rect 12198 34444 12204 34446
rect 12268 34444 12274 34508
rect 14365 34506 14431 34509
rect 18965 34506 19031 34509
rect 14365 34504 19031 34506
rect 14365 34448 14370 34504
rect 14426 34448 18970 34504
rect 19026 34448 19031 34504
rect 14365 34446 19031 34448
rect 14365 34443 14431 34446
rect 18965 34443 19031 34446
rect -300 34310 2790 34370
rect -300 34280 160 34310
rect 4838 34308 4844 34372
rect 4908 34370 4914 34372
rect 7414 34370 7420 34372
rect 4908 34310 7420 34370
rect 4908 34308 4914 34310
rect 7414 34308 7420 34310
rect 7484 34308 7490 34372
rect 20437 34370 20503 34373
rect 21840 34370 22300 34400
rect 20437 34368 22300 34370
rect 20437 34312 20442 34368
rect 20498 34312 22300 34368
rect 20437 34310 22300 34312
rect 20437 34307 20503 34310
rect 3418 34304 3734 34305
rect 3418 34240 3424 34304
rect 3488 34240 3504 34304
rect 3568 34240 3584 34304
rect 3648 34240 3664 34304
rect 3728 34240 3734 34304
rect 3418 34239 3734 34240
rect 8363 34304 8679 34305
rect 8363 34240 8369 34304
rect 8433 34240 8449 34304
rect 8513 34240 8529 34304
rect 8593 34240 8609 34304
rect 8673 34240 8679 34304
rect 8363 34239 8679 34240
rect 13308 34304 13624 34305
rect 13308 34240 13314 34304
rect 13378 34240 13394 34304
rect 13458 34240 13474 34304
rect 13538 34240 13554 34304
rect 13618 34240 13624 34304
rect 13308 34239 13624 34240
rect 18253 34304 18569 34305
rect 18253 34240 18259 34304
rect 18323 34240 18339 34304
rect 18403 34240 18419 34304
rect 18483 34240 18499 34304
rect 18563 34240 18569 34304
rect 21840 34280 22300 34310
rect 18253 34239 18569 34240
rect 4102 34172 4108 34236
rect 4172 34234 4178 34236
rect 6545 34234 6611 34237
rect 4172 34232 6611 34234
rect 4172 34176 6550 34232
rect 6606 34176 6611 34232
rect 4172 34174 6611 34176
rect 4172 34172 4178 34174
rect 6545 34171 6611 34174
rect 7097 34234 7163 34237
rect 7414 34234 7420 34236
rect 7097 34232 7420 34234
rect 7097 34176 7102 34232
rect 7158 34176 7420 34232
rect 7097 34174 7420 34176
rect 7097 34171 7163 34174
rect 7414 34172 7420 34174
rect 7484 34172 7490 34236
rect 7598 34172 7604 34236
rect 7668 34234 7674 34236
rect 7925 34234 7991 34237
rect 7668 34232 7991 34234
rect 7668 34176 7930 34232
rect 7986 34176 7991 34232
rect 7668 34174 7991 34176
rect 7668 34172 7674 34174
rect 7925 34171 7991 34174
rect 13721 34234 13787 34237
rect 14457 34234 14523 34237
rect 14733 34234 14799 34237
rect 13721 34232 14799 34234
rect 13721 34176 13726 34232
rect 13782 34176 14462 34232
rect 14518 34176 14738 34232
rect 14794 34176 14799 34232
rect 13721 34174 14799 34176
rect 13721 34171 13787 34174
rect 14457 34171 14523 34174
rect 14733 34171 14799 34174
rect 15193 34234 15259 34237
rect 17350 34234 17356 34236
rect 15193 34232 17356 34234
rect 15193 34176 15198 34232
rect 15254 34176 17356 34232
rect 15193 34174 17356 34176
rect 15193 34171 15259 34174
rect 17350 34172 17356 34174
rect 17420 34172 17426 34236
rect -300 34098 160 34128
rect 3325 34098 3391 34101
rect -300 34096 3391 34098
rect -300 34040 3330 34096
rect 3386 34040 3391 34096
rect -300 34038 3391 34040
rect -300 34008 160 34038
rect 3325 34035 3391 34038
rect 4061 34098 4127 34101
rect 18781 34098 18847 34101
rect 19425 34100 19491 34101
rect 19374 34098 19380 34100
rect 4061 34096 18847 34098
rect 4061 34040 4066 34096
rect 4122 34040 18786 34096
rect 18842 34040 18847 34096
rect 4061 34038 18847 34040
rect 19334 34038 19380 34098
rect 19444 34096 19491 34100
rect 19486 34040 19491 34096
rect 4061 34035 4127 34038
rect 18781 34035 18847 34038
rect 19374 34036 19380 34038
rect 19444 34036 19491 34040
rect 19425 34035 19491 34036
rect 2998 33900 3004 33964
rect 3068 33962 3074 33964
rect 4064 33962 4124 34035
rect 3068 33902 4124 33962
rect 5257 33962 5323 33965
rect 6494 33962 6500 33964
rect 5257 33960 6500 33962
rect 5257 33904 5262 33960
rect 5318 33904 6500 33960
rect 5257 33902 6500 33904
rect 3068 33900 3074 33902
rect 5257 33899 5323 33902
rect 6494 33900 6500 33902
rect 6564 33900 6570 33964
rect 8569 33962 8635 33965
rect 9305 33962 9371 33965
rect 8569 33960 9371 33962
rect 8569 33904 8574 33960
rect 8630 33904 9310 33960
rect 9366 33904 9371 33960
rect 8569 33902 9371 33904
rect 8569 33899 8635 33902
rect 9305 33899 9371 33902
rect 11053 33962 11119 33965
rect 16614 33962 16620 33964
rect 11053 33960 16620 33962
rect 11053 33904 11058 33960
rect 11114 33904 16620 33960
rect 11053 33902 16620 33904
rect 11053 33899 11119 33902
rect 16614 33900 16620 33902
rect 16684 33900 16690 33964
rect 18505 33962 18571 33965
rect 19701 33962 19767 33965
rect 18505 33960 19767 33962
rect 18505 33904 18510 33960
rect 18566 33904 19706 33960
rect 19762 33904 19767 33960
rect 18505 33902 19767 33904
rect 18505 33899 18571 33902
rect 19701 33899 19767 33902
rect -300 33826 160 33856
rect 2773 33826 2839 33829
rect -300 33824 2839 33826
rect -300 33768 2778 33824
rect 2834 33768 2839 33824
rect -300 33766 2839 33768
rect -300 33736 160 33766
rect 2773 33763 2839 33766
rect 6310 33764 6316 33828
rect 6380 33826 6386 33828
rect 6729 33826 6795 33829
rect 6380 33824 6795 33826
rect 6380 33768 6734 33824
rect 6790 33768 6795 33824
rect 6380 33766 6795 33768
rect 6380 33764 6386 33766
rect 6729 33763 6795 33766
rect 9029 33826 9095 33829
rect 9949 33826 10015 33829
rect 9029 33824 10015 33826
rect 9029 33768 9034 33824
rect 9090 33768 9954 33824
rect 10010 33768 10015 33824
rect 9029 33766 10015 33768
rect 9029 33763 9095 33766
rect 9949 33763 10015 33766
rect 13813 33826 13879 33829
rect 15009 33826 15075 33829
rect 13813 33824 15075 33826
rect 13813 33768 13818 33824
rect 13874 33768 15014 33824
rect 15070 33768 15075 33824
rect 13813 33766 15075 33768
rect 13813 33763 13879 33766
rect 15009 33763 15075 33766
rect 19517 33826 19583 33829
rect 19742 33826 19748 33828
rect 19517 33824 19748 33826
rect 19517 33768 19522 33824
rect 19578 33768 19748 33824
rect 19517 33766 19748 33768
rect 19517 33763 19583 33766
rect 19742 33764 19748 33766
rect 19812 33764 19818 33828
rect 21173 33826 21239 33829
rect 21840 33826 22300 33856
rect 21173 33824 22300 33826
rect 21173 33768 21178 33824
rect 21234 33768 22300 33824
rect 21173 33766 22300 33768
rect 21173 33763 21239 33766
rect 5890 33760 6206 33761
rect 5890 33696 5896 33760
rect 5960 33696 5976 33760
rect 6040 33696 6056 33760
rect 6120 33696 6136 33760
rect 6200 33696 6206 33760
rect 5890 33695 6206 33696
rect 10835 33760 11151 33761
rect 10835 33696 10841 33760
rect 10905 33696 10921 33760
rect 10985 33696 11001 33760
rect 11065 33696 11081 33760
rect 11145 33696 11151 33760
rect 10835 33695 11151 33696
rect 15780 33760 16096 33761
rect 15780 33696 15786 33760
rect 15850 33696 15866 33760
rect 15930 33696 15946 33760
rect 16010 33696 16026 33760
rect 16090 33696 16096 33760
rect 15780 33695 16096 33696
rect 20725 33760 21041 33761
rect 20725 33696 20731 33760
rect 20795 33696 20811 33760
rect 20875 33696 20891 33760
rect 20955 33696 20971 33760
rect 21035 33696 21041 33760
rect 21840 33736 22300 33766
rect 20725 33695 21041 33696
rect 13813 33690 13879 33693
rect 15653 33690 15719 33693
rect 13813 33688 15719 33690
rect 13813 33632 13818 33688
rect 13874 33632 15658 33688
rect 15714 33632 15719 33688
rect 13813 33630 15719 33632
rect 13813 33627 13879 33630
rect 15653 33627 15719 33630
rect -300 33554 160 33584
rect 1301 33554 1367 33557
rect -300 33552 1367 33554
rect -300 33496 1306 33552
rect 1362 33496 1367 33552
rect -300 33494 1367 33496
rect -300 33464 160 33494
rect 1301 33491 1367 33494
rect 3693 33554 3759 33557
rect 4470 33554 4476 33556
rect 3693 33552 4476 33554
rect 3693 33496 3698 33552
rect 3754 33496 4476 33552
rect 3693 33494 4476 33496
rect 3693 33491 3759 33494
rect 4470 33492 4476 33494
rect 4540 33492 4546 33556
rect 8845 33554 8911 33557
rect 18137 33554 18203 33557
rect 7054 33552 18203 33554
rect 7054 33496 8850 33552
rect 8906 33496 18142 33552
rect 18198 33496 18203 33552
rect 7054 33494 18203 33496
rect 422 33356 428 33420
rect 492 33418 498 33420
rect 4153 33418 4219 33421
rect 492 33416 4219 33418
rect 492 33360 4158 33416
rect 4214 33360 4219 33416
rect 492 33358 4219 33360
rect 492 33356 498 33358
rect 4153 33355 4219 33358
rect 4286 33356 4292 33420
rect 4356 33418 4362 33420
rect 4429 33418 4495 33421
rect 4356 33416 4495 33418
rect 4356 33360 4434 33416
rect 4490 33360 4495 33416
rect 4356 33358 4495 33360
rect 4356 33356 4362 33358
rect 4429 33355 4495 33358
rect -300 33282 160 33312
rect 1945 33282 2011 33285
rect -300 33280 2011 33282
rect -300 33224 1950 33280
rect 2006 33224 2011 33280
rect -300 33222 2011 33224
rect -300 33192 160 33222
rect 1945 33219 2011 33222
rect 3418 33216 3734 33217
rect 3418 33152 3424 33216
rect 3488 33152 3504 33216
rect 3568 33152 3584 33216
rect 3648 33152 3664 33216
rect 3728 33152 3734 33216
rect 3418 33151 3734 33152
rect 1209 33146 1275 33149
rect 798 33144 1275 33146
rect 798 33088 1214 33144
rect 1270 33088 1275 33144
rect 798 33086 1275 33088
rect -300 33010 160 33040
rect 798 33010 858 33086
rect 1209 33083 1275 33086
rect 4245 33146 4311 33149
rect 7054 33146 7114 33494
rect 8845 33491 8911 33494
rect 18137 33491 18203 33494
rect 18689 33554 18755 33557
rect 19057 33554 19123 33557
rect 18689 33552 19123 33554
rect 18689 33496 18694 33552
rect 18750 33496 19062 33552
rect 19118 33496 19123 33552
rect 18689 33494 19123 33496
rect 18689 33491 18755 33494
rect 19057 33491 19123 33494
rect 17125 33418 17191 33421
rect 20253 33418 20319 33421
rect 17125 33416 20319 33418
rect 17125 33360 17130 33416
rect 17186 33360 20258 33416
rect 20314 33360 20319 33416
rect 17125 33358 20319 33360
rect 17125 33355 17191 33358
rect 20253 33355 20319 33358
rect 19333 33284 19399 33285
rect 19701 33284 19767 33285
rect 18822 33220 18828 33284
rect 18892 33282 18898 33284
rect 18892 33222 19258 33282
rect 18892 33220 18898 33222
rect 8363 33216 8679 33217
rect 8363 33152 8369 33216
rect 8433 33152 8449 33216
rect 8513 33152 8529 33216
rect 8593 33152 8609 33216
rect 8673 33152 8679 33216
rect 8363 33151 8679 33152
rect 13308 33216 13624 33217
rect 13308 33152 13314 33216
rect 13378 33152 13394 33216
rect 13458 33152 13474 33216
rect 13538 33152 13554 33216
rect 13618 33152 13624 33216
rect 13308 33151 13624 33152
rect 18253 33216 18569 33217
rect 18253 33152 18259 33216
rect 18323 33152 18339 33216
rect 18403 33152 18419 33216
rect 18483 33152 18499 33216
rect 18563 33152 18569 33216
rect 18253 33151 18569 33152
rect 4245 33144 7114 33146
rect 4245 33088 4250 33144
rect 4306 33088 7114 33144
rect 4245 33086 7114 33088
rect 8845 33146 8911 33149
rect 11237 33146 11303 33149
rect 8845 33144 11303 33146
rect 8845 33088 8850 33144
rect 8906 33088 11242 33144
rect 11298 33088 11303 33144
rect 8845 33086 11303 33088
rect 4245 33083 4311 33086
rect 8845 33083 8911 33086
rect 11237 33083 11303 33086
rect -300 32950 858 33010
rect 5165 33010 5231 33013
rect 8569 33010 8635 33013
rect 5165 33008 8635 33010
rect 5165 32952 5170 33008
rect 5226 32952 8574 33008
rect 8630 32952 8635 33008
rect 5165 32950 8635 32952
rect -300 32920 160 32950
rect 5165 32947 5231 32950
rect 8569 32947 8635 32950
rect 9029 33010 9095 33013
rect 9581 33010 9647 33013
rect 11973 33010 12039 33013
rect 9029 33008 12039 33010
rect 9029 32952 9034 33008
rect 9090 32952 9586 33008
rect 9642 32952 11978 33008
rect 12034 32952 12039 33008
rect 9029 32950 12039 32952
rect 9029 32947 9095 32950
rect 9581 32947 9647 32950
rect 11973 32947 12039 32950
rect 13169 33010 13235 33013
rect 16205 33010 16271 33013
rect 13169 33008 16271 33010
rect 13169 32952 13174 33008
rect 13230 32952 16210 33008
rect 16266 32952 16271 33008
rect 13169 32950 16271 32952
rect 13169 32947 13235 32950
rect 16205 32947 16271 32950
rect 18689 33010 18755 33013
rect 18822 33010 18828 33012
rect 18689 33008 18828 33010
rect 18689 32952 18694 33008
rect 18750 32952 18828 33008
rect 18689 32950 18828 32952
rect 18689 32947 18755 32950
rect 18822 32948 18828 32950
rect 18892 32948 18898 33012
rect 19198 33010 19258 33222
rect 19333 33280 19380 33284
rect 19444 33282 19450 33284
rect 19701 33282 19748 33284
rect 19333 33224 19338 33280
rect 19333 33220 19380 33224
rect 19444 33222 19490 33282
rect 19656 33280 19748 33282
rect 19656 33224 19706 33280
rect 19656 33222 19748 33224
rect 19444 33220 19450 33222
rect 19701 33220 19748 33222
rect 19812 33220 19818 33284
rect 20437 33282 20503 33285
rect 21840 33282 22300 33312
rect 20437 33280 22300 33282
rect 20437 33224 20442 33280
rect 20498 33224 22300 33280
rect 20437 33222 22300 33224
rect 19333 33219 19399 33220
rect 19701 33219 19767 33220
rect 20437 33219 20503 33222
rect 21840 33192 22300 33222
rect 19374 33010 19380 33012
rect 19198 32950 19380 33010
rect 19374 32948 19380 32950
rect 19444 32948 19450 33012
rect 473 32874 539 32877
rect 2446 32874 2452 32876
rect 473 32872 2452 32874
rect 473 32816 478 32872
rect 534 32816 2452 32872
rect 473 32814 2452 32816
rect 473 32811 539 32814
rect 2446 32812 2452 32814
rect 2516 32812 2522 32876
rect 3877 32874 3943 32877
rect 6310 32874 6316 32876
rect 3877 32872 6316 32874
rect 3877 32816 3882 32872
rect 3938 32816 6316 32872
rect 3877 32814 6316 32816
rect 3877 32811 3943 32814
rect 6310 32812 6316 32814
rect 6380 32812 6386 32876
rect 8886 32812 8892 32876
rect 8956 32874 8962 32876
rect 9029 32874 9095 32877
rect 8956 32872 9095 32874
rect 8956 32816 9034 32872
rect 9090 32816 9095 32872
rect 8956 32814 9095 32816
rect 8956 32812 8962 32814
rect 9029 32811 9095 32814
rect 14825 32874 14891 32877
rect 18689 32874 18755 32877
rect 20345 32874 20411 32877
rect 14825 32872 17786 32874
rect 14825 32816 14830 32872
rect 14886 32816 17786 32872
rect 14825 32814 17786 32816
rect 14825 32811 14891 32814
rect -300 32738 160 32768
rect 2773 32738 2839 32741
rect -300 32736 2839 32738
rect -300 32680 2778 32736
rect 2834 32680 2839 32736
rect -300 32678 2839 32680
rect -300 32648 160 32678
rect 2773 32675 2839 32678
rect 5890 32672 6206 32673
rect 5890 32608 5896 32672
rect 5960 32608 5976 32672
rect 6040 32608 6056 32672
rect 6120 32608 6136 32672
rect 6200 32608 6206 32672
rect 5890 32607 6206 32608
rect 10835 32672 11151 32673
rect 10835 32608 10841 32672
rect 10905 32608 10921 32672
rect 10985 32608 11001 32672
rect 11065 32608 11081 32672
rect 11145 32608 11151 32672
rect 10835 32607 11151 32608
rect 15780 32672 16096 32673
rect 15780 32608 15786 32672
rect 15850 32608 15866 32672
rect 15930 32608 15946 32672
rect 16010 32608 16026 32672
rect 16090 32608 16096 32672
rect 15780 32607 16096 32608
rect 1393 32600 1459 32605
rect 1393 32544 1398 32600
rect 1454 32544 1459 32600
rect 1393 32539 1459 32544
rect 2589 32602 2655 32605
rect 2773 32602 2839 32605
rect 5441 32602 5507 32605
rect 2589 32600 5507 32602
rect 2589 32544 2594 32600
rect 2650 32544 2778 32600
rect 2834 32544 5446 32600
rect 5502 32544 5507 32600
rect 2589 32542 5507 32544
rect 2589 32539 2655 32542
rect 2773 32539 2839 32542
rect 5441 32539 5507 32542
rect 13077 32604 13143 32605
rect 17726 32604 17786 32814
rect 18689 32872 20411 32874
rect 18689 32816 18694 32872
rect 18750 32816 20350 32872
rect 20406 32816 20411 32872
rect 18689 32814 20411 32816
rect 18689 32811 18755 32814
rect 20345 32811 20411 32814
rect 19425 32738 19491 32741
rect 20069 32738 20135 32741
rect 19425 32736 20135 32738
rect 19425 32680 19430 32736
rect 19486 32680 20074 32736
rect 20130 32680 20135 32736
rect 19425 32678 20135 32680
rect 19425 32675 19491 32678
rect 20069 32675 20135 32678
rect 21265 32738 21331 32741
rect 21840 32738 22300 32768
rect 21265 32736 22300 32738
rect 21265 32680 21270 32736
rect 21326 32680 22300 32736
rect 21265 32678 22300 32680
rect 21265 32675 21331 32678
rect 20725 32672 21041 32673
rect 20725 32608 20731 32672
rect 20795 32608 20811 32672
rect 20875 32608 20891 32672
rect 20955 32608 20971 32672
rect 21035 32608 21041 32672
rect 21840 32648 22300 32678
rect 20725 32607 21041 32608
rect 13077 32600 13124 32604
rect 13188 32602 13194 32604
rect 13077 32544 13082 32600
rect 13077 32540 13124 32544
rect 13188 32542 13234 32602
rect 13188 32540 13194 32542
rect 17718 32540 17724 32604
rect 17788 32540 17794 32604
rect 13077 32539 13143 32540
rect -300 32466 160 32496
rect 1396 32466 1456 32539
rect -300 32406 1456 32466
rect 4337 32466 4403 32469
rect 7373 32466 7439 32469
rect 17125 32466 17191 32469
rect 4337 32464 17191 32466
rect 4337 32408 4342 32464
rect 4398 32408 7378 32464
rect 7434 32408 17130 32464
rect 17186 32408 17191 32464
rect 4337 32406 17191 32408
rect -300 32376 160 32406
rect 4337 32403 4403 32406
rect 7373 32403 7439 32406
rect 17125 32403 17191 32406
rect 18045 32466 18111 32469
rect 19425 32466 19491 32469
rect 18045 32464 19491 32466
rect 18045 32408 18050 32464
rect 18106 32408 19430 32464
rect 19486 32408 19491 32464
rect 18045 32406 19491 32408
rect 18045 32403 18111 32406
rect 19425 32403 19491 32406
rect 3509 32330 3575 32333
rect 18229 32330 18295 32333
rect 3509 32328 18295 32330
rect 3509 32272 3514 32328
rect 3570 32272 18234 32328
rect 18290 32272 18295 32328
rect 3509 32270 18295 32272
rect 3509 32267 3575 32270
rect 18229 32267 18295 32270
rect -300 32194 160 32224
rect 1301 32194 1367 32197
rect -300 32192 1367 32194
rect -300 32136 1306 32192
rect 1362 32136 1367 32192
rect -300 32134 1367 32136
rect -300 32104 160 32134
rect 1301 32131 1367 32134
rect 4654 32132 4660 32196
rect 4724 32194 4730 32196
rect 4797 32194 4863 32197
rect 4724 32192 4863 32194
rect 4724 32136 4802 32192
rect 4858 32136 4863 32192
rect 4724 32134 4863 32136
rect 4724 32132 4730 32134
rect 4797 32131 4863 32134
rect 9673 32194 9739 32197
rect 11053 32194 11119 32197
rect 9673 32192 11119 32194
rect 9673 32136 9678 32192
rect 9734 32136 11058 32192
rect 11114 32136 11119 32192
rect 9673 32134 11119 32136
rect 9673 32131 9739 32134
rect 11053 32131 11119 32134
rect 20529 32194 20595 32197
rect 21840 32194 22300 32224
rect 20529 32192 22300 32194
rect 20529 32136 20534 32192
rect 20590 32136 22300 32192
rect 20529 32134 22300 32136
rect 20529 32131 20595 32134
rect 3418 32128 3734 32129
rect 3418 32064 3424 32128
rect 3488 32064 3504 32128
rect 3568 32064 3584 32128
rect 3648 32064 3664 32128
rect 3728 32064 3734 32128
rect 3418 32063 3734 32064
rect 8363 32128 8679 32129
rect 8363 32064 8369 32128
rect 8433 32064 8449 32128
rect 8513 32064 8529 32128
rect 8593 32064 8609 32128
rect 8673 32064 8679 32128
rect 8363 32063 8679 32064
rect 13308 32128 13624 32129
rect 13308 32064 13314 32128
rect 13378 32064 13394 32128
rect 13458 32064 13474 32128
rect 13538 32064 13554 32128
rect 13618 32064 13624 32128
rect 13308 32063 13624 32064
rect 18253 32128 18569 32129
rect 18253 32064 18259 32128
rect 18323 32064 18339 32128
rect 18403 32064 18419 32128
rect 18483 32064 18499 32128
rect 18563 32064 18569 32128
rect 21840 32104 22300 32134
rect 18253 32063 18569 32064
rect 4613 32058 4679 32061
rect 6269 32058 6335 32061
rect 4613 32056 6335 32058
rect 4613 32000 4618 32056
rect 4674 32000 6274 32056
rect 6330 32000 6335 32056
rect 4613 31998 6335 32000
rect 4613 31995 4679 31998
rect 6269 31995 6335 31998
rect 9949 32058 10015 32061
rect 10225 32058 10291 32061
rect 9949 32056 10291 32058
rect 9949 32000 9954 32056
rect 10010 32000 10230 32056
rect 10286 32000 10291 32056
rect 9949 31998 10291 32000
rect 9949 31995 10015 31998
rect 10225 31995 10291 31998
rect 14733 32056 14799 32061
rect 14733 32000 14738 32056
rect 14794 32000 14799 32056
rect 14733 31995 14799 32000
rect -300 31922 160 31952
rect 749 31922 815 31925
rect -300 31920 815 31922
rect -300 31864 754 31920
rect 810 31864 815 31920
rect -300 31862 815 31864
rect -300 31832 160 31862
rect 749 31859 815 31862
rect 1761 31922 1827 31925
rect 5022 31922 5028 31924
rect 1761 31920 5028 31922
rect 1761 31864 1766 31920
rect 1822 31864 5028 31920
rect 1761 31862 5028 31864
rect 1761 31859 1827 31862
rect 5022 31860 5028 31862
rect 5092 31860 5098 31924
rect 7005 31922 7071 31925
rect 9397 31922 9463 31925
rect 7005 31920 9463 31922
rect 7005 31864 7010 31920
rect 7066 31864 9402 31920
rect 9458 31864 9463 31920
rect 7005 31862 9463 31864
rect 7005 31859 7071 31862
rect 9397 31859 9463 31862
rect 12065 31922 12131 31925
rect 14736 31922 14796 31995
rect 15101 31922 15167 31925
rect 12065 31920 15167 31922
rect 12065 31864 12070 31920
rect 12126 31864 15106 31920
rect 15162 31864 15167 31920
rect 12065 31862 15167 31864
rect 12065 31859 12131 31862
rect 15101 31859 15167 31862
rect 17401 31922 17467 31925
rect 19057 31922 19123 31925
rect 17401 31920 19123 31922
rect 17401 31864 17406 31920
rect 17462 31864 19062 31920
rect 19118 31864 19123 31920
rect 17401 31862 19123 31864
rect 17401 31859 17467 31862
rect 19057 31859 19123 31862
rect 2221 31786 2287 31789
rect 8017 31786 8083 31789
rect 8937 31786 9003 31789
rect 614 31726 1594 31786
rect -300 31650 160 31680
rect 614 31650 674 31726
rect 1393 31650 1459 31653
rect -300 31590 674 31650
rect 752 31648 1459 31650
rect 752 31592 1398 31648
rect 1454 31592 1459 31648
rect 752 31590 1459 31592
rect 1534 31650 1594 31726
rect 2221 31784 9003 31786
rect 2221 31728 2226 31784
rect 2282 31728 8022 31784
rect 8078 31728 8942 31784
rect 8998 31728 9003 31784
rect 2221 31726 9003 31728
rect 2221 31723 2287 31726
rect 8017 31723 8083 31726
rect 8937 31723 9003 31726
rect 14273 31786 14339 31789
rect 15009 31786 15075 31789
rect 14273 31784 15075 31786
rect 14273 31728 14278 31784
rect 14334 31728 15014 31784
rect 15070 31728 15075 31784
rect 14273 31726 15075 31728
rect 14273 31723 14339 31726
rect 15009 31723 15075 31726
rect 18229 31786 18295 31789
rect 19885 31786 19951 31789
rect 18229 31784 19951 31786
rect 18229 31728 18234 31784
rect 18290 31728 19890 31784
rect 19946 31728 19951 31784
rect 18229 31726 19951 31728
rect 18229 31723 18295 31726
rect 19885 31723 19951 31726
rect 3785 31650 3851 31653
rect 1534 31648 3851 31650
rect 1534 31592 3790 31648
rect 3846 31592 3851 31648
rect 1534 31590 3851 31592
rect -300 31560 160 31590
rect -300 31378 160 31408
rect 752 31378 812 31590
rect 1393 31587 1459 31590
rect 3785 31587 3851 31590
rect 6862 31588 6868 31652
rect 6932 31650 6938 31652
rect 7005 31650 7071 31653
rect 6932 31648 7071 31650
rect 6932 31592 7010 31648
rect 7066 31592 7071 31648
rect 6932 31590 7071 31592
rect 6932 31588 6938 31590
rect 7005 31587 7071 31590
rect 7230 31588 7236 31652
rect 7300 31650 7306 31652
rect 7373 31650 7439 31653
rect 7300 31648 7439 31650
rect 7300 31592 7378 31648
rect 7434 31592 7439 31648
rect 7300 31590 7439 31592
rect 7300 31588 7306 31590
rect 7373 31587 7439 31590
rect 9397 31650 9463 31653
rect 9806 31650 9812 31652
rect 9397 31648 9812 31650
rect 9397 31592 9402 31648
rect 9458 31592 9812 31648
rect 9397 31590 9812 31592
rect 9397 31587 9463 31590
rect 9806 31588 9812 31590
rect 9876 31588 9882 31652
rect 13169 31650 13235 31653
rect 14733 31650 14799 31653
rect 21840 31650 22300 31680
rect 13169 31648 14799 31650
rect 13169 31592 13174 31648
rect 13230 31592 14738 31648
rect 14794 31592 14799 31648
rect 13169 31590 14799 31592
rect 13169 31587 13235 31590
rect 14733 31587 14799 31590
rect 21176 31590 22300 31650
rect 5890 31584 6206 31585
rect 5890 31520 5896 31584
rect 5960 31520 5976 31584
rect 6040 31520 6056 31584
rect 6120 31520 6136 31584
rect 6200 31520 6206 31584
rect 5890 31519 6206 31520
rect 10835 31584 11151 31585
rect 10835 31520 10841 31584
rect 10905 31520 10921 31584
rect 10985 31520 11001 31584
rect 11065 31520 11081 31584
rect 11145 31520 11151 31584
rect 10835 31519 11151 31520
rect 15780 31584 16096 31585
rect 15780 31520 15786 31584
rect 15850 31520 15866 31584
rect 15930 31520 15946 31584
rect 16010 31520 16026 31584
rect 16090 31520 16096 31584
rect 15780 31519 16096 31520
rect 20725 31584 21041 31585
rect 20725 31520 20731 31584
rect 20795 31520 20811 31584
rect 20875 31520 20891 31584
rect 20955 31520 20971 31584
rect 21035 31520 21041 31584
rect 20725 31519 21041 31520
rect 1945 31514 2011 31517
rect 5165 31514 5231 31517
rect 1945 31512 5231 31514
rect 1945 31456 1950 31512
rect 2006 31456 5170 31512
rect 5226 31456 5231 31512
rect 1945 31454 5231 31456
rect 1945 31451 2011 31454
rect 5165 31451 5231 31454
rect 8109 31514 8175 31517
rect 10409 31514 10475 31517
rect 8109 31512 10475 31514
rect 8109 31456 8114 31512
rect 8170 31456 10414 31512
rect 10470 31456 10475 31512
rect 8109 31454 10475 31456
rect 8109 31451 8175 31454
rect 10409 31451 10475 31454
rect 16430 31452 16436 31516
rect 16500 31514 16506 31516
rect 19742 31514 19748 31516
rect 16500 31454 19748 31514
rect 16500 31452 16506 31454
rect 19742 31452 19748 31454
rect 19812 31452 19818 31516
rect -300 31318 812 31378
rect -300 31288 160 31318
rect 2262 31316 2268 31380
rect 2332 31378 2338 31380
rect 2957 31378 3023 31381
rect 6269 31378 6335 31381
rect 2332 31376 6335 31378
rect 2332 31320 2962 31376
rect 3018 31320 6274 31376
rect 6330 31320 6335 31376
rect 2332 31318 6335 31320
rect 2332 31316 2338 31318
rect 2957 31315 3023 31318
rect 6269 31315 6335 31318
rect 8201 31378 8267 31381
rect 10777 31378 10843 31381
rect 15469 31378 15535 31381
rect 8201 31376 10843 31378
rect 8201 31320 8206 31376
rect 8262 31320 10782 31376
rect 10838 31320 10843 31376
rect 8201 31318 10843 31320
rect 8201 31315 8267 31318
rect 10777 31315 10843 31318
rect 11792 31376 15535 31378
rect 11792 31320 15474 31376
rect 15530 31320 15535 31376
rect 11792 31318 15535 31320
rect 11792 31245 11852 31318
rect 15469 31315 15535 31318
rect 15653 31378 15719 31381
rect 16430 31378 16436 31380
rect 15653 31376 16436 31378
rect 15653 31320 15658 31376
rect 15714 31320 16436 31376
rect 15653 31318 16436 31320
rect 15653 31315 15719 31318
rect 16430 31316 16436 31318
rect 16500 31316 16506 31380
rect 16941 31378 17007 31381
rect 18086 31378 18092 31380
rect 16941 31376 18092 31378
rect 16941 31320 16946 31376
rect 17002 31320 18092 31376
rect 16941 31318 18092 31320
rect 16941 31315 17007 31318
rect 18086 31316 18092 31318
rect 18156 31316 18162 31380
rect 18413 31378 18479 31381
rect 21176 31378 21236 31590
rect 21840 31560 22300 31590
rect 18413 31376 21236 31378
rect 18413 31320 18418 31376
rect 18474 31320 21236 31376
rect 18413 31318 21236 31320
rect 18413 31315 18479 31318
rect 2497 31242 2563 31245
rect 6913 31242 6979 31245
rect 2497 31240 6979 31242
rect 2497 31184 2502 31240
rect 2558 31184 6918 31240
rect 6974 31184 6979 31240
rect 2497 31182 6979 31184
rect 2497 31179 2563 31182
rect 6913 31179 6979 31182
rect 7097 31242 7163 31245
rect 7414 31242 7420 31244
rect 7097 31240 7420 31242
rect 7097 31184 7102 31240
rect 7158 31184 7420 31240
rect 7097 31182 7420 31184
rect 7097 31179 7163 31182
rect 7414 31180 7420 31182
rect 7484 31242 7490 31244
rect 11053 31242 11119 31245
rect 7484 31240 11119 31242
rect 7484 31184 11058 31240
rect 11114 31184 11119 31240
rect 7484 31182 11119 31184
rect 7484 31180 7490 31182
rect 11053 31179 11119 31182
rect 11278 31180 11284 31244
rect 11348 31242 11354 31244
rect 11789 31242 11855 31245
rect 18137 31242 18203 31245
rect 11348 31240 11855 31242
rect 11348 31184 11794 31240
rect 11850 31184 11855 31240
rect 11348 31182 11855 31184
rect 11348 31180 11354 31182
rect 11789 31179 11855 31182
rect 12390 31240 18203 31242
rect 12390 31184 18142 31240
rect 18198 31184 18203 31240
rect 12390 31182 18203 31184
rect -300 31106 160 31136
rect 1393 31106 1459 31109
rect 2865 31106 2931 31109
rect -300 31104 1459 31106
rect -300 31048 1398 31104
rect 1454 31048 1459 31104
rect -300 31046 1459 31048
rect -300 31016 160 31046
rect 1393 31043 1459 31046
rect 2730 31104 2931 31106
rect 2730 31048 2870 31104
rect 2926 31048 2931 31104
rect 2730 31046 2931 31048
rect -300 30834 160 30864
rect 2730 30834 2790 31046
rect 2865 31043 2931 31046
rect 4654 31044 4660 31108
rect 4724 31106 4730 31108
rect 5206 31106 5212 31108
rect 4724 31046 5212 31106
rect 4724 31044 4730 31046
rect 5206 31044 5212 31046
rect 5276 31044 5282 31108
rect 5390 31044 5396 31108
rect 5460 31106 5466 31108
rect 5809 31106 5875 31109
rect 12390 31106 12450 31182
rect 18137 31179 18203 31182
rect 18321 31242 18387 31245
rect 18321 31240 19304 31242
rect 18321 31184 18326 31240
rect 18382 31184 19304 31240
rect 18321 31182 19304 31184
rect 18321 31179 18387 31182
rect 19244 31109 19304 31182
rect 19926 31180 19932 31244
rect 19996 31242 20002 31244
rect 20621 31242 20687 31245
rect 19996 31240 20687 31242
rect 19996 31184 20626 31240
rect 20682 31184 20687 31240
rect 19996 31182 20687 31184
rect 19996 31180 20002 31182
rect 20621 31179 20687 31182
rect 5460 31104 5875 31106
rect 5460 31048 5814 31104
rect 5870 31048 5875 31104
rect 5460 31046 5875 31048
rect 5460 31044 5466 31046
rect 5809 31043 5875 31046
rect 10550 31046 12450 31106
rect 16297 31106 16363 31109
rect 16798 31106 16804 31108
rect 16297 31104 16804 31106
rect 16297 31048 16302 31104
rect 16358 31048 16804 31104
rect 16297 31046 16804 31048
rect 3418 31040 3734 31041
rect 3418 30976 3424 31040
rect 3488 30976 3504 31040
rect 3568 30976 3584 31040
rect 3648 30976 3664 31040
rect 3728 30976 3734 31040
rect 3418 30975 3734 30976
rect 8363 31040 8679 31041
rect 8363 30976 8369 31040
rect 8433 30976 8449 31040
rect 8513 30976 8529 31040
rect 8593 30976 8609 31040
rect 8673 30976 8679 31040
rect 8363 30975 8679 30976
rect 8109 30970 8175 30973
rect 5030 30968 8175 30970
rect 5030 30912 8114 30968
rect 8170 30912 8175 30968
rect 5030 30910 8175 30912
rect -300 30774 2790 30834
rect 3601 30834 3667 30837
rect 5030 30834 5090 30910
rect 8109 30907 8175 30910
rect 3601 30832 5090 30834
rect 3601 30776 3606 30832
rect 3662 30776 5090 30832
rect 3601 30774 5090 30776
rect -300 30744 160 30774
rect 3601 30771 3667 30774
rect 5206 30772 5212 30836
rect 5276 30834 5282 30836
rect 9765 30834 9831 30837
rect 5276 30832 9831 30834
rect 5276 30776 9770 30832
rect 9826 30776 9831 30832
rect 5276 30774 9831 30776
rect 5276 30772 5282 30774
rect 9765 30771 9831 30774
rect 1853 30698 1919 30701
rect 7189 30698 7255 30701
rect 8201 30700 8267 30701
rect 1853 30696 7255 30698
rect 1853 30640 1858 30696
rect 1914 30640 7194 30696
rect 7250 30640 7255 30696
rect 1853 30638 7255 30640
rect 1853 30635 1919 30638
rect 7189 30635 7255 30638
rect 8150 30636 8156 30700
rect 8220 30698 8267 30700
rect 8220 30696 8312 30698
rect 8262 30640 8312 30696
rect 8220 30638 8312 30640
rect 8220 30636 8267 30638
rect 8201 30635 8267 30636
rect -300 30562 160 30592
rect 2773 30562 2839 30565
rect -300 30560 2839 30562
rect -300 30504 2778 30560
rect 2834 30504 2839 30560
rect -300 30502 2839 30504
rect -300 30472 160 30502
rect 2773 30499 2839 30502
rect 5890 30496 6206 30497
rect 5890 30432 5896 30496
rect 5960 30432 5976 30496
rect 6040 30432 6056 30496
rect 6120 30432 6136 30496
rect 6200 30432 6206 30496
rect 5890 30431 6206 30432
rect 2497 30426 2563 30429
rect 5349 30426 5415 30429
rect 2497 30424 5415 30426
rect 2497 30368 2502 30424
rect 2558 30368 5354 30424
rect 5410 30368 5415 30424
rect 2497 30366 5415 30368
rect 2497 30363 2563 30366
rect 5349 30363 5415 30366
rect 7557 30426 7623 30429
rect 10550 30426 10610 31046
rect 16297 31043 16363 31046
rect 16798 31044 16804 31046
rect 16868 31044 16874 31108
rect 18689 31106 18755 31109
rect 19057 31106 19123 31109
rect 18689 31104 19123 31106
rect 18689 31048 18694 31104
rect 18750 31048 19062 31104
rect 19118 31048 19123 31104
rect 18689 31046 19123 31048
rect 18689 31043 18755 31046
rect 19057 31043 19123 31046
rect 19241 31104 19307 31109
rect 19241 31048 19246 31104
rect 19302 31048 19307 31104
rect 19241 31043 19307 31048
rect 20437 31106 20503 31109
rect 21840 31106 22300 31136
rect 20437 31104 22300 31106
rect 20437 31048 20442 31104
rect 20498 31048 22300 31104
rect 20437 31046 22300 31048
rect 20437 31043 20503 31046
rect 13308 31040 13624 31041
rect 13308 30976 13314 31040
rect 13378 30976 13394 31040
rect 13458 30976 13474 31040
rect 13538 30976 13554 31040
rect 13618 30976 13624 31040
rect 13308 30975 13624 30976
rect 18253 31040 18569 31041
rect 18253 30976 18259 31040
rect 18323 30976 18339 31040
rect 18403 30976 18419 31040
rect 18483 30976 18499 31040
rect 18563 30976 18569 31040
rect 21840 31016 22300 31046
rect 18253 30975 18569 30976
rect 14641 30970 14707 30973
rect 13862 30968 14707 30970
rect 13862 30912 14646 30968
rect 14702 30912 14707 30968
rect 13862 30910 14707 30912
rect 13862 30837 13922 30910
rect 14641 30907 14707 30910
rect 18781 30970 18847 30973
rect 19793 30970 19859 30973
rect 18781 30968 19859 30970
rect 18781 30912 18786 30968
rect 18842 30912 19798 30968
rect 19854 30912 19859 30968
rect 18781 30910 19859 30912
rect 18781 30907 18847 30910
rect 19793 30907 19859 30910
rect 13813 30832 13922 30837
rect 13813 30776 13818 30832
rect 13874 30776 13922 30832
rect 13813 30774 13922 30776
rect 14089 30834 14155 30837
rect 17125 30834 17191 30837
rect 19149 30834 19215 30837
rect 14089 30832 14290 30834
rect 14089 30776 14094 30832
rect 14150 30776 14290 30832
rect 14089 30774 14290 30776
rect 13813 30771 13879 30774
rect 14089 30771 14155 30774
rect 10777 30698 10843 30701
rect 14089 30698 14155 30701
rect 10777 30696 14155 30698
rect 10777 30640 10782 30696
rect 10838 30640 14094 30696
rect 14150 30640 14155 30696
rect 10777 30638 14155 30640
rect 10777 30635 10843 30638
rect 14089 30635 14155 30638
rect 12433 30562 12499 30565
rect 14038 30562 14044 30564
rect 12433 30560 14044 30562
rect 12433 30504 12438 30560
rect 12494 30504 14044 30560
rect 12433 30502 14044 30504
rect 12433 30499 12499 30502
rect 14038 30500 14044 30502
rect 14108 30500 14114 30564
rect 10835 30496 11151 30497
rect 10835 30432 10841 30496
rect 10905 30432 10921 30496
rect 10985 30432 11001 30496
rect 11065 30432 11081 30496
rect 11145 30432 11151 30496
rect 10835 30431 11151 30432
rect 7557 30424 10610 30426
rect 7557 30368 7562 30424
rect 7618 30368 10610 30424
rect 7557 30366 10610 30368
rect 7557 30363 7623 30366
rect -300 30290 160 30320
rect 3417 30290 3483 30293
rect -300 30288 3483 30290
rect -300 30232 3422 30288
rect 3478 30232 3483 30288
rect -300 30230 3483 30232
rect -300 30200 160 30230
rect 3417 30227 3483 30230
rect 4797 30290 4863 30293
rect 5073 30290 5139 30293
rect 4797 30288 5139 30290
rect 4797 30232 4802 30288
rect 4858 30232 5078 30288
rect 5134 30232 5139 30288
rect 4797 30230 5139 30232
rect 4797 30227 4863 30230
rect 5073 30227 5139 30230
rect 5533 30290 5599 30293
rect 6545 30290 6611 30293
rect 5533 30288 6611 30290
rect 5533 30232 5538 30288
rect 5594 30232 6550 30288
rect 6606 30232 6611 30288
rect 5533 30230 6611 30232
rect 14230 30290 14290 30774
rect 17125 30832 19215 30834
rect 17125 30776 17130 30832
rect 17186 30776 19154 30832
rect 19210 30776 19215 30832
rect 17125 30774 19215 30776
rect 17125 30771 17191 30774
rect 19149 30771 19215 30774
rect 15653 30698 15719 30701
rect 16614 30698 16620 30700
rect 15653 30696 16620 30698
rect 15653 30640 15658 30696
rect 15714 30640 16620 30696
rect 15653 30638 16620 30640
rect 15653 30635 15719 30638
rect 16614 30636 16620 30638
rect 16684 30636 16690 30700
rect 19006 30562 19012 30564
rect 17174 30502 19012 30562
rect 15780 30496 16096 30497
rect 15780 30432 15786 30496
rect 15850 30432 15866 30496
rect 15930 30432 15946 30496
rect 16010 30432 16026 30496
rect 16090 30432 16096 30496
rect 15780 30431 16096 30432
rect 16205 30426 16271 30429
rect 17174 30426 17234 30502
rect 19006 30500 19012 30502
rect 19076 30500 19082 30564
rect 21265 30562 21331 30565
rect 21840 30562 22300 30592
rect 21265 30560 22300 30562
rect 21265 30504 21270 30560
rect 21326 30504 22300 30560
rect 21265 30502 22300 30504
rect 21265 30499 21331 30502
rect 20725 30496 21041 30497
rect 20725 30432 20731 30496
rect 20795 30432 20811 30496
rect 20875 30432 20891 30496
rect 20955 30432 20971 30496
rect 21035 30432 21041 30496
rect 21840 30472 22300 30502
rect 20725 30431 21041 30432
rect 16205 30424 17234 30426
rect 16205 30368 16210 30424
rect 16266 30368 17234 30424
rect 16205 30366 17234 30368
rect 16205 30363 16271 30366
rect 17350 30364 17356 30428
rect 17420 30426 17426 30428
rect 19006 30426 19012 30428
rect 17420 30366 19012 30426
rect 17420 30364 17426 30366
rect 19006 30364 19012 30366
rect 19076 30364 19082 30428
rect 14230 30230 16866 30290
rect 5533 30227 5599 30230
rect 6545 30227 6611 30230
rect 1025 30156 1091 30157
rect 974 30154 980 30156
rect 934 30094 980 30154
rect 1044 30152 1091 30156
rect 1761 30154 1827 30157
rect 1086 30096 1091 30152
rect 974 30092 980 30094
rect 1044 30092 1091 30096
rect 1025 30091 1091 30092
rect 1718 30152 1827 30154
rect 1718 30096 1766 30152
rect 1822 30096 1827 30152
rect 1718 30091 1827 30096
rect 2078 30092 2084 30156
rect 2148 30154 2154 30156
rect 4429 30154 4495 30157
rect 2148 30152 4495 30154
rect 2148 30096 4434 30152
rect 4490 30096 4495 30152
rect 2148 30094 4495 30096
rect 2148 30092 2154 30094
rect 4429 30091 4495 30094
rect 5441 30154 5507 30157
rect 9121 30154 9187 30157
rect 5441 30152 9187 30154
rect 5441 30096 5446 30152
rect 5502 30096 9126 30152
rect 9182 30096 9187 30152
rect 5441 30094 9187 30096
rect 5441 30091 5507 30094
rect 9121 30091 9187 30094
rect 11697 30154 11763 30157
rect 15469 30154 15535 30157
rect 16806 30156 16866 30230
rect 11697 30152 15535 30154
rect 11697 30096 11702 30152
rect 11758 30096 15474 30152
rect 15530 30096 15535 30152
rect 11697 30094 15535 30096
rect 11697 30091 11763 30094
rect 15469 30091 15535 30094
rect 16798 30092 16804 30156
rect 16868 30092 16874 30156
rect 18229 30154 18295 30157
rect 19241 30154 19307 30157
rect 18229 30152 19307 30154
rect 18229 30096 18234 30152
rect 18290 30096 19246 30152
rect 19302 30096 19307 30152
rect 18229 30094 19307 30096
rect 18229 30091 18295 30094
rect 19241 30091 19307 30094
rect -300 30018 160 30048
rect 1718 30018 1778 30091
rect 3969 30020 4035 30021
rect -300 29958 1778 30018
rect -300 29928 160 29958
rect 3918 29956 3924 30020
rect 3988 30018 4035 30020
rect 20437 30018 20503 30021
rect 21840 30018 22300 30048
rect 3988 30016 4080 30018
rect 4030 29960 4080 30016
rect 3988 29958 4080 29960
rect 20437 30016 22300 30018
rect 20437 29960 20442 30016
rect 20498 29960 22300 30016
rect 20437 29958 22300 29960
rect 3988 29956 4035 29958
rect 3969 29955 4035 29956
rect 20437 29955 20503 29958
rect 3418 29952 3734 29953
rect 3418 29888 3424 29952
rect 3488 29888 3504 29952
rect 3568 29888 3584 29952
rect 3648 29888 3664 29952
rect 3728 29888 3734 29952
rect 3418 29887 3734 29888
rect 8363 29952 8679 29953
rect 8363 29888 8369 29952
rect 8433 29888 8449 29952
rect 8513 29888 8529 29952
rect 8593 29888 8609 29952
rect 8673 29888 8679 29952
rect 8363 29887 8679 29888
rect 13308 29952 13624 29953
rect 13308 29888 13314 29952
rect 13378 29888 13394 29952
rect 13458 29888 13474 29952
rect 13538 29888 13554 29952
rect 13618 29888 13624 29952
rect 13308 29887 13624 29888
rect 18253 29952 18569 29953
rect 18253 29888 18259 29952
rect 18323 29888 18339 29952
rect 18403 29888 18419 29952
rect 18483 29888 18499 29952
rect 18563 29888 18569 29952
rect 21840 29928 22300 29958
rect 18253 29887 18569 29888
rect 2773 29880 2839 29885
rect 2773 29824 2778 29880
rect 2834 29824 2839 29880
rect 2773 29819 2839 29824
rect 4153 29882 4219 29885
rect 4286 29882 4292 29884
rect 4153 29880 4292 29882
rect 4153 29824 4158 29880
rect 4214 29824 4292 29880
rect 4153 29822 4292 29824
rect 4153 29819 4219 29822
rect 4286 29820 4292 29822
rect 4356 29882 4362 29884
rect 7414 29882 7420 29884
rect 4356 29822 7420 29882
rect 4356 29820 4362 29822
rect 7414 29820 7420 29822
rect 7484 29820 7490 29884
rect -300 29746 160 29776
rect 1209 29746 1275 29749
rect -300 29744 1275 29746
rect -300 29688 1214 29744
rect 1270 29688 1275 29744
rect -300 29686 1275 29688
rect 2776 29746 2836 29819
rect 3325 29746 3391 29749
rect 2776 29744 3391 29746
rect 2776 29688 3330 29744
rect 3386 29688 3391 29744
rect 2776 29686 3391 29688
rect -300 29656 160 29686
rect 1209 29683 1275 29686
rect 3325 29683 3391 29686
rect 3969 29746 4035 29749
rect 5206 29746 5212 29748
rect 3969 29744 5212 29746
rect 3969 29688 3974 29744
rect 4030 29688 5212 29744
rect 3969 29686 5212 29688
rect 3969 29683 4035 29686
rect 5206 29684 5212 29686
rect 5276 29684 5282 29748
rect 7373 29746 7439 29749
rect 11697 29746 11763 29749
rect 7373 29744 11763 29746
rect 7373 29688 7378 29744
rect 7434 29688 11702 29744
rect 11758 29688 11763 29744
rect 7373 29686 11763 29688
rect 7373 29683 7439 29686
rect 11697 29683 11763 29686
rect 14222 29684 14228 29748
rect 14292 29746 14298 29748
rect 15101 29746 15167 29749
rect 14292 29744 15167 29746
rect 14292 29688 15106 29744
rect 15162 29688 15167 29744
rect 14292 29686 15167 29688
rect 14292 29684 14298 29686
rect 15101 29683 15167 29686
rect 1669 29610 1735 29613
rect 1669 29608 11714 29610
rect 1669 29552 1674 29608
rect 1730 29552 11714 29608
rect 1669 29550 11714 29552
rect 1669 29547 1735 29550
rect -300 29474 160 29504
rect 565 29474 631 29477
rect -300 29472 631 29474
rect -300 29416 570 29472
rect 626 29416 631 29472
rect -300 29414 631 29416
rect -300 29384 160 29414
rect 565 29411 631 29414
rect 2957 29474 3023 29477
rect 4337 29474 4403 29477
rect 2957 29472 4403 29474
rect 2957 29416 2962 29472
rect 3018 29416 4342 29472
rect 4398 29416 4403 29472
rect 2957 29414 4403 29416
rect 2957 29411 3023 29414
rect 4337 29411 4403 29414
rect 6269 29474 6335 29477
rect 7782 29474 7788 29476
rect 6269 29472 7788 29474
rect 6269 29416 6274 29472
rect 6330 29416 7788 29472
rect 6269 29414 7788 29416
rect 6269 29411 6335 29414
rect 7782 29412 7788 29414
rect 7852 29412 7858 29476
rect 5890 29408 6206 29409
rect 5890 29344 5896 29408
rect 5960 29344 5976 29408
rect 6040 29344 6056 29408
rect 6120 29344 6136 29408
rect 6200 29344 6206 29408
rect 5890 29343 6206 29344
rect 10835 29408 11151 29409
rect 10835 29344 10841 29408
rect 10905 29344 10921 29408
rect 10985 29344 11001 29408
rect 11065 29344 11081 29408
rect 11145 29344 11151 29408
rect 10835 29343 11151 29344
rect 2773 29338 2839 29341
rect 2998 29338 3004 29340
rect 2773 29336 3004 29338
rect 2773 29280 2778 29336
rect 2834 29280 3004 29336
rect 2773 29278 3004 29280
rect 2773 29275 2839 29278
rect 2998 29276 3004 29278
rect 3068 29276 3074 29340
rect 3417 29338 3483 29341
rect 4654 29338 4660 29340
rect 3417 29336 4660 29338
rect 3417 29280 3422 29336
rect 3478 29280 4660 29336
rect 3417 29278 4660 29280
rect 3417 29275 3483 29278
rect 4654 29276 4660 29278
rect 4724 29276 4730 29340
rect 5022 29276 5028 29340
rect 5092 29338 5098 29340
rect 5441 29338 5507 29341
rect 11654 29338 11714 29550
rect 19374 29548 19380 29612
rect 19444 29610 19450 29612
rect 19517 29610 19583 29613
rect 19444 29608 19583 29610
rect 19444 29552 19522 29608
rect 19578 29552 19583 29608
rect 19444 29550 19583 29552
rect 19444 29548 19450 29550
rect 19517 29547 19583 29550
rect 13813 29474 13879 29477
rect 12390 29472 13879 29474
rect 12390 29416 13818 29472
rect 13874 29416 13879 29472
rect 12390 29414 13879 29416
rect 12390 29338 12450 29414
rect 13813 29411 13879 29414
rect 21265 29474 21331 29477
rect 21840 29474 22300 29504
rect 21265 29472 22300 29474
rect 21265 29416 21270 29472
rect 21326 29416 22300 29472
rect 21265 29414 22300 29416
rect 21265 29411 21331 29414
rect 15780 29408 16096 29409
rect 15780 29344 15786 29408
rect 15850 29344 15866 29408
rect 15930 29344 15946 29408
rect 16010 29344 16026 29408
rect 16090 29344 16096 29408
rect 15780 29343 16096 29344
rect 20725 29408 21041 29409
rect 20725 29344 20731 29408
rect 20795 29344 20811 29408
rect 20875 29344 20891 29408
rect 20955 29344 20971 29408
rect 21035 29344 21041 29408
rect 21840 29384 22300 29414
rect 20725 29343 21041 29344
rect 5092 29336 5780 29338
rect 5092 29280 5446 29336
rect 5502 29280 5780 29336
rect 5092 29278 5780 29280
rect 5092 29276 5098 29278
rect 5441 29275 5507 29278
rect -300 29202 160 29232
rect 1577 29202 1643 29205
rect 5533 29202 5599 29205
rect -300 29200 1643 29202
rect -300 29144 1582 29200
rect 1638 29144 1643 29200
rect -300 29142 1643 29144
rect -300 29112 160 29142
rect 1577 29139 1643 29142
rect 4294 29200 5599 29202
rect 4294 29144 5538 29200
rect 5594 29144 5599 29200
rect 4294 29142 5599 29144
rect 5720 29202 5780 29278
rect 7606 29278 9690 29338
rect 11654 29278 12450 29338
rect 12709 29338 12775 29341
rect 13118 29338 13124 29340
rect 12709 29336 13124 29338
rect 12709 29280 12714 29336
rect 12770 29280 13124 29336
rect 12709 29278 13124 29280
rect 7606 29202 7666 29278
rect 5720 29142 7666 29202
rect 7741 29202 7807 29205
rect 9438 29202 9444 29204
rect 7741 29200 9444 29202
rect 7741 29144 7746 29200
rect 7802 29144 9444 29200
rect 7741 29142 9444 29144
rect 1158 29004 1164 29068
rect 1228 29066 1234 29068
rect 1301 29066 1367 29069
rect 1228 29064 1367 29066
rect 1228 29008 1306 29064
rect 1362 29008 1367 29064
rect 1228 29006 1367 29008
rect 1228 29004 1234 29006
rect 1301 29003 1367 29006
rect 1526 29004 1532 29068
rect 1596 29066 1602 29068
rect 2405 29066 2471 29069
rect 4294 29066 4354 29142
rect 5533 29139 5599 29142
rect 7741 29139 7807 29142
rect 9438 29140 9444 29142
rect 9508 29140 9514 29204
rect 9630 29202 9690 29278
rect 12709 29275 12775 29278
rect 13118 29276 13124 29278
rect 13188 29276 13194 29340
rect 14222 29202 14228 29204
rect 9630 29142 14228 29202
rect 14222 29140 14228 29142
rect 14292 29140 14298 29204
rect 16430 29140 16436 29204
rect 16500 29202 16506 29204
rect 17033 29202 17099 29205
rect 16500 29200 17099 29202
rect 16500 29144 17038 29200
rect 17094 29144 17099 29200
rect 16500 29142 17099 29144
rect 16500 29140 16506 29142
rect 17033 29139 17099 29142
rect 18638 29140 18644 29204
rect 18708 29202 18714 29204
rect 19057 29202 19123 29205
rect 18708 29200 19123 29202
rect 18708 29144 19062 29200
rect 19118 29144 19123 29200
rect 18708 29142 19123 29144
rect 18708 29140 18714 29142
rect 19057 29139 19123 29142
rect 19241 29202 19307 29205
rect 21265 29202 21331 29205
rect 19241 29200 21331 29202
rect 19241 29144 19246 29200
rect 19302 29144 21270 29200
rect 21326 29144 21331 29200
rect 19241 29142 21331 29144
rect 19241 29139 19307 29142
rect 21265 29139 21331 29142
rect 1596 29064 2471 29066
rect 1596 29008 2410 29064
rect 2466 29008 2471 29064
rect 1596 29006 2471 29008
rect 1596 29004 1602 29006
rect 2405 29003 2471 29006
rect 2730 29006 4354 29066
rect 4797 29066 4863 29069
rect 8293 29066 8359 29069
rect 9397 29068 9463 29069
rect 4797 29064 8359 29066
rect 4797 29008 4802 29064
rect 4858 29008 8298 29064
rect 8354 29008 8359 29064
rect 4797 29006 8359 29008
rect -300 28930 160 28960
rect 749 28930 815 28933
rect -300 28928 815 28930
rect -300 28872 754 28928
rect 810 28872 815 28928
rect -300 28870 815 28872
rect -300 28840 160 28870
rect 749 28867 815 28870
rect 1894 28868 1900 28932
rect 1964 28930 1970 28932
rect 2730 28930 2790 29006
rect 4797 29003 4863 29006
rect 8293 29003 8359 29006
rect 9254 29004 9260 29068
rect 9324 29004 9330 29068
rect 9397 29064 9444 29068
rect 9508 29066 9514 29068
rect 10317 29066 10383 29069
rect 10542 29066 10548 29068
rect 9397 29008 9402 29064
rect 9397 29004 9444 29008
rect 9508 29006 9554 29066
rect 10317 29064 10548 29066
rect 10317 29008 10322 29064
rect 10378 29008 10548 29064
rect 10317 29006 10548 29008
rect 9508 29004 9514 29006
rect 3233 28930 3299 28933
rect 1964 28870 2790 28930
rect 3190 28928 3299 28930
rect 3190 28872 3238 28928
rect 3294 28872 3299 28928
rect 1964 28868 1970 28870
rect 3190 28867 3299 28872
rect 9262 28930 9322 29004
rect 9397 29003 9463 29004
rect 10317 29003 10383 29006
rect 10542 29004 10548 29006
rect 10612 29066 10618 29068
rect 11237 29066 11303 29069
rect 10612 29064 11303 29066
rect 10612 29008 11242 29064
rect 11298 29008 11303 29064
rect 10612 29006 11303 29008
rect 10612 29004 10618 29006
rect 11237 29003 11303 29006
rect 12157 29066 12223 29069
rect 15193 29068 15259 29069
rect 14406 29066 14412 29068
rect 12157 29064 14412 29066
rect 12157 29008 12162 29064
rect 12218 29008 14412 29064
rect 12157 29006 14412 29008
rect 12157 29003 12223 29006
rect 14406 29004 14412 29006
rect 14476 29004 14482 29068
rect 15142 29066 15148 29068
rect 15102 29006 15148 29066
rect 15212 29064 15259 29068
rect 15254 29008 15259 29064
rect 15142 29004 15148 29006
rect 15212 29004 15259 29008
rect 16982 29004 16988 29068
rect 17052 29066 17058 29068
rect 17401 29066 17467 29069
rect 17052 29064 17467 29066
rect 17052 29008 17406 29064
rect 17462 29008 17467 29064
rect 17052 29006 17467 29008
rect 17052 29004 17058 29006
rect 15193 29003 15259 29004
rect 17401 29003 17467 29006
rect 17585 29066 17651 29069
rect 17718 29066 17724 29068
rect 17585 29064 17724 29066
rect 17585 29008 17590 29064
rect 17646 29008 17724 29064
rect 17585 29006 17724 29008
rect 17585 29003 17651 29006
rect 17718 29004 17724 29006
rect 17788 29004 17794 29068
rect 9857 28930 9923 28933
rect 12709 28932 12775 28933
rect 12709 28930 12756 28932
rect 9262 28928 9923 28930
rect 9262 28872 9862 28928
rect 9918 28872 9923 28928
rect 9262 28870 9923 28872
rect 12664 28928 12756 28930
rect 12664 28872 12714 28928
rect 12664 28870 12756 28872
rect 9857 28867 9923 28870
rect 12709 28868 12756 28870
rect 12820 28868 12826 28932
rect 12934 28868 12940 28932
rect 13004 28930 13010 28932
rect 13169 28930 13235 28933
rect 13004 28928 13235 28930
rect 13004 28872 13174 28928
rect 13230 28872 13235 28928
rect 13004 28870 13235 28872
rect 13004 28868 13010 28870
rect 12709 28867 12775 28868
rect 13169 28867 13235 28870
rect 20437 28930 20503 28933
rect 21840 28930 22300 28960
rect 20437 28928 22300 28930
rect 20437 28872 20442 28928
rect 20498 28872 22300 28928
rect 20437 28870 22300 28872
rect 20437 28867 20503 28870
rect 1025 28794 1091 28797
rect 3190 28794 3250 28867
rect 3418 28864 3734 28865
rect 3418 28800 3424 28864
rect 3488 28800 3504 28864
rect 3568 28800 3584 28864
rect 3648 28800 3664 28864
rect 3728 28800 3734 28864
rect 3418 28799 3734 28800
rect 8363 28864 8679 28865
rect 8363 28800 8369 28864
rect 8433 28800 8449 28864
rect 8513 28800 8529 28864
rect 8593 28800 8609 28864
rect 8673 28800 8679 28864
rect 8363 28799 8679 28800
rect 13308 28864 13624 28865
rect 13308 28800 13314 28864
rect 13378 28800 13394 28864
rect 13458 28800 13474 28864
rect 13538 28800 13554 28864
rect 13618 28800 13624 28864
rect 13308 28799 13624 28800
rect 18253 28864 18569 28865
rect 18253 28800 18259 28864
rect 18323 28800 18339 28864
rect 18403 28800 18419 28864
rect 18483 28800 18499 28864
rect 18563 28800 18569 28864
rect 21840 28840 22300 28870
rect 18253 28799 18569 28800
rect 1025 28792 3250 28794
rect 1025 28736 1030 28792
rect 1086 28736 3250 28792
rect 1025 28734 3250 28736
rect 6453 28794 6519 28797
rect 7414 28794 7420 28796
rect 6453 28792 7420 28794
rect 6453 28736 6458 28792
rect 6514 28736 7420 28792
rect 6453 28734 7420 28736
rect 1025 28731 1091 28734
rect 6453 28731 6519 28734
rect 7414 28732 7420 28734
rect 7484 28732 7490 28796
rect -300 28658 160 28688
rect 1485 28658 1551 28661
rect -300 28656 1551 28658
rect -300 28600 1490 28656
rect 1546 28600 1551 28656
rect -300 28598 1551 28600
rect -300 28568 160 28598
rect 1485 28595 1551 28598
rect 1669 28658 1735 28661
rect 2262 28658 2268 28660
rect 1669 28656 2268 28658
rect 1669 28600 1674 28656
rect 1730 28600 2268 28656
rect 1669 28598 2268 28600
rect 1669 28595 1735 28598
rect 2262 28596 2268 28598
rect 2332 28596 2338 28660
rect 2589 28658 2655 28661
rect 8293 28658 8359 28661
rect 2589 28656 8359 28658
rect 2589 28600 2594 28656
rect 2650 28600 8298 28656
rect 8354 28600 8359 28656
rect 2589 28598 8359 28600
rect 2589 28595 2655 28598
rect 8293 28595 8359 28598
rect 9581 28658 9647 28661
rect 10317 28658 10383 28661
rect 9581 28656 10383 28658
rect 9581 28600 9586 28656
rect 9642 28600 10322 28656
rect 10378 28600 10383 28656
rect 9581 28598 10383 28600
rect 9581 28595 9647 28598
rect 10317 28595 10383 28598
rect 11789 28656 11855 28661
rect 11789 28600 11794 28656
rect 11850 28600 11855 28656
rect 11789 28595 11855 28600
rect 13813 28658 13879 28661
rect 14038 28658 14044 28660
rect 13813 28656 14044 28658
rect 13813 28600 13818 28656
rect 13874 28600 14044 28656
rect 13813 28598 14044 28600
rect 13813 28595 13879 28598
rect 14038 28596 14044 28598
rect 14108 28658 14114 28660
rect 15193 28658 15259 28661
rect 14108 28656 15259 28658
rect 14108 28600 15198 28656
rect 15254 28600 15259 28656
rect 14108 28598 15259 28600
rect 14108 28596 14114 28598
rect 15193 28595 15259 28598
rect 1669 28522 1735 28525
rect 8109 28522 8175 28525
rect 10685 28522 10751 28525
rect 1669 28520 8034 28522
rect 1669 28464 1674 28520
rect 1730 28464 8034 28520
rect 1669 28462 8034 28464
rect 1669 28459 1735 28462
rect -300 28386 160 28416
rect 4613 28386 4679 28389
rect -300 28384 4679 28386
rect -300 28328 4618 28384
rect 4674 28328 4679 28384
rect -300 28326 4679 28328
rect 7974 28386 8034 28462
rect 8109 28520 10751 28522
rect 8109 28464 8114 28520
rect 8170 28464 10690 28520
rect 10746 28464 10751 28520
rect 8109 28462 10751 28464
rect 8109 28459 8175 28462
rect 10685 28459 10751 28462
rect 10041 28386 10107 28389
rect 7974 28384 10107 28386
rect 7974 28328 10046 28384
rect 10102 28328 10107 28384
rect 7974 28326 10107 28328
rect -300 28296 160 28326
rect 4613 28323 4679 28326
rect 10041 28323 10107 28326
rect 5890 28320 6206 28321
rect 5890 28256 5896 28320
rect 5960 28256 5976 28320
rect 6040 28256 6056 28320
rect 6120 28256 6136 28320
rect 6200 28256 6206 28320
rect 5890 28255 6206 28256
rect 10835 28320 11151 28321
rect 10835 28256 10841 28320
rect 10905 28256 10921 28320
rect 10985 28256 11001 28320
rect 11065 28256 11081 28320
rect 11145 28256 11151 28320
rect 10835 28255 11151 28256
rect 2078 28188 2084 28252
rect 2148 28250 2154 28252
rect 2405 28250 2471 28253
rect 2148 28248 2471 28250
rect 2148 28192 2410 28248
rect 2466 28192 2471 28248
rect 2148 28190 2471 28192
rect 2148 28188 2154 28190
rect 2405 28187 2471 28190
rect 2814 28188 2820 28252
rect 2884 28250 2890 28252
rect 3049 28250 3115 28253
rect 2884 28248 3115 28250
rect 2884 28192 3054 28248
rect 3110 28192 3115 28248
rect 2884 28190 3115 28192
rect 2884 28188 2890 28190
rect 3049 28187 3115 28190
rect 5073 28248 5139 28253
rect 5073 28192 5078 28248
rect 5134 28192 5139 28248
rect 5073 28187 5139 28192
rect -300 28114 160 28144
rect 3785 28114 3851 28117
rect 5076 28116 5136 28187
rect 11792 28117 11852 28595
rect 12750 28460 12756 28524
rect 12820 28522 12826 28524
rect 14089 28522 14155 28525
rect 12820 28520 14155 28522
rect 12820 28464 14094 28520
rect 14150 28464 14155 28520
rect 12820 28462 14155 28464
rect 12820 28460 12826 28462
rect 14089 28459 14155 28462
rect 20486 28462 21282 28522
rect 20486 28389 20546 28462
rect 12433 28386 12499 28389
rect 13537 28386 13603 28389
rect 12433 28384 13140 28386
rect 12433 28328 12438 28384
rect 12494 28328 13140 28384
rect 12433 28326 13140 28328
rect 12433 28323 12499 28326
rect -300 28112 3851 28114
rect -300 28056 3790 28112
rect 3846 28056 3851 28112
rect -300 28054 3851 28056
rect -300 28024 160 28054
rect 3785 28051 3851 28054
rect 5022 28052 5028 28116
rect 5092 28114 5136 28116
rect 5901 28114 5967 28117
rect 5092 28112 5967 28114
rect 5092 28056 5906 28112
rect 5962 28056 5967 28112
rect 5092 28054 5967 28056
rect 5092 28052 5098 28054
rect 5901 28051 5967 28054
rect 11789 28112 11855 28117
rect 11789 28056 11794 28112
rect 11850 28056 11855 28112
rect 11789 28051 11855 28056
rect 289 27978 355 27981
rect 2221 27978 2287 27981
rect 2630 27978 2636 27980
rect 289 27976 1548 27978
rect 289 27920 294 27976
rect 350 27920 1548 27976
rect 289 27918 1548 27920
rect 289 27915 355 27918
rect -300 27842 160 27872
rect 1301 27842 1367 27845
rect -300 27840 1367 27842
rect -300 27784 1306 27840
rect 1362 27784 1367 27840
rect -300 27782 1367 27784
rect 1488 27842 1548 27918
rect 2221 27976 2636 27978
rect 2221 27920 2226 27976
rect 2282 27920 2636 27976
rect 2221 27918 2636 27920
rect 2221 27915 2287 27918
rect 2630 27916 2636 27918
rect 2700 27916 2706 27980
rect 3049 27978 3115 27981
rect 12893 27978 12959 27981
rect 3049 27976 12959 27978
rect 3049 27920 3054 27976
rect 3110 27920 12898 27976
rect 12954 27920 12959 27976
rect 3049 27918 12959 27920
rect 13080 27978 13140 28326
rect 13537 28384 15210 28386
rect 13537 28328 13542 28384
rect 13598 28328 15210 28384
rect 13537 28326 15210 28328
rect 13537 28323 13603 28326
rect 15150 28252 15210 28326
rect 20437 28384 20546 28389
rect 20437 28328 20442 28384
rect 20498 28328 20546 28384
rect 20437 28326 20546 28328
rect 21222 28386 21282 28462
rect 21840 28386 22300 28416
rect 21222 28326 22300 28386
rect 20437 28323 20503 28326
rect 15780 28320 16096 28321
rect 15780 28256 15786 28320
rect 15850 28256 15866 28320
rect 15930 28256 15946 28320
rect 16010 28256 16026 28320
rect 16090 28256 16096 28320
rect 15780 28255 16096 28256
rect 20725 28320 21041 28321
rect 20725 28256 20731 28320
rect 20795 28256 20811 28320
rect 20875 28256 20891 28320
rect 20955 28256 20971 28320
rect 21035 28256 21041 28320
rect 21840 28296 22300 28326
rect 20725 28255 21041 28256
rect 15142 28188 15148 28252
rect 15212 28188 15218 28252
rect 19241 28250 19307 28253
rect 19374 28250 19380 28252
rect 19241 28248 19380 28250
rect 19241 28192 19246 28248
rect 19302 28192 19380 28248
rect 19241 28190 19380 28192
rect 19241 28187 19307 28190
rect 19374 28188 19380 28190
rect 19444 28188 19450 28252
rect 13813 28114 13879 28117
rect 17769 28114 17835 28117
rect 13813 28112 17835 28114
rect 13813 28056 13818 28112
rect 13874 28056 17774 28112
rect 17830 28056 17835 28112
rect 13813 28054 17835 28056
rect 13813 28051 13879 28054
rect 17769 28051 17835 28054
rect 19241 28114 19307 28117
rect 21817 28114 21883 28117
rect 19241 28112 21883 28114
rect 19241 28056 19246 28112
rect 19302 28056 21822 28112
rect 21878 28056 21883 28112
rect 19241 28054 21883 28056
rect 19241 28051 19307 28054
rect 21817 28051 21883 28054
rect 13080 27918 18890 27978
rect 3049 27915 3115 27918
rect 12893 27915 12959 27918
rect 2262 27842 2268 27844
rect 1488 27782 2268 27842
rect -300 27752 160 27782
rect 1301 27779 1367 27782
rect 2262 27780 2268 27782
rect 2332 27780 2338 27844
rect 2446 27780 2452 27844
rect 2516 27842 2522 27844
rect 3049 27842 3115 27845
rect 2516 27840 3115 27842
rect 2516 27784 3054 27840
rect 3110 27784 3115 27840
rect 2516 27782 3115 27784
rect 2516 27780 2522 27782
rect 3049 27779 3115 27782
rect 3418 27776 3734 27777
rect 3418 27712 3424 27776
rect 3488 27712 3504 27776
rect 3568 27712 3584 27776
rect 3648 27712 3664 27776
rect 3728 27712 3734 27776
rect 3418 27711 3734 27712
rect 8363 27776 8679 27777
rect 8363 27712 8369 27776
rect 8433 27712 8449 27776
rect 8513 27712 8529 27776
rect 8593 27712 8609 27776
rect 8673 27712 8679 27776
rect 8363 27711 8679 27712
rect 13308 27776 13624 27777
rect 13308 27712 13314 27776
rect 13378 27712 13394 27776
rect 13458 27712 13474 27776
rect 13538 27712 13554 27776
rect 13618 27712 13624 27776
rect 13308 27711 13624 27712
rect 18253 27776 18569 27777
rect 18253 27712 18259 27776
rect 18323 27712 18339 27776
rect 18403 27712 18419 27776
rect 18483 27712 18499 27776
rect 18563 27712 18569 27776
rect 18253 27711 18569 27712
rect 2037 27706 2103 27709
rect 3969 27708 4035 27709
rect 2998 27706 3004 27708
rect 2037 27704 3004 27706
rect 2037 27648 2042 27704
rect 2098 27648 3004 27704
rect 2037 27646 3004 27648
rect 2037 27643 2103 27646
rect 2998 27644 3004 27646
rect 3068 27644 3074 27708
rect 3918 27706 3924 27708
rect 3878 27646 3924 27706
rect 3988 27704 4035 27708
rect 4030 27648 4035 27704
rect 3918 27644 3924 27646
rect 3988 27644 4035 27648
rect 3969 27643 4035 27644
rect 6361 27706 6427 27709
rect 7189 27706 7255 27709
rect 6361 27704 7255 27706
rect 6361 27648 6366 27704
rect 6422 27648 7194 27704
rect 7250 27648 7255 27704
rect 6361 27646 7255 27648
rect 6361 27643 6427 27646
rect 7189 27643 7255 27646
rect 12341 27706 12407 27709
rect 13077 27706 13143 27709
rect 12341 27704 13143 27706
rect 12341 27648 12346 27704
rect 12402 27648 13082 27704
rect 13138 27648 13143 27704
rect 12341 27646 13143 27648
rect 12341 27643 12407 27646
rect 13077 27643 13143 27646
rect 14958 27644 14964 27708
rect 15028 27706 15034 27708
rect 15653 27706 15719 27709
rect 15028 27704 15719 27706
rect 15028 27648 15658 27704
rect 15714 27648 15719 27704
rect 15028 27646 15719 27648
rect 15028 27644 15034 27646
rect 15653 27643 15719 27646
rect -300 27570 160 27600
rect 3233 27570 3299 27573
rect -300 27568 3299 27570
rect -300 27512 3238 27568
rect 3294 27512 3299 27568
rect -300 27510 3299 27512
rect -300 27480 160 27510
rect 3233 27507 3299 27510
rect 3969 27570 4035 27573
rect 4102 27570 4108 27572
rect 3969 27568 4108 27570
rect 3969 27512 3974 27568
rect 4030 27512 4108 27568
rect 3969 27510 4108 27512
rect 3969 27507 4035 27510
rect 4102 27508 4108 27510
rect 4172 27508 4178 27572
rect 13905 27570 13971 27573
rect 12390 27568 13971 27570
rect 12390 27512 13910 27568
rect 13966 27512 13971 27568
rect 12390 27510 13971 27512
rect 18830 27570 18890 27918
rect 20437 27842 20503 27845
rect 21840 27842 22300 27872
rect 20437 27840 22300 27842
rect 20437 27784 20442 27840
rect 20498 27784 22300 27840
rect 20437 27782 22300 27784
rect 20437 27779 20503 27782
rect 21840 27752 22300 27782
rect 19190 27644 19196 27708
rect 19260 27706 19266 27708
rect 19701 27706 19767 27709
rect 19260 27704 19767 27706
rect 19260 27648 19706 27704
rect 19762 27648 19767 27704
rect 19260 27646 19767 27648
rect 19260 27644 19266 27646
rect 19701 27643 19767 27646
rect 20621 27570 20687 27573
rect 18830 27568 20687 27570
rect 18830 27512 20626 27568
rect 20682 27512 20687 27568
rect 18830 27510 20687 27512
rect 289 27434 355 27437
rect 1342 27434 1348 27436
rect 289 27432 1348 27434
rect 289 27376 294 27432
rect 350 27376 1348 27432
rect 289 27374 1348 27376
rect 289 27371 355 27374
rect 1342 27372 1348 27374
rect 1412 27372 1418 27436
rect 3693 27434 3759 27437
rect 12390 27434 12450 27510
rect 13905 27507 13971 27510
rect 20621 27507 20687 27510
rect 3693 27432 12450 27434
rect 3693 27376 3698 27432
rect 3754 27376 12450 27432
rect 3693 27374 12450 27376
rect 3693 27371 3759 27374
rect -300 27298 160 27328
rect 1301 27298 1367 27301
rect -300 27296 1367 27298
rect -300 27240 1306 27296
rect 1362 27240 1367 27296
rect -300 27238 1367 27240
rect -300 27208 160 27238
rect 1301 27235 1367 27238
rect 3325 27298 3391 27301
rect 4286 27298 4292 27300
rect 3325 27296 4292 27298
rect 3325 27240 3330 27296
rect 3386 27240 4292 27296
rect 3325 27238 4292 27240
rect 3325 27235 3391 27238
rect 4286 27236 4292 27238
rect 4356 27236 4362 27300
rect 21265 27298 21331 27301
rect 21840 27298 22300 27328
rect 21265 27296 22300 27298
rect 21265 27240 21270 27296
rect 21326 27240 22300 27296
rect 21265 27238 22300 27240
rect 21265 27235 21331 27238
rect 5890 27232 6206 27233
rect 5890 27168 5896 27232
rect 5960 27168 5976 27232
rect 6040 27168 6056 27232
rect 6120 27168 6136 27232
rect 6200 27168 6206 27232
rect 5890 27167 6206 27168
rect 10835 27232 11151 27233
rect 10835 27168 10841 27232
rect 10905 27168 10921 27232
rect 10985 27168 11001 27232
rect 11065 27168 11081 27232
rect 11145 27168 11151 27232
rect 10835 27167 11151 27168
rect 15780 27232 16096 27233
rect 15780 27168 15786 27232
rect 15850 27168 15866 27232
rect 15930 27168 15946 27232
rect 16010 27168 16026 27232
rect 16090 27168 16096 27232
rect 15780 27167 16096 27168
rect 20725 27232 21041 27233
rect 20725 27168 20731 27232
rect 20795 27168 20811 27232
rect 20875 27168 20891 27232
rect 20955 27168 20971 27232
rect 21035 27168 21041 27232
rect 21840 27208 22300 27238
rect 20725 27167 21041 27168
rect 1710 27100 1716 27164
rect 1780 27162 1786 27164
rect 2405 27162 2471 27165
rect 3141 27162 3207 27165
rect 6729 27162 6795 27165
rect 9622 27162 9628 27164
rect 1780 27160 2790 27162
rect 1780 27104 2410 27160
rect 2466 27104 2790 27160
rect 1780 27102 2790 27104
rect 1780 27100 1786 27102
rect 2405 27099 2471 27102
rect -300 27026 160 27056
rect 1117 27026 1183 27029
rect -300 27024 1183 27026
rect -300 26968 1122 27024
rect 1178 26968 1183 27024
rect -300 26966 1183 26968
rect -300 26936 160 26966
rect 1117 26963 1183 26966
rect 2730 26890 2790 27102
rect 3141 27160 4492 27162
rect 3141 27104 3146 27160
rect 3202 27104 4492 27160
rect 3141 27102 4492 27104
rect 3141 27099 3207 27102
rect 3601 27026 3667 27029
rect 4245 27026 4311 27029
rect 3601 27024 4311 27026
rect 3601 26968 3606 27024
rect 3662 26968 4250 27024
rect 4306 26968 4311 27024
rect 3601 26966 4311 26968
rect 4432 27026 4492 27102
rect 6729 27160 9628 27162
rect 6729 27104 6734 27160
rect 6790 27104 9628 27160
rect 6729 27102 9628 27104
rect 6729 27099 6795 27102
rect 9622 27100 9628 27102
rect 9692 27100 9698 27164
rect 7281 27026 7347 27029
rect 8201 27028 8267 27029
rect 8150 27026 8156 27028
rect 4432 27024 7347 27026
rect 4432 26968 7286 27024
rect 7342 26968 7347 27024
rect 4432 26966 7347 26968
rect 8110 26966 8156 27026
rect 8220 27026 8267 27028
rect 9121 27026 9187 27029
rect 8220 27024 9187 27026
rect 8262 26968 9126 27024
rect 9182 26968 9187 27024
rect 3601 26963 3667 26966
rect 4245 26963 4311 26966
rect 7281 26963 7347 26966
rect 8150 26964 8156 26966
rect 8220 26966 9187 26968
rect 8220 26964 8267 26966
rect 8201 26963 8267 26964
rect 9121 26963 9187 26966
rect 9806 26964 9812 27028
rect 9876 27026 9882 27028
rect 10961 27026 11027 27029
rect 12341 27028 12407 27029
rect 12341 27026 12388 27028
rect 9876 27024 11027 27026
rect 9876 26968 10966 27024
rect 11022 26968 11027 27024
rect 9876 26966 11027 26968
rect 12296 27024 12388 27026
rect 12296 26968 12346 27024
rect 12296 26966 12388 26968
rect 9876 26964 9882 26966
rect 10961 26963 11027 26966
rect 12341 26964 12388 26966
rect 12452 26964 12458 27028
rect 17718 26964 17724 27028
rect 17788 27026 17794 27028
rect 18597 27026 18663 27029
rect 17788 27024 18663 27026
rect 17788 26968 18602 27024
rect 18658 26968 18663 27024
rect 17788 26966 18663 26968
rect 17788 26964 17794 26966
rect 12341 26963 12407 26964
rect 18597 26963 18663 26966
rect 4705 26890 4771 26893
rect 2730 26888 4771 26890
rect 2730 26832 4710 26888
rect 4766 26832 4771 26888
rect 2730 26830 4771 26832
rect 4705 26827 4771 26830
rect 5349 26890 5415 26893
rect 18873 26890 18939 26893
rect 5349 26888 18939 26890
rect 5349 26832 5354 26888
rect 5410 26832 18878 26888
rect 18934 26832 18939 26888
rect 5349 26830 18939 26832
rect 5349 26827 5415 26830
rect 18873 26827 18939 26830
rect -300 26754 160 26784
rect 1301 26754 1367 26757
rect -300 26752 1367 26754
rect -300 26696 1306 26752
rect 1362 26696 1367 26752
rect -300 26694 1367 26696
rect -300 26664 160 26694
rect 1301 26691 1367 26694
rect 11789 26754 11855 26757
rect 12341 26754 12407 26757
rect 11789 26752 12407 26754
rect 11789 26696 11794 26752
rect 11850 26696 12346 26752
rect 12402 26696 12407 26752
rect 11789 26694 12407 26696
rect 11789 26691 11855 26694
rect 12341 26691 12407 26694
rect 14733 26754 14799 26757
rect 17309 26754 17375 26757
rect 14733 26752 17375 26754
rect 14733 26696 14738 26752
rect 14794 26696 17314 26752
rect 17370 26696 17375 26752
rect 14733 26694 17375 26696
rect 14733 26691 14799 26694
rect 17309 26691 17375 26694
rect 20529 26754 20595 26757
rect 21840 26754 22300 26784
rect 20529 26752 22300 26754
rect 20529 26696 20534 26752
rect 20590 26696 22300 26752
rect 20529 26694 22300 26696
rect 20529 26691 20595 26694
rect 3418 26688 3734 26689
rect 3418 26624 3424 26688
rect 3488 26624 3504 26688
rect 3568 26624 3584 26688
rect 3648 26624 3664 26688
rect 3728 26624 3734 26688
rect 3418 26623 3734 26624
rect 8363 26688 8679 26689
rect 8363 26624 8369 26688
rect 8433 26624 8449 26688
rect 8513 26624 8529 26688
rect 8593 26624 8609 26688
rect 8673 26624 8679 26688
rect 8363 26623 8679 26624
rect 13308 26688 13624 26689
rect 13308 26624 13314 26688
rect 13378 26624 13394 26688
rect 13458 26624 13474 26688
rect 13538 26624 13554 26688
rect 13618 26624 13624 26688
rect 13308 26623 13624 26624
rect 18253 26688 18569 26689
rect 18253 26624 18259 26688
rect 18323 26624 18339 26688
rect 18403 26624 18419 26688
rect 18483 26624 18499 26688
rect 18563 26624 18569 26688
rect 21840 26664 22300 26694
rect 18253 26623 18569 26624
rect 9806 26556 9812 26620
rect 9876 26618 9882 26620
rect 12157 26618 12223 26621
rect 9876 26616 12223 26618
rect 9876 26560 12162 26616
rect 12218 26560 12223 26616
rect 9876 26558 12223 26560
rect 9876 26556 9882 26558
rect 12157 26555 12223 26558
rect 12893 26618 12959 26621
rect 13118 26618 13124 26620
rect 12893 26616 13124 26618
rect 12893 26560 12898 26616
rect 12954 26560 13124 26616
rect 12893 26558 13124 26560
rect 12893 26555 12959 26558
rect 13118 26556 13124 26558
rect 13188 26556 13194 26620
rect 16614 26556 16620 26620
rect 16684 26618 16690 26620
rect 16849 26618 16915 26621
rect 16684 26616 16915 26618
rect 16684 26560 16854 26616
rect 16910 26560 16915 26616
rect 16684 26558 16915 26560
rect 16684 26556 16690 26558
rect 16849 26555 16915 26558
rect -300 26482 160 26512
rect 1209 26482 1275 26485
rect -300 26480 1275 26482
rect -300 26424 1214 26480
rect 1270 26424 1275 26480
rect -300 26422 1275 26424
rect -300 26392 160 26422
rect 1209 26419 1275 26422
rect 1761 26482 1827 26485
rect 19333 26482 19399 26485
rect 20253 26482 20319 26485
rect 1761 26480 14106 26482
rect 1761 26424 1766 26480
rect 1822 26424 14106 26480
rect 1761 26422 14106 26424
rect 1761 26419 1827 26422
rect 1209 26346 1275 26349
rect 3049 26346 3115 26349
rect 1209 26344 3115 26346
rect 1209 26288 1214 26344
rect 1270 26288 3054 26344
rect 3110 26288 3115 26344
rect 1209 26286 3115 26288
rect 1209 26283 1275 26286
rect 3049 26283 3115 26286
rect 4102 26284 4108 26348
rect 4172 26346 4178 26348
rect 4981 26346 5047 26349
rect 8109 26346 8175 26349
rect 4172 26344 8175 26346
rect 4172 26288 4986 26344
rect 5042 26288 8114 26344
rect 8170 26288 8175 26344
rect 4172 26286 8175 26288
rect 4172 26284 4178 26286
rect 4981 26283 5047 26286
rect 8109 26283 8175 26286
rect 8569 26346 8635 26349
rect 9949 26346 10015 26349
rect 8569 26344 10015 26346
rect 8569 26288 8574 26344
rect 8630 26288 9954 26344
rect 10010 26288 10015 26344
rect 8569 26286 10015 26288
rect 8569 26283 8635 26286
rect 9949 26283 10015 26286
rect 11973 26346 12039 26349
rect 11973 26344 12818 26346
rect 11973 26288 11978 26344
rect 12034 26288 12818 26344
rect 11973 26286 12818 26288
rect 11973 26283 12039 26286
rect -300 26210 160 26240
rect 3601 26210 3667 26213
rect -300 26208 3667 26210
rect -300 26152 3606 26208
rect 3662 26152 3667 26208
rect -300 26150 3667 26152
rect -300 26120 160 26150
rect 3601 26147 3667 26150
rect 6269 26210 6335 26213
rect 6862 26210 6868 26212
rect 6269 26208 6868 26210
rect 6269 26152 6274 26208
rect 6330 26152 6868 26208
rect 6269 26150 6868 26152
rect 6269 26147 6335 26150
rect 6862 26148 6868 26150
rect 6932 26148 6938 26212
rect 7833 26210 7899 26213
rect 10317 26210 10383 26213
rect 7833 26208 10383 26210
rect 7833 26152 7838 26208
rect 7894 26152 10322 26208
rect 10378 26152 10383 26208
rect 7833 26150 10383 26152
rect 7833 26147 7899 26150
rect 10317 26147 10383 26150
rect 11421 26210 11487 26213
rect 11646 26210 11652 26212
rect 11421 26208 11652 26210
rect 11421 26152 11426 26208
rect 11482 26152 11652 26208
rect 11421 26150 11652 26152
rect 11421 26147 11487 26150
rect 11646 26148 11652 26150
rect 11716 26148 11722 26212
rect 5890 26144 6206 26145
rect 5890 26080 5896 26144
rect 5960 26080 5976 26144
rect 6040 26080 6056 26144
rect 6120 26080 6136 26144
rect 6200 26080 6206 26144
rect 5890 26079 6206 26080
rect 10835 26144 11151 26145
rect 10835 26080 10841 26144
rect 10905 26080 10921 26144
rect 10985 26080 11001 26144
rect 11065 26080 11081 26144
rect 11145 26080 11151 26144
rect 10835 26079 11151 26080
rect 1945 26074 2011 26077
rect 6913 26074 6979 26077
rect 1945 26072 5596 26074
rect 1945 26016 1950 26072
rect 2006 26016 5596 26072
rect 1945 26014 5596 26016
rect 1945 26011 2011 26014
rect -300 25938 160 25968
rect 3141 25938 3207 25941
rect -300 25936 3207 25938
rect -300 25880 3146 25936
rect 3202 25880 3207 25936
rect -300 25878 3207 25880
rect -300 25848 160 25878
rect 3141 25875 3207 25878
rect 5165 25938 5231 25941
rect 5390 25938 5396 25940
rect 5165 25936 5396 25938
rect 5165 25880 5170 25936
rect 5226 25880 5396 25936
rect 5165 25878 5396 25880
rect 5165 25875 5231 25878
rect 5390 25876 5396 25878
rect 5460 25876 5466 25940
rect 5536 25938 5596 26014
rect 6272 26072 6979 26074
rect 6272 26016 6918 26072
rect 6974 26016 6979 26072
rect 6272 26014 6979 26016
rect 6272 25938 6332 26014
rect 6913 26011 6979 26014
rect 9857 26074 9923 26077
rect 10133 26074 10199 26077
rect 9857 26072 10199 26074
rect 9857 26016 9862 26072
rect 9918 26016 10138 26072
rect 10194 26016 10199 26072
rect 9857 26014 10199 26016
rect 12758 26074 12818 26286
rect 12758 26014 13968 26074
rect 9857 26011 9923 26014
rect 10133 26011 10199 26014
rect 13908 25941 13968 26014
rect 7281 25938 7347 25941
rect 12709 25938 12775 25941
rect 13537 25938 13603 25941
rect 5536 25878 6332 25938
rect 6686 25936 10794 25938
rect 6686 25880 7286 25936
rect 7342 25880 10794 25936
rect 6686 25878 10794 25880
rect 1393 25802 1459 25805
rect 752 25800 1459 25802
rect 752 25744 1398 25800
rect 1454 25744 1459 25800
rect 752 25742 1459 25744
rect -300 25666 160 25696
rect 752 25666 812 25742
rect 1393 25739 1459 25742
rect 2998 25740 3004 25804
rect 3068 25802 3074 25804
rect 3693 25802 3759 25805
rect 4245 25802 4311 25805
rect 6494 25802 6500 25804
rect 3068 25800 3986 25802
rect 3068 25744 3698 25800
rect 3754 25744 3986 25800
rect 3068 25742 3986 25744
rect 3068 25740 3074 25742
rect 3693 25739 3759 25742
rect -300 25606 812 25666
rect 1117 25666 1183 25669
rect 2446 25666 2452 25668
rect 1117 25664 2452 25666
rect 1117 25608 1122 25664
rect 1178 25608 2452 25664
rect 1117 25606 2452 25608
rect -300 25576 160 25606
rect 1117 25603 1183 25606
rect 2446 25604 2452 25606
rect 2516 25604 2522 25668
rect 3926 25666 3986 25742
rect 4245 25800 6500 25802
rect 4245 25744 4250 25800
rect 4306 25744 6500 25800
rect 4245 25742 6500 25744
rect 4245 25739 4311 25742
rect 6494 25740 6500 25742
rect 6564 25740 6570 25804
rect 6686 25666 6746 25878
rect 7281 25875 7347 25878
rect 7557 25802 7623 25805
rect 10041 25802 10107 25805
rect 7557 25800 10107 25802
rect 7557 25744 7562 25800
rect 7618 25744 10046 25800
rect 10102 25744 10107 25800
rect 7557 25742 10107 25744
rect 10734 25802 10794 25878
rect 12709 25936 13603 25938
rect 12709 25880 12714 25936
rect 12770 25880 13542 25936
rect 13598 25880 13603 25936
rect 12709 25878 13603 25880
rect 12709 25875 12775 25878
rect 13537 25875 13603 25878
rect 13905 25936 13971 25941
rect 13905 25880 13910 25936
rect 13966 25880 13971 25936
rect 13905 25875 13971 25880
rect 14046 25938 14106 26422
rect 19333 26480 20319 26482
rect 19333 26424 19338 26480
rect 19394 26424 20258 26480
rect 20314 26424 20319 26480
rect 19333 26422 20319 26424
rect 19333 26419 19399 26422
rect 20253 26419 20319 26422
rect 16205 26210 16271 26213
rect 19057 26210 19123 26213
rect 16205 26208 19123 26210
rect 16205 26152 16210 26208
rect 16266 26152 19062 26208
rect 19118 26152 19123 26208
rect 16205 26150 19123 26152
rect 16205 26147 16271 26150
rect 19057 26147 19123 26150
rect 21265 26210 21331 26213
rect 21840 26210 22300 26240
rect 21265 26208 22300 26210
rect 21265 26152 21270 26208
rect 21326 26152 22300 26208
rect 21265 26150 22300 26152
rect 21265 26147 21331 26150
rect 15780 26144 16096 26145
rect 15780 26080 15786 26144
rect 15850 26080 15866 26144
rect 15930 26080 15946 26144
rect 16010 26080 16026 26144
rect 16090 26080 16096 26144
rect 15780 26079 16096 26080
rect 20725 26144 21041 26145
rect 20725 26080 20731 26144
rect 20795 26080 20811 26144
rect 20875 26080 20891 26144
rect 20955 26080 20971 26144
rect 21035 26080 21041 26144
rect 21840 26120 22300 26150
rect 20725 26079 21041 26080
rect 14181 25938 14247 25941
rect 18505 25938 18571 25941
rect 14046 25936 18571 25938
rect 14046 25880 14186 25936
rect 14242 25880 18510 25936
rect 18566 25880 18571 25936
rect 14046 25878 18571 25880
rect 14181 25875 14247 25878
rect 18505 25875 18571 25878
rect 11329 25802 11395 25805
rect 10734 25800 11395 25802
rect 10734 25744 11334 25800
rect 11390 25744 11395 25800
rect 10734 25742 11395 25744
rect 7557 25739 7623 25742
rect 10041 25739 10107 25742
rect 11329 25739 11395 25742
rect 13537 25802 13603 25805
rect 13537 25800 16682 25802
rect 13537 25744 13542 25800
rect 13598 25744 16682 25800
rect 13537 25742 16682 25744
rect 13537 25739 13603 25742
rect 3926 25606 6746 25666
rect 12065 25666 12131 25669
rect 12709 25666 12775 25669
rect 12065 25664 12775 25666
rect 12065 25608 12070 25664
rect 12126 25608 12714 25664
rect 12770 25608 12775 25664
rect 12065 25606 12775 25608
rect 12065 25603 12131 25606
rect 12709 25603 12775 25606
rect 3418 25600 3734 25601
rect 3418 25536 3424 25600
rect 3488 25536 3504 25600
rect 3568 25536 3584 25600
rect 3648 25536 3664 25600
rect 3728 25536 3734 25600
rect 3418 25535 3734 25536
rect 8363 25600 8679 25601
rect 8363 25536 8369 25600
rect 8433 25536 8449 25600
rect 8513 25536 8529 25600
rect 8593 25536 8609 25600
rect 8673 25536 8679 25600
rect 8363 25535 8679 25536
rect 13308 25600 13624 25601
rect 13308 25536 13314 25600
rect 13378 25536 13394 25600
rect 13458 25536 13474 25600
rect 13538 25536 13554 25600
rect 13618 25536 13624 25600
rect 13308 25535 13624 25536
rect 790 25468 796 25532
rect 860 25530 866 25532
rect 1117 25530 1183 25533
rect 860 25528 1183 25530
rect 860 25472 1122 25528
rect 1178 25472 1183 25528
rect 860 25470 1183 25472
rect 860 25468 866 25470
rect 1117 25467 1183 25470
rect 1485 25530 1551 25533
rect 4245 25530 4311 25533
rect 5022 25530 5028 25532
rect 1485 25528 3296 25530
rect 1485 25472 1490 25528
rect 1546 25472 3296 25528
rect 1485 25470 3296 25472
rect 1485 25467 1551 25470
rect -300 25394 160 25424
rect 1209 25394 1275 25397
rect 2865 25396 2931 25397
rect -300 25392 1275 25394
rect -300 25336 1214 25392
rect 1270 25336 1275 25392
rect -300 25334 1275 25336
rect -300 25304 160 25334
rect 1209 25331 1275 25334
rect 2814 25332 2820 25396
rect 2884 25394 2931 25396
rect 3236 25394 3296 25470
rect 4245 25528 5028 25530
rect 4245 25472 4250 25528
rect 4306 25472 5028 25528
rect 4245 25470 5028 25472
rect 4245 25467 4311 25470
rect 5022 25468 5028 25470
rect 5092 25530 5098 25532
rect 6729 25530 6795 25533
rect 5092 25528 6795 25530
rect 5092 25472 6734 25528
rect 6790 25472 6795 25528
rect 5092 25470 6795 25472
rect 5092 25468 5098 25470
rect 6729 25467 6795 25470
rect 9029 25530 9095 25533
rect 9254 25530 9260 25532
rect 9029 25528 9260 25530
rect 9029 25472 9034 25528
rect 9090 25472 9260 25528
rect 9029 25470 9260 25472
rect 9029 25467 9095 25470
rect 9254 25468 9260 25470
rect 9324 25468 9330 25532
rect 9622 25468 9628 25532
rect 9692 25530 9698 25532
rect 11513 25530 11579 25533
rect 9692 25528 11579 25530
rect 9692 25472 11518 25528
rect 11574 25472 11579 25528
rect 9692 25470 11579 25472
rect 9692 25468 9698 25470
rect 11513 25467 11579 25470
rect 4153 25394 4219 25397
rect 10133 25394 10199 25397
rect 2884 25392 2976 25394
rect 2926 25336 2976 25392
rect 2884 25334 2976 25336
rect 3236 25392 4219 25394
rect 3236 25336 4158 25392
rect 4214 25336 4219 25392
rect 3236 25334 4219 25336
rect 2884 25332 2931 25334
rect 2865 25331 2931 25332
rect 4153 25331 4219 25334
rect 5030 25392 10199 25394
rect 5030 25336 10138 25392
rect 10194 25336 10199 25392
rect 5030 25334 10199 25336
rect 1853 25258 1919 25261
rect 5030 25258 5090 25334
rect 10133 25331 10199 25334
rect 10501 25394 10567 25397
rect 10501 25392 16498 25394
rect 10501 25336 10506 25392
rect 10562 25336 16498 25392
rect 10501 25334 16498 25336
rect 10501 25331 10567 25334
rect 1853 25256 5090 25258
rect 1853 25200 1858 25256
rect 1914 25200 5090 25256
rect 1853 25198 5090 25200
rect 5257 25258 5323 25261
rect 16205 25258 16271 25261
rect 5257 25256 16271 25258
rect 5257 25200 5262 25256
rect 5318 25200 16210 25256
rect 16266 25200 16271 25256
rect 5257 25198 16271 25200
rect 1853 25195 1919 25198
rect 5257 25195 5323 25198
rect 16205 25195 16271 25198
rect -300 25122 160 25152
rect 1301 25122 1367 25125
rect -300 25120 1367 25122
rect -300 25064 1306 25120
rect 1362 25064 1367 25120
rect -300 25062 1367 25064
rect -300 25032 160 25062
rect 1301 25059 1367 25062
rect 7833 25122 7899 25125
rect 9305 25122 9371 25125
rect 7833 25120 9371 25122
rect 7833 25064 7838 25120
rect 7894 25064 9310 25120
rect 9366 25064 9371 25120
rect 7833 25062 9371 25064
rect 7833 25059 7899 25062
rect 9305 25059 9371 25062
rect 9765 25122 9831 25125
rect 9765 25120 9874 25122
rect 9765 25064 9770 25120
rect 9826 25064 9874 25120
rect 9765 25059 9874 25064
rect 12934 25060 12940 25124
rect 13004 25122 13010 25124
rect 14457 25122 14523 25125
rect 15561 25124 15627 25125
rect 13004 25120 14523 25122
rect 13004 25064 14462 25120
rect 14518 25064 14523 25120
rect 13004 25062 14523 25064
rect 13004 25060 13010 25062
rect 14457 25059 14523 25062
rect 15510 25060 15516 25124
rect 15580 25122 15627 25124
rect 15580 25120 15672 25122
rect 15622 25064 15672 25120
rect 15580 25062 15672 25064
rect 15580 25060 15627 25062
rect 15561 25059 15627 25060
rect 5890 25056 6206 25057
rect 5890 24992 5896 25056
rect 5960 24992 5976 25056
rect 6040 24992 6056 25056
rect 6120 24992 6136 25056
rect 6200 24992 6206 25056
rect 5890 24991 6206 24992
rect 2129 24986 2195 24989
rect 2681 24986 2747 24989
rect 7741 24986 7807 24989
rect 2129 24984 2330 24986
rect 2129 24928 2134 24984
rect 2190 24928 2330 24984
rect 2129 24926 2330 24928
rect 2129 24923 2195 24926
rect -300 24850 160 24880
rect 749 24850 815 24853
rect -300 24848 815 24850
rect -300 24792 754 24848
rect 810 24792 815 24848
rect -300 24790 815 24792
rect 2270 24850 2330 24926
rect 2681 24984 5826 24986
rect 2681 24928 2686 24984
rect 2742 24928 5826 24984
rect 2681 24926 5826 24928
rect 2681 24923 2747 24926
rect 5533 24850 5599 24853
rect 2270 24848 5599 24850
rect 2270 24792 5538 24848
rect 5594 24792 5599 24848
rect 2270 24790 5599 24792
rect 5766 24850 5826 24926
rect 6548 24984 7807 24986
rect 6548 24928 7746 24984
rect 7802 24928 7807 24984
rect 6548 24926 7807 24928
rect 6548 24850 6608 24926
rect 7741 24923 7807 24926
rect 8753 24986 8819 24989
rect 8886 24986 8892 24988
rect 8753 24984 8892 24986
rect 8753 24928 8758 24984
rect 8814 24928 8892 24984
rect 8753 24926 8892 24928
rect 8753 24923 8819 24926
rect 8886 24924 8892 24926
rect 8956 24924 8962 24988
rect 9814 24853 9874 25059
rect 10835 25056 11151 25057
rect 10835 24992 10841 25056
rect 10905 24992 10921 25056
rect 10985 24992 11001 25056
rect 11065 24992 11081 25056
rect 11145 24992 11151 25056
rect 10835 24991 11151 24992
rect 15780 25056 16096 25057
rect 15780 24992 15786 25056
rect 15850 24992 15866 25056
rect 15930 24992 15946 25056
rect 16010 24992 16026 25056
rect 16090 24992 16096 25056
rect 15780 24991 16096 24992
rect 11278 24924 11284 24988
rect 11348 24986 11354 24988
rect 11881 24986 11947 24989
rect 11348 24984 11947 24986
rect 11348 24928 11886 24984
rect 11942 24928 11947 24984
rect 11348 24926 11947 24928
rect 11348 24924 11354 24926
rect 11881 24923 11947 24926
rect 13813 24984 13879 24989
rect 13813 24928 13818 24984
rect 13874 24928 13879 24984
rect 13813 24923 13879 24928
rect 6729 24852 6795 24853
rect 5766 24790 6608 24850
rect -300 24760 160 24790
rect 749 24787 815 24790
rect 5533 24787 5599 24790
rect 6678 24788 6684 24852
rect 6748 24850 6795 24852
rect 6748 24848 6840 24850
rect 6790 24792 6840 24848
rect 6748 24790 6840 24792
rect 9765 24848 9874 24853
rect 9765 24792 9770 24848
rect 9826 24792 9874 24848
rect 9765 24790 9874 24792
rect 10041 24850 10107 24853
rect 10409 24850 10475 24853
rect 10041 24848 10475 24850
rect 10041 24792 10046 24848
rect 10102 24792 10414 24848
rect 10470 24792 10475 24848
rect 10041 24790 10475 24792
rect 6748 24788 6795 24790
rect 6729 24787 6795 24788
rect 9765 24787 9831 24790
rect 10041 24787 10107 24790
rect 10409 24787 10475 24790
rect 11053 24850 11119 24853
rect 13816 24850 13876 24923
rect 11053 24848 13876 24850
rect 11053 24792 11058 24848
rect 11114 24792 13876 24848
rect 11053 24790 13876 24792
rect 16438 24850 16498 25334
rect 16622 25258 16682 25742
rect 19885 25666 19951 25669
rect 21840 25666 22300 25696
rect 19885 25664 22300 25666
rect 19885 25608 19890 25664
rect 19946 25608 22300 25664
rect 19885 25606 22300 25608
rect 19885 25603 19951 25606
rect 18253 25600 18569 25601
rect 18253 25536 18259 25600
rect 18323 25536 18339 25600
rect 18403 25536 18419 25600
rect 18483 25536 18499 25600
rect 18563 25536 18569 25600
rect 21840 25576 22300 25606
rect 18253 25535 18569 25536
rect 20621 25394 20687 25397
rect 20486 25392 20687 25394
rect 20486 25336 20626 25392
rect 20682 25336 20687 25392
rect 20486 25334 20687 25336
rect 16757 25258 16823 25261
rect 17861 25258 17927 25261
rect 16622 25256 17927 25258
rect 16622 25200 16762 25256
rect 16818 25200 17866 25256
rect 17922 25200 17927 25256
rect 16622 25198 17927 25200
rect 20486 25258 20546 25334
rect 20621 25331 20687 25334
rect 20486 25198 21282 25258
rect 16757 25195 16823 25198
rect 17861 25195 17927 25198
rect 19241 25122 19307 25125
rect 19558 25122 19564 25124
rect 19241 25120 19564 25122
rect 19241 25064 19246 25120
rect 19302 25064 19564 25120
rect 19241 25062 19564 25064
rect 19241 25059 19307 25062
rect 19558 25060 19564 25062
rect 19628 25060 19634 25124
rect 21222 25122 21282 25198
rect 21840 25122 22300 25152
rect 21222 25062 22300 25122
rect 20725 25056 21041 25057
rect 20725 24992 20731 25056
rect 20795 24992 20811 25056
rect 20875 24992 20891 25056
rect 20955 24992 20971 25056
rect 21035 24992 21041 25056
rect 21840 25032 22300 25062
rect 20725 24991 21041 24992
rect 16941 24850 17007 24853
rect 16438 24848 17007 24850
rect 16438 24792 16946 24848
rect 17002 24792 17007 24848
rect 16438 24790 17007 24792
rect 11053 24787 11119 24790
rect 16941 24787 17007 24790
rect 19190 24788 19196 24852
rect 19260 24850 19266 24852
rect 19609 24850 19675 24853
rect 19260 24848 19675 24850
rect 19260 24792 19614 24848
rect 19670 24792 19675 24848
rect 19260 24790 19675 24792
rect 19260 24788 19266 24790
rect 19609 24787 19675 24790
rect 2497 24714 2563 24717
rect 12985 24714 13051 24717
rect 2497 24712 13051 24714
rect 2497 24656 2502 24712
rect 2558 24656 12990 24712
rect 13046 24656 13051 24712
rect 2497 24654 13051 24656
rect 2497 24651 2563 24654
rect 12985 24651 13051 24654
rect -300 24578 160 24608
rect 1301 24578 1367 24581
rect -300 24576 1367 24578
rect -300 24520 1306 24576
rect 1362 24520 1367 24576
rect -300 24518 1367 24520
rect -300 24488 160 24518
rect 1301 24515 1367 24518
rect 6310 24516 6316 24580
rect 6380 24578 6386 24580
rect 6453 24578 6519 24581
rect 6380 24576 6519 24578
rect 6380 24520 6458 24576
rect 6514 24520 6519 24576
rect 6380 24518 6519 24520
rect 6380 24516 6386 24518
rect 6453 24515 6519 24518
rect 9622 24516 9628 24580
rect 9692 24578 9698 24580
rect 9949 24578 10015 24581
rect 9692 24576 10015 24578
rect 9692 24520 9954 24576
rect 10010 24520 10015 24576
rect 9692 24518 10015 24520
rect 9692 24516 9698 24518
rect 9949 24515 10015 24518
rect 20253 24578 20319 24581
rect 21840 24578 22300 24608
rect 20253 24576 22300 24578
rect 20253 24520 20258 24576
rect 20314 24520 22300 24576
rect 20253 24518 22300 24520
rect 20253 24515 20319 24518
rect 3418 24512 3734 24513
rect 3418 24448 3424 24512
rect 3488 24448 3504 24512
rect 3568 24448 3584 24512
rect 3648 24448 3664 24512
rect 3728 24448 3734 24512
rect 3418 24447 3734 24448
rect 8363 24512 8679 24513
rect 8363 24448 8369 24512
rect 8433 24448 8449 24512
rect 8513 24448 8529 24512
rect 8593 24448 8609 24512
rect 8673 24448 8679 24512
rect 8363 24447 8679 24448
rect 13308 24512 13624 24513
rect 13308 24448 13314 24512
rect 13378 24448 13394 24512
rect 13458 24448 13474 24512
rect 13538 24448 13554 24512
rect 13618 24448 13624 24512
rect 13308 24447 13624 24448
rect 18253 24512 18569 24513
rect 18253 24448 18259 24512
rect 18323 24448 18339 24512
rect 18403 24448 18419 24512
rect 18483 24448 18499 24512
rect 18563 24448 18569 24512
rect 21840 24488 22300 24518
rect 18253 24447 18569 24448
rect 4153 24442 4219 24445
rect 7649 24442 7715 24445
rect 11881 24442 11947 24445
rect 4153 24440 7715 24442
rect 4153 24384 4158 24440
rect 4214 24384 7654 24440
rect 7710 24384 7715 24440
rect 4153 24382 7715 24384
rect 4153 24379 4219 24382
rect 7649 24379 7715 24382
rect 9630 24440 11947 24442
rect 9630 24384 11886 24440
rect 11942 24384 11947 24440
rect 9630 24382 11947 24384
rect -300 24306 160 24336
rect 1209 24306 1275 24309
rect -300 24304 1275 24306
rect -300 24248 1214 24304
rect 1270 24248 1275 24304
rect -300 24246 1275 24248
rect -300 24216 160 24246
rect 1209 24243 1275 24246
rect 2497 24306 2563 24309
rect 4613 24308 4679 24309
rect 4102 24306 4108 24308
rect 2497 24304 4108 24306
rect 2497 24248 2502 24304
rect 2558 24248 4108 24304
rect 2497 24246 4108 24248
rect 2497 24243 2563 24246
rect 4102 24244 4108 24246
rect 4172 24244 4178 24308
rect 4613 24306 4660 24308
rect 4568 24304 4660 24306
rect 4568 24248 4618 24304
rect 4568 24246 4660 24248
rect 4613 24244 4660 24246
rect 4724 24244 4730 24308
rect 5533 24306 5599 24309
rect 6310 24306 6316 24308
rect 5533 24304 6316 24306
rect 5533 24248 5538 24304
rect 5594 24248 6316 24304
rect 5533 24246 6316 24248
rect 4613 24243 4679 24244
rect 5533 24243 5599 24246
rect 6310 24244 6316 24246
rect 6380 24306 6386 24308
rect 9630 24306 9690 24382
rect 11881 24379 11947 24382
rect 11053 24306 11119 24309
rect 6380 24246 9690 24306
rect 10412 24304 11119 24306
rect 10412 24248 11058 24304
rect 11114 24248 11119 24304
rect 10412 24246 11119 24248
rect 6380 24244 6386 24246
rect 1710 24108 1716 24172
rect 1780 24170 1786 24172
rect 2630 24170 2636 24172
rect 1780 24110 2636 24170
rect 1780 24108 1786 24110
rect 2630 24108 2636 24110
rect 2700 24170 2706 24172
rect 10412 24170 10472 24246
rect 11053 24243 11119 24246
rect 11421 24306 11487 24309
rect 14457 24306 14523 24309
rect 11421 24304 14523 24306
rect 11421 24248 11426 24304
rect 11482 24248 14462 24304
rect 14518 24248 14523 24304
rect 11421 24246 14523 24248
rect 11421 24243 11487 24246
rect 14457 24243 14523 24246
rect 15009 24170 15075 24173
rect 2700 24110 10472 24170
rect 10550 24168 15075 24170
rect 10550 24112 15014 24168
rect 15070 24112 15075 24168
rect 10550 24110 15075 24112
rect 2700 24108 2706 24110
rect -300 24034 160 24064
rect 657 24034 723 24037
rect -300 24032 723 24034
rect -300 23976 662 24032
rect 718 23976 723 24032
rect -300 23974 723 23976
rect -300 23944 160 23974
rect 657 23971 723 23974
rect 1761 24034 1827 24037
rect 5165 24034 5231 24037
rect 1761 24032 5231 24034
rect 1761 23976 1766 24032
rect 1822 23976 5170 24032
rect 5226 23976 5231 24032
rect 1761 23974 5231 23976
rect 1761 23971 1827 23974
rect 5165 23971 5231 23974
rect 8201 24034 8267 24037
rect 10550 24034 10610 24110
rect 15009 24107 15075 24110
rect 15377 24170 15443 24173
rect 16614 24170 16620 24172
rect 15377 24168 16620 24170
rect 15377 24112 15382 24168
rect 15438 24112 16620 24168
rect 15377 24110 16620 24112
rect 15377 24107 15443 24110
rect 16614 24108 16620 24110
rect 16684 24108 16690 24172
rect 20437 24170 20503 24173
rect 20437 24168 21282 24170
rect 20437 24112 20442 24168
rect 20498 24112 21282 24168
rect 20437 24110 21282 24112
rect 20437 24107 20503 24110
rect 8201 24032 10610 24034
rect 8201 23976 8206 24032
rect 8262 23976 10610 24032
rect 8201 23974 10610 23976
rect 12341 24034 12407 24037
rect 12566 24034 12572 24036
rect 12341 24032 12572 24034
rect 12341 23976 12346 24032
rect 12402 23976 12572 24032
rect 12341 23974 12572 23976
rect 8201 23971 8267 23974
rect 12341 23971 12407 23974
rect 12566 23972 12572 23974
rect 12636 23972 12642 24036
rect 21222 24034 21282 24110
rect 21840 24034 22300 24064
rect 21222 23974 22300 24034
rect 5890 23968 6206 23969
rect 5890 23904 5896 23968
rect 5960 23904 5976 23968
rect 6040 23904 6056 23968
rect 6120 23904 6136 23968
rect 6200 23904 6206 23968
rect 5890 23903 6206 23904
rect 10835 23968 11151 23969
rect 10835 23904 10841 23968
rect 10905 23904 10921 23968
rect 10985 23904 11001 23968
rect 11065 23904 11081 23968
rect 11145 23904 11151 23968
rect 10835 23903 11151 23904
rect 15780 23968 16096 23969
rect 15780 23904 15786 23968
rect 15850 23904 15866 23968
rect 15930 23904 15946 23968
rect 16010 23904 16026 23968
rect 16090 23904 16096 23968
rect 15780 23903 16096 23904
rect 20725 23968 21041 23969
rect 20725 23904 20731 23968
rect 20795 23904 20811 23968
rect 20875 23904 20891 23968
rect 20955 23904 20971 23968
rect 21035 23904 21041 23968
rect 21840 23944 22300 23974
rect 20725 23903 21041 23904
rect 5165 23900 5231 23901
rect 1158 23836 1164 23900
rect 1228 23898 1234 23900
rect 5022 23898 5028 23900
rect 1228 23838 5028 23898
rect 1228 23836 1234 23838
rect 5022 23836 5028 23838
rect 5092 23836 5098 23900
rect 5165 23896 5212 23900
rect 5276 23898 5282 23900
rect 7097 23898 7163 23901
rect 7414 23898 7420 23900
rect 5165 23840 5170 23896
rect 5165 23836 5212 23840
rect 5276 23838 5322 23898
rect 7097 23896 7420 23898
rect 7097 23840 7102 23896
rect 7158 23840 7420 23896
rect 7097 23838 7420 23840
rect 5276 23836 5282 23838
rect 5165 23835 5231 23836
rect 7097 23835 7163 23838
rect 7414 23836 7420 23838
rect 7484 23836 7490 23900
rect 9622 23836 9628 23900
rect 9692 23898 9698 23900
rect 9949 23898 10015 23901
rect 12750 23898 12756 23900
rect 9692 23896 10015 23898
rect 9692 23840 9954 23896
rect 10010 23840 10015 23896
rect 9692 23838 10015 23840
rect 9692 23836 9698 23838
rect 9949 23835 10015 23838
rect 11286 23838 12756 23898
rect -300 23762 160 23792
rect 1301 23762 1367 23765
rect -300 23760 1367 23762
rect -300 23704 1306 23760
rect 1362 23704 1367 23760
rect -300 23702 1367 23704
rect -300 23672 160 23702
rect 1301 23699 1367 23702
rect 2129 23762 2195 23765
rect 7465 23762 7531 23765
rect 9806 23762 9812 23764
rect 2129 23760 7531 23762
rect 2129 23704 2134 23760
rect 2190 23704 7470 23760
rect 7526 23704 7531 23760
rect 2129 23702 7531 23704
rect 2129 23699 2195 23702
rect 7465 23699 7531 23702
rect 7606 23702 9812 23762
rect 1301 23626 1367 23629
rect 4838 23626 4844 23628
rect 1301 23624 4844 23626
rect 1301 23568 1306 23624
rect 1362 23568 4844 23624
rect 1301 23566 4844 23568
rect 1301 23563 1367 23566
rect 4838 23564 4844 23566
rect 4908 23564 4914 23628
rect 5206 23564 5212 23628
rect 5276 23626 5282 23628
rect 7606 23626 7666 23702
rect 9806 23700 9812 23702
rect 9876 23700 9882 23764
rect 5276 23566 7666 23626
rect 7925 23626 7991 23629
rect 9213 23628 9279 23629
rect 9213 23626 9260 23628
rect 7925 23624 8954 23626
rect 7925 23568 7930 23624
rect 7986 23568 8954 23624
rect 7925 23566 8954 23568
rect 9168 23624 9260 23626
rect 9168 23568 9218 23624
rect 9168 23566 9260 23568
rect 5276 23564 5282 23566
rect 7925 23563 8034 23566
rect -300 23490 160 23520
rect 749 23490 815 23493
rect -300 23488 815 23490
rect -300 23432 754 23488
rect 810 23432 815 23488
rect -300 23430 815 23432
rect -300 23400 160 23430
rect 749 23427 815 23430
rect 1485 23490 1551 23493
rect 1894 23490 1900 23492
rect 1485 23488 1900 23490
rect 1485 23432 1490 23488
rect 1546 23432 1900 23488
rect 1485 23430 1900 23432
rect 1485 23427 1551 23430
rect 1894 23428 1900 23430
rect 1964 23428 1970 23492
rect 5993 23490 6059 23493
rect 7046 23490 7052 23492
rect 5993 23488 7052 23490
rect 5993 23432 5998 23488
rect 6054 23432 7052 23488
rect 5993 23430 7052 23432
rect 5993 23427 6059 23430
rect 7046 23428 7052 23430
rect 7116 23428 7122 23492
rect 3418 23424 3734 23425
rect 3418 23360 3424 23424
rect 3488 23360 3504 23424
rect 3568 23360 3584 23424
rect 3648 23360 3664 23424
rect 3728 23360 3734 23424
rect 3418 23359 3734 23360
rect 4061 23354 4127 23357
rect 4654 23354 4660 23356
rect 4061 23352 4660 23354
rect 4061 23296 4066 23352
rect 4122 23296 4660 23352
rect 4061 23294 4660 23296
rect 4061 23291 4127 23294
rect 4654 23292 4660 23294
rect 4724 23354 4730 23356
rect 7974 23354 8034 23563
rect 8363 23424 8679 23425
rect 8363 23360 8369 23424
rect 8433 23360 8449 23424
rect 8513 23360 8529 23424
rect 8593 23360 8609 23424
rect 8673 23360 8679 23424
rect 8363 23359 8679 23360
rect 4724 23294 8034 23354
rect 8894 23354 8954 23566
rect 9213 23564 9260 23566
rect 9324 23564 9330 23628
rect 9806 23564 9812 23628
rect 9876 23626 9882 23628
rect 11286 23626 11346 23838
rect 12750 23836 12756 23838
rect 12820 23836 12826 23900
rect 12433 23762 12499 23765
rect 12566 23762 12572 23764
rect 12433 23760 12572 23762
rect 12433 23704 12438 23760
rect 12494 23704 12572 23760
rect 12433 23702 12572 23704
rect 12433 23699 12499 23702
rect 12566 23700 12572 23702
rect 12636 23700 12642 23764
rect 12801 23762 12867 23765
rect 13169 23762 13235 23765
rect 12801 23760 13235 23762
rect 12801 23704 12806 23760
rect 12862 23704 13174 23760
rect 13230 23704 13235 23760
rect 12801 23702 13235 23704
rect 12801 23699 12867 23702
rect 13169 23699 13235 23702
rect 9876 23566 11346 23626
rect 11881 23626 11947 23629
rect 12525 23626 12591 23629
rect 14089 23626 14155 23629
rect 11881 23624 14155 23626
rect 11881 23568 11886 23624
rect 11942 23568 12530 23624
rect 12586 23568 14094 23624
rect 14150 23568 14155 23624
rect 11881 23566 14155 23568
rect 9876 23564 9882 23566
rect 9213 23563 9279 23564
rect 11881 23563 11947 23566
rect 12525 23563 12591 23566
rect 14089 23563 14155 23566
rect 14590 23564 14596 23628
rect 14660 23626 14666 23628
rect 14733 23626 14799 23629
rect 14660 23624 14799 23626
rect 14660 23568 14738 23624
rect 14794 23568 14799 23624
rect 14660 23566 14799 23568
rect 14660 23564 14666 23566
rect 14733 23563 14799 23566
rect 15193 23626 15259 23629
rect 15745 23626 15811 23629
rect 15193 23624 15811 23626
rect 15193 23568 15198 23624
rect 15254 23568 15750 23624
rect 15806 23568 15811 23624
rect 15193 23566 15811 23568
rect 15193 23563 15259 23566
rect 15745 23563 15811 23566
rect 17534 23564 17540 23628
rect 17604 23626 17610 23628
rect 17604 23566 19258 23626
rect 17604 23564 17610 23566
rect 9305 23490 9371 23493
rect 9622 23490 9628 23492
rect 9305 23488 9628 23490
rect 9305 23432 9310 23488
rect 9366 23432 9628 23488
rect 9305 23430 9628 23432
rect 9305 23427 9371 23430
rect 9622 23428 9628 23430
rect 9692 23428 9698 23492
rect 9765 23490 9831 23493
rect 11237 23490 11303 23493
rect 9765 23488 11303 23490
rect 9765 23432 9770 23488
rect 9826 23432 11242 23488
rect 11298 23432 11303 23488
rect 9765 23430 11303 23432
rect 9765 23427 9831 23430
rect 11237 23427 11303 23430
rect 16246 23428 16252 23492
rect 16316 23490 16322 23492
rect 17350 23490 17356 23492
rect 16316 23430 17356 23490
rect 16316 23428 16322 23430
rect 17350 23428 17356 23430
rect 17420 23428 17426 23492
rect 13308 23424 13624 23425
rect 13308 23360 13314 23424
rect 13378 23360 13394 23424
rect 13458 23360 13474 23424
rect 13538 23360 13554 23424
rect 13618 23360 13624 23424
rect 13308 23359 13624 23360
rect 18253 23424 18569 23425
rect 18253 23360 18259 23424
rect 18323 23360 18339 23424
rect 18403 23360 18419 23424
rect 18483 23360 18499 23424
rect 18563 23360 18569 23424
rect 18253 23359 18569 23360
rect 10317 23354 10383 23357
rect 8894 23352 10383 23354
rect 8894 23296 10322 23352
rect 10378 23296 10383 23352
rect 8894 23294 10383 23296
rect 4724 23292 4730 23294
rect 10317 23291 10383 23294
rect 16573 23354 16639 23357
rect 17769 23354 17835 23357
rect 16573 23352 17835 23354
rect 16573 23296 16578 23352
rect 16634 23296 17774 23352
rect 17830 23296 17835 23352
rect 16573 23294 17835 23296
rect 19198 23354 19258 23566
rect 20437 23490 20503 23493
rect 21840 23490 22300 23520
rect 20437 23488 22300 23490
rect 20437 23432 20442 23488
rect 20498 23432 22300 23488
rect 20437 23430 22300 23432
rect 20437 23427 20503 23430
rect 21840 23400 22300 23430
rect 19333 23354 19399 23357
rect 19198 23352 19399 23354
rect 19198 23296 19338 23352
rect 19394 23296 19399 23352
rect 19198 23294 19399 23296
rect 16573 23291 16639 23294
rect 17769 23291 17835 23294
rect 19333 23291 19399 23294
rect -300 23218 160 23248
rect 1669 23218 1735 23221
rect -300 23216 1735 23218
rect -300 23160 1674 23216
rect 1730 23160 1735 23216
rect -300 23158 1735 23160
rect -300 23128 160 23158
rect 1669 23155 1735 23158
rect 2957 23218 3023 23221
rect 3141 23218 3207 23221
rect 2957 23216 3207 23218
rect 2957 23160 2962 23216
rect 3018 23160 3146 23216
rect 3202 23160 3207 23216
rect 2957 23158 3207 23160
rect 2957 23155 3023 23158
rect 3141 23155 3207 23158
rect 3969 23218 4035 23221
rect 13905 23218 13971 23221
rect 3969 23216 13971 23218
rect 3969 23160 3974 23216
rect 4030 23160 13910 23216
rect 13966 23160 13971 23216
rect 3969 23158 13971 23160
rect 3969 23155 4035 23158
rect 13905 23155 13971 23158
rect 3182 23020 3188 23084
rect 3252 23082 3258 23084
rect 3325 23082 3391 23085
rect 3252 23080 3391 23082
rect 3252 23024 3330 23080
rect 3386 23024 3391 23080
rect 3252 23022 3391 23024
rect 3252 23020 3258 23022
rect 3325 23019 3391 23022
rect 4838 23020 4844 23084
rect 4908 23082 4914 23084
rect 9029 23082 9095 23085
rect 4908 23080 9095 23082
rect 4908 23024 9034 23080
rect 9090 23024 9095 23080
rect 4908 23022 9095 23024
rect 4908 23020 4914 23022
rect 9029 23019 9095 23022
rect 9254 23020 9260 23084
rect 9324 23082 9330 23084
rect 10777 23082 10843 23085
rect 12065 23084 12131 23085
rect 12014 23082 12020 23084
rect 9324 23080 10843 23082
rect 9324 23024 10782 23080
rect 10838 23024 10843 23080
rect 9324 23022 10843 23024
rect 11974 23022 12020 23082
rect 12084 23080 12131 23084
rect 12126 23024 12131 23080
rect 9324 23020 9330 23022
rect 10777 23019 10843 23022
rect 12014 23020 12020 23022
rect 12084 23020 12131 23024
rect 12065 23019 12131 23020
rect -300 22946 160 22976
rect 749 22946 815 22949
rect -300 22944 815 22946
rect -300 22888 754 22944
rect 810 22888 815 22944
rect -300 22886 815 22888
rect -300 22856 160 22886
rect 749 22883 815 22886
rect 2773 22946 2839 22949
rect 4521 22946 4587 22949
rect 2773 22944 4587 22946
rect 2773 22888 2778 22944
rect 2834 22888 4526 22944
rect 4582 22888 4587 22944
rect 2773 22886 4587 22888
rect 2773 22883 2839 22886
rect 4521 22883 4587 22886
rect 6269 22946 6335 22949
rect 10174 22946 10180 22948
rect 6269 22944 10180 22946
rect 6269 22888 6274 22944
rect 6330 22888 10180 22944
rect 6269 22886 10180 22888
rect 6269 22883 6335 22886
rect 10174 22884 10180 22886
rect 10244 22884 10250 22948
rect 21265 22946 21331 22949
rect 21840 22946 22300 22976
rect 21265 22944 22300 22946
rect 21265 22888 21270 22944
rect 21326 22888 22300 22944
rect 21265 22886 22300 22888
rect 21265 22883 21331 22886
rect 5890 22880 6206 22881
rect 5890 22816 5896 22880
rect 5960 22816 5976 22880
rect 6040 22816 6056 22880
rect 6120 22816 6136 22880
rect 6200 22816 6206 22880
rect 5890 22815 6206 22816
rect 10835 22880 11151 22881
rect 10835 22816 10841 22880
rect 10905 22816 10921 22880
rect 10985 22816 11001 22880
rect 11065 22816 11081 22880
rect 11145 22816 11151 22880
rect 10835 22815 11151 22816
rect 15780 22880 16096 22881
rect 15780 22816 15786 22880
rect 15850 22816 15866 22880
rect 15930 22816 15946 22880
rect 16010 22816 16026 22880
rect 16090 22816 16096 22880
rect 15780 22815 16096 22816
rect 20725 22880 21041 22881
rect 20725 22816 20731 22880
rect 20795 22816 20811 22880
rect 20875 22816 20891 22880
rect 20955 22816 20971 22880
rect 21035 22816 21041 22880
rect 21840 22856 22300 22886
rect 20725 22815 21041 22816
rect 2814 22748 2820 22812
rect 2884 22810 2890 22812
rect 3969 22810 4035 22813
rect 5574 22810 5580 22812
rect 2884 22808 5580 22810
rect 2884 22752 3974 22808
rect 4030 22752 5580 22808
rect 2884 22750 5580 22752
rect 2884 22748 2890 22750
rect 3969 22747 4035 22750
rect 5574 22748 5580 22750
rect 5644 22748 5650 22812
rect 7230 22748 7236 22812
rect 7300 22810 7306 22812
rect 9070 22810 9076 22812
rect 7300 22750 9076 22810
rect 7300 22748 7306 22750
rect 9070 22748 9076 22750
rect 9140 22748 9146 22812
rect 9213 22810 9279 22813
rect 10593 22812 10659 22813
rect 10542 22810 10548 22812
rect 9213 22808 10548 22810
rect 10612 22808 10659 22812
rect 9213 22752 9218 22808
rect 9274 22752 10548 22808
rect 10654 22752 10659 22808
rect 9213 22750 10548 22752
rect 9213 22747 9279 22750
rect 10542 22748 10548 22750
rect 10612 22748 10659 22752
rect 10593 22747 10659 22748
rect -300 22674 160 22704
rect 1393 22674 1459 22677
rect -300 22672 1459 22674
rect -300 22616 1398 22672
rect 1454 22616 1459 22672
rect -300 22614 1459 22616
rect -300 22584 160 22614
rect 1393 22611 1459 22614
rect 1577 22674 1643 22677
rect 9029 22674 9095 22677
rect 1577 22672 9095 22674
rect 1577 22616 1582 22672
rect 1638 22616 9034 22672
rect 9090 22616 9095 22672
rect 1577 22614 9095 22616
rect 1577 22611 1643 22614
rect 9029 22611 9095 22614
rect 9857 22674 9923 22677
rect 14641 22676 14707 22677
rect 9990 22674 9996 22676
rect 9857 22672 9996 22674
rect 9857 22616 9862 22672
rect 9918 22616 9996 22672
rect 9857 22614 9996 22616
rect 9857 22611 9923 22614
rect 9990 22612 9996 22614
rect 10060 22612 10066 22676
rect 12198 22612 12204 22676
rect 12268 22612 12274 22676
rect 14590 22674 14596 22676
rect 14550 22614 14596 22674
rect 14660 22672 14707 22676
rect 14702 22616 14707 22672
rect 14590 22612 14596 22614
rect 14660 22612 14707 22616
rect 14774 22612 14780 22676
rect 14844 22674 14850 22676
rect 19926 22674 19932 22676
rect 14844 22614 19932 22674
rect 14844 22612 14850 22614
rect 19926 22612 19932 22614
rect 19996 22612 20002 22676
rect 3601 22538 3667 22541
rect 7649 22538 7715 22541
rect 3601 22536 7715 22538
rect 3601 22480 3606 22536
rect 3662 22480 7654 22536
rect 7710 22480 7715 22536
rect 3601 22478 7715 22480
rect 3601 22475 3667 22478
rect 7649 22475 7715 22478
rect 9029 22538 9095 22541
rect 12206 22538 12266 22612
rect 14641 22611 14707 22612
rect 9029 22536 12266 22538
rect 9029 22480 9034 22536
rect 9090 22480 12266 22536
rect 9029 22478 12266 22480
rect 12985 22538 13051 22541
rect 17125 22538 17191 22541
rect 12985 22536 17191 22538
rect 12985 22480 12990 22536
rect 13046 22480 17130 22536
rect 17186 22480 17191 22536
rect 12985 22478 17191 22480
rect 9029 22475 9095 22478
rect 12985 22475 13051 22478
rect 17125 22475 17191 22478
rect 18086 22476 18092 22540
rect 18156 22538 18162 22540
rect 19517 22538 19583 22541
rect 18156 22536 19583 22538
rect 18156 22480 19522 22536
rect 19578 22480 19583 22536
rect 18156 22478 19583 22480
rect 18156 22476 18162 22478
rect 19517 22475 19583 22478
rect 19701 22540 19767 22541
rect 19701 22536 19748 22540
rect 19812 22538 19818 22540
rect 19701 22480 19706 22536
rect 19701 22476 19748 22480
rect 19812 22478 19858 22538
rect 19812 22476 19818 22478
rect 19701 22475 19767 22476
rect -300 22402 160 22432
rect 749 22402 815 22405
rect -300 22400 815 22402
rect -300 22344 754 22400
rect 810 22344 815 22400
rect -300 22342 815 22344
rect -300 22312 160 22342
rect 749 22339 815 22342
rect 4153 22402 4219 22405
rect 4705 22402 4771 22405
rect 4153 22400 4771 22402
rect 4153 22344 4158 22400
rect 4214 22344 4710 22400
rect 4766 22344 4771 22400
rect 4153 22342 4771 22344
rect 4153 22339 4219 22342
rect 4705 22339 4771 22342
rect 13905 22402 13971 22405
rect 15510 22402 15516 22404
rect 13905 22400 15516 22402
rect 13905 22344 13910 22400
rect 13966 22344 15516 22400
rect 13905 22342 15516 22344
rect 13905 22339 13971 22342
rect 15510 22340 15516 22342
rect 15580 22402 15586 22404
rect 16246 22402 16252 22404
rect 15580 22342 16252 22402
rect 15580 22340 15586 22342
rect 16246 22340 16252 22342
rect 16316 22340 16322 22404
rect 19374 22340 19380 22404
rect 19444 22402 19450 22404
rect 19517 22402 19583 22405
rect 19444 22400 19583 22402
rect 19444 22344 19522 22400
rect 19578 22344 19583 22400
rect 19444 22342 19583 22344
rect 19444 22340 19450 22342
rect 19517 22339 19583 22342
rect 20437 22402 20503 22405
rect 21840 22402 22300 22432
rect 20437 22400 22300 22402
rect 20437 22344 20442 22400
rect 20498 22344 22300 22400
rect 20437 22342 22300 22344
rect 20437 22339 20503 22342
rect 3418 22336 3734 22337
rect 3418 22272 3424 22336
rect 3488 22272 3504 22336
rect 3568 22272 3584 22336
rect 3648 22272 3664 22336
rect 3728 22272 3734 22336
rect 3418 22271 3734 22272
rect 8363 22336 8679 22337
rect 8363 22272 8369 22336
rect 8433 22272 8449 22336
rect 8513 22272 8529 22336
rect 8593 22272 8609 22336
rect 8673 22272 8679 22336
rect 8363 22271 8679 22272
rect 13308 22336 13624 22337
rect 13308 22272 13314 22336
rect 13378 22272 13394 22336
rect 13458 22272 13474 22336
rect 13538 22272 13554 22336
rect 13618 22272 13624 22336
rect 13308 22271 13624 22272
rect 18253 22336 18569 22337
rect 18253 22272 18259 22336
rect 18323 22272 18339 22336
rect 18403 22272 18419 22336
rect 18483 22272 18499 22336
rect 18563 22272 18569 22336
rect 21840 22312 22300 22342
rect 18253 22271 18569 22272
rect 2957 22266 3023 22269
rect 7465 22268 7531 22269
rect 4286 22266 4292 22268
rect 2730 22264 3023 22266
rect 2730 22208 2962 22264
rect 3018 22208 3023 22264
rect 2730 22206 3023 22208
rect -300 22130 160 22160
rect 1393 22130 1459 22133
rect -300 22128 1459 22130
rect -300 22072 1398 22128
rect 1454 22072 1459 22128
rect -300 22070 1459 22072
rect -300 22040 160 22070
rect 1393 22067 1459 22070
rect 2129 22130 2195 22133
rect 2730 22130 2790 22206
rect 2957 22203 3023 22206
rect 3972 22206 4292 22266
rect 3972 22133 4032 22206
rect 4286 22204 4292 22206
rect 4356 22204 4362 22268
rect 7414 22266 7420 22268
rect 7374 22206 7420 22266
rect 7484 22264 7531 22268
rect 7526 22208 7531 22264
rect 7414 22204 7420 22206
rect 7484 22204 7531 22208
rect 7465 22203 7531 22204
rect 10501 22268 10567 22269
rect 10501 22264 10548 22268
rect 10612 22266 10618 22268
rect 16849 22266 16915 22269
rect 10501 22208 10506 22264
rect 10501 22204 10548 22208
rect 10612 22206 10658 22266
rect 16849 22264 17188 22266
rect 16849 22208 16854 22264
rect 16910 22208 17188 22264
rect 16849 22206 17188 22208
rect 10612 22204 10618 22206
rect 10501 22203 10567 22204
rect 16849 22203 16915 22206
rect 2129 22128 2790 22130
rect 2129 22072 2134 22128
rect 2190 22072 2790 22128
rect 2129 22070 2790 22072
rect 3969 22128 4035 22133
rect 3969 22072 3974 22128
rect 4030 22072 4035 22128
rect 2129 22067 2195 22070
rect 3969 22067 4035 22072
rect 4102 22068 4108 22132
rect 4172 22130 4178 22132
rect 6361 22130 6427 22133
rect 4172 22128 6427 22130
rect 4172 22072 6366 22128
rect 6422 22072 6427 22128
rect 4172 22070 6427 22072
rect 4172 22068 4178 22070
rect 6361 22067 6427 22070
rect 8017 22130 8083 22133
rect 13169 22130 13235 22133
rect 8017 22128 13235 22130
rect 8017 22072 8022 22128
rect 8078 22072 13174 22128
rect 13230 22072 13235 22128
rect 8017 22070 13235 22072
rect 8017 22067 8083 22070
rect 13169 22067 13235 22070
rect 14733 22130 14799 22133
rect 15326 22130 15332 22132
rect 14733 22128 15332 22130
rect 14733 22072 14738 22128
rect 14794 22072 15332 22128
rect 14733 22070 15332 22072
rect 14733 22067 14799 22070
rect 15326 22068 15332 22070
rect 15396 22068 15402 22132
rect 17128 21997 17188 22206
rect 1209 21994 1275 21997
rect 1894 21994 1900 21996
rect 1209 21992 1900 21994
rect 1209 21936 1214 21992
rect 1270 21936 1900 21992
rect 1209 21934 1900 21936
rect 1209 21931 1275 21934
rect 1894 21932 1900 21934
rect 1964 21932 1970 21996
rect 3601 21994 3667 21997
rect 8109 21994 8175 21997
rect 3601 21992 8175 21994
rect 3601 21936 3606 21992
rect 3662 21936 8114 21992
rect 8170 21936 8175 21992
rect 3601 21934 8175 21936
rect 3601 21931 3667 21934
rect 8109 21931 8175 21934
rect 10225 21994 10291 21997
rect 11830 21994 11836 21996
rect 10225 21992 11836 21994
rect 10225 21936 10230 21992
rect 10286 21936 11836 21992
rect 10225 21934 11836 21936
rect 10225 21931 10291 21934
rect 11830 21932 11836 21934
rect 11900 21932 11906 21996
rect 13629 21994 13695 21997
rect 14641 21994 14707 21997
rect 13629 21992 14707 21994
rect 13629 21936 13634 21992
rect 13690 21936 14646 21992
rect 14702 21936 14707 21992
rect 13629 21934 14707 21936
rect 13629 21931 13695 21934
rect 14641 21931 14707 21934
rect 17125 21992 17191 21997
rect 17125 21936 17130 21992
rect 17186 21936 17191 21992
rect 17125 21931 17191 21936
rect -300 21858 160 21888
rect 841 21858 907 21861
rect -300 21856 907 21858
rect -300 21800 846 21856
rect 902 21800 907 21856
rect -300 21798 907 21800
rect -300 21768 160 21798
rect 841 21795 907 21798
rect 9765 21858 9831 21861
rect 10409 21858 10475 21861
rect 9765 21856 10475 21858
rect 9765 21800 9770 21856
rect 9826 21800 10414 21856
rect 10470 21800 10475 21856
rect 9765 21798 10475 21800
rect 9765 21795 9831 21798
rect 10409 21795 10475 21798
rect 21265 21858 21331 21861
rect 21840 21858 22300 21888
rect 21265 21856 22300 21858
rect 21265 21800 21270 21856
rect 21326 21800 22300 21856
rect 21265 21798 22300 21800
rect 21265 21795 21331 21798
rect 5890 21792 6206 21793
rect 5890 21728 5896 21792
rect 5960 21728 5976 21792
rect 6040 21728 6056 21792
rect 6120 21728 6136 21792
rect 6200 21728 6206 21792
rect 5890 21727 6206 21728
rect 10835 21792 11151 21793
rect 10835 21728 10841 21792
rect 10905 21728 10921 21792
rect 10985 21728 11001 21792
rect 11065 21728 11081 21792
rect 11145 21728 11151 21792
rect 10835 21727 11151 21728
rect 15780 21792 16096 21793
rect 15780 21728 15786 21792
rect 15850 21728 15866 21792
rect 15930 21728 15946 21792
rect 16010 21728 16026 21792
rect 16090 21728 16096 21792
rect 15780 21727 16096 21728
rect 20725 21792 21041 21793
rect 20725 21728 20731 21792
rect 20795 21728 20811 21792
rect 20875 21728 20891 21792
rect 20955 21728 20971 21792
rect 21035 21728 21041 21792
rect 21840 21768 22300 21798
rect 20725 21727 21041 21728
rect 2998 21660 3004 21724
rect 3068 21722 3074 21724
rect 3233 21722 3299 21725
rect 3068 21720 3299 21722
rect 3068 21664 3238 21720
rect 3294 21664 3299 21720
rect 3068 21662 3299 21664
rect 3068 21660 3074 21662
rect 3233 21659 3299 21662
rect 4521 21722 4587 21725
rect 5574 21722 5580 21724
rect 4521 21720 5580 21722
rect 4521 21664 4526 21720
rect 4582 21664 5580 21720
rect 4521 21662 5580 21664
rect 4521 21659 4587 21662
rect 5574 21660 5580 21662
rect 5644 21660 5650 21724
rect 6678 21660 6684 21724
rect 6748 21722 6754 21724
rect 9029 21722 9095 21725
rect 15009 21722 15075 21725
rect 6748 21720 9095 21722
rect 6748 21664 9034 21720
rect 9090 21664 9095 21720
rect 6748 21662 9095 21664
rect 6748 21660 6754 21662
rect 9029 21659 9095 21662
rect 14230 21720 15075 21722
rect 14230 21664 15014 21720
rect 15070 21664 15075 21720
rect 14230 21662 15075 21664
rect -300 21586 160 21616
rect 933 21586 999 21589
rect -300 21584 999 21586
rect -300 21528 938 21584
rect 994 21528 999 21584
rect -300 21526 999 21528
rect -300 21496 160 21526
rect 933 21523 999 21526
rect 1117 21586 1183 21589
rect 3417 21586 3483 21589
rect 1117 21584 3483 21586
rect 1117 21528 1122 21584
rect 1178 21528 3422 21584
rect 3478 21528 3483 21584
rect 1117 21526 3483 21528
rect 1117 21523 1183 21526
rect 3417 21523 3483 21526
rect 4061 21586 4127 21589
rect 11697 21586 11763 21589
rect 12065 21586 12131 21589
rect 14230 21588 14290 21662
rect 15009 21659 15075 21662
rect 4061 21584 12131 21586
rect 4061 21528 4066 21584
rect 4122 21528 11702 21584
rect 11758 21528 12070 21584
rect 12126 21528 12131 21584
rect 4061 21526 12131 21528
rect 4061 21523 4127 21526
rect 11697 21523 11763 21526
rect 12065 21523 12131 21526
rect 14222 21524 14228 21588
rect 14292 21524 14298 21588
rect 790 21388 796 21452
rect 860 21450 866 21452
rect 9305 21450 9371 21453
rect 860 21448 9371 21450
rect 860 21392 9310 21448
rect 9366 21392 9371 21448
rect 860 21390 9371 21392
rect 860 21388 866 21390
rect 9305 21387 9371 21390
rect 10133 21450 10199 21453
rect 16481 21450 16547 21453
rect 10133 21448 16547 21450
rect 10133 21392 10138 21448
rect 10194 21392 16486 21448
rect 16542 21392 16547 21448
rect 10133 21390 16547 21392
rect 10133 21387 10199 21390
rect 16481 21387 16547 21390
rect 17769 21450 17835 21453
rect 19057 21450 19123 21453
rect 17769 21448 19123 21450
rect 17769 21392 17774 21448
rect 17830 21392 19062 21448
rect 19118 21392 19123 21448
rect 17769 21390 19123 21392
rect 17769 21387 17835 21390
rect 19057 21387 19123 21390
rect -300 21314 160 21344
rect 1945 21314 2011 21317
rect -300 21312 2011 21314
rect -300 21256 1950 21312
rect 2006 21256 2011 21312
rect -300 21254 2011 21256
rect -300 21224 160 21254
rect 1945 21251 2011 21254
rect 4705 21314 4771 21317
rect 5901 21314 5967 21317
rect 4705 21312 5967 21314
rect 4705 21256 4710 21312
rect 4766 21256 5906 21312
rect 5962 21256 5967 21312
rect 4705 21254 5967 21256
rect 4705 21251 4771 21254
rect 5901 21251 5967 21254
rect 13813 21312 13879 21317
rect 13813 21256 13818 21312
rect 13874 21256 13879 21312
rect 13813 21251 13879 21256
rect 19885 21314 19951 21317
rect 21840 21314 22300 21344
rect 19885 21312 22300 21314
rect 19885 21256 19890 21312
rect 19946 21256 22300 21312
rect 19885 21254 22300 21256
rect 19885 21251 19951 21254
rect 3418 21248 3734 21249
rect 3418 21184 3424 21248
rect 3488 21184 3504 21248
rect 3568 21184 3584 21248
rect 3648 21184 3664 21248
rect 3728 21184 3734 21248
rect 3418 21183 3734 21184
rect 8363 21248 8679 21249
rect 8363 21184 8369 21248
rect 8433 21184 8449 21248
rect 8513 21184 8529 21248
rect 8593 21184 8609 21248
rect 8673 21184 8679 21248
rect 8363 21183 8679 21184
rect 13308 21248 13624 21249
rect 13308 21184 13314 21248
rect 13378 21184 13394 21248
rect 13458 21184 13474 21248
rect 13538 21184 13554 21248
rect 13618 21184 13624 21248
rect 13308 21183 13624 21184
rect 933 21178 999 21181
rect 2078 21178 2084 21180
rect 933 21176 2084 21178
rect 933 21120 938 21176
rect 994 21120 2084 21176
rect 933 21118 2084 21120
rect 933 21115 999 21118
rect 2078 21116 2084 21118
rect 2148 21116 2154 21180
rect 3969 21178 4035 21181
rect 5390 21178 5396 21180
rect 3969 21176 5396 21178
rect 3969 21120 3974 21176
rect 4030 21120 5396 21176
rect 3969 21118 5396 21120
rect 3969 21115 4035 21118
rect 5390 21116 5396 21118
rect 5460 21116 5466 21180
rect -300 21042 160 21072
rect 1117 21042 1183 21045
rect -300 21040 1183 21042
rect -300 20984 1122 21040
rect 1178 20984 1183 21040
rect -300 20982 1183 20984
rect -300 20952 160 20982
rect 1117 20979 1183 20982
rect 1669 21042 1735 21045
rect 10225 21042 10291 21045
rect 1669 21040 10291 21042
rect 1669 20984 1674 21040
rect 1730 20984 10230 21040
rect 10286 20984 10291 21040
rect 1669 20982 10291 20984
rect 1669 20979 1735 20982
rect 10225 20979 10291 20982
rect 12382 20980 12388 21044
rect 12452 21042 12458 21044
rect 12985 21042 13051 21045
rect 12452 21040 13051 21042
rect 12452 20984 12990 21040
rect 13046 20984 13051 21040
rect 12452 20982 13051 20984
rect 12452 20980 12458 20982
rect 12985 20979 13051 20982
rect 13537 21042 13603 21045
rect 13816 21042 13876 21251
rect 18253 21248 18569 21249
rect 18253 21184 18259 21248
rect 18323 21184 18339 21248
rect 18403 21184 18419 21248
rect 18483 21184 18499 21248
rect 18563 21184 18569 21248
rect 21840 21224 22300 21254
rect 18253 21183 18569 21184
rect 15510 21116 15516 21180
rect 15580 21178 15586 21180
rect 16430 21178 16436 21180
rect 15580 21118 16436 21178
rect 15580 21116 15586 21118
rect 16430 21116 16436 21118
rect 16500 21116 16506 21180
rect 13537 21040 13876 21042
rect 13537 20984 13542 21040
rect 13598 20984 13876 21040
rect 13537 20982 13876 20984
rect 16297 21042 16363 21045
rect 18965 21042 19031 21045
rect 16297 21040 19031 21042
rect 16297 20984 16302 21040
rect 16358 20984 18970 21040
rect 19026 20984 19031 21040
rect 16297 20982 19031 20984
rect 13537 20979 13603 20982
rect 16297 20979 16363 20982
rect 18965 20979 19031 20982
rect 2773 20906 2839 20909
rect 2730 20904 2839 20906
rect 2730 20848 2778 20904
rect 2834 20848 2839 20904
rect 2730 20843 2839 20848
rect 3325 20906 3391 20909
rect 6637 20906 6703 20909
rect 3325 20904 6703 20906
rect 3325 20848 3330 20904
rect 3386 20848 6642 20904
rect 6698 20848 6703 20904
rect 3325 20846 6703 20848
rect 3325 20843 3391 20846
rect 6637 20843 6703 20846
rect 6862 20844 6868 20908
rect 6932 20906 6938 20908
rect 7782 20906 7788 20908
rect 6932 20846 7788 20906
rect 6932 20844 6938 20846
rect 7782 20844 7788 20846
rect 7852 20844 7858 20908
rect 8661 20906 8727 20909
rect 11973 20906 12039 20909
rect 13118 20906 13124 20908
rect 8661 20904 13124 20906
rect 8661 20848 8666 20904
rect 8722 20848 11978 20904
rect 12034 20848 13124 20904
rect 8661 20846 13124 20848
rect 8661 20843 8727 20846
rect 11973 20843 12039 20846
rect 13118 20844 13124 20846
rect 13188 20906 13194 20908
rect 14917 20906 14983 20909
rect 13188 20904 14983 20906
rect 13188 20848 14922 20904
rect 14978 20848 14983 20904
rect 13188 20846 14983 20848
rect 13188 20844 13194 20846
rect 14917 20843 14983 20846
rect 19006 20844 19012 20908
rect 19076 20906 19082 20908
rect 21725 20906 21791 20909
rect 19076 20904 21791 20906
rect 19076 20848 21730 20904
rect 21786 20848 21791 20904
rect 19076 20846 21791 20848
rect 19076 20844 19082 20846
rect 21725 20843 21791 20846
rect -300 20770 160 20800
rect 2730 20770 2790 20843
rect -300 20710 2790 20770
rect -300 20680 160 20710
rect 4838 20708 4844 20772
rect 4908 20770 4914 20772
rect 5717 20770 5783 20773
rect 4908 20768 5783 20770
rect 4908 20712 5722 20768
rect 5778 20712 5783 20768
rect 4908 20710 5783 20712
rect 4908 20708 4914 20710
rect 5717 20707 5783 20710
rect 6361 20770 6427 20773
rect 6494 20770 6500 20772
rect 6361 20768 6500 20770
rect 6361 20712 6366 20768
rect 6422 20712 6500 20768
rect 6361 20710 6500 20712
rect 6361 20707 6427 20710
rect 6494 20708 6500 20710
rect 6564 20708 6570 20772
rect 6862 20708 6868 20772
rect 6932 20770 6938 20772
rect 7465 20770 7531 20773
rect 6932 20768 7531 20770
rect 6932 20712 7470 20768
rect 7526 20712 7531 20768
rect 6932 20710 7531 20712
rect 6932 20708 6938 20710
rect 7465 20707 7531 20710
rect 7966 20708 7972 20772
rect 8036 20770 8042 20772
rect 10133 20770 10199 20773
rect 8036 20768 10199 20770
rect 8036 20712 10138 20768
rect 10194 20712 10199 20768
rect 8036 20710 10199 20712
rect 8036 20708 8042 20710
rect 10133 20707 10199 20710
rect 13537 20770 13603 20773
rect 16481 20772 16547 20773
rect 14958 20770 14964 20772
rect 13537 20768 14964 20770
rect 13537 20712 13542 20768
rect 13598 20712 14964 20768
rect 13537 20710 14964 20712
rect 13537 20707 13603 20710
rect 14958 20708 14964 20710
rect 15028 20708 15034 20772
rect 16430 20770 16436 20772
rect 16390 20710 16436 20770
rect 16500 20768 16547 20772
rect 16542 20712 16547 20768
rect 16430 20708 16436 20710
rect 16500 20708 16547 20712
rect 16481 20707 16547 20708
rect 21265 20770 21331 20773
rect 21840 20770 22300 20800
rect 21265 20768 22300 20770
rect 21265 20712 21270 20768
rect 21326 20712 22300 20768
rect 21265 20710 22300 20712
rect 21265 20707 21331 20710
rect 5890 20704 6206 20705
rect 5890 20640 5896 20704
rect 5960 20640 5976 20704
rect 6040 20640 6056 20704
rect 6120 20640 6136 20704
rect 6200 20640 6206 20704
rect 5890 20639 6206 20640
rect 10835 20704 11151 20705
rect 10835 20640 10841 20704
rect 10905 20640 10921 20704
rect 10985 20640 11001 20704
rect 11065 20640 11081 20704
rect 11145 20640 11151 20704
rect 10835 20639 11151 20640
rect 15780 20704 16096 20705
rect 15780 20640 15786 20704
rect 15850 20640 15866 20704
rect 15930 20640 15946 20704
rect 16010 20640 16026 20704
rect 16090 20640 16096 20704
rect 15780 20639 16096 20640
rect 20725 20704 21041 20705
rect 20725 20640 20731 20704
rect 20795 20640 20811 20704
rect 20875 20640 20891 20704
rect 20955 20640 20971 20704
rect 21035 20640 21041 20704
rect 21840 20680 22300 20710
rect 20725 20639 21041 20640
rect 1945 20634 2011 20637
rect 4981 20634 5047 20637
rect 1945 20632 5047 20634
rect 1945 20576 1950 20632
rect 2006 20576 4986 20632
rect 5042 20576 5047 20632
rect 1945 20574 5047 20576
rect 1945 20571 2011 20574
rect 4981 20571 5047 20574
rect 7281 20634 7347 20637
rect 9949 20634 10015 20637
rect 7281 20632 10015 20634
rect 7281 20576 7286 20632
rect 7342 20576 9954 20632
rect 10010 20576 10015 20632
rect 7281 20574 10015 20576
rect 7281 20571 7347 20574
rect 9949 20571 10015 20574
rect 16481 20634 16547 20637
rect 18086 20634 18092 20636
rect 16481 20632 18092 20634
rect 16481 20576 16486 20632
rect 16542 20576 18092 20632
rect 16481 20574 18092 20576
rect 16481 20571 16547 20574
rect 18086 20572 18092 20574
rect 18156 20572 18162 20636
rect -300 20498 160 20528
rect 749 20498 815 20501
rect -300 20496 815 20498
rect -300 20440 754 20496
rect 810 20440 815 20496
rect -300 20438 815 20440
rect -300 20408 160 20438
rect 749 20435 815 20438
rect 2957 20498 3023 20501
rect 5206 20498 5212 20500
rect 2957 20496 5212 20498
rect 2957 20440 2962 20496
rect 3018 20440 5212 20496
rect 2957 20438 5212 20440
rect 2957 20435 3023 20438
rect 5206 20436 5212 20438
rect 5276 20436 5282 20500
rect 5441 20498 5507 20501
rect 5574 20498 5580 20500
rect 5441 20496 5580 20498
rect 5441 20440 5446 20496
rect 5502 20440 5580 20496
rect 5441 20438 5580 20440
rect 5441 20435 5507 20438
rect 5574 20436 5580 20438
rect 5644 20498 5650 20500
rect 12065 20498 12131 20501
rect 5644 20496 12131 20498
rect 5644 20440 12070 20496
rect 12126 20440 12131 20496
rect 5644 20438 12131 20440
rect 5644 20436 5650 20438
rect 12065 20435 12131 20438
rect 12750 20436 12756 20500
rect 12820 20498 12826 20500
rect 14774 20498 14780 20500
rect 12820 20438 14780 20498
rect 12820 20436 12826 20438
rect 14774 20436 14780 20438
rect 14844 20436 14850 20500
rect 3509 20362 3575 20365
rect 2730 20360 3575 20362
rect 2730 20304 3514 20360
rect 3570 20304 3575 20360
rect 2730 20302 3575 20304
rect -300 20226 160 20256
rect 2730 20226 2790 20302
rect 3509 20299 3575 20302
rect 3693 20362 3759 20365
rect 7373 20362 7439 20365
rect 8150 20362 8156 20364
rect 3693 20360 5090 20362
rect 3693 20304 3698 20360
rect 3754 20304 5090 20360
rect 3693 20302 5090 20304
rect 3693 20299 3759 20302
rect 5030 20229 5090 20302
rect 7373 20360 8156 20362
rect 7373 20304 7378 20360
rect 7434 20304 8156 20360
rect 7373 20302 8156 20304
rect 7373 20299 7439 20302
rect 8150 20300 8156 20302
rect 8220 20362 8226 20364
rect 17217 20362 17283 20365
rect 8220 20360 17283 20362
rect 8220 20304 17222 20360
rect 17278 20304 17283 20360
rect 8220 20302 17283 20304
rect 8220 20300 8226 20302
rect 17217 20299 17283 20302
rect 3233 20228 3299 20229
rect 3182 20226 3188 20228
rect -300 20166 2790 20226
rect 3142 20166 3188 20226
rect 3252 20224 3299 20228
rect 3294 20168 3299 20224
rect -300 20136 160 20166
rect 3182 20164 3188 20166
rect 3252 20164 3299 20168
rect 5030 20224 5139 20229
rect 5030 20168 5078 20224
rect 5134 20168 5139 20224
rect 5030 20166 5139 20168
rect 3233 20163 3299 20164
rect 5073 20163 5139 20166
rect 10542 20164 10548 20228
rect 10612 20226 10618 20228
rect 12709 20226 12775 20229
rect 13997 20228 14063 20229
rect 13997 20226 14044 20228
rect 10612 20224 12775 20226
rect 10612 20168 12714 20224
rect 12770 20168 12775 20224
rect 10612 20166 12775 20168
rect 13952 20224 14044 20226
rect 13952 20168 14002 20224
rect 13952 20166 14044 20168
rect 10612 20164 10618 20166
rect 12709 20163 12775 20166
rect 13997 20164 14044 20166
rect 14108 20164 14114 20228
rect 21541 20226 21607 20229
rect 21840 20226 22300 20256
rect 21541 20224 22300 20226
rect 21541 20168 21546 20224
rect 21602 20168 22300 20224
rect 21541 20166 22300 20168
rect 13997 20163 14063 20164
rect 21541 20163 21607 20166
rect 3418 20160 3734 20161
rect 3418 20096 3424 20160
rect 3488 20096 3504 20160
rect 3568 20096 3584 20160
rect 3648 20096 3664 20160
rect 3728 20096 3734 20160
rect 3418 20095 3734 20096
rect 8363 20160 8679 20161
rect 8363 20096 8369 20160
rect 8433 20096 8449 20160
rect 8513 20096 8529 20160
rect 8593 20096 8609 20160
rect 8673 20096 8679 20160
rect 8363 20095 8679 20096
rect 13308 20160 13624 20161
rect 13308 20096 13314 20160
rect 13378 20096 13394 20160
rect 13458 20096 13474 20160
rect 13538 20096 13554 20160
rect 13618 20096 13624 20160
rect 13308 20095 13624 20096
rect 18253 20160 18569 20161
rect 18253 20096 18259 20160
rect 18323 20096 18339 20160
rect 18403 20096 18419 20160
rect 18483 20096 18499 20160
rect 18563 20096 18569 20160
rect 21840 20136 22300 20166
rect 18253 20095 18569 20096
rect 2221 20090 2287 20093
rect 2221 20088 2330 20090
rect 2221 20032 2226 20088
rect 2282 20032 2330 20088
rect 2221 20027 2330 20032
rect 2814 20028 2820 20092
rect 2884 20090 2890 20092
rect 3233 20090 3299 20093
rect 2884 20088 3299 20090
rect 2884 20032 3238 20088
rect 3294 20032 3299 20088
rect 2884 20030 3299 20032
rect 2884 20028 2890 20030
rect 3233 20027 3299 20030
rect 5257 20090 5323 20093
rect 5390 20090 5396 20092
rect 5257 20088 5396 20090
rect 5257 20032 5262 20088
rect 5318 20032 5396 20088
rect 5257 20030 5396 20032
rect 5257 20027 5323 20030
rect 5390 20028 5396 20030
rect 5460 20028 5466 20092
rect -300 19954 160 19984
rect 1853 19954 1919 19957
rect -300 19952 1919 19954
rect -300 19896 1858 19952
rect 1914 19896 1919 19952
rect -300 19894 1919 19896
rect -300 19864 160 19894
rect 1853 19891 1919 19894
rect 2270 19954 2330 20027
rect 4981 19954 5047 19957
rect 7373 19954 7439 19957
rect 2270 19952 7439 19954
rect 2270 19896 4986 19952
rect 5042 19896 7378 19952
rect 7434 19896 7439 19952
rect 2270 19894 7439 19896
rect 2129 19818 2195 19821
rect 2270 19818 2330 19894
rect 4981 19891 5047 19894
rect 7373 19891 7439 19894
rect 12014 19892 12020 19956
rect 12084 19954 12090 19956
rect 13854 19954 13860 19956
rect 12084 19894 13860 19954
rect 12084 19892 12090 19894
rect 13854 19892 13860 19894
rect 13924 19892 13930 19956
rect 14917 19954 14983 19957
rect 17769 19954 17835 19957
rect 14917 19952 17835 19954
rect 14917 19896 14922 19952
rect 14978 19896 17774 19952
rect 17830 19896 17835 19952
rect 14917 19894 17835 19896
rect 14917 19891 14983 19894
rect 17769 19891 17835 19894
rect 2129 19816 2330 19818
rect 2129 19760 2134 19816
rect 2190 19760 2330 19816
rect 2129 19758 2330 19760
rect 4153 19818 4219 19821
rect 7373 19818 7439 19821
rect 4153 19816 7439 19818
rect 4153 19760 4158 19816
rect 4214 19760 7378 19816
rect 7434 19760 7439 19816
rect 4153 19758 7439 19760
rect 2129 19755 2195 19758
rect 4153 19755 4219 19758
rect 7373 19755 7439 19758
rect 10225 19816 10291 19821
rect 10225 19760 10230 19816
rect 10286 19760 10291 19816
rect 10225 19755 10291 19760
rect 10869 19818 10935 19821
rect 15285 19818 15351 19821
rect 10869 19816 15351 19818
rect 10869 19760 10874 19816
rect 10930 19760 15290 19816
rect 15346 19760 15351 19816
rect 10869 19758 15351 19760
rect 10869 19755 10935 19758
rect 15285 19755 15351 19758
rect 15469 19818 15535 19821
rect 17718 19818 17724 19820
rect 15469 19816 17724 19818
rect 15469 19760 15474 19816
rect 15530 19760 17724 19816
rect 15469 19758 17724 19760
rect 15469 19755 15535 19758
rect 17718 19756 17724 19758
rect 17788 19756 17794 19820
rect -300 19682 160 19712
rect 3141 19682 3207 19685
rect 5257 19682 5323 19685
rect -300 19622 1410 19682
rect -300 19592 160 19622
rect -300 19410 160 19440
rect 1209 19410 1275 19413
rect -300 19408 1275 19410
rect -300 19352 1214 19408
rect 1270 19352 1275 19408
rect -300 19350 1275 19352
rect 1350 19410 1410 19622
rect 3141 19680 5323 19682
rect 3141 19624 3146 19680
rect 3202 19624 5262 19680
rect 5318 19624 5323 19680
rect 3141 19622 5323 19624
rect 3141 19619 3207 19622
rect 5257 19619 5323 19622
rect 8150 19620 8156 19684
rect 8220 19682 8226 19684
rect 10228 19682 10288 19755
rect 8220 19622 10288 19682
rect 21541 19682 21607 19685
rect 21840 19682 22300 19712
rect 21541 19680 22300 19682
rect 21541 19624 21546 19680
rect 21602 19624 22300 19680
rect 21541 19622 22300 19624
rect 8220 19620 8226 19622
rect 21541 19619 21607 19622
rect 5890 19616 6206 19617
rect 5890 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6206 19616
rect 5890 19551 6206 19552
rect 10835 19616 11151 19617
rect 10835 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11151 19616
rect 10835 19551 11151 19552
rect 15780 19616 16096 19617
rect 15780 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16096 19616
rect 15780 19551 16096 19552
rect 20725 19616 21041 19617
rect 20725 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21041 19616
rect 21840 19592 22300 19622
rect 20725 19551 21041 19552
rect 2681 19546 2747 19549
rect 2681 19544 3848 19546
rect 2681 19488 2686 19544
rect 2742 19488 3848 19544
rect 2681 19486 3848 19488
rect 2681 19483 2747 19486
rect 2681 19410 2747 19413
rect 1350 19408 2747 19410
rect 1350 19352 2686 19408
rect 2742 19352 2747 19408
rect 1350 19350 2747 19352
rect -300 19320 160 19350
rect 1209 19347 1275 19350
rect 2681 19347 2747 19350
rect 3182 19348 3188 19412
rect 3252 19410 3258 19412
rect 3325 19410 3391 19413
rect 3252 19408 3391 19410
rect 3252 19352 3330 19408
rect 3386 19352 3391 19408
rect 3252 19350 3391 19352
rect 3788 19410 3848 19486
rect 3918 19484 3924 19548
rect 3988 19546 3994 19548
rect 5533 19546 5599 19549
rect 3988 19544 5599 19546
rect 3988 19488 5538 19544
rect 5594 19488 5599 19544
rect 3988 19486 5599 19488
rect 3988 19484 3994 19486
rect 5533 19483 5599 19486
rect 6545 19546 6611 19549
rect 6545 19544 9506 19546
rect 6545 19488 6550 19544
rect 6606 19488 9506 19544
rect 6545 19486 9506 19488
rect 6545 19483 6611 19486
rect 6361 19410 6427 19413
rect 3788 19408 6427 19410
rect 3788 19352 6366 19408
rect 6422 19352 6427 19408
rect 3788 19350 6427 19352
rect 3252 19348 3258 19350
rect 3325 19347 3391 19350
rect 6361 19347 6427 19350
rect 8937 19410 9003 19413
rect 9254 19410 9260 19412
rect 8937 19408 9260 19410
rect 8937 19352 8942 19408
rect 8998 19352 9260 19408
rect 8937 19350 9260 19352
rect 8937 19347 9003 19350
rect 9254 19348 9260 19350
rect 9324 19348 9330 19412
rect 9446 19410 9506 19486
rect 10358 19484 10364 19548
rect 10428 19546 10434 19548
rect 10501 19546 10567 19549
rect 10428 19544 10567 19546
rect 10428 19488 10506 19544
rect 10562 19488 10567 19544
rect 10428 19486 10567 19488
rect 10428 19484 10434 19486
rect 10501 19483 10567 19486
rect 11646 19484 11652 19548
rect 11716 19546 11722 19548
rect 11881 19546 11947 19549
rect 13353 19546 13419 19549
rect 11716 19544 11947 19546
rect 11716 19488 11886 19544
rect 11942 19488 11947 19544
rect 11716 19486 11947 19488
rect 11716 19484 11722 19486
rect 11881 19483 11947 19486
rect 12988 19544 13419 19546
rect 12988 19488 13358 19544
rect 13414 19488 13419 19544
rect 12988 19486 13419 19488
rect 11278 19410 11284 19412
rect 9446 19350 11284 19410
rect 11278 19348 11284 19350
rect 11348 19410 11354 19412
rect 12988 19410 13048 19486
rect 13353 19483 13419 19486
rect 11348 19350 13048 19410
rect 11348 19348 11354 19350
rect 1669 19274 1735 19277
rect 10409 19274 10475 19277
rect 1669 19272 6194 19274
rect 1669 19216 1674 19272
rect 1730 19216 6194 19272
rect 1669 19214 6194 19216
rect 1669 19211 1735 19214
rect -300 19138 160 19168
rect 6134 19138 6194 19214
rect 8158 19272 10475 19274
rect 8158 19216 10414 19272
rect 10470 19216 10475 19272
rect 8158 19214 10475 19216
rect 8158 19138 8218 19214
rect 10409 19211 10475 19214
rect 10542 19212 10548 19276
rect 10612 19274 10618 19276
rect 10685 19274 10751 19277
rect 13997 19274 14063 19277
rect 10612 19272 10751 19274
rect 10612 19216 10690 19272
rect 10746 19216 10751 19272
rect 10612 19214 10751 19216
rect 10612 19212 10618 19214
rect 10685 19211 10751 19214
rect 13172 19272 14063 19274
rect 13172 19216 14002 19272
rect 14058 19216 14063 19272
rect 13172 19214 14063 19216
rect -300 19078 1962 19138
rect 6134 19078 8218 19138
rect 9765 19136 9831 19141
rect 9765 19080 9770 19136
rect 9826 19080 9831 19136
rect -300 19048 160 19078
rect 381 19002 447 19005
rect 1761 19002 1827 19005
rect 381 19000 1827 19002
rect 381 18944 386 19000
rect 442 18944 1766 19000
rect 1822 18944 1827 19000
rect 381 18942 1827 18944
rect 381 18939 447 18942
rect 1761 18939 1827 18942
rect -300 18866 160 18896
rect 749 18866 815 18869
rect -300 18864 815 18866
rect -300 18808 754 18864
rect 810 18808 815 18864
rect -300 18806 815 18808
rect -300 18776 160 18806
rect 749 18803 815 18806
rect -300 18594 160 18624
rect 749 18594 815 18597
rect -300 18592 815 18594
rect -300 18536 754 18592
rect 810 18536 815 18592
rect -300 18534 815 18536
rect 1902 18594 1962 19078
rect 9765 19075 9831 19080
rect 9949 19138 10015 19141
rect 13172 19138 13232 19214
rect 13997 19211 14063 19214
rect 9949 19136 13232 19138
rect 9949 19080 9954 19136
rect 10010 19080 13232 19136
rect 9949 19078 13232 19080
rect 20069 19138 20135 19141
rect 21840 19138 22300 19168
rect 20069 19136 22300 19138
rect 20069 19080 20074 19136
rect 20130 19080 22300 19136
rect 20069 19078 22300 19080
rect 9949 19075 10015 19078
rect 20069 19075 20135 19078
rect 3418 19072 3734 19073
rect 3418 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3734 19072
rect 3418 19007 3734 19008
rect 8363 19072 8679 19073
rect 8363 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8679 19072
rect 8363 19007 8679 19008
rect 9397 19002 9463 19005
rect 9768 19002 9828 19075
rect 13308 19072 13624 19073
rect 13308 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13624 19072
rect 13308 19007 13624 19008
rect 18253 19072 18569 19073
rect 18253 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18569 19072
rect 21840 19048 22300 19078
rect 18253 19007 18569 19008
rect 12341 19004 12407 19005
rect 12341 19002 12388 19004
rect 9397 19000 9828 19002
rect 9397 18944 9402 19000
rect 9458 18944 9828 19000
rect 9397 18942 9828 18944
rect 12296 19000 12388 19002
rect 12296 18944 12346 19000
rect 12296 18942 12388 18944
rect 9397 18939 9463 18942
rect 12341 18940 12388 18942
rect 12452 18940 12458 19004
rect 12341 18939 12407 18940
rect 2589 18866 2655 18869
rect 6678 18866 6684 18868
rect 2589 18864 6684 18866
rect 2589 18808 2594 18864
rect 2650 18808 6684 18864
rect 2589 18806 6684 18808
rect 2589 18803 2655 18806
rect 6678 18804 6684 18806
rect 6748 18804 6754 18868
rect 7281 18866 7347 18869
rect 7414 18866 7420 18868
rect 7281 18864 7420 18866
rect 7281 18808 7286 18864
rect 7342 18808 7420 18864
rect 7281 18806 7420 18808
rect 7281 18803 7347 18806
rect 7414 18804 7420 18806
rect 7484 18804 7490 18868
rect 7833 18866 7899 18869
rect 7966 18866 7972 18868
rect 7833 18864 7972 18866
rect 7833 18808 7838 18864
rect 7894 18808 7972 18864
rect 7833 18806 7972 18808
rect 7833 18803 7899 18806
rect 7966 18804 7972 18806
rect 8036 18804 8042 18868
rect 9254 18804 9260 18868
rect 9324 18866 9330 18868
rect 10041 18866 10107 18869
rect 9324 18864 10107 18866
rect 9324 18808 10046 18864
rect 10102 18808 10107 18864
rect 9324 18806 10107 18808
rect 9324 18804 9330 18806
rect 10041 18803 10107 18806
rect 10501 18866 10567 18869
rect 14590 18866 14596 18868
rect 10501 18864 14596 18866
rect 10501 18808 10506 18864
rect 10562 18808 14596 18864
rect 10501 18806 14596 18808
rect 10501 18803 10567 18806
rect 14590 18804 14596 18806
rect 14660 18866 14666 18868
rect 14917 18866 14983 18869
rect 14660 18864 14983 18866
rect 14660 18808 14922 18864
rect 14978 18808 14983 18864
rect 14660 18806 14983 18808
rect 14660 18804 14666 18806
rect 14917 18803 14983 18806
rect 2037 18730 2103 18733
rect 11830 18730 11836 18732
rect 2037 18728 11836 18730
rect 2037 18672 2042 18728
rect 2098 18672 11836 18728
rect 2037 18670 11836 18672
rect 2037 18667 2103 18670
rect 11830 18668 11836 18670
rect 11900 18668 11906 18732
rect 12341 18730 12407 18733
rect 21449 18730 21515 18733
rect 12341 18728 21515 18730
rect 12341 18672 12346 18728
rect 12402 18672 21454 18728
rect 21510 18672 21515 18728
rect 12341 18670 21515 18672
rect 12341 18667 12407 18670
rect 21449 18667 21515 18670
rect 3049 18594 3115 18597
rect 1902 18592 3115 18594
rect 1902 18536 3054 18592
rect 3110 18536 3115 18592
rect 1902 18534 3115 18536
rect -300 18504 160 18534
rect 749 18531 815 18534
rect 3049 18531 3115 18534
rect 21265 18594 21331 18597
rect 21840 18594 22300 18624
rect 21265 18592 22300 18594
rect 21265 18536 21270 18592
rect 21326 18536 22300 18592
rect 21265 18534 22300 18536
rect 21265 18531 21331 18534
rect 5890 18528 6206 18529
rect 5890 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6206 18528
rect 5890 18463 6206 18464
rect 10835 18528 11151 18529
rect 10835 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11151 18528
rect 10835 18463 11151 18464
rect 15780 18528 16096 18529
rect 15780 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16096 18528
rect 15780 18463 16096 18464
rect 20725 18528 21041 18529
rect 20725 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21041 18528
rect 21840 18504 22300 18534
rect 20725 18463 21041 18464
rect 1485 18458 1551 18461
rect 2446 18458 2452 18460
rect 1485 18456 2452 18458
rect 1485 18400 1490 18456
rect 1546 18400 2452 18456
rect 1485 18398 2452 18400
rect 1485 18395 1551 18398
rect 2446 18396 2452 18398
rect 2516 18396 2522 18460
rect 2630 18396 2636 18460
rect 2700 18458 2706 18460
rect 2865 18458 2931 18461
rect 3049 18460 3115 18461
rect 2700 18456 2931 18458
rect 2700 18400 2870 18456
rect 2926 18400 2931 18456
rect 2700 18398 2931 18400
rect 2700 18396 2706 18398
rect 2865 18395 2931 18398
rect 2998 18396 3004 18460
rect 3068 18458 3115 18460
rect 3601 18458 3667 18461
rect 5574 18458 5580 18460
rect 3068 18456 3160 18458
rect 3110 18400 3160 18456
rect 3068 18398 3160 18400
rect 3601 18456 5580 18458
rect 3601 18400 3606 18456
rect 3662 18400 5580 18456
rect 3601 18398 5580 18400
rect 3068 18396 3115 18398
rect 3049 18395 3115 18396
rect 3601 18395 3667 18398
rect 5574 18396 5580 18398
rect 5644 18396 5650 18460
rect 14273 18458 14339 18461
rect 14406 18458 14412 18460
rect 14273 18456 14412 18458
rect 14273 18400 14278 18456
rect 14334 18400 14412 18456
rect 14273 18398 14412 18400
rect 14273 18395 14339 18398
rect 14406 18396 14412 18398
rect 14476 18396 14482 18460
rect -300 18322 160 18352
rect 1209 18322 1275 18325
rect -300 18320 1275 18322
rect -300 18264 1214 18320
rect 1270 18264 1275 18320
rect -300 18262 1275 18264
rect -300 18232 160 18262
rect 1209 18259 1275 18262
rect 1577 18322 1643 18325
rect 2262 18322 2268 18324
rect 1577 18320 2268 18322
rect 1577 18264 1582 18320
rect 1638 18264 2268 18320
rect 1577 18262 2268 18264
rect 1577 18259 1643 18262
rect 2262 18260 2268 18262
rect 2332 18260 2338 18324
rect 5901 18322 5967 18325
rect 3604 18320 5967 18322
rect 3604 18264 5906 18320
rect 5962 18264 5967 18320
rect 3604 18262 5967 18264
rect 749 18188 815 18189
rect 749 18186 796 18188
rect 704 18184 796 18186
rect 704 18128 754 18184
rect 704 18126 796 18128
rect 749 18124 796 18126
rect 860 18124 866 18188
rect 1117 18186 1183 18189
rect 3604 18186 3664 18262
rect 5901 18259 5967 18262
rect 6310 18260 6316 18324
rect 6380 18322 6386 18324
rect 7465 18322 7531 18325
rect 13629 18322 13695 18325
rect 16941 18322 17007 18325
rect 6380 18320 17007 18322
rect 6380 18264 7470 18320
rect 7526 18264 13634 18320
rect 13690 18264 16946 18320
rect 17002 18264 17007 18320
rect 6380 18262 17007 18264
rect 6380 18260 6386 18262
rect 7465 18259 7531 18262
rect 13629 18259 13695 18262
rect 16941 18259 17007 18262
rect 19190 18260 19196 18324
rect 19260 18322 19266 18324
rect 21817 18322 21883 18325
rect 19260 18320 21883 18322
rect 19260 18264 21822 18320
rect 21878 18264 21883 18320
rect 19260 18262 21883 18264
rect 19260 18260 19266 18262
rect 21817 18259 21883 18262
rect 1117 18184 3664 18186
rect 1117 18128 1122 18184
rect 1178 18128 3664 18184
rect 1117 18126 3664 18128
rect 3785 18186 3851 18189
rect 4245 18186 4311 18189
rect 3785 18184 4311 18186
rect 3785 18128 3790 18184
rect 3846 18128 4250 18184
rect 4306 18128 4311 18184
rect 3785 18126 4311 18128
rect 749 18123 815 18124
rect 1117 18123 1183 18126
rect 3785 18123 3851 18126
rect 4245 18123 4311 18126
rect 6678 18124 6684 18188
rect 6748 18186 6754 18188
rect 9305 18186 9371 18189
rect 6748 18184 9371 18186
rect 6748 18128 9310 18184
rect 9366 18128 9371 18184
rect 6748 18126 9371 18128
rect 6748 18124 6754 18126
rect 9305 18123 9371 18126
rect 9622 18124 9628 18188
rect 9692 18186 9698 18188
rect 10685 18186 10751 18189
rect 9692 18184 10751 18186
rect 9692 18128 10690 18184
rect 10746 18128 10751 18184
rect 9692 18126 10751 18128
rect 9692 18124 9698 18126
rect 10685 18123 10751 18126
rect 13118 18124 13124 18188
rect 13188 18186 13194 18188
rect 15469 18186 15535 18189
rect 13188 18184 15535 18186
rect 13188 18128 15474 18184
rect 15530 18128 15535 18184
rect 13188 18126 15535 18128
rect 13188 18124 13194 18126
rect 15469 18123 15535 18126
rect 16573 18186 16639 18189
rect 20110 18186 20116 18188
rect 16573 18184 20116 18186
rect 16573 18128 16578 18184
rect 16634 18128 20116 18184
rect 16573 18126 20116 18128
rect 16573 18123 16639 18126
rect 20110 18124 20116 18126
rect 20180 18124 20186 18188
rect -300 18050 160 18080
rect 1485 18050 1551 18053
rect 12341 18050 12407 18053
rect -300 18048 1551 18050
rect -300 17992 1490 18048
rect 1546 17992 1551 18048
rect -300 17990 1551 17992
rect -300 17960 160 17990
rect 1485 17987 1551 17990
rect 8756 18048 12407 18050
rect 8756 17992 12346 18048
rect 12402 17992 12407 18048
rect 8756 17990 12407 17992
rect 3418 17984 3734 17985
rect 3418 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3734 17984
rect 3418 17919 3734 17920
rect 8363 17984 8679 17985
rect 8363 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8679 17984
rect 8363 17919 8679 17920
rect 4102 17852 4108 17916
rect 4172 17914 4178 17916
rect 4245 17914 4311 17917
rect 4172 17912 4311 17914
rect 4172 17856 4250 17912
rect 4306 17856 4311 17912
rect 4172 17854 4311 17856
rect 4172 17852 4178 17854
rect 4245 17851 4311 17854
rect -300 17778 160 17808
rect 2681 17778 2747 17781
rect -300 17776 2747 17778
rect -300 17720 2686 17776
rect 2742 17720 2747 17776
rect -300 17718 2747 17720
rect -300 17688 160 17718
rect 2681 17715 2747 17718
rect 3509 17778 3575 17781
rect 5441 17778 5507 17781
rect 8756 17778 8816 17990
rect 12341 17987 12407 17990
rect 20989 18050 21055 18053
rect 21840 18050 22300 18080
rect 20989 18048 22300 18050
rect 20989 17992 20994 18048
rect 21050 17992 22300 18048
rect 20989 17990 22300 17992
rect 20989 17987 21055 17990
rect 13308 17984 13624 17985
rect 13308 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13624 17984
rect 13308 17919 13624 17920
rect 18253 17984 18569 17985
rect 18253 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18569 17984
rect 21840 17960 22300 17990
rect 18253 17919 18569 17920
rect 9489 17912 9555 17917
rect 9489 17856 9494 17912
rect 9550 17856 9555 17912
rect 9489 17851 9555 17856
rect 3509 17776 5507 17778
rect 3509 17720 3514 17776
rect 3570 17720 5446 17776
rect 5502 17720 5507 17776
rect 3509 17718 5507 17720
rect 3509 17715 3575 17718
rect 5441 17715 5507 17718
rect 5720 17718 8816 17778
rect 9492 17778 9552 17851
rect 14222 17778 14228 17780
rect 9492 17718 14228 17778
rect 1894 17580 1900 17644
rect 1964 17642 1970 17644
rect 5720 17642 5780 17718
rect 14222 17716 14228 17718
rect 14292 17716 14298 17780
rect 1964 17582 5780 17642
rect 9581 17642 9647 17645
rect 9806 17642 9812 17644
rect 9581 17640 9812 17642
rect 9581 17584 9586 17640
rect 9642 17584 9812 17640
rect 9581 17582 9812 17584
rect 1964 17580 1970 17582
rect 9581 17579 9647 17582
rect 9806 17580 9812 17582
rect 9876 17580 9882 17644
rect 17585 17642 17651 17645
rect 11286 17640 17651 17642
rect 11286 17584 17590 17640
rect 17646 17584 17651 17640
rect 11286 17582 17651 17584
rect -300 17506 160 17536
rect 1577 17506 1643 17509
rect -300 17504 1643 17506
rect -300 17448 1582 17504
rect 1638 17448 1643 17504
rect -300 17446 1643 17448
rect -300 17416 160 17446
rect 1577 17443 1643 17446
rect 4654 17444 4660 17508
rect 4724 17506 4730 17508
rect 5073 17506 5139 17509
rect 4724 17504 5139 17506
rect 4724 17448 5078 17504
rect 5134 17448 5139 17504
rect 4724 17446 5139 17448
rect 4724 17444 4730 17446
rect 2313 17370 2379 17373
rect 4662 17370 4722 17444
rect 5073 17443 5139 17446
rect 7833 17506 7899 17509
rect 7833 17504 10426 17506
rect 7833 17448 7838 17504
rect 7894 17448 10426 17504
rect 7833 17446 10426 17448
rect 7833 17443 7899 17446
rect 5890 17440 6206 17441
rect 5890 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6206 17440
rect 5890 17375 6206 17376
rect 2313 17368 4722 17370
rect 2313 17312 2318 17368
rect 2374 17312 4722 17368
rect 2313 17310 4722 17312
rect 10133 17370 10199 17373
rect 10133 17368 10242 17370
rect 10133 17312 10138 17368
rect 10194 17312 10242 17368
rect 2313 17307 2379 17310
rect 10133 17307 10242 17312
rect -300 17234 160 17264
rect 2129 17234 2195 17237
rect 9857 17234 9923 17237
rect 10182 17236 10242 17307
rect -300 17232 2195 17234
rect -300 17176 2134 17232
rect 2190 17176 2195 17232
rect -300 17174 2195 17176
rect -300 17144 160 17174
rect 2129 17171 2195 17174
rect 9814 17232 9923 17234
rect 9814 17176 9862 17232
rect 9918 17176 9923 17232
rect 9814 17171 9923 17176
rect 10174 17172 10180 17236
rect 10244 17172 10250 17236
rect 10366 17234 10426 17446
rect 10835 17440 11151 17441
rect 10835 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11151 17440
rect 10835 17375 11151 17376
rect 11286 17372 11346 17582
rect 17585 17579 17651 17582
rect 21265 17506 21331 17509
rect 21840 17506 22300 17536
rect 21265 17504 22300 17506
rect 21265 17448 21270 17504
rect 21326 17448 22300 17504
rect 21265 17446 22300 17448
rect 21265 17443 21331 17446
rect 15780 17440 16096 17441
rect 15780 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16096 17440
rect 15780 17375 16096 17376
rect 20725 17440 21041 17441
rect 20725 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21041 17440
rect 21840 17416 22300 17446
rect 20725 17375 21041 17376
rect 11278 17308 11284 17372
rect 11348 17308 11354 17372
rect 10366 17174 17418 17234
rect 4337 17098 4403 17101
rect 9305 17098 9371 17101
rect 9814 17100 9874 17171
rect 4337 17096 9371 17098
rect 4337 17040 4342 17096
rect 4398 17040 9310 17096
rect 9366 17040 9371 17096
rect 4337 17038 9371 17040
rect 4337 17035 4403 17038
rect 9305 17035 9371 17038
rect 9806 17036 9812 17100
rect 9876 17036 9882 17100
rect 9949 17098 10015 17101
rect 10409 17098 10475 17101
rect 11789 17100 11855 17101
rect 11789 17098 11836 17100
rect 9949 17096 10475 17098
rect 9949 17040 9954 17096
rect 10010 17040 10414 17096
rect 10470 17040 10475 17096
rect 9949 17038 10475 17040
rect 11744 17096 11836 17098
rect 11744 17040 11794 17096
rect 11744 17038 11836 17040
rect 9949 17035 10015 17038
rect 10409 17035 10475 17038
rect 11789 17036 11836 17038
rect 11900 17036 11906 17100
rect 12065 17098 12131 17101
rect 12617 17098 12683 17101
rect 15377 17098 15443 17101
rect 12065 17096 12683 17098
rect 12065 17040 12070 17096
rect 12126 17040 12622 17096
rect 12678 17040 12683 17096
rect 12065 17038 12683 17040
rect 11789 17035 11855 17036
rect 12065 17035 12131 17038
rect 12617 17035 12683 17038
rect 13172 17096 15443 17098
rect 13172 17040 15382 17096
rect 15438 17040 15443 17096
rect 13172 17038 15443 17040
rect 17358 17098 17418 17174
rect 18045 17098 18111 17101
rect 17358 17096 18111 17098
rect 17358 17040 18050 17096
rect 18106 17040 18111 17096
rect 17358 17038 18111 17040
rect -300 16962 160 16992
rect 1577 16962 1643 16965
rect -300 16960 1643 16962
rect -300 16904 1582 16960
rect 1638 16904 1643 16960
rect -300 16902 1643 16904
rect -300 16872 160 16902
rect 1577 16899 1643 16902
rect 1761 16962 1827 16965
rect 2589 16962 2655 16965
rect 1761 16960 2655 16962
rect 1761 16904 1766 16960
rect 1822 16904 2594 16960
rect 2650 16904 2655 16960
rect 1761 16902 2655 16904
rect 1761 16899 1827 16902
rect 2589 16899 2655 16902
rect 5022 16900 5028 16964
rect 5092 16962 5098 16964
rect 5901 16962 5967 16965
rect 5092 16960 5967 16962
rect 5092 16904 5906 16960
rect 5962 16904 5967 16960
rect 5092 16902 5967 16904
rect 5092 16900 5098 16902
rect 5901 16899 5967 16902
rect 9765 16962 9831 16965
rect 13172 16962 13232 17038
rect 15377 17035 15443 17038
rect 18045 17035 18111 17038
rect 19793 17098 19859 17101
rect 19977 17098 20043 17101
rect 19793 17096 20043 17098
rect 19793 17040 19798 17096
rect 19854 17040 19982 17096
rect 20038 17040 20043 17096
rect 19793 17038 20043 17040
rect 19793 17035 19859 17038
rect 19977 17035 20043 17038
rect 9765 16960 13232 16962
rect 9765 16904 9770 16960
rect 9826 16904 13232 16960
rect 9765 16902 13232 16904
rect 20897 16962 20963 16965
rect 21840 16962 22300 16992
rect 20897 16960 22300 16962
rect 20897 16904 20902 16960
rect 20958 16904 22300 16960
rect 20897 16902 22300 16904
rect 9765 16899 9831 16902
rect 20897 16899 20963 16902
rect 3418 16896 3734 16897
rect 3418 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3734 16896
rect 3418 16831 3734 16832
rect 8363 16896 8679 16897
rect 8363 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8679 16896
rect 8363 16831 8679 16832
rect 13308 16896 13624 16897
rect 13308 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13624 16896
rect 13308 16831 13624 16832
rect 18253 16896 18569 16897
rect 18253 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18569 16896
rect 21840 16872 22300 16902
rect 18253 16831 18569 16832
rect 1669 16826 1735 16829
rect 3049 16826 3115 16829
rect 1669 16824 3115 16826
rect 1669 16768 1674 16824
rect 1730 16768 3054 16824
rect 3110 16768 3115 16824
rect 1669 16766 3115 16768
rect 1669 16763 1735 16766
rect 3049 16763 3115 16766
rect 4153 16826 4219 16829
rect 7097 16826 7163 16829
rect 4153 16824 7163 16826
rect 4153 16768 4158 16824
rect 4214 16768 7102 16824
rect 7158 16768 7163 16824
rect 4153 16766 7163 16768
rect 4153 16763 4219 16766
rect 7097 16763 7163 16766
rect 9213 16826 9279 16829
rect 9622 16826 9628 16828
rect 9213 16824 9628 16826
rect 9213 16768 9218 16824
rect 9274 16768 9628 16824
rect 9213 16766 9628 16768
rect 9213 16763 9279 16766
rect 9622 16764 9628 16766
rect 9692 16764 9698 16828
rect 9857 16826 9923 16829
rect 11789 16826 11855 16829
rect 9857 16824 11855 16826
rect 9857 16768 9862 16824
rect 9918 16768 11794 16824
rect 11850 16768 11855 16824
rect 9857 16766 11855 16768
rect 9857 16763 9923 16766
rect 11789 16763 11855 16766
rect 14038 16764 14044 16828
rect 14108 16826 14114 16828
rect 16481 16826 16547 16829
rect 14108 16824 16547 16826
rect 14108 16768 16486 16824
rect 16542 16768 16547 16824
rect 14108 16766 16547 16768
rect 14108 16764 14114 16766
rect 16481 16763 16547 16766
rect -300 16690 160 16720
rect 1761 16690 1827 16693
rect -300 16688 1827 16690
rect -300 16632 1766 16688
rect 1822 16632 1827 16688
rect -300 16630 1827 16632
rect -300 16600 160 16630
rect 1761 16627 1827 16630
rect 2681 16690 2747 16693
rect 16021 16690 16087 16693
rect 2681 16688 16087 16690
rect 2681 16632 2686 16688
rect 2742 16632 16026 16688
rect 16082 16632 16087 16688
rect 2681 16630 16087 16632
rect 2681 16627 2747 16630
rect 16021 16627 16087 16630
rect 19742 16628 19748 16692
rect 19812 16690 19818 16692
rect 21725 16690 21791 16693
rect 19812 16688 21791 16690
rect 19812 16632 21730 16688
rect 21786 16632 21791 16688
rect 19812 16630 21791 16632
rect 19812 16628 19818 16630
rect 21725 16627 21791 16630
rect 749 16554 815 16557
rect 2078 16554 2084 16556
rect 749 16552 2084 16554
rect 749 16496 754 16552
rect 810 16496 2084 16552
rect 749 16494 2084 16496
rect 749 16491 815 16494
rect 2078 16492 2084 16494
rect 2148 16492 2154 16556
rect 2497 16554 2563 16557
rect 3417 16554 3483 16557
rect 2497 16552 3483 16554
rect 2497 16496 2502 16552
rect 2558 16496 3422 16552
rect 3478 16496 3483 16552
rect 2497 16494 3483 16496
rect 2497 16491 2563 16494
rect 3417 16491 3483 16494
rect 3969 16554 4035 16557
rect 15193 16554 15259 16557
rect 16481 16554 16547 16557
rect 18045 16556 18111 16557
rect 17350 16554 17356 16556
rect 3969 16552 15259 16554
rect 3969 16496 3974 16552
rect 4030 16496 15198 16552
rect 15254 16496 15259 16552
rect 3969 16494 15259 16496
rect 3969 16491 4035 16494
rect 15193 16491 15259 16494
rect 15334 16494 16268 16554
rect -300 16418 160 16448
rect 657 16418 723 16421
rect -300 16416 723 16418
rect -300 16360 662 16416
rect 718 16360 723 16416
rect -300 16358 723 16360
rect -300 16328 160 16358
rect 657 16355 723 16358
rect 2221 16418 2287 16421
rect 3785 16418 3851 16421
rect 2221 16416 3851 16418
rect 2221 16360 2226 16416
rect 2282 16360 3790 16416
rect 3846 16360 3851 16416
rect 2221 16358 3851 16360
rect 2221 16355 2287 16358
rect 3785 16355 3851 16358
rect 4102 16356 4108 16420
rect 4172 16418 4178 16420
rect 4889 16418 4955 16421
rect 4172 16416 4955 16418
rect 4172 16360 4894 16416
rect 4950 16360 4955 16416
rect 4172 16358 4955 16360
rect 4172 16356 4178 16358
rect 4889 16355 4955 16358
rect 6494 16356 6500 16420
rect 6564 16418 6570 16420
rect 7833 16418 7899 16421
rect 6564 16416 7899 16418
rect 6564 16360 7838 16416
rect 7894 16360 7899 16416
rect 6564 16358 7899 16360
rect 6564 16356 6570 16358
rect 7833 16355 7899 16358
rect 12157 16418 12223 16421
rect 15334 16418 15394 16494
rect 12157 16416 15394 16418
rect 12157 16360 12162 16416
rect 12218 16360 15394 16416
rect 12157 16358 15394 16360
rect 16208 16418 16268 16494
rect 16481 16552 17356 16554
rect 16481 16496 16486 16552
rect 16542 16496 17356 16552
rect 16481 16494 17356 16496
rect 16481 16491 16547 16494
rect 17350 16492 17356 16494
rect 17420 16492 17426 16556
rect 18045 16552 18092 16556
rect 18156 16554 18162 16556
rect 20437 16554 20503 16557
rect 18045 16496 18050 16552
rect 18045 16492 18092 16496
rect 18156 16494 18202 16554
rect 20437 16552 21282 16554
rect 20437 16496 20442 16552
rect 20498 16496 21282 16552
rect 20437 16494 21282 16496
rect 18156 16492 18162 16494
rect 18045 16491 18111 16492
rect 20437 16491 20503 16494
rect 19374 16418 19380 16420
rect 16208 16358 19380 16418
rect 12157 16355 12223 16358
rect 19374 16356 19380 16358
rect 19444 16356 19450 16420
rect 21222 16418 21282 16494
rect 21840 16418 22300 16448
rect 21222 16358 22300 16418
rect 5890 16352 6206 16353
rect 5890 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6206 16352
rect 5890 16287 6206 16288
rect 10835 16352 11151 16353
rect 10835 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11151 16352
rect 10835 16287 11151 16288
rect 15780 16352 16096 16353
rect 15780 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16096 16352
rect 15780 16287 16096 16288
rect 20725 16352 21041 16353
rect 20725 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21041 16352
rect 21840 16328 22300 16358
rect 20725 16287 21041 16288
rect 3918 16282 3924 16284
rect 3052 16222 3924 16282
rect -300 16146 160 16176
rect 841 16146 907 16149
rect -300 16144 907 16146
rect -300 16088 846 16144
rect 902 16088 907 16144
rect -300 16086 907 16088
rect -300 16056 160 16086
rect 841 16083 907 16086
rect 2865 16146 2931 16149
rect 3052 16146 3112 16222
rect 3918 16220 3924 16222
rect 3988 16220 3994 16284
rect 4337 16282 4403 16285
rect 9673 16282 9739 16285
rect 4110 16280 4403 16282
rect 4110 16224 4342 16280
rect 4398 16224 4403 16280
rect 4110 16222 4403 16224
rect 2865 16144 3112 16146
rect 2865 16088 2870 16144
rect 2926 16088 3112 16144
rect 2865 16086 3112 16088
rect 2865 16083 2931 16086
rect 3182 16084 3188 16148
rect 3252 16146 3258 16148
rect 4110 16146 4170 16222
rect 4337 16219 4403 16222
rect 8572 16280 9739 16282
rect 8572 16224 9678 16280
rect 9734 16224 9739 16280
rect 8572 16222 9739 16224
rect 3252 16086 4170 16146
rect 5441 16146 5507 16149
rect 6310 16146 6316 16148
rect 5441 16144 6316 16146
rect 5441 16088 5446 16144
rect 5502 16088 6316 16144
rect 5441 16086 6316 16088
rect 3252 16084 3258 16086
rect 5441 16083 5507 16086
rect 6310 16084 6316 16086
rect 6380 16084 6386 16148
rect 7598 16084 7604 16148
rect 7668 16146 7674 16148
rect 8109 16146 8175 16149
rect 8572 16146 8632 16222
rect 9673 16219 9739 16222
rect 11646 16220 11652 16284
rect 11716 16282 11722 16284
rect 15510 16282 15516 16284
rect 11716 16222 15516 16282
rect 11716 16220 11722 16222
rect 15510 16220 15516 16222
rect 15580 16220 15586 16284
rect 7668 16144 8632 16146
rect 7668 16088 8114 16144
rect 8170 16088 8632 16144
rect 7668 16086 8632 16088
rect 8753 16146 8819 16149
rect 11053 16146 11119 16149
rect 8753 16144 11119 16146
rect 8753 16088 8758 16144
rect 8814 16088 11058 16144
rect 11114 16088 11119 16144
rect 8753 16086 11119 16088
rect 7668 16084 7674 16086
rect 8109 16083 8175 16086
rect 8753 16083 8819 16086
rect 11053 16083 11119 16086
rect 14457 16146 14523 16149
rect 15510 16146 15516 16148
rect 14457 16144 15516 16146
rect 14457 16088 14462 16144
rect 14518 16088 15516 16144
rect 14457 16086 15516 16088
rect 14457 16083 14523 16086
rect 15510 16084 15516 16086
rect 15580 16084 15586 16148
rect 16941 16146 17007 16149
rect 18689 16146 18755 16149
rect 16941 16144 18755 16146
rect 16941 16088 16946 16144
rect 17002 16088 18694 16144
rect 18750 16088 18755 16144
rect 16941 16086 18755 16088
rect 16941 16083 17007 16086
rect 18689 16083 18755 16086
rect 1761 16012 1827 16013
rect 1710 16010 1716 16012
rect 1670 15950 1716 16010
rect 1780 16008 1827 16012
rect 1822 15952 1827 16008
rect 1710 15948 1716 15950
rect 1780 15948 1827 15952
rect 1761 15947 1827 15948
rect 2037 16010 2103 16013
rect 17769 16010 17835 16013
rect 2037 16008 17835 16010
rect 2037 15952 2042 16008
rect 2098 15952 17774 16008
rect 17830 15952 17835 16008
rect 2037 15950 17835 15952
rect 2037 15947 2103 15950
rect 17769 15947 17835 15950
rect 17902 15948 17908 16012
rect 17972 16010 17978 16012
rect 19517 16010 19583 16013
rect 17972 16008 19583 16010
rect 17972 15952 19522 16008
rect 19578 15952 19583 16008
rect 17972 15950 19583 15952
rect 17972 15948 17978 15950
rect 19517 15947 19583 15950
rect -300 15874 160 15904
rect 1669 15874 1735 15877
rect -300 15872 1735 15874
rect -300 15816 1674 15872
rect 1730 15816 1735 15872
rect -300 15814 1735 15816
rect -300 15784 160 15814
rect 1669 15811 1735 15814
rect 3877 15874 3943 15877
rect 5901 15874 5967 15877
rect 3877 15872 5967 15874
rect 3877 15816 3882 15872
rect 3938 15816 5906 15872
rect 5962 15816 5967 15872
rect 3877 15814 5967 15816
rect 3877 15811 3943 15814
rect 5901 15811 5967 15814
rect 9305 15874 9371 15877
rect 11830 15874 11836 15876
rect 9305 15872 11836 15874
rect 9305 15816 9310 15872
rect 9366 15816 11836 15872
rect 9305 15814 11836 15816
rect 9305 15811 9371 15814
rect 11830 15812 11836 15814
rect 11900 15874 11906 15876
rect 11900 15814 12588 15874
rect 11900 15812 11906 15814
rect 3418 15808 3734 15809
rect 3418 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3734 15808
rect 3418 15743 3734 15744
rect 8363 15808 8679 15809
rect 8363 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8679 15808
rect 8363 15743 8679 15744
rect 6729 15738 6795 15741
rect 7005 15738 7071 15741
rect 6729 15736 7071 15738
rect 6729 15680 6734 15736
rect 6790 15680 7010 15736
rect 7066 15680 7071 15736
rect 6729 15678 7071 15680
rect 6729 15675 6795 15678
rect 7005 15675 7071 15678
rect 9121 15738 9187 15741
rect 9305 15738 9371 15741
rect 11605 15738 11671 15741
rect 9121 15736 11671 15738
rect 9121 15680 9126 15736
rect 9182 15680 9310 15736
rect 9366 15680 11610 15736
rect 11666 15680 11671 15736
rect 9121 15678 11671 15680
rect 9121 15675 9187 15678
rect 9305 15675 9371 15678
rect 11605 15675 11671 15678
rect -300 15602 160 15632
rect 2129 15602 2195 15605
rect -300 15600 2195 15602
rect -300 15544 2134 15600
rect 2190 15544 2195 15600
rect -300 15542 2195 15544
rect -300 15512 160 15542
rect 2129 15539 2195 15542
rect 4838 15540 4844 15604
rect 4908 15602 4914 15604
rect 5441 15602 5507 15605
rect 5574 15602 5580 15604
rect 4908 15600 5580 15602
rect 4908 15544 5446 15600
rect 5502 15544 5580 15600
rect 4908 15542 5580 15544
rect 4908 15540 4914 15542
rect 5441 15539 5507 15542
rect 5574 15540 5580 15542
rect 5644 15540 5650 15604
rect 6637 15602 6703 15605
rect 6862 15602 6868 15604
rect 6637 15600 6868 15602
rect 6637 15544 6642 15600
rect 6698 15544 6868 15600
rect 6637 15542 6868 15544
rect 6637 15539 6703 15542
rect 6862 15540 6868 15542
rect 6932 15540 6938 15604
rect 7465 15602 7531 15605
rect 12341 15602 12407 15605
rect 7465 15600 12407 15602
rect 7465 15544 7470 15600
rect 7526 15544 12346 15600
rect 12402 15544 12407 15600
rect 7465 15542 12407 15544
rect 12528 15602 12588 15814
rect 12934 15812 12940 15876
rect 13004 15874 13010 15876
rect 13169 15874 13235 15877
rect 13004 15872 13235 15874
rect 13004 15816 13174 15872
rect 13230 15816 13235 15872
rect 13004 15814 13235 15816
rect 13004 15812 13010 15814
rect 13169 15811 13235 15814
rect 20437 15874 20503 15877
rect 21840 15874 22300 15904
rect 20437 15872 22300 15874
rect 20437 15816 20442 15872
rect 20498 15816 22300 15872
rect 20437 15814 22300 15816
rect 20437 15811 20503 15814
rect 13308 15808 13624 15809
rect 13308 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13624 15808
rect 13308 15743 13624 15744
rect 18253 15808 18569 15809
rect 18253 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18569 15808
rect 21840 15784 22300 15814
rect 18253 15743 18569 15744
rect 16665 15738 16731 15741
rect 13724 15736 16731 15738
rect 13724 15680 16670 15736
rect 16726 15680 16731 15736
rect 13724 15678 16731 15680
rect 13724 15602 13784 15678
rect 16665 15675 16731 15678
rect 12528 15542 13784 15602
rect 7465 15539 7531 15542
rect 12341 15539 12407 15542
rect 14958 15540 14964 15604
rect 15028 15602 15034 15604
rect 18413 15602 18479 15605
rect 15028 15600 18479 15602
rect 15028 15544 18418 15600
rect 18474 15544 18479 15600
rect 15028 15542 18479 15544
rect 15028 15540 15034 15542
rect 18413 15539 18479 15542
rect 238 15404 244 15468
rect 308 15466 314 15468
rect 6821 15466 6887 15469
rect 15561 15466 15627 15469
rect 308 15406 6378 15466
rect 308 15404 314 15406
rect -300 15330 160 15360
rect 1577 15330 1643 15333
rect -300 15328 1643 15330
rect -300 15272 1582 15328
rect 1638 15272 1643 15328
rect -300 15270 1643 15272
rect -300 15240 160 15270
rect 1577 15267 1643 15270
rect 5533 15332 5599 15333
rect 5533 15328 5580 15332
rect 5644 15330 5650 15332
rect 6318 15330 6378 15406
rect 6821 15464 15627 15466
rect 6821 15408 6826 15464
rect 6882 15408 15566 15464
rect 15622 15408 15627 15464
rect 6821 15406 15627 15408
rect 6821 15403 6887 15406
rect 15561 15403 15627 15406
rect 16798 15404 16804 15468
rect 16868 15466 16874 15468
rect 16941 15466 17007 15469
rect 16868 15464 17007 15466
rect 16868 15408 16946 15464
rect 17002 15408 17007 15464
rect 16868 15406 17007 15408
rect 16868 15404 16874 15406
rect 16941 15403 17007 15406
rect 8661 15330 8727 15333
rect 9581 15330 9647 15333
rect 5533 15272 5538 15328
rect 5533 15268 5580 15272
rect 5644 15270 5690 15330
rect 6318 15270 7068 15330
rect 5644 15268 5650 15270
rect 5533 15267 5599 15268
rect 5890 15264 6206 15265
rect 5890 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6206 15264
rect 5890 15199 6206 15200
rect 289 15194 355 15197
rect 790 15194 796 15196
rect 289 15192 796 15194
rect 289 15136 294 15192
rect 350 15136 796 15192
rect 289 15134 796 15136
rect 289 15131 355 15134
rect 790 15132 796 15134
rect 860 15132 866 15196
rect 6545 15194 6611 15197
rect 6862 15194 6868 15196
rect 6545 15192 6868 15194
rect 6545 15136 6550 15192
rect 6606 15136 6868 15192
rect 6545 15134 6868 15136
rect 6545 15131 6611 15134
rect 6862 15132 6868 15134
rect 6932 15132 6938 15196
rect 7008 15194 7068 15270
rect 8661 15328 9647 15330
rect 8661 15272 8666 15328
rect 8722 15272 9586 15328
rect 9642 15272 9647 15328
rect 8661 15270 9647 15272
rect 8661 15267 8727 15270
rect 9581 15267 9647 15270
rect 9949 15330 10015 15333
rect 10358 15330 10364 15332
rect 9949 15328 10364 15330
rect 9949 15272 9954 15328
rect 10010 15272 10364 15328
rect 9949 15270 10364 15272
rect 9949 15267 10015 15270
rect 10358 15268 10364 15270
rect 10428 15268 10434 15332
rect 14549 15330 14615 15333
rect 14917 15330 14983 15333
rect 14549 15328 14983 15330
rect 14549 15272 14554 15328
rect 14610 15272 14922 15328
rect 14978 15272 14983 15328
rect 14549 15270 14983 15272
rect 14549 15267 14615 15270
rect 14917 15267 14983 15270
rect 21265 15330 21331 15333
rect 21840 15330 22300 15360
rect 21265 15328 22300 15330
rect 21265 15272 21270 15328
rect 21326 15272 22300 15328
rect 21265 15270 22300 15272
rect 21265 15267 21331 15270
rect 10835 15264 11151 15265
rect 10835 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11151 15264
rect 10835 15199 11151 15200
rect 15780 15264 16096 15265
rect 15780 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16096 15264
rect 15780 15199 16096 15200
rect 20725 15264 21041 15265
rect 20725 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21041 15264
rect 21840 15240 22300 15270
rect 20725 15199 21041 15200
rect 12157 15194 12223 15197
rect 7008 15134 9322 15194
rect -300 15058 160 15088
rect 1945 15058 2011 15061
rect -300 15056 2011 15058
rect -300 15000 1950 15056
rect 2006 15000 2011 15056
rect -300 14998 2011 15000
rect -300 14968 160 14998
rect 1945 14995 2011 14998
rect 6545 15058 6611 15061
rect 6821 15058 6887 15061
rect 6545 15056 6887 15058
rect 6545 15000 6550 15056
rect 6606 15000 6826 15056
rect 6882 15000 6887 15056
rect 6545 14998 6887 15000
rect 6545 14995 6611 14998
rect 6821 14995 6887 14998
rect 7741 15058 7807 15061
rect 9121 15058 9187 15061
rect 7741 15056 9187 15058
rect 7741 15000 7746 15056
rect 7802 15000 9126 15056
rect 9182 15000 9187 15056
rect 7741 14998 9187 15000
rect 9262 15058 9322 15134
rect 11240 15192 12223 15194
rect 11240 15136 12162 15192
rect 12218 15136 12223 15192
rect 11240 15134 12223 15136
rect 11240 15058 11300 15134
rect 12157 15131 12223 15134
rect 14273 15194 14339 15197
rect 15193 15194 15259 15197
rect 14273 15192 15259 15194
rect 14273 15136 14278 15192
rect 14334 15136 15198 15192
rect 15254 15136 15259 15192
rect 14273 15134 15259 15136
rect 14273 15131 14339 15134
rect 15193 15131 15259 15134
rect 18689 15194 18755 15197
rect 18822 15194 18828 15196
rect 18689 15192 18828 15194
rect 18689 15136 18694 15192
rect 18750 15136 18828 15192
rect 18689 15134 18828 15136
rect 18689 15131 18755 15134
rect 18822 15132 18828 15134
rect 18892 15132 18898 15196
rect 12157 15060 12223 15061
rect 12157 15058 12204 15060
rect 9262 14998 11300 15058
rect 12112 15056 12204 15058
rect 12112 15000 12162 15056
rect 12112 14998 12204 15000
rect 7741 14995 7807 14998
rect 9121 14995 9187 14998
rect 12157 14996 12204 14998
rect 12268 14996 12274 15060
rect 13854 14996 13860 15060
rect 13924 15058 13930 15060
rect 16982 15058 16988 15060
rect 13924 14998 16988 15058
rect 13924 14996 13930 14998
rect 16982 14996 16988 14998
rect 17052 14996 17058 15060
rect 17350 14996 17356 15060
rect 17420 15058 17426 15060
rect 18638 15058 18644 15060
rect 17420 14998 18644 15058
rect 17420 14996 17426 14998
rect 18638 14996 18644 14998
rect 18708 14996 18714 15060
rect 12157 14995 12223 14996
rect 473 14922 539 14925
rect 1894 14922 1900 14924
rect 473 14920 1900 14922
rect 473 14864 478 14920
rect 534 14864 1900 14920
rect 473 14862 1900 14864
rect 473 14859 539 14862
rect 1894 14860 1900 14862
rect 1964 14860 1970 14924
rect 3325 14922 3391 14925
rect 4613 14922 4679 14925
rect 3325 14920 4679 14922
rect 3325 14864 3330 14920
rect 3386 14864 4618 14920
rect 4674 14864 4679 14920
rect 3325 14862 4679 14864
rect 3325 14859 3391 14862
rect 4613 14859 4679 14862
rect 7649 14922 7715 14925
rect 8017 14922 8083 14925
rect 8569 14922 8635 14925
rect 10593 14922 10659 14925
rect 12893 14922 12959 14925
rect 17401 14922 17467 14925
rect 18638 14922 18644 14924
rect 7649 14920 10426 14922
rect 7649 14864 7654 14920
rect 7710 14864 8022 14920
rect 8078 14864 8574 14920
rect 8630 14864 10426 14920
rect 7649 14862 10426 14864
rect 7649 14859 7715 14862
rect 8017 14859 8083 14862
rect 8569 14859 8635 14862
rect -300 14786 160 14816
rect 841 14786 907 14789
rect -300 14784 907 14786
rect -300 14728 846 14784
rect 902 14728 907 14784
rect -300 14726 907 14728
rect -300 14696 160 14726
rect 841 14723 907 14726
rect 5390 14724 5396 14788
rect 5460 14786 5466 14788
rect 6177 14786 6243 14789
rect 5460 14784 6243 14786
rect 5460 14728 6182 14784
rect 6238 14728 6243 14784
rect 5460 14726 6243 14728
rect 10366 14786 10426 14862
rect 10593 14920 12959 14922
rect 10593 14864 10598 14920
rect 10654 14864 12898 14920
rect 12954 14864 12959 14920
rect 10593 14862 12959 14864
rect 10593 14859 10659 14862
rect 12893 14859 12959 14862
rect 13080 14862 13784 14922
rect 11053 14786 11119 14789
rect 13080 14786 13140 14862
rect 10366 14784 11119 14786
rect 10366 14728 11058 14784
rect 11114 14728 11119 14784
rect 10366 14726 11119 14728
rect 5460 14724 5466 14726
rect 6177 14723 6243 14726
rect 11053 14723 11119 14726
rect 11240 14726 13140 14786
rect 13724 14786 13784 14862
rect 17401 14920 18644 14922
rect 17401 14864 17406 14920
rect 17462 14864 18644 14920
rect 17401 14862 18644 14864
rect 17401 14859 17467 14862
rect 18638 14860 18644 14862
rect 18708 14860 18714 14924
rect 20437 14786 20503 14789
rect 21840 14786 22300 14816
rect 13724 14726 17602 14786
rect 3418 14720 3734 14721
rect 3418 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3734 14720
rect 3418 14655 3734 14656
rect 8363 14720 8679 14721
rect 8363 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8679 14720
rect 8363 14655 8679 14656
rect 2681 14652 2747 14653
rect 2630 14650 2636 14652
rect 2554 14590 2636 14650
rect 2700 14650 2747 14652
rect 2998 14650 3004 14652
rect 2700 14648 3004 14650
rect 2742 14592 3004 14648
rect 2630 14588 2636 14590
rect 2700 14590 3004 14592
rect 2700 14588 2747 14590
rect 2998 14588 3004 14590
rect 3068 14588 3074 14652
rect 5206 14588 5212 14652
rect 5276 14650 5282 14652
rect 6269 14650 6335 14653
rect 11240 14650 11300 14726
rect 13308 14720 13624 14721
rect 13308 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13624 14720
rect 13308 14655 13624 14656
rect 5276 14648 6335 14650
rect 5276 14592 6274 14648
rect 6330 14592 6335 14648
rect 5276 14590 6335 14592
rect 5276 14588 5282 14590
rect 2681 14587 2747 14588
rect 6269 14587 6335 14590
rect 9216 14590 11300 14650
rect 12065 14650 12131 14653
rect 12617 14650 12683 14653
rect 12065 14648 12683 14650
rect 12065 14592 12070 14648
rect 12126 14592 12622 14648
rect 12678 14592 12683 14648
rect 12065 14590 12683 14592
rect -300 14514 160 14544
rect 565 14516 631 14517
rect 565 14514 612 14516
rect -300 14454 306 14514
rect 520 14512 612 14514
rect 520 14456 570 14512
rect 520 14454 612 14456
rect -300 14424 160 14454
rect 246 14378 306 14454
rect 565 14452 612 14454
rect 676 14452 682 14516
rect 1158 14452 1164 14516
rect 1228 14514 1234 14516
rect 1393 14514 1459 14517
rect 1228 14512 1459 14514
rect 1228 14456 1398 14512
rect 1454 14456 1459 14512
rect 1228 14454 1459 14456
rect 1228 14452 1234 14454
rect 565 14451 631 14452
rect 1393 14451 1459 14454
rect 4286 14452 4292 14516
rect 4356 14514 4362 14516
rect 4705 14514 4771 14517
rect 7281 14514 7347 14517
rect 7925 14514 7991 14517
rect 4356 14512 7991 14514
rect 4356 14456 4710 14512
rect 4766 14456 7286 14512
rect 7342 14456 7930 14512
rect 7986 14456 7991 14512
rect 4356 14454 7991 14456
rect 4356 14452 4362 14454
rect 4705 14451 4771 14454
rect 7281 14451 7347 14454
rect 7925 14451 7991 14454
rect 933 14378 999 14381
rect 246 14376 999 14378
rect 246 14320 938 14376
rect 994 14320 999 14376
rect 246 14318 999 14320
rect 933 14315 999 14318
rect 4797 14378 4863 14381
rect 9216 14378 9276 14590
rect 12065 14587 12131 14590
rect 12617 14587 12683 14590
rect 14222 14588 14228 14652
rect 14292 14650 14298 14652
rect 16205 14650 16271 14653
rect 17542 14652 17602 14726
rect 20437 14784 22300 14786
rect 20437 14728 20442 14784
rect 20498 14728 22300 14784
rect 20437 14726 22300 14728
rect 20437 14723 20503 14726
rect 18253 14720 18569 14721
rect 18253 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18569 14720
rect 21840 14696 22300 14726
rect 18253 14655 18569 14656
rect 14292 14648 16271 14650
rect 14292 14592 16210 14648
rect 16266 14592 16271 14648
rect 14292 14590 16271 14592
rect 14292 14588 14298 14590
rect 16205 14587 16271 14590
rect 17534 14588 17540 14652
rect 17604 14588 17610 14652
rect 9857 14514 9923 14517
rect 11513 14514 11579 14517
rect 15009 14514 15075 14517
rect 9857 14512 15075 14514
rect 9857 14456 9862 14512
rect 9918 14456 11518 14512
rect 11574 14456 15014 14512
rect 15070 14456 15075 14512
rect 9857 14454 15075 14456
rect 9857 14451 9923 14454
rect 11513 14451 11579 14454
rect 15009 14451 15075 14454
rect 15142 14452 15148 14516
rect 15212 14514 15218 14516
rect 19190 14514 19196 14516
rect 15212 14454 19196 14514
rect 15212 14452 15218 14454
rect 19190 14452 19196 14454
rect 19260 14452 19266 14516
rect 4797 14376 9276 14378
rect 4797 14320 4802 14376
rect 4858 14320 9276 14376
rect 4797 14318 9276 14320
rect 4797 14315 4863 14318
rect 9622 14316 9628 14380
rect 9692 14378 9698 14380
rect 14273 14378 14339 14381
rect 9692 14376 14339 14378
rect 9692 14320 14278 14376
rect 14334 14320 14339 14376
rect 9692 14318 14339 14320
rect 9692 14316 9698 14318
rect 14273 14315 14339 14318
rect 14406 14316 14412 14380
rect 14476 14378 14482 14380
rect 14825 14378 14891 14381
rect 14476 14376 14891 14378
rect 14476 14320 14830 14376
rect 14886 14320 14891 14376
rect 14476 14318 14891 14320
rect 14476 14316 14482 14318
rect 14825 14315 14891 14318
rect 15101 14380 15167 14381
rect 15101 14376 15148 14380
rect 15212 14378 15218 14380
rect 16297 14378 16363 14381
rect 15101 14320 15106 14376
rect 15101 14316 15148 14320
rect 15212 14318 15258 14378
rect 15656 14376 16363 14378
rect 15656 14320 16302 14376
rect 16358 14320 16363 14376
rect 15656 14318 16363 14320
rect 15212 14316 15218 14318
rect 15101 14315 15167 14316
rect -300 14242 160 14272
rect -300 14182 306 14242
rect -300 14152 160 14182
rect 246 14106 306 14182
rect 1342 14180 1348 14244
rect 1412 14242 1418 14244
rect 4102 14242 4108 14244
rect 1412 14182 4108 14242
rect 1412 14180 1418 14182
rect 4102 14180 4108 14182
rect 4172 14180 4178 14244
rect 7741 14242 7807 14245
rect 8753 14242 8819 14245
rect 7741 14240 8819 14242
rect 7741 14184 7746 14240
rect 7802 14184 8758 14240
rect 8814 14184 8819 14240
rect 7741 14182 8819 14184
rect 7741 14179 7807 14182
rect 8753 14179 8819 14182
rect 13118 14180 13124 14244
rect 13188 14242 13194 14244
rect 15656 14242 15716 14318
rect 16297 14315 16363 14318
rect 17677 14378 17743 14381
rect 18229 14378 18295 14381
rect 17677 14376 18295 14378
rect 17677 14320 17682 14376
rect 17738 14320 18234 14376
rect 18290 14320 18295 14376
rect 17677 14318 18295 14320
rect 17677 14315 17743 14318
rect 18229 14315 18295 14318
rect 13188 14182 15716 14242
rect 21265 14242 21331 14245
rect 21840 14242 22300 14272
rect 21265 14240 22300 14242
rect 21265 14184 21270 14240
rect 21326 14184 22300 14240
rect 21265 14182 22300 14184
rect 13188 14180 13194 14182
rect 21265 14179 21331 14182
rect 5890 14176 6206 14177
rect 5890 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6206 14176
rect 5890 14111 6206 14112
rect 10835 14176 11151 14177
rect 10835 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11151 14176
rect 10835 14111 11151 14112
rect 15780 14176 16096 14177
rect 15780 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16096 14176
rect 15780 14111 16096 14112
rect 20725 14176 21041 14177
rect 20725 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21041 14176
rect 21840 14152 22300 14182
rect 20725 14111 21041 14112
rect 2589 14106 2655 14109
rect 246 14104 2655 14106
rect 246 14048 2594 14104
rect 2650 14048 2655 14104
rect 246 14046 2655 14048
rect 2589 14043 2655 14046
rect 4061 14104 4127 14109
rect 6361 14108 6427 14109
rect 4061 14048 4066 14104
rect 4122 14048 4127 14104
rect 4061 14043 4127 14048
rect 6310 14044 6316 14108
rect 6380 14106 6427 14108
rect 7281 14106 7347 14109
rect 7414 14106 7420 14108
rect 6380 14104 6472 14106
rect 6422 14048 6472 14104
rect 6380 14046 6472 14048
rect 7281 14104 7420 14106
rect 7281 14048 7286 14104
rect 7342 14048 7420 14104
rect 7281 14046 7420 14048
rect 6380 14044 6427 14046
rect 6361 14043 6427 14044
rect 7281 14043 7347 14046
rect 7414 14044 7420 14046
rect 7484 14044 7490 14108
rect 9949 14106 10015 14109
rect 10685 14106 10751 14109
rect 9949 14104 10751 14106
rect 9949 14048 9954 14104
rect 10010 14048 10690 14104
rect 10746 14048 10751 14104
rect 9949 14046 10751 14048
rect 9949 14043 10015 14046
rect 10685 14043 10751 14046
rect 12065 14106 12131 14109
rect 14774 14106 14780 14108
rect 12065 14104 14780 14106
rect 12065 14048 12070 14104
rect 12126 14048 14780 14104
rect 12065 14046 14780 14048
rect 12065 14043 12131 14046
rect 14774 14044 14780 14046
rect 14844 14044 14850 14108
rect 15469 14106 15535 14109
rect 15150 14104 15535 14106
rect 15150 14048 15474 14104
rect 15530 14048 15535 14104
rect 15150 14046 15535 14048
rect -300 13970 160 14000
rect 2037 13970 2103 13973
rect 4064 13970 4124 14043
rect -300 13968 2103 13970
rect -300 13912 2042 13968
rect 2098 13912 2103 13968
rect -300 13910 2103 13912
rect -300 13880 160 13910
rect 2037 13907 2103 13910
rect 2270 13910 4124 13970
rect 4429 13970 4495 13973
rect 15150 13970 15210 14046
rect 15469 14043 15535 14046
rect 4429 13968 15210 13970
rect 4429 13912 4434 13968
rect 4490 13912 15210 13968
rect 4429 13910 15210 13912
rect 289 13834 355 13837
rect 2270 13834 2330 13910
rect 4429 13907 4495 13910
rect 15326 13908 15332 13972
rect 15396 13970 15402 13972
rect 20110 13970 20116 13972
rect 15396 13910 20116 13970
rect 15396 13908 15402 13910
rect 20110 13908 20116 13910
rect 20180 13908 20186 13972
rect 289 13832 2330 13834
rect 289 13776 294 13832
rect 350 13776 2330 13832
rect 289 13774 2330 13776
rect 3877 13834 3943 13837
rect 7189 13834 7255 13837
rect 3877 13832 7255 13834
rect 3877 13776 3882 13832
rect 3938 13776 7194 13832
rect 7250 13776 7255 13832
rect 3877 13774 7255 13776
rect 289 13771 355 13774
rect 3877 13771 3943 13774
rect 7189 13771 7255 13774
rect 7925 13834 7991 13837
rect 8201 13834 8267 13837
rect 7925 13832 8267 13834
rect 7925 13776 7930 13832
rect 7986 13776 8206 13832
rect 8262 13776 8267 13832
rect 7925 13774 8267 13776
rect 7925 13771 7991 13774
rect 8201 13771 8267 13774
rect 9029 13834 9095 13837
rect 9673 13834 9739 13837
rect 9029 13832 9739 13834
rect 9029 13776 9034 13832
rect 9090 13776 9678 13832
rect 9734 13776 9739 13832
rect 9029 13774 9739 13776
rect 9029 13771 9095 13774
rect 9673 13771 9739 13774
rect 10593 13834 10659 13837
rect 10593 13832 14704 13834
rect 10593 13776 10598 13832
rect 10654 13776 14704 13832
rect 10593 13774 14704 13776
rect 10593 13771 10659 13774
rect -300 13698 160 13728
rect 1485 13698 1551 13701
rect -300 13696 1551 13698
rect -300 13640 1490 13696
rect 1546 13640 1551 13696
rect -300 13638 1551 13640
rect -300 13608 160 13638
rect 1485 13635 1551 13638
rect 4102 13636 4108 13700
rect 4172 13698 4178 13700
rect 5533 13698 5599 13701
rect 4172 13696 5599 13698
rect 4172 13640 5538 13696
rect 5594 13640 5599 13696
rect 4172 13638 5599 13640
rect 4172 13636 4178 13638
rect 5533 13635 5599 13638
rect 7281 13698 7347 13701
rect 7414 13698 7420 13700
rect 7281 13696 7420 13698
rect 7281 13640 7286 13696
rect 7342 13640 7420 13696
rect 7281 13638 7420 13640
rect 7281 13635 7347 13638
rect 7414 13636 7420 13638
rect 7484 13636 7490 13700
rect 14644 13698 14704 13774
rect 14774 13772 14780 13836
rect 14844 13834 14850 13836
rect 17309 13834 17375 13837
rect 14844 13832 17375 13834
rect 14844 13776 17314 13832
rect 17370 13776 17375 13832
rect 14844 13774 17375 13776
rect 14844 13772 14850 13774
rect 17309 13771 17375 13774
rect 16941 13698 17007 13701
rect 14644 13696 17007 13698
rect 14644 13640 16946 13696
rect 17002 13640 17007 13696
rect 14644 13638 17007 13640
rect 16941 13635 17007 13638
rect 19517 13698 19583 13701
rect 21840 13698 22300 13728
rect 19517 13696 22300 13698
rect 19517 13640 19522 13696
rect 19578 13640 22300 13696
rect 19517 13638 22300 13640
rect 19517 13635 19583 13638
rect 3418 13632 3734 13633
rect 3418 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3734 13632
rect 3418 13567 3734 13568
rect 8363 13632 8679 13633
rect 8363 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8679 13632
rect 8363 13567 8679 13568
rect 13308 13632 13624 13633
rect 13308 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13624 13632
rect 13308 13567 13624 13568
rect 18253 13632 18569 13633
rect 18253 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18569 13632
rect 21840 13608 22300 13638
rect 18253 13567 18569 13568
rect 5993 13562 6059 13565
rect 7373 13562 7439 13565
rect 5993 13560 7439 13562
rect 5993 13504 5998 13560
rect 6054 13504 7378 13560
rect 7434 13504 7439 13560
rect 5993 13502 7439 13504
rect 5993 13499 6059 13502
rect 7373 13499 7439 13502
rect 9990 13500 9996 13564
rect 10060 13562 10066 13564
rect 12709 13562 12775 13565
rect 16430 13562 16436 13564
rect 10060 13560 12775 13562
rect 10060 13504 12714 13560
rect 12770 13504 12775 13560
rect 10060 13502 12775 13504
rect 10060 13500 10066 13502
rect 12709 13499 12775 13502
rect 14460 13502 16436 13562
rect -300 13426 160 13456
rect 3969 13426 4035 13429
rect -300 13424 4035 13426
rect -300 13368 3974 13424
rect 4030 13368 4035 13424
rect -300 13366 4035 13368
rect -300 13336 160 13366
rect 3969 13363 4035 13366
rect 5574 13364 5580 13428
rect 5644 13426 5650 13428
rect 5809 13426 5875 13429
rect 5644 13424 5875 13426
rect 5644 13368 5814 13424
rect 5870 13368 5875 13424
rect 5644 13366 5875 13368
rect 5644 13364 5650 13366
rect 5809 13363 5875 13366
rect 6913 13426 6979 13429
rect 8661 13426 8727 13429
rect 6913 13424 8727 13426
rect 6913 13368 6918 13424
rect 6974 13368 8666 13424
rect 8722 13368 8727 13424
rect 6913 13366 8727 13368
rect 6913 13363 6979 13366
rect 8661 13363 8727 13366
rect 9581 13426 9647 13429
rect 11462 13426 11468 13428
rect 9581 13424 11468 13426
rect 9581 13368 9586 13424
rect 9642 13368 11468 13424
rect 9581 13366 11468 13368
rect 9581 13363 9647 13366
rect 11462 13364 11468 13366
rect 11532 13364 11538 13428
rect 12566 13364 12572 13428
rect 12636 13426 12642 13428
rect 14460 13426 14520 13502
rect 16430 13500 16436 13502
rect 16500 13500 16506 13564
rect 17585 13562 17651 13565
rect 17718 13562 17724 13564
rect 17585 13560 17724 13562
rect 17585 13504 17590 13560
rect 17646 13504 17724 13560
rect 17585 13502 17724 13504
rect 17585 13499 17651 13502
rect 17718 13500 17724 13502
rect 17788 13500 17794 13564
rect 12636 13366 14520 13426
rect 12636 13364 12642 13366
rect 14590 13364 14596 13428
rect 14660 13426 14666 13428
rect 16614 13426 16620 13428
rect 14660 13366 16620 13426
rect 14660 13364 14666 13366
rect 16614 13364 16620 13366
rect 16684 13364 16690 13428
rect 2497 13290 2563 13293
rect 2630 13290 2636 13292
rect 2497 13288 2636 13290
rect 2497 13232 2502 13288
rect 2558 13232 2636 13288
rect 2497 13230 2636 13232
rect 2497 13227 2563 13230
rect 2630 13228 2636 13230
rect 2700 13228 2706 13292
rect 3969 13290 4035 13293
rect 4981 13292 5047 13293
rect 4102 13290 4108 13292
rect 3969 13288 4108 13290
rect 3969 13232 3974 13288
rect 4030 13232 4108 13288
rect 3969 13230 4108 13232
rect 3969 13227 4035 13230
rect 4102 13228 4108 13230
rect 4172 13228 4178 13292
rect 4981 13290 5028 13292
rect 4936 13288 5028 13290
rect 4936 13232 4986 13288
rect 4936 13230 5028 13232
rect 4981 13228 5028 13230
rect 5092 13228 5098 13292
rect 15929 13290 15995 13293
rect 5490 13288 15995 13290
rect 5490 13232 15934 13288
rect 15990 13232 15995 13288
rect 5490 13230 15995 13232
rect 4981 13227 5047 13228
rect -300 13154 160 13184
rect 1761 13154 1827 13157
rect 5490 13154 5550 13230
rect 15929 13227 15995 13230
rect 16246 13228 16252 13292
rect 16316 13290 16322 13292
rect 16665 13290 16731 13293
rect 16316 13288 16731 13290
rect 16316 13232 16670 13288
rect 16726 13232 16731 13288
rect 16316 13230 16731 13232
rect 16316 13228 16322 13230
rect 16665 13227 16731 13230
rect -300 13152 1827 13154
rect -300 13096 1766 13152
rect 1822 13096 1827 13152
rect -300 13094 1827 13096
rect -300 13064 160 13094
rect 1761 13091 1827 13094
rect 2776 13094 5550 13154
rect 6453 13154 6519 13157
rect 6729 13154 6795 13157
rect 6453 13152 6795 13154
rect 6453 13096 6458 13152
rect 6514 13096 6734 13152
rect 6790 13096 6795 13152
rect 6453 13094 6795 13096
rect 1301 13018 1367 13021
rect 2776 13018 2836 13094
rect 6453 13091 6519 13094
rect 6729 13091 6795 13094
rect 8293 13154 8359 13157
rect 10133 13154 10199 13157
rect 10409 13156 10475 13157
rect 10358 13154 10364 13156
rect 8293 13152 10199 13154
rect 8293 13096 8298 13152
rect 8354 13096 10138 13152
rect 10194 13096 10199 13152
rect 8293 13094 10199 13096
rect 10318 13094 10364 13154
rect 10428 13152 10475 13156
rect 10470 13096 10475 13152
rect 8293 13091 8359 13094
rect 10133 13091 10199 13094
rect 10358 13092 10364 13094
rect 10428 13092 10475 13096
rect 10409 13091 10475 13092
rect 11237 13154 11303 13157
rect 15101 13156 15167 13157
rect 14406 13154 14412 13156
rect 11237 13152 14412 13154
rect 11237 13096 11242 13152
rect 11298 13096 14412 13152
rect 11237 13094 14412 13096
rect 11237 13091 11303 13094
rect 14406 13092 14412 13094
rect 14476 13092 14482 13156
rect 15101 13154 15148 13156
rect 15056 13152 15148 13154
rect 15056 13096 15106 13152
rect 15056 13094 15148 13096
rect 15101 13092 15148 13094
rect 15212 13092 15218 13156
rect 15510 13092 15516 13156
rect 15580 13092 15586 13156
rect 21265 13154 21331 13157
rect 21840 13154 22300 13184
rect 21265 13152 22300 13154
rect 21265 13096 21270 13152
rect 21326 13096 22300 13152
rect 21265 13094 22300 13096
rect 15101 13091 15167 13092
rect 5890 13088 6206 13089
rect 5890 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6206 13088
rect 5890 13023 6206 13024
rect 10835 13088 11151 13089
rect 10835 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11151 13088
rect 10835 13023 11151 13024
rect 1301 13016 2836 13018
rect 1301 12960 1306 13016
rect 1362 12960 2836 13016
rect 1301 12958 2836 12960
rect 3233 13018 3299 13021
rect 3233 13016 4308 13018
rect 3233 12960 3238 13016
rect 3294 12960 4308 13016
rect 3233 12958 4308 12960
rect 1301 12955 1367 12958
rect 3233 12955 3299 12958
rect -300 12882 160 12912
rect 4061 12882 4127 12885
rect -300 12880 4127 12882
rect -300 12824 4066 12880
rect 4122 12824 4127 12880
rect -300 12822 4127 12824
rect 4248 12882 4308 12958
rect 4838 12956 4844 13020
rect 4908 13018 4914 13020
rect 4981 13018 5047 13021
rect 4908 13016 5047 13018
rect 4908 12960 4986 13016
rect 5042 12960 5047 13016
rect 4908 12958 5047 12960
rect 4908 12956 4914 12958
rect 4981 12955 5047 12958
rect 6361 13018 6427 13021
rect 7005 13018 7071 13021
rect 6361 13016 7071 13018
rect 6361 12960 6366 13016
rect 6422 12960 7010 13016
rect 7066 12960 7071 13016
rect 6361 12958 7071 12960
rect 6361 12955 6427 12958
rect 7005 12955 7071 12958
rect 11605 13018 11671 13021
rect 15518 13018 15578 13092
rect 21265 13091 21331 13094
rect 15780 13088 16096 13089
rect 15780 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16096 13088
rect 15780 13023 16096 13024
rect 20725 13088 21041 13089
rect 20725 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21041 13088
rect 21840 13064 22300 13094
rect 20725 13023 21041 13024
rect 11605 13016 15578 13018
rect 11605 12960 11610 13016
rect 11666 12960 15578 13016
rect 11605 12958 15578 12960
rect 11605 12955 11671 12958
rect 17677 12882 17743 12885
rect 4248 12880 17786 12882
rect 4248 12824 17682 12880
rect 17738 12824 17786 12880
rect 4248 12822 17786 12824
rect -300 12792 160 12822
rect 4061 12819 4127 12822
rect 17677 12819 17786 12822
rect 2262 12684 2268 12748
rect 2332 12746 2338 12748
rect 6361 12746 6427 12749
rect 2332 12744 6427 12746
rect 2332 12688 6366 12744
rect 6422 12688 6427 12744
rect 2332 12686 6427 12688
rect 2332 12684 2338 12686
rect 6361 12683 6427 12686
rect 8661 12746 8727 12749
rect 11421 12746 11487 12749
rect 16113 12746 16179 12749
rect 8661 12744 11487 12746
rect 8661 12688 8666 12744
rect 8722 12688 11426 12744
rect 11482 12688 11487 12744
rect 8661 12686 11487 12688
rect 8661 12683 8727 12686
rect 11421 12683 11487 12686
rect 11654 12744 16179 12746
rect 11654 12688 16118 12744
rect 16174 12688 16179 12744
rect 11654 12686 16179 12688
rect -300 12610 160 12640
rect 3877 12610 3943 12613
rect 4981 12610 5047 12613
rect -300 12550 2146 12610
rect -300 12520 160 12550
rect -300 12338 160 12368
rect 1669 12338 1735 12341
rect -300 12336 1735 12338
rect -300 12280 1674 12336
rect 1730 12280 1735 12336
rect -300 12278 1735 12280
rect -300 12248 160 12278
rect 1669 12275 1735 12278
rect -300 12066 160 12096
rect 1577 12066 1643 12069
rect -300 12064 1643 12066
rect -300 12008 1582 12064
rect 1638 12008 1643 12064
rect -300 12006 1643 12008
rect -300 11976 160 12006
rect 1577 12003 1643 12006
rect 2086 11930 2146 12550
rect 3877 12608 5047 12610
rect 3877 12552 3882 12608
rect 3938 12552 4986 12608
rect 5042 12552 5047 12608
rect 3877 12550 5047 12552
rect 3877 12547 3943 12550
rect 4981 12547 5047 12550
rect 5390 12548 5396 12612
rect 5460 12610 5466 12612
rect 5625 12610 5691 12613
rect 5460 12608 5691 12610
rect 5460 12552 5630 12608
rect 5686 12552 5691 12608
rect 5460 12550 5691 12552
rect 5460 12548 5466 12550
rect 5625 12547 5691 12550
rect 3418 12544 3734 12545
rect 3418 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3734 12544
rect 3418 12479 3734 12480
rect 8363 12544 8679 12545
rect 8363 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8679 12544
rect 8363 12479 8679 12480
rect 3785 12440 3851 12443
rect 3926 12440 4170 12474
rect 3785 12438 4170 12440
rect 3785 12382 3790 12438
rect 3846 12414 4170 12438
rect 3846 12382 3986 12414
rect 3785 12380 3986 12382
rect 3785 12377 3851 12380
rect 4110 12338 4170 12414
rect 5712 12412 5718 12476
rect 5782 12474 5788 12476
rect 10593 12474 10659 12477
rect 5782 12414 8264 12474
rect 5782 12412 5788 12414
rect 4889 12338 4955 12341
rect 4110 12336 4955 12338
rect 3742 12244 3986 12304
rect 4110 12280 4894 12336
rect 4950 12280 4955 12336
rect 4110 12278 4955 12280
rect 4889 12275 4955 12278
rect 5574 12276 5580 12340
rect 5644 12338 5650 12340
rect 7557 12338 7623 12341
rect 5644 12336 7623 12338
rect 5644 12280 7562 12336
rect 7618 12280 7623 12336
rect 5644 12278 7623 12280
rect 8204 12338 8264 12414
rect 10228 12472 10659 12474
rect 10228 12416 10598 12472
rect 10654 12416 10659 12472
rect 10228 12414 10659 12416
rect 10228 12338 10288 12414
rect 10593 12411 10659 12414
rect 11654 12338 11714 12686
rect 16113 12683 16179 12686
rect 16665 12746 16731 12749
rect 16798 12746 16804 12748
rect 16665 12744 16804 12746
rect 16665 12688 16670 12744
rect 16726 12688 16804 12744
rect 16665 12686 16804 12688
rect 16665 12683 16731 12686
rect 16798 12684 16804 12686
rect 16868 12684 16874 12748
rect 14733 12610 14799 12613
rect 16297 12610 16363 12613
rect 16941 12610 17007 12613
rect 14733 12608 17007 12610
rect 14733 12552 14738 12608
rect 14794 12552 16302 12608
rect 16358 12552 16946 12608
rect 17002 12552 17007 12608
rect 14733 12550 17007 12552
rect 14733 12547 14799 12550
rect 16297 12547 16363 12550
rect 16941 12547 17007 12550
rect 13308 12544 13624 12545
rect 13308 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13624 12544
rect 13308 12479 13624 12480
rect 13813 12474 13879 12477
rect 15285 12474 15351 12477
rect 13813 12472 15351 12474
rect 13813 12416 13818 12472
rect 13874 12416 15290 12472
rect 15346 12416 15351 12472
rect 13813 12414 15351 12416
rect 13813 12411 13879 12414
rect 15285 12411 15351 12414
rect 15653 12472 15719 12477
rect 16297 12476 16363 12477
rect 15653 12416 15658 12472
rect 15714 12416 15719 12472
rect 15653 12411 15719 12416
rect 16246 12412 16252 12476
rect 16316 12474 16363 12476
rect 17726 12474 17786 12819
rect 20294 12684 20300 12748
rect 20364 12746 20370 12748
rect 21633 12746 21699 12749
rect 20364 12744 21699 12746
rect 20364 12688 21638 12744
rect 21694 12688 21699 12744
rect 20364 12686 21699 12688
rect 20364 12684 20370 12686
rect 21633 12683 21699 12686
rect 19057 12610 19123 12613
rect 21840 12610 22300 12640
rect 19057 12608 22300 12610
rect 19057 12552 19062 12608
rect 19118 12552 22300 12608
rect 19057 12550 22300 12552
rect 19057 12547 19123 12550
rect 18253 12544 18569 12545
rect 18253 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18569 12544
rect 21840 12520 22300 12550
rect 18253 12479 18569 12480
rect 16316 12472 16408 12474
rect 16358 12416 16408 12472
rect 16316 12414 16408 12416
rect 17726 12414 18154 12474
rect 16316 12412 16363 12414
rect 16297 12411 16363 12412
rect 8204 12278 10288 12338
rect 10366 12278 11714 12338
rect 14089 12338 14155 12341
rect 15656 12338 15716 12411
rect 14089 12336 15716 12338
rect 14089 12280 14094 12336
rect 14150 12280 15716 12336
rect 14089 12278 15716 12280
rect 5644 12276 5650 12278
rect 7557 12275 7623 12278
rect 2589 12202 2655 12205
rect 3742 12202 3802 12244
rect 2589 12200 3802 12202
rect 2589 12144 2594 12200
rect 2650 12144 3802 12200
rect 2589 12142 3802 12144
rect 3926 12202 3986 12244
rect 10366 12202 10426 12278
rect 14089 12275 14155 12278
rect 17534 12276 17540 12340
rect 17604 12338 17610 12340
rect 17677 12338 17743 12341
rect 17604 12336 17743 12338
rect 17604 12280 17682 12336
rect 17738 12280 17743 12336
rect 17604 12278 17743 12280
rect 17604 12276 17610 12278
rect 17677 12275 17743 12278
rect 11053 12202 11119 12205
rect 3926 12142 10426 12202
rect 10504 12200 11119 12202
rect 10504 12144 11058 12200
rect 11114 12144 11119 12200
rect 10504 12142 11119 12144
rect 2589 12139 2655 12142
rect 2865 12066 2931 12069
rect 4429 12066 4495 12069
rect 2865 12064 4495 12066
rect 2865 12008 2870 12064
rect 2926 12008 4434 12064
rect 4490 12008 4495 12064
rect 2865 12006 4495 12008
rect 2865 12003 2931 12006
rect 4429 12003 4495 12006
rect 4838 12004 4844 12068
rect 4908 12066 4914 12068
rect 5349 12066 5415 12069
rect 4908 12064 5415 12066
rect 4908 12008 5354 12064
rect 5410 12008 5415 12064
rect 4908 12006 5415 12008
rect 4908 12004 4914 12006
rect 5349 12003 5415 12006
rect 5533 12066 5599 12069
rect 5717 12066 5783 12069
rect 5533 12064 5783 12066
rect 5533 12008 5538 12064
rect 5594 12008 5722 12064
rect 5778 12008 5783 12064
rect 5533 12006 5783 12008
rect 5533 12003 5599 12006
rect 5717 12003 5783 12006
rect 7598 12004 7604 12068
rect 7668 12066 7674 12068
rect 8569 12066 8635 12069
rect 10504 12066 10564 12142
rect 11053 12139 11119 12142
rect 11237 12202 11303 12205
rect 17309 12202 17375 12205
rect 11237 12200 17375 12202
rect 11237 12144 11242 12200
rect 11298 12144 17314 12200
rect 17370 12144 17375 12200
rect 11237 12142 17375 12144
rect 18094 12202 18154 12414
rect 19333 12202 19399 12205
rect 18094 12200 19399 12202
rect 18094 12144 19338 12200
rect 19394 12144 19399 12200
rect 18094 12142 19399 12144
rect 11237 12139 11303 12142
rect 17309 12139 17375 12142
rect 19333 12139 19399 12142
rect 19885 12202 19951 12205
rect 19885 12200 21282 12202
rect 19885 12144 19890 12200
rect 19946 12144 21282 12200
rect 19885 12142 21282 12144
rect 19885 12139 19951 12142
rect 7668 12064 10564 12066
rect 7668 12008 8574 12064
rect 8630 12008 10564 12064
rect 7668 12006 10564 12008
rect 7668 12004 7674 12006
rect 8569 12003 8635 12006
rect 11462 12004 11468 12068
rect 11532 12066 11538 12068
rect 13854 12066 13860 12068
rect 11532 12006 13860 12066
rect 11532 12004 11538 12006
rect 13854 12004 13860 12006
rect 13924 12004 13930 12068
rect 14406 12004 14412 12068
rect 14476 12066 14482 12068
rect 15285 12066 15351 12069
rect 14476 12064 15351 12066
rect 14476 12008 15290 12064
rect 15346 12008 15351 12064
rect 14476 12006 15351 12008
rect 14476 12004 14482 12006
rect 15285 12003 15351 12006
rect 16297 12066 16363 12069
rect 19558 12066 19564 12068
rect 16297 12064 19564 12066
rect 16297 12008 16302 12064
rect 16358 12008 19564 12064
rect 16297 12006 19564 12008
rect 16297 12003 16363 12006
rect 19558 12004 19564 12006
rect 19628 12004 19634 12068
rect 21222 12066 21282 12142
rect 21840 12066 22300 12096
rect 21222 12006 22300 12066
rect 5890 12000 6206 12001
rect 5890 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6206 12000
rect 5890 11935 6206 11936
rect 10835 12000 11151 12001
rect 10835 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11151 12000
rect 10835 11935 11151 11936
rect 15780 12000 16096 12001
rect 15780 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16096 12000
rect 15780 11935 16096 11936
rect 20725 12000 21041 12001
rect 20725 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21041 12000
rect 21840 11976 22300 12006
rect 20725 11935 21041 11936
rect 5533 11930 5599 11933
rect 11881 11930 11947 11933
rect 13261 11930 13327 11933
rect 2086 11928 5599 11930
rect 2086 11872 5538 11928
rect 5594 11872 5599 11928
rect 2086 11870 5599 11872
rect 5533 11867 5599 11870
rect 6686 11870 10610 11930
rect -300 11794 160 11824
rect 1853 11794 1919 11797
rect -300 11792 1919 11794
rect -300 11736 1858 11792
rect 1914 11736 1919 11792
rect -300 11734 1919 11736
rect -300 11704 160 11734
rect 1853 11731 1919 11734
rect 2446 11732 2452 11796
rect 2516 11794 2522 11796
rect 4061 11794 4127 11797
rect 5390 11794 5396 11796
rect 2516 11734 3848 11794
rect 2516 11732 2522 11734
rect 3788 11692 3848 11734
rect 4061 11792 5396 11794
rect 4061 11736 4066 11792
rect 4122 11736 5396 11792
rect 4061 11734 5396 11736
rect 4061 11731 4127 11734
rect 5390 11732 5396 11734
rect 5460 11732 5466 11796
rect 6177 11794 6243 11797
rect 6686 11794 6746 11870
rect 6177 11792 6746 11794
rect 6177 11736 6182 11792
rect 6238 11736 6746 11792
rect 6177 11734 6746 11736
rect 6821 11796 6887 11797
rect 6821 11792 6868 11796
rect 6932 11794 6938 11796
rect 9765 11794 9831 11797
rect 6821 11736 6826 11792
rect 6177 11731 6243 11734
rect 6821 11732 6868 11736
rect 6932 11734 6978 11794
rect 7606 11792 9831 11794
rect 7606 11736 9770 11792
rect 9826 11736 9831 11792
rect 7606 11734 9831 11736
rect 10550 11794 10610 11870
rect 11881 11928 13327 11930
rect 11881 11872 11886 11928
rect 11942 11872 13266 11928
rect 13322 11872 13327 11928
rect 11881 11870 13327 11872
rect 11881 11867 11947 11870
rect 13261 11867 13327 11870
rect 13905 11930 13971 11933
rect 14222 11930 14228 11932
rect 13905 11928 14228 11930
rect 13905 11872 13910 11928
rect 13966 11872 14228 11928
rect 13905 11870 14228 11872
rect 13905 11867 13971 11870
rect 14222 11868 14228 11870
rect 14292 11868 14298 11932
rect 17166 11868 17172 11932
rect 17236 11930 17242 11932
rect 17861 11930 17927 11933
rect 17236 11928 17927 11930
rect 17236 11872 17866 11928
rect 17922 11872 17927 11928
rect 17236 11870 17927 11872
rect 17236 11868 17242 11870
rect 17861 11867 17927 11870
rect 14641 11794 14707 11797
rect 10550 11792 14707 11794
rect 10550 11736 14646 11792
rect 14702 11736 14707 11792
rect 10550 11734 14707 11736
rect 6932 11732 6938 11734
rect 6821 11731 6887 11732
rect 3788 11658 3986 11692
rect 7414 11658 7420 11660
rect 3788 11632 7420 11658
rect 3926 11598 7420 11632
rect 7414 11596 7420 11598
rect 7484 11596 7490 11660
rect -300 11522 160 11552
rect 1945 11522 2011 11525
rect -300 11520 2011 11522
rect -300 11464 1950 11520
rect 2006 11464 2011 11520
rect -300 11462 2011 11464
rect -300 11432 160 11462
rect 1945 11459 2011 11462
rect 4153 11522 4219 11525
rect 4286 11522 4292 11524
rect 4153 11520 4292 11522
rect 4153 11464 4158 11520
rect 4214 11464 4292 11520
rect 4153 11462 4292 11464
rect 4153 11459 4219 11462
rect 4286 11460 4292 11462
rect 4356 11460 4362 11524
rect 4521 11522 4587 11525
rect 4889 11522 4955 11525
rect 7606 11522 7666 11734
rect 9765 11731 9831 11734
rect 14641 11731 14707 11734
rect 14958 11732 14964 11796
rect 15028 11794 15034 11796
rect 15101 11794 15167 11797
rect 15377 11796 15443 11797
rect 15326 11794 15332 11796
rect 15028 11792 15167 11794
rect 15028 11736 15106 11792
rect 15162 11736 15167 11792
rect 15028 11734 15167 11736
rect 15286 11734 15332 11794
rect 15396 11792 15443 11796
rect 15438 11736 15443 11792
rect 15028 11732 15034 11734
rect 15101 11731 15167 11734
rect 15326 11732 15332 11734
rect 15396 11732 15443 11736
rect 15510 11732 15516 11796
rect 15580 11794 15586 11796
rect 15580 11734 19350 11794
rect 15580 11732 15586 11734
rect 15377 11731 15443 11732
rect 8017 11658 8083 11661
rect 10225 11658 10291 11661
rect 8017 11656 10291 11658
rect 8017 11600 8022 11656
rect 8078 11600 10230 11656
rect 10286 11600 10291 11656
rect 8017 11598 10291 11600
rect 8017 11595 8083 11598
rect 10225 11595 10291 11598
rect 11881 11658 11947 11661
rect 17769 11658 17835 11661
rect 11881 11656 17835 11658
rect 11881 11600 11886 11656
rect 11942 11600 17774 11656
rect 17830 11600 17835 11656
rect 11881 11598 17835 11600
rect 19290 11658 19350 11734
rect 19793 11658 19859 11661
rect 19290 11656 19859 11658
rect 19290 11600 19798 11656
rect 19854 11600 19859 11656
rect 19290 11598 19859 11600
rect 11881 11595 11947 11598
rect 17769 11595 17835 11598
rect 19793 11595 19859 11598
rect 4521 11520 4955 11522
rect 4521 11464 4526 11520
rect 4582 11464 4894 11520
rect 4950 11464 4955 11520
rect 4521 11462 4955 11464
rect 4521 11459 4587 11462
rect 4889 11459 4955 11462
rect 5582 11462 7666 11522
rect 13721 11522 13787 11525
rect 16246 11522 16252 11524
rect 13721 11520 16252 11522
rect 13721 11464 13726 11520
rect 13782 11464 16252 11520
rect 13721 11462 16252 11464
rect 3418 11456 3734 11457
rect 3418 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3734 11456
rect 3418 11391 3734 11392
rect 4889 11386 4955 11389
rect 5441 11386 5507 11389
rect 4889 11384 5507 11386
rect 4889 11328 4894 11384
rect 4950 11328 5446 11384
rect 5502 11328 5507 11384
rect 4889 11326 5507 11328
rect 4889 11323 4955 11326
rect 5441 11323 5507 11326
rect -300 11250 160 11280
rect 4061 11250 4127 11253
rect -300 11248 4127 11250
rect -300 11192 4066 11248
rect 4122 11192 4127 11248
rect -300 11190 4127 11192
rect -300 11160 160 11190
rect 4061 11187 4127 11190
rect 4521 11250 4587 11253
rect 5582 11250 5642 11462
rect 13721 11459 13787 11462
rect 16246 11460 16252 11462
rect 16316 11460 16322 11524
rect 16614 11460 16620 11524
rect 16684 11522 16690 11524
rect 17217 11522 17283 11525
rect 16684 11520 17283 11522
rect 16684 11464 17222 11520
rect 17278 11464 17283 11520
rect 16684 11462 17283 11464
rect 16684 11460 16690 11462
rect 17217 11459 17283 11462
rect 19425 11522 19491 11525
rect 21840 11522 22300 11552
rect 19425 11520 22300 11522
rect 19425 11464 19430 11520
rect 19486 11464 22300 11520
rect 19425 11462 22300 11464
rect 19425 11459 19491 11462
rect 8363 11456 8679 11457
rect 8363 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8679 11456
rect 8363 11391 8679 11392
rect 13308 11456 13624 11457
rect 13308 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13624 11456
rect 13308 11391 13624 11392
rect 18253 11456 18569 11457
rect 18253 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18569 11456
rect 21840 11432 22300 11462
rect 18253 11391 18569 11392
rect 6085 11386 6151 11389
rect 7005 11386 7071 11389
rect 6085 11384 7071 11386
rect 6085 11328 6090 11384
rect 6146 11328 7010 11384
rect 7066 11328 7071 11384
rect 6085 11326 7071 11328
rect 6085 11323 6151 11326
rect 7005 11323 7071 11326
rect 8748 11324 8754 11388
rect 8818 11386 8824 11388
rect 13077 11386 13143 11389
rect 8818 11384 13143 11386
rect 8818 11328 13082 11384
rect 13138 11328 13143 11384
rect 8818 11326 13143 11328
rect 8818 11324 8824 11326
rect 13077 11323 13143 11326
rect 14089 11386 14155 11389
rect 17953 11386 18019 11389
rect 14089 11384 18019 11386
rect 14089 11328 14094 11384
rect 14150 11328 17958 11384
rect 18014 11328 18019 11384
rect 14089 11326 18019 11328
rect 14089 11323 14155 11326
rect 17953 11323 18019 11326
rect 9213 11250 9279 11253
rect 4521 11248 5642 11250
rect 4521 11192 4526 11248
rect 4582 11192 5642 11248
rect 4521 11190 5642 11192
rect 5766 11248 9279 11250
rect 5766 11192 9218 11248
rect 9274 11192 9279 11248
rect 5766 11190 9279 11192
rect 4521 11187 4587 11190
rect 2037 11114 2103 11117
rect 2497 11116 2563 11117
rect 2262 11114 2268 11116
rect 2037 11112 2268 11114
rect 2037 11056 2042 11112
rect 2098 11056 2268 11112
rect 2037 11054 2268 11056
rect 2037 11051 2103 11054
rect 2262 11052 2268 11054
rect 2332 11052 2338 11116
rect 2446 11052 2452 11116
rect 2516 11114 2563 11116
rect 4797 11116 4863 11117
rect 4797 11114 4844 11116
rect 2516 11112 2608 11114
rect 2558 11056 2608 11112
rect 2516 11054 2608 11056
rect 4752 11112 4844 11114
rect 4752 11056 4802 11112
rect 4752 11054 4844 11056
rect 2516 11052 2563 11054
rect 2497 11051 2563 11052
rect 4797 11052 4844 11054
rect 4908 11052 4914 11116
rect 5165 11114 5231 11117
rect 5441 11114 5507 11117
rect 5165 11112 5507 11114
rect 5165 11056 5170 11112
rect 5226 11056 5446 11112
rect 5502 11056 5507 11112
rect 5165 11054 5507 11056
rect 4797 11051 4863 11052
rect 5165 11051 5231 11054
rect 5441 11051 5507 11054
rect -300 10978 160 11008
rect 841 10978 907 10981
rect -300 10976 907 10978
rect -300 10920 846 10976
rect 902 10920 907 10976
rect -300 10918 907 10920
rect -300 10888 160 10918
rect 841 10915 907 10918
rect 1393 10978 1459 10981
rect 1526 10978 1532 10980
rect 1393 10976 1532 10978
rect 1393 10920 1398 10976
rect 1454 10920 1532 10976
rect 1393 10918 1532 10920
rect 1393 10915 1459 10918
rect 1526 10916 1532 10918
rect 1596 10916 1602 10980
rect 2497 10978 2563 10981
rect 2497 10976 4170 10978
rect 2497 10920 2502 10976
rect 2558 10920 4170 10976
rect 2497 10918 4170 10920
rect 2497 10915 2563 10918
rect 2221 10842 2287 10845
rect 2086 10840 2287 10842
rect 2086 10784 2226 10840
rect 2282 10784 2287 10840
rect 2086 10782 2287 10784
rect 4110 10842 4170 10918
rect 4286 10916 4292 10980
rect 4356 10978 4362 10980
rect 4521 10978 4587 10981
rect 4889 10980 4955 10981
rect 4356 10976 4587 10978
rect 4356 10920 4526 10976
rect 4582 10920 4587 10976
rect 4356 10918 4587 10920
rect 4356 10916 4362 10918
rect 4521 10915 4587 10918
rect 4838 10916 4844 10980
rect 4908 10978 4955 10980
rect 4908 10976 5000 10978
rect 4950 10920 5000 10976
rect 4908 10918 5000 10920
rect 4908 10916 4955 10918
rect 4889 10915 4955 10916
rect 5766 10842 5826 11190
rect 9213 11187 9279 11190
rect 12014 11188 12020 11252
rect 12084 11250 12090 11252
rect 18965 11250 19031 11253
rect 12084 11248 19031 11250
rect 12084 11192 18970 11248
rect 19026 11192 19031 11248
rect 12084 11190 19031 11192
rect 12084 11188 12090 11190
rect 18965 11187 19031 11190
rect 6361 11114 6427 11117
rect 6545 11114 6611 11117
rect 6361 11112 6611 11114
rect 6361 11056 6366 11112
rect 6422 11056 6550 11112
rect 6606 11056 6611 11112
rect 6361 11054 6611 11056
rect 6361 11051 6427 11054
rect 6545 11051 6611 11054
rect 6862 11052 6868 11116
rect 6932 11114 6938 11116
rect 10409 11114 10475 11117
rect 12065 11114 12131 11117
rect 19057 11114 19123 11117
rect 6932 11112 10475 11114
rect 6932 11056 10414 11112
rect 10470 11056 10475 11112
rect 6932 11054 10475 11056
rect 6932 11052 6938 11054
rect 10409 11051 10475 11054
rect 10550 11054 11346 11114
rect 7097 10978 7163 10981
rect 7649 10978 7715 10981
rect 10550 10978 10610 11054
rect 7097 10976 10610 10978
rect 7097 10920 7102 10976
rect 7158 10920 7654 10976
rect 7710 10920 10610 10976
rect 7097 10918 10610 10920
rect 11286 10978 11346 11054
rect 12065 11112 19123 11114
rect 12065 11056 12070 11112
rect 12126 11056 19062 11112
rect 19118 11056 19123 11112
rect 12065 11054 19123 11056
rect 12065 11051 12131 11054
rect 19057 11051 19123 11054
rect 14089 10978 14155 10981
rect 15653 10978 15719 10981
rect 18781 10980 18847 10981
rect 18781 10978 18828 10980
rect 11286 10918 13922 10978
rect 7097 10915 7163 10918
rect 7649 10915 7715 10918
rect 5890 10912 6206 10913
rect 5890 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6206 10912
rect 5890 10847 6206 10848
rect 10835 10912 11151 10913
rect 10835 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11151 10912
rect 10835 10847 11151 10848
rect 4110 10782 5826 10842
rect 7649 10842 7715 10845
rect 10685 10842 10751 10845
rect 11605 10844 11671 10845
rect 13862 10844 13922 10918
rect 14089 10976 15719 10978
rect 14089 10920 14094 10976
rect 14150 10920 15658 10976
rect 15714 10920 15719 10976
rect 14089 10918 15719 10920
rect 18736 10976 18828 10978
rect 18736 10920 18786 10976
rect 18736 10918 18828 10920
rect 14089 10915 14155 10918
rect 15653 10915 15719 10918
rect 18781 10916 18828 10918
rect 18892 10916 18898 10980
rect 21265 10978 21331 10981
rect 21840 10978 22300 11008
rect 21265 10976 22300 10978
rect 21265 10920 21270 10976
rect 21326 10920 22300 10976
rect 21265 10918 22300 10920
rect 18781 10915 18847 10916
rect 21265 10915 21331 10918
rect 15780 10912 16096 10913
rect 15780 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16096 10912
rect 15780 10847 16096 10848
rect 20725 10912 21041 10913
rect 20725 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21041 10912
rect 21840 10888 22300 10918
rect 20725 10847 21041 10848
rect 11605 10842 11652 10844
rect 7649 10840 10751 10842
rect 7649 10784 7654 10840
rect 7710 10784 10690 10840
rect 10746 10784 10751 10840
rect 7649 10782 10751 10784
rect 11560 10840 11652 10842
rect 11560 10784 11610 10840
rect 11560 10782 11652 10784
rect -300 10706 160 10736
rect 1025 10706 1091 10709
rect -300 10704 1091 10706
rect -300 10648 1030 10704
rect 1086 10648 1091 10704
rect -300 10646 1091 10648
rect -300 10616 160 10646
rect 1025 10643 1091 10646
rect 2086 10570 2146 10782
rect 2221 10779 2287 10782
rect 7649 10779 7715 10782
rect 10685 10779 10751 10782
rect 11605 10780 11652 10782
rect 11716 10780 11722 10844
rect 13854 10780 13860 10844
rect 13924 10780 13930 10844
rect 14089 10842 14155 10845
rect 15285 10842 15351 10845
rect 14089 10840 15351 10842
rect 14089 10784 14094 10840
rect 14150 10784 15290 10840
rect 15346 10784 15351 10840
rect 14089 10782 15351 10784
rect 11605 10779 11671 10780
rect 14089 10779 14155 10782
rect 15285 10779 15351 10782
rect 16205 10842 16271 10845
rect 16205 10840 17602 10842
rect 16205 10784 16210 10840
rect 16266 10784 17602 10840
rect 16205 10782 17602 10784
rect 16205 10779 16271 10782
rect 3969 10708 4035 10709
rect 2262 10644 2268 10708
rect 2332 10706 2338 10708
rect 2998 10706 3004 10708
rect 2332 10646 3004 10706
rect 2332 10644 2338 10646
rect 2998 10644 3004 10646
rect 3068 10644 3074 10708
rect 3918 10706 3924 10708
rect 3878 10646 3924 10706
rect 3988 10704 4035 10708
rect 4030 10648 4035 10704
rect 3918 10644 3924 10646
rect 3988 10644 4035 10648
rect 5022 10644 5028 10708
rect 5092 10706 5098 10708
rect 8017 10706 8083 10709
rect 5092 10704 8083 10706
rect 5092 10648 8022 10704
rect 8078 10648 8083 10704
rect 5092 10646 8083 10648
rect 5092 10644 5098 10646
rect 3969 10643 4035 10644
rect 8017 10643 8083 10646
rect 10041 10706 10107 10709
rect 11462 10706 11468 10708
rect 10041 10704 11468 10706
rect 10041 10648 10046 10704
rect 10102 10648 11468 10704
rect 10041 10646 11468 10648
rect 10041 10643 10107 10646
rect 11462 10644 11468 10646
rect 11532 10644 11538 10708
rect 11789 10706 11855 10709
rect 17033 10706 17099 10709
rect 17542 10708 17602 10782
rect 11789 10704 17099 10706
rect 11789 10648 11794 10704
rect 11850 10648 17038 10704
rect 17094 10648 17099 10704
rect 11789 10646 17099 10648
rect 11789 10643 11855 10646
rect 17033 10643 17099 10646
rect 17534 10644 17540 10708
rect 17604 10644 17610 10708
rect 2221 10570 2287 10573
rect 2086 10568 2287 10570
rect 2086 10512 2226 10568
rect 2282 10512 2287 10568
rect 2086 10510 2287 10512
rect 2221 10507 2287 10510
rect 2998 10508 3004 10572
rect 3068 10570 3074 10572
rect 11237 10570 11303 10573
rect 3068 10568 11303 10570
rect 3068 10512 11242 10568
rect 11298 10512 11303 10568
rect 3068 10510 11303 10512
rect 3068 10508 3074 10510
rect 11237 10507 11303 10510
rect 11830 10508 11836 10572
rect 11900 10570 11906 10572
rect 14038 10570 14044 10572
rect 11900 10510 14044 10570
rect 11900 10508 11906 10510
rect 14038 10508 14044 10510
rect 14108 10508 14114 10572
rect 14406 10508 14412 10572
rect 14476 10570 14482 10572
rect 15510 10570 15516 10572
rect 14476 10510 15516 10570
rect 14476 10508 14482 10510
rect 15510 10508 15516 10510
rect 15580 10508 15586 10572
rect 16297 10570 16363 10573
rect 20161 10570 20227 10573
rect 16297 10568 20227 10570
rect 16297 10512 16302 10568
rect 16358 10512 20166 10568
rect 20222 10512 20227 10568
rect 16297 10510 20227 10512
rect 16297 10507 16363 10510
rect 20161 10507 20227 10510
rect -300 10434 160 10464
rect 2313 10434 2379 10437
rect -300 10432 2379 10434
rect -300 10376 2318 10432
rect 2374 10376 2379 10432
rect -300 10374 2379 10376
rect -300 10344 160 10374
rect 2313 10371 2379 10374
rect 5533 10436 5599 10437
rect 5533 10432 5580 10436
rect 5644 10434 5650 10436
rect 6821 10434 6887 10437
rect 7189 10434 7255 10437
rect 8017 10436 8083 10437
rect 7966 10434 7972 10436
rect 5533 10376 5538 10432
rect 5533 10372 5580 10376
rect 5644 10374 5690 10434
rect 6821 10432 7255 10434
rect 6821 10376 6826 10432
rect 6882 10376 7194 10432
rect 7250 10376 7255 10432
rect 6821 10374 7255 10376
rect 7926 10374 7972 10434
rect 8036 10432 8083 10436
rect 8078 10376 8083 10432
rect 5644 10372 5650 10374
rect 5533 10371 5599 10372
rect 6821 10371 6887 10374
rect 7189 10371 7255 10374
rect 7966 10372 7972 10374
rect 8036 10372 8083 10376
rect 8886 10372 8892 10436
rect 8956 10434 8962 10436
rect 9121 10434 9187 10437
rect 9438 10434 9444 10436
rect 8956 10432 9187 10434
rect 8956 10376 9126 10432
rect 9182 10376 9187 10432
rect 8956 10374 9187 10376
rect 8956 10372 8962 10374
rect 8017 10371 8083 10372
rect 9121 10371 9187 10374
rect 9262 10374 9444 10434
rect 3418 10368 3734 10369
rect 3418 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3734 10368
rect 3418 10303 3734 10304
rect 8363 10368 8679 10369
rect 8363 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8679 10368
rect 8363 10303 8679 10304
rect 2589 10300 2655 10301
rect 2589 10298 2636 10300
rect 2544 10296 2636 10298
rect 2544 10240 2594 10296
rect 2544 10238 2636 10240
rect 2589 10236 2636 10238
rect 2700 10236 2706 10300
rect 3969 10298 4035 10301
rect 4102 10298 4108 10300
rect 3969 10296 4108 10298
rect 3969 10240 3974 10296
rect 4030 10240 4108 10296
rect 3969 10238 4108 10240
rect 2589 10235 2655 10236
rect 3969 10235 4035 10238
rect 4102 10236 4108 10238
rect 4172 10236 4178 10300
rect 5390 10236 5396 10300
rect 5460 10298 5466 10300
rect 5460 10238 8218 10298
rect 5460 10236 5466 10238
rect -300 10162 160 10192
rect -300 10102 4170 10162
rect -300 10072 160 10102
rect 1894 9964 1900 10028
rect 1964 10026 1970 10028
rect 4110 10026 4170 10102
rect 4521 10026 4587 10029
rect 7649 10026 7715 10029
rect 7966 10026 7972 10028
rect 1964 9966 2330 10026
rect 4110 10024 4587 10026
rect 4110 9968 4526 10024
rect 4582 9968 4587 10024
rect 4110 9966 4587 9968
rect 1964 9964 1970 9966
rect -300 9890 160 9920
rect 2270 9890 2330 9966
rect 4521 9963 4587 9966
rect 5628 9966 6378 10026
rect 4705 9890 4771 9893
rect -300 9830 2146 9890
rect 2270 9888 4771 9890
rect 2270 9832 4710 9888
rect 4766 9832 4771 9888
rect 2270 9830 4771 9832
rect -300 9800 160 9830
rect 2086 9754 2146 9830
rect 4705 9827 4771 9830
rect 4061 9754 4127 9757
rect 5628 9754 5688 9966
rect 6318 9890 6378 9966
rect 7649 10024 7972 10026
rect 7649 9968 7654 10024
rect 7710 9968 7972 10024
rect 7649 9966 7972 9968
rect 7649 9963 7715 9966
rect 7966 9964 7972 9966
rect 8036 9964 8042 10028
rect 8158 10026 8218 10238
rect 8886 10236 8892 10300
rect 8956 10236 8962 10300
rect 9070 10236 9076 10300
rect 9140 10298 9146 10300
rect 9262 10298 9322 10374
rect 9438 10372 9444 10374
rect 9508 10372 9514 10436
rect 10680 10372 10686 10436
rect 10750 10434 10756 10436
rect 11237 10434 11303 10437
rect 10750 10432 11303 10434
rect 10750 10376 11242 10432
rect 11298 10376 11303 10432
rect 10750 10374 11303 10376
rect 10750 10372 10756 10374
rect 11237 10371 11303 10374
rect 11462 10372 11468 10436
rect 11532 10434 11538 10436
rect 12801 10434 12867 10437
rect 11532 10432 12867 10434
rect 11532 10376 12806 10432
rect 12862 10376 12867 10432
rect 11532 10374 12867 10376
rect 11532 10372 11538 10374
rect 12801 10371 12867 10374
rect 13721 10434 13787 10437
rect 17769 10434 17835 10437
rect 20529 10434 20595 10437
rect 21840 10434 22300 10464
rect 13721 10432 17970 10434
rect 13721 10376 13726 10432
rect 13782 10376 17774 10432
rect 17830 10376 17970 10432
rect 13721 10374 17970 10376
rect 13721 10371 13787 10374
rect 17769 10371 17835 10374
rect 13308 10368 13624 10369
rect 13308 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13624 10368
rect 13308 10303 13624 10304
rect 9140 10238 9322 10298
rect 9140 10236 9146 10238
rect 9438 10236 9444 10300
rect 9508 10298 9514 10300
rect 12750 10298 12756 10300
rect 9508 10238 12756 10298
rect 9508 10236 9514 10238
rect 12750 10236 12756 10238
rect 12820 10236 12826 10300
rect 17033 10298 17099 10301
rect 13862 10296 17099 10298
rect 13862 10240 17038 10296
rect 17094 10240 17099 10296
rect 13862 10238 17099 10240
rect 8753 10162 8819 10165
rect 8894 10162 8954 10236
rect 8753 10160 8954 10162
rect 8753 10104 8758 10160
rect 8814 10104 8954 10160
rect 8753 10102 8954 10104
rect 9765 10162 9831 10165
rect 13862 10162 13922 10238
rect 17033 10235 17099 10238
rect 14457 10164 14523 10165
rect 14406 10162 14412 10164
rect 9765 10160 13922 10162
rect 9765 10104 9770 10160
rect 9826 10104 13922 10160
rect 9765 10102 13922 10104
rect 14366 10102 14412 10162
rect 14476 10160 14523 10164
rect 14518 10104 14523 10160
rect 8753 10099 8819 10102
rect 9765 10099 9831 10102
rect 14406 10100 14412 10102
rect 14476 10100 14523 10104
rect 14457 10099 14523 10100
rect 14641 10162 14707 10165
rect 17166 10162 17172 10164
rect 14641 10160 17172 10162
rect 14641 10104 14646 10160
rect 14702 10104 17172 10160
rect 14641 10102 17172 10104
rect 14641 10099 14707 10102
rect 17166 10100 17172 10102
rect 17236 10100 17242 10164
rect 17910 10162 17970 10374
rect 20529 10432 22300 10434
rect 20529 10376 20534 10432
rect 20590 10376 22300 10432
rect 20529 10374 22300 10376
rect 20529 10371 20595 10374
rect 18253 10368 18569 10369
rect 18253 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18569 10368
rect 21840 10344 22300 10374
rect 18253 10303 18569 10304
rect 18822 10162 18828 10164
rect 17910 10102 18828 10162
rect 18822 10100 18828 10102
rect 18892 10100 18898 10164
rect 17677 10026 17743 10029
rect 17861 10028 17927 10029
rect 17861 10026 17908 10028
rect 8158 10024 17743 10026
rect 8158 9968 17682 10024
rect 17738 9968 17743 10024
rect 8158 9966 17743 9968
rect 17816 10024 17908 10026
rect 17816 9968 17866 10024
rect 17816 9966 17908 9968
rect 17677 9963 17743 9966
rect 17861 9964 17908 9966
rect 17972 9964 17978 10028
rect 18086 9964 18092 10028
rect 18156 10026 18162 10028
rect 18505 10026 18571 10029
rect 18156 10024 18571 10026
rect 18156 9968 18510 10024
rect 18566 9968 18571 10024
rect 18156 9966 18571 9968
rect 18156 9964 18162 9966
rect 17861 9963 17927 9964
rect 18505 9963 18571 9966
rect 18689 10026 18755 10029
rect 18689 10024 21282 10026
rect 18689 9968 18694 10024
rect 18750 9968 21282 10024
rect 18689 9966 21282 9968
rect 18689 9963 18755 9966
rect 8201 9890 8267 9893
rect 10133 9890 10199 9893
rect 6318 9888 8267 9890
rect 6318 9832 8206 9888
rect 8262 9832 8267 9888
rect 6318 9830 8267 9832
rect 8201 9827 8267 9830
rect 8342 9888 10199 9890
rect 8342 9832 10138 9888
rect 10194 9832 10199 9888
rect 8342 9830 10199 9832
rect 5890 9824 6206 9825
rect 5890 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6206 9824
rect 5890 9759 6206 9760
rect 8342 9757 8402 9830
rect 10133 9827 10199 9830
rect 11237 9890 11303 9893
rect 12525 9890 12591 9893
rect 12801 9892 12867 9893
rect 12750 9890 12756 9892
rect 11237 9888 12591 9890
rect 11237 9832 11242 9888
rect 11298 9832 12530 9888
rect 12586 9832 12591 9888
rect 11237 9830 12591 9832
rect 12710 9830 12756 9890
rect 12820 9888 12867 9892
rect 12862 9832 12867 9888
rect 11237 9827 11303 9830
rect 12525 9827 12591 9830
rect 12750 9828 12756 9830
rect 12820 9828 12867 9832
rect 12801 9827 12867 9828
rect 13077 9890 13143 9893
rect 15653 9890 15719 9893
rect 13077 9888 15719 9890
rect 13077 9832 13082 9888
rect 13138 9832 15658 9888
rect 15714 9832 15719 9888
rect 13077 9830 15719 9832
rect 13077 9827 13143 9830
rect 15653 9827 15719 9830
rect 16297 9890 16363 9893
rect 19701 9890 19767 9893
rect 16297 9888 19767 9890
rect 16297 9832 16302 9888
rect 16358 9832 19706 9888
rect 19762 9832 19767 9888
rect 16297 9830 19767 9832
rect 21222 9890 21282 9966
rect 21840 9890 22300 9920
rect 21222 9830 22300 9890
rect 16297 9827 16363 9830
rect 19701 9827 19767 9830
rect 10835 9824 11151 9825
rect 10835 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11151 9824
rect 10835 9759 11151 9760
rect 15780 9824 16096 9825
rect 15780 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16096 9824
rect 15780 9759 16096 9760
rect 20725 9824 21041 9825
rect 20725 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21041 9824
rect 21840 9800 22300 9830
rect 20725 9759 21041 9760
rect 2086 9752 4127 9754
rect 2086 9696 4066 9752
rect 4122 9696 4127 9752
rect 2086 9694 4127 9696
rect 4061 9691 4127 9694
rect 5352 9694 5688 9754
rect 7189 9754 7255 9757
rect 7649 9754 7715 9757
rect 8109 9756 8175 9757
rect 8109 9754 8156 9756
rect 7189 9752 7715 9754
rect 7189 9696 7194 9752
rect 7250 9696 7654 9752
rect 7710 9696 7715 9752
rect 7189 9694 7715 9696
rect 8064 9752 8156 9754
rect 8064 9696 8114 9752
rect 8064 9694 8156 9696
rect -300 9618 160 9648
rect 5352 9621 5412 9694
rect 7189 9691 7255 9694
rect 7649 9691 7715 9694
rect 8109 9692 8156 9694
rect 8220 9692 8226 9756
rect 8293 9752 8402 9757
rect 8293 9696 8298 9752
rect 8354 9696 8402 9752
rect 8293 9694 8402 9696
rect 8661 9754 8727 9757
rect 10317 9754 10383 9757
rect 8661 9752 10383 9754
rect 8661 9696 8666 9752
rect 8722 9696 10322 9752
rect 10378 9696 10383 9752
rect 8661 9694 10383 9696
rect 8109 9691 8175 9692
rect 8293 9691 8359 9694
rect 8661 9691 8727 9694
rect 10317 9691 10383 9694
rect 11646 9692 11652 9756
rect 11716 9754 11722 9756
rect 19425 9754 19491 9757
rect 11716 9694 15716 9754
rect 11716 9692 11722 9694
rect 1301 9618 1367 9621
rect -300 9616 1367 9618
rect -300 9560 1306 9616
rect 1362 9560 1367 9616
rect -300 9558 1367 9560
rect -300 9528 160 9558
rect 1301 9555 1367 9558
rect 2630 9556 2636 9620
rect 2700 9618 2706 9620
rect 2773 9618 2839 9621
rect 3325 9618 3391 9621
rect 2700 9616 2839 9618
rect 2700 9560 2778 9616
rect 2834 9560 2839 9616
rect 2700 9558 2839 9560
rect 2700 9556 2706 9558
rect 2773 9555 2839 9558
rect 3006 9616 3391 9618
rect 3006 9560 3330 9616
rect 3386 9560 3391 9616
rect 3006 9558 3391 9560
rect 1342 9420 1348 9484
rect 1412 9482 1418 9484
rect 3006 9482 3066 9558
rect 3325 9555 3391 9558
rect 4153 9618 4219 9621
rect 4470 9618 4476 9620
rect 4153 9616 4476 9618
rect 4153 9560 4158 9616
rect 4214 9560 4476 9616
rect 4153 9558 4476 9560
rect 4153 9555 4219 9558
rect 4470 9556 4476 9558
rect 4540 9556 4546 9620
rect 5349 9616 5415 9621
rect 5349 9560 5354 9616
rect 5410 9560 5415 9616
rect 5349 9555 5415 9560
rect 6177 9618 6243 9621
rect 6913 9618 6979 9621
rect 10501 9618 10567 9621
rect 6177 9616 10567 9618
rect 6177 9560 6182 9616
rect 6238 9560 6918 9616
rect 6974 9560 10506 9616
rect 10562 9560 10567 9616
rect 6177 9558 10567 9560
rect 6177 9555 6243 9558
rect 6913 9555 6979 9558
rect 10501 9555 10567 9558
rect 10961 9618 11027 9621
rect 15285 9618 15351 9621
rect 10961 9616 15351 9618
rect 10961 9560 10966 9616
rect 11022 9560 15290 9616
rect 15346 9560 15351 9616
rect 10961 9558 15351 9560
rect 15656 9618 15716 9694
rect 19290 9752 19491 9754
rect 19290 9696 19430 9752
rect 19486 9696 19491 9752
rect 19290 9694 19491 9696
rect 19290 9618 19350 9694
rect 19425 9691 19491 9694
rect 15656 9558 19350 9618
rect 10961 9555 11027 9558
rect 15285 9555 15351 9558
rect 5073 9484 5139 9485
rect 1412 9422 3066 9482
rect 1412 9420 1418 9422
rect 3182 9420 3188 9484
rect 3252 9482 3258 9484
rect 3252 9422 4170 9482
rect 3252 9420 3258 9422
rect -300 9346 160 9376
rect 1577 9346 1643 9349
rect -300 9344 1643 9346
rect -300 9288 1582 9344
rect 1638 9288 1643 9344
rect -300 9286 1643 9288
rect -300 9256 160 9286
rect 1577 9283 1643 9286
rect 2814 9284 2820 9348
rect 2884 9346 2890 9348
rect 3233 9346 3299 9349
rect 2884 9344 3299 9346
rect 2884 9288 3238 9344
rect 3294 9288 3299 9344
rect 2884 9286 3299 9288
rect 4110 9346 4170 9422
rect 5022 9420 5028 9484
rect 5092 9482 5139 9484
rect 5993 9482 6059 9485
rect 7281 9482 7347 9485
rect 5092 9480 5184 9482
rect 5134 9424 5184 9480
rect 5092 9422 5184 9424
rect 5993 9480 7347 9482
rect 5993 9424 5998 9480
rect 6054 9424 7286 9480
rect 7342 9424 7347 9480
rect 5993 9422 7347 9424
rect 5092 9420 5139 9422
rect 5073 9419 5139 9420
rect 5993 9419 6059 9422
rect 7281 9419 7347 9422
rect 7465 9482 7531 9485
rect 7782 9482 7788 9484
rect 7465 9480 7788 9482
rect 7465 9424 7470 9480
rect 7526 9424 7788 9480
rect 7465 9422 7788 9424
rect 7465 9419 7531 9422
rect 7782 9420 7788 9422
rect 7852 9420 7858 9484
rect 14181 9482 14247 9485
rect 15142 9482 15148 9484
rect 8158 9422 14060 9482
rect 5022 9346 5028 9348
rect 4110 9286 5028 9346
rect 2884 9284 2890 9286
rect 3233 9283 3299 9286
rect 5022 9284 5028 9286
rect 5092 9284 5098 9348
rect 5349 9346 5415 9349
rect 8158 9346 8218 9422
rect 14000 9349 14060 9422
rect 14181 9480 15148 9482
rect 14181 9424 14186 9480
rect 14242 9424 15148 9480
rect 14181 9422 15148 9424
rect 14181 9419 14247 9422
rect 15142 9420 15148 9422
rect 15212 9420 15218 9484
rect 15653 9482 15719 9485
rect 19885 9482 19951 9485
rect 15653 9480 19951 9482
rect 15653 9424 15658 9480
rect 15714 9424 19890 9480
rect 19946 9424 19951 9480
rect 15653 9422 19951 9424
rect 15653 9419 15719 9422
rect 19885 9419 19951 9422
rect 5349 9344 8218 9346
rect 5349 9288 5354 9344
rect 5410 9288 8218 9344
rect 5349 9286 8218 9288
rect 9949 9346 10015 9349
rect 10358 9346 10364 9348
rect 9949 9344 10364 9346
rect 9949 9288 9954 9344
rect 10010 9288 10364 9344
rect 9949 9286 10364 9288
rect 5349 9283 5415 9286
rect 9949 9283 10015 9286
rect 10358 9284 10364 9286
rect 10428 9284 10434 9348
rect 10501 9346 10567 9349
rect 12341 9346 12407 9349
rect 10501 9344 12407 9346
rect 10501 9288 10506 9344
rect 10562 9288 12346 9344
rect 12402 9288 12407 9344
rect 10501 9286 12407 9288
rect 10501 9283 10567 9286
rect 12341 9283 12407 9286
rect 12934 9284 12940 9348
rect 13004 9284 13010 9348
rect 13997 9344 14063 9349
rect 13997 9288 14002 9344
rect 14058 9288 14063 9344
rect 3418 9280 3734 9281
rect 3418 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3734 9280
rect 3418 9215 3734 9216
rect 8363 9280 8679 9281
rect 8363 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8679 9280
rect 8363 9215 8679 9216
rect 4061 9210 4127 9213
rect 6177 9210 6243 9213
rect 8201 9212 8267 9213
rect 8150 9210 8156 9212
rect 4061 9208 6243 9210
rect 4061 9152 4066 9208
rect 4122 9152 6182 9208
rect 6238 9152 6243 9208
rect 4061 9150 6243 9152
rect 8110 9150 8156 9210
rect 8220 9208 8267 9212
rect 8262 9152 8267 9208
rect 4061 9147 4127 9150
rect 6177 9147 6243 9150
rect 8150 9148 8156 9150
rect 8220 9148 8267 9152
rect 8886 9148 8892 9212
rect 8956 9210 8962 9212
rect 11881 9210 11947 9213
rect 8956 9208 11947 9210
rect 8956 9152 11886 9208
rect 11942 9152 11947 9208
rect 8956 9150 11947 9152
rect 8956 9148 8962 9150
rect 8201 9147 8267 9148
rect 11881 9147 11947 9150
rect 12198 9148 12204 9212
rect 12268 9210 12274 9212
rect 12341 9210 12407 9213
rect 12268 9208 12407 9210
rect 12268 9152 12346 9208
rect 12402 9152 12407 9208
rect 12268 9150 12407 9152
rect 12268 9148 12274 9150
rect 12341 9147 12407 9150
rect -300 9074 160 9104
rect 1761 9074 1827 9077
rect -300 9072 1827 9074
rect -300 9016 1766 9072
rect 1822 9016 1827 9072
rect -300 9014 1827 9016
rect -300 8984 160 9014
rect 1761 9011 1827 9014
rect 1894 9012 1900 9076
rect 1964 9074 1970 9076
rect 2262 9074 2268 9076
rect 1964 9014 2268 9074
rect 1964 9012 1970 9014
rect 2262 9012 2268 9014
rect 2332 9012 2338 9076
rect 3969 9074 4035 9077
rect 4102 9074 4108 9076
rect 3969 9072 4108 9074
rect 3969 9016 3974 9072
rect 4030 9016 4108 9072
rect 3969 9014 4108 9016
rect 3969 9011 4035 9014
rect 4102 9012 4108 9014
rect 4172 9012 4178 9076
rect 4705 9074 4771 9077
rect 4340 9072 4771 9074
rect 4340 9016 4710 9072
rect 4766 9016 4771 9072
rect 4340 9014 4771 9016
rect 1710 8876 1716 8940
rect 1780 8938 1786 8940
rect 2262 8938 2268 8940
rect 1780 8878 2268 8938
rect 1780 8876 1786 8878
rect 2262 8876 2268 8878
rect 2332 8876 2338 8940
rect 2630 8876 2636 8940
rect 2700 8938 2706 8940
rect 4340 8938 4400 9014
rect 4705 9011 4771 9014
rect 5390 9012 5396 9076
rect 5460 9074 5466 9076
rect 6913 9074 6979 9077
rect 5460 9072 6979 9074
rect 5460 9016 6918 9072
rect 6974 9016 6979 9072
rect 5460 9014 6979 9016
rect 5460 9012 5466 9014
rect 6913 9011 6979 9014
rect 7833 9074 7899 9077
rect 8201 9074 8267 9077
rect 7833 9072 8267 9074
rect 7833 9016 7838 9072
rect 7894 9016 8206 9072
rect 8262 9016 8267 9072
rect 7833 9014 8267 9016
rect 7833 9011 7899 9014
rect 8201 9011 8267 9014
rect 8569 9074 8635 9077
rect 9806 9074 9812 9076
rect 8569 9072 9812 9074
rect 8569 9016 8574 9072
rect 8630 9016 9812 9072
rect 8569 9014 9812 9016
rect 8569 9011 8635 9014
rect 9806 9012 9812 9014
rect 9876 9012 9882 9076
rect 10358 9012 10364 9076
rect 10428 9074 10434 9076
rect 12942 9074 13002 9284
rect 13997 9283 14063 9288
rect 14273 9346 14339 9349
rect 16798 9346 16804 9348
rect 14273 9344 16804 9346
rect 14273 9288 14278 9344
rect 14334 9288 16804 9344
rect 14273 9286 16804 9288
rect 14273 9283 14339 9286
rect 16798 9284 16804 9286
rect 16868 9284 16874 9348
rect 17033 9346 17099 9349
rect 19333 9348 19399 9349
rect 18086 9346 18092 9348
rect 17033 9344 18092 9346
rect 17033 9288 17038 9344
rect 17094 9288 18092 9344
rect 17033 9286 18092 9288
rect 17033 9283 17099 9286
rect 18086 9284 18092 9286
rect 18156 9284 18162 9348
rect 19333 9344 19380 9348
rect 19444 9346 19450 9348
rect 20345 9346 20411 9349
rect 21840 9346 22300 9376
rect 19333 9288 19338 9344
rect 19333 9284 19380 9288
rect 19444 9286 19490 9346
rect 20345 9344 22300 9346
rect 20345 9288 20350 9344
rect 20406 9288 22300 9344
rect 20345 9286 22300 9288
rect 19444 9284 19450 9286
rect 19333 9283 19399 9284
rect 20345 9283 20411 9286
rect 13308 9280 13624 9281
rect 13308 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13624 9280
rect 13308 9215 13624 9216
rect 18253 9280 18569 9281
rect 18253 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18569 9280
rect 21840 9256 22300 9286
rect 18253 9215 18569 9216
rect 13905 9210 13971 9213
rect 14549 9210 14615 9213
rect 13905 9208 14615 9210
rect 13905 9152 13910 9208
rect 13966 9152 14554 9208
rect 14610 9152 14615 9208
rect 13905 9150 14615 9152
rect 13905 9147 13971 9150
rect 14549 9147 14615 9150
rect 14917 9212 14983 9213
rect 14917 9208 14964 9212
rect 15028 9210 15034 9212
rect 15745 9210 15811 9213
rect 18045 9210 18111 9213
rect 14917 9152 14922 9208
rect 14917 9148 14964 9152
rect 15028 9150 15074 9210
rect 15745 9208 18111 9210
rect 15745 9152 15750 9208
rect 15806 9152 18050 9208
rect 18106 9152 18111 9208
rect 15745 9150 18111 9152
rect 15028 9148 15034 9150
rect 14917 9147 14983 9148
rect 15745 9147 15811 9150
rect 18045 9147 18111 9150
rect 18689 9210 18755 9213
rect 18822 9210 18828 9212
rect 18689 9208 18828 9210
rect 18689 9152 18694 9208
rect 18750 9152 18828 9208
rect 18689 9150 18828 9152
rect 18689 9147 18755 9150
rect 18822 9148 18828 9150
rect 18892 9148 18898 9212
rect 19149 9210 19215 9213
rect 20294 9210 20300 9212
rect 19149 9208 20300 9210
rect 19149 9152 19154 9208
rect 19210 9152 20300 9208
rect 19149 9150 20300 9152
rect 19149 9147 19215 9150
rect 20294 9148 20300 9150
rect 20364 9148 20370 9212
rect 18873 9074 18939 9077
rect 10428 9014 13002 9074
rect 13080 9072 18939 9074
rect 13080 9016 18878 9072
rect 18934 9016 18939 9072
rect 13080 9014 18939 9016
rect 10428 9012 10434 9014
rect 2700 8878 4400 8938
rect 2700 8876 2706 8878
rect 4470 8876 4476 8940
rect 4540 8938 4546 8940
rect 4705 8938 4771 8941
rect 12893 8938 12959 8941
rect 13080 8938 13140 9014
rect 18873 9011 18939 9014
rect 19517 9074 19583 9077
rect 19926 9074 19932 9076
rect 19517 9072 19932 9074
rect 19517 9016 19522 9072
rect 19578 9016 19932 9072
rect 19517 9014 19932 9016
rect 19517 9011 19583 9014
rect 19926 9012 19932 9014
rect 19996 9012 20002 9076
rect 15469 8938 15535 8941
rect 16389 8938 16455 8941
rect 16982 8938 16988 8940
rect 4540 8936 13140 8938
rect 4540 8880 4710 8936
rect 4766 8880 12898 8936
rect 12954 8880 13140 8936
rect 4540 8878 13140 8880
rect 13724 8936 15535 8938
rect 13724 8880 15474 8936
rect 15530 8880 15535 8936
rect 13724 8878 15535 8880
rect 4540 8876 4546 8878
rect 4705 8875 4771 8878
rect 12893 8875 12959 8878
rect -300 8802 160 8832
rect 2313 8802 2379 8805
rect -300 8800 2379 8802
rect -300 8744 2318 8800
rect 2374 8744 2379 8800
rect -300 8742 2379 8744
rect -300 8712 160 8742
rect 2313 8739 2379 8742
rect 7189 8802 7255 8805
rect 7557 8802 7623 8805
rect 7189 8800 7623 8802
rect 7189 8744 7194 8800
rect 7250 8744 7562 8800
rect 7618 8744 7623 8800
rect 7189 8742 7623 8744
rect 7189 8739 7255 8742
rect 7557 8739 7623 8742
rect 7782 8740 7788 8804
rect 7852 8802 7858 8804
rect 10358 8802 10364 8804
rect 7852 8742 10364 8802
rect 7852 8740 7858 8742
rect 10358 8740 10364 8742
rect 10428 8740 10434 8804
rect 10542 8740 10548 8804
rect 10612 8740 10618 8804
rect 11513 8802 11579 8805
rect 11973 8802 12039 8805
rect 11513 8800 12039 8802
rect 11513 8744 11518 8800
rect 11574 8744 11978 8800
rect 12034 8744 12039 8800
rect 11513 8742 12039 8744
rect 5890 8736 6206 8737
rect 5890 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6206 8736
rect 5890 8671 6206 8672
rect 2037 8666 2103 8669
rect 4797 8666 4863 8669
rect 2037 8664 4863 8666
rect 2037 8608 2042 8664
rect 2098 8608 4802 8664
rect 4858 8608 4863 8664
rect 2037 8606 4863 8608
rect 2037 8603 2103 8606
rect 4797 8603 4863 8606
rect 6545 8666 6611 8669
rect 8477 8666 8543 8669
rect 6545 8664 8543 8666
rect 6545 8608 6550 8664
rect 6606 8608 8482 8664
rect 8538 8608 8543 8664
rect 6545 8606 8543 8608
rect 6545 8603 6611 8606
rect 8477 8603 8543 8606
rect 10041 8666 10107 8669
rect 10550 8666 10610 8740
rect 11513 8739 11579 8742
rect 11973 8739 12039 8742
rect 12382 8740 12388 8804
rect 12452 8802 12458 8804
rect 13724 8802 13784 8878
rect 15469 8875 15535 8878
rect 15656 8878 16268 8938
rect 12452 8742 13784 8802
rect 12452 8740 12458 8742
rect 13854 8740 13860 8804
rect 13924 8802 13930 8804
rect 15656 8802 15716 8878
rect 13924 8742 15716 8802
rect 16208 8802 16268 8878
rect 16389 8936 16988 8938
rect 16389 8880 16394 8936
rect 16450 8880 16988 8936
rect 16389 8878 16988 8880
rect 16389 8875 16455 8878
rect 16982 8876 16988 8878
rect 17052 8876 17058 8940
rect 18321 8938 18387 8941
rect 18321 8936 21282 8938
rect 18321 8880 18326 8936
rect 18382 8880 21282 8936
rect 18321 8878 21282 8880
rect 18321 8875 18387 8878
rect 19241 8802 19307 8805
rect 16208 8800 19307 8802
rect 16208 8744 19246 8800
rect 19302 8744 19307 8800
rect 16208 8742 19307 8744
rect 21222 8802 21282 8878
rect 21840 8802 22300 8832
rect 21222 8742 22300 8802
rect 13924 8740 13930 8742
rect 19241 8739 19307 8742
rect 10835 8736 11151 8737
rect 10835 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11151 8736
rect 10835 8671 11151 8672
rect 15780 8736 16096 8737
rect 15780 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16096 8736
rect 15780 8671 16096 8672
rect 20725 8736 21041 8737
rect 20725 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21041 8736
rect 21840 8712 22300 8742
rect 20725 8671 21041 8672
rect 15285 8666 15351 8669
rect 10041 8664 10610 8666
rect 10041 8608 10046 8664
rect 10102 8608 10610 8664
rect 10041 8606 10610 8608
rect 11286 8664 15351 8666
rect 11286 8608 15290 8664
rect 15346 8608 15351 8664
rect 11286 8606 15351 8608
rect 10041 8603 10107 8606
rect -300 8530 160 8560
rect 1209 8530 1275 8533
rect -300 8528 1275 8530
rect -300 8472 1214 8528
rect 1270 8472 1275 8528
rect -300 8470 1275 8472
rect -300 8440 160 8470
rect 1209 8467 1275 8470
rect 2221 8530 2287 8533
rect 2998 8530 3004 8532
rect 2221 8528 3004 8530
rect 2221 8472 2226 8528
rect 2282 8472 3004 8528
rect 2221 8470 3004 8472
rect 2221 8467 2287 8470
rect 2998 8468 3004 8470
rect 3068 8468 3074 8532
rect 3182 8468 3188 8532
rect 3252 8530 3258 8532
rect 3417 8530 3483 8533
rect 3252 8528 3483 8530
rect 3252 8472 3422 8528
rect 3478 8472 3483 8528
rect 3252 8470 3483 8472
rect 3252 8468 3258 8470
rect 3417 8467 3483 8470
rect 4429 8530 4495 8533
rect 6085 8530 6151 8533
rect 4429 8528 6151 8530
rect 4429 8472 4434 8528
rect 4490 8472 6090 8528
rect 6146 8472 6151 8528
rect 4429 8470 6151 8472
rect 4429 8467 4495 8470
rect 6085 8467 6151 8470
rect 7557 8530 7623 8533
rect 11286 8530 11346 8606
rect 15285 8603 15351 8606
rect 16205 8666 16271 8669
rect 19425 8666 19491 8669
rect 16205 8664 19491 8666
rect 16205 8608 16210 8664
rect 16266 8608 19430 8664
rect 19486 8608 19491 8664
rect 16205 8606 19491 8608
rect 16205 8603 16271 8606
rect 19425 8603 19491 8606
rect 7557 8528 11346 8530
rect 7557 8472 7562 8528
rect 7618 8472 11346 8528
rect 7557 8470 11346 8472
rect 12249 8530 12315 8533
rect 12801 8530 12867 8533
rect 12249 8528 12867 8530
rect 12249 8472 12254 8528
rect 12310 8472 12806 8528
rect 12862 8472 12867 8528
rect 12249 8470 12867 8472
rect 7557 8467 7623 8470
rect 12249 8467 12315 8470
rect 12801 8467 12867 8470
rect 12985 8530 13051 8533
rect 18689 8530 18755 8533
rect 12985 8528 18755 8530
rect 12985 8472 12990 8528
rect 13046 8472 18694 8528
rect 18750 8472 18755 8528
rect 12985 8470 18755 8472
rect 12985 8467 13051 8470
rect 18689 8467 18755 8470
rect 841 8394 907 8397
rect 1669 8394 1735 8397
rect 841 8392 1735 8394
rect 841 8336 846 8392
rect 902 8336 1674 8392
rect 1730 8336 1735 8392
rect 841 8334 1735 8336
rect 841 8331 907 8334
rect 1669 8331 1735 8334
rect 2405 8396 2471 8397
rect 2405 8392 2452 8396
rect 2516 8394 2522 8396
rect 2957 8394 3023 8397
rect 8385 8394 8451 8397
rect 20069 8394 20135 8397
rect 2405 8336 2410 8392
rect 2405 8332 2452 8336
rect 2516 8334 2562 8394
rect 2957 8392 8451 8394
rect 2957 8336 2962 8392
rect 3018 8336 8390 8392
rect 8446 8336 8451 8392
rect 2957 8334 8451 8336
rect 2516 8332 2522 8334
rect 2405 8331 2471 8332
rect 2957 8331 3023 8334
rect 8385 8331 8451 8334
rect 10366 8392 20135 8394
rect 10366 8336 20074 8392
rect 20130 8336 20135 8392
rect 10366 8334 20135 8336
rect -300 8258 160 8288
rect 3141 8258 3207 8261
rect -300 8256 3207 8258
rect -300 8200 3146 8256
rect 3202 8200 3207 8256
rect -300 8198 3207 8200
rect -300 8168 160 8198
rect 3141 8195 3207 8198
rect 5390 8196 5396 8260
rect 5460 8258 5466 8260
rect 5717 8258 5783 8261
rect 5460 8256 5783 8258
rect 5460 8200 5722 8256
rect 5778 8200 5783 8256
rect 5460 8198 5783 8200
rect 5460 8196 5466 8198
rect 5717 8195 5783 8198
rect 5993 8258 6059 8261
rect 6494 8258 6500 8260
rect 5993 8256 6500 8258
rect 5993 8200 5998 8256
rect 6054 8200 6500 8256
rect 5993 8198 6500 8200
rect 5993 8195 6059 8198
rect 6494 8196 6500 8198
rect 6564 8196 6570 8260
rect 3418 8192 3734 8193
rect 3418 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3734 8192
rect 3418 8127 3734 8128
rect 8363 8192 8679 8193
rect 8363 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8679 8192
rect 8363 8127 8679 8128
rect 841 8122 907 8125
rect 4061 8124 4127 8125
rect 1710 8122 1716 8124
rect 841 8120 1716 8122
rect 841 8064 846 8120
rect 902 8064 1716 8120
rect 841 8062 1716 8064
rect 841 8059 907 8062
rect 1710 8060 1716 8062
rect 1780 8060 1786 8124
rect 4061 8120 4108 8124
rect 4172 8122 4178 8124
rect 5809 8122 5875 8125
rect 6177 8122 6243 8125
rect 4061 8064 4066 8120
rect 4061 8060 4108 8064
rect 4172 8062 4218 8122
rect 5809 8120 6243 8122
rect 5809 8064 5814 8120
rect 5870 8064 6182 8120
rect 6238 8064 6243 8120
rect 5809 8062 6243 8064
rect 4172 8060 4178 8062
rect 4061 8059 4127 8060
rect 5809 8059 5875 8062
rect 6177 8059 6243 8062
rect 7465 8122 7531 8125
rect 7741 8122 7807 8125
rect 7465 8120 7807 8122
rect 7465 8064 7470 8120
rect 7526 8064 7746 8120
rect 7802 8064 7807 8120
rect 7465 8062 7807 8064
rect 7465 8059 7531 8062
rect 7741 8059 7807 8062
rect -300 7986 160 8016
rect 4061 7986 4127 7989
rect -300 7984 4127 7986
rect -300 7928 4066 7984
rect 4122 7928 4127 7984
rect -300 7926 4127 7928
rect -300 7896 160 7926
rect 4061 7923 4127 7926
rect 5257 7986 5323 7989
rect 10366 7986 10426 8334
rect 20069 8331 20135 8334
rect 10869 8258 10935 8261
rect 12341 8258 12407 8261
rect 10869 8256 12407 8258
rect 10869 8200 10874 8256
rect 10930 8200 12346 8256
rect 12402 8200 12407 8256
rect 10869 8198 12407 8200
rect 10869 8195 10935 8198
rect 12341 8195 12407 8198
rect 13997 8258 14063 8261
rect 18045 8258 18111 8261
rect 21840 8258 22300 8288
rect 13997 8256 18111 8258
rect 13997 8200 14002 8256
rect 14058 8200 18050 8256
rect 18106 8200 18111 8256
rect 13997 8198 18111 8200
rect 13997 8195 14063 8198
rect 18045 8195 18111 8198
rect 19198 8198 22300 8258
rect 13308 8192 13624 8193
rect 13308 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13624 8192
rect 13308 8127 13624 8128
rect 18253 8192 18569 8193
rect 18253 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18569 8192
rect 18253 8127 18569 8128
rect 10542 8060 10548 8124
rect 10612 8122 10618 8124
rect 12525 8122 12591 8125
rect 10612 8120 12591 8122
rect 10612 8064 12530 8120
rect 12586 8064 12591 8120
rect 10612 8062 12591 8064
rect 10612 8060 10618 8062
rect 12525 8059 12591 8062
rect 13997 8122 14063 8125
rect 16205 8122 16271 8125
rect 13997 8120 16271 8122
rect 13997 8064 14002 8120
rect 14058 8064 16210 8120
rect 16266 8064 16271 8120
rect 13997 8062 16271 8064
rect 13997 8059 14063 8062
rect 16205 8059 16271 8062
rect 16665 8120 16731 8125
rect 16665 8064 16670 8120
rect 16726 8064 16731 8120
rect 16665 8059 16731 8064
rect 16798 8060 16804 8124
rect 16868 8122 16874 8124
rect 17309 8122 17375 8125
rect 16868 8120 17375 8122
rect 16868 8064 17314 8120
rect 17370 8064 17375 8120
rect 16868 8062 17375 8064
rect 16868 8060 16874 8062
rect 17309 8059 17375 8062
rect 5257 7984 10426 7986
rect 5257 7928 5262 7984
rect 5318 7928 10426 7984
rect 5257 7926 10426 7928
rect 5257 7923 5323 7926
rect 10542 7924 10548 7988
rect 10612 7986 10618 7988
rect 13854 7986 13860 7988
rect 10612 7926 13860 7986
rect 10612 7924 10618 7926
rect 13854 7924 13860 7926
rect 13924 7924 13930 7988
rect 14273 7986 14339 7989
rect 16389 7986 16455 7989
rect 14273 7984 16455 7986
rect 14273 7928 14278 7984
rect 14334 7928 16394 7984
rect 16450 7928 16455 7984
rect 14273 7926 16455 7928
rect 16668 7986 16728 8059
rect 19198 7986 19258 8198
rect 21840 8168 22300 8198
rect 19333 8122 19399 8125
rect 19558 8122 19564 8124
rect 19333 8120 19564 8122
rect 19333 8064 19338 8120
rect 19394 8064 19564 8120
rect 19333 8062 19564 8064
rect 19333 8059 19399 8062
rect 19558 8060 19564 8062
rect 19628 8060 19634 8124
rect 16668 7926 19258 7986
rect 14273 7923 14339 7926
rect 16389 7923 16455 7926
rect 1393 7852 1459 7853
rect 1342 7788 1348 7852
rect 1412 7850 1459 7852
rect 1853 7852 1919 7853
rect 1412 7848 1504 7850
rect 1454 7792 1504 7848
rect 1412 7790 1504 7792
rect 1853 7848 1900 7852
rect 1964 7850 1970 7852
rect 1853 7792 1858 7848
rect 1412 7788 1459 7790
rect 1393 7787 1459 7788
rect 1853 7788 1900 7792
rect 1964 7790 2010 7850
rect 1964 7788 1970 7790
rect 2814 7788 2820 7852
rect 2884 7850 2890 7852
rect 3693 7850 3759 7853
rect 2884 7848 3759 7850
rect 2884 7792 3698 7848
rect 3754 7792 3759 7848
rect 2884 7790 3759 7792
rect 2884 7788 2890 7790
rect 1853 7787 1919 7788
rect 3693 7787 3759 7790
rect 3918 7788 3924 7852
rect 3988 7850 3994 7852
rect 4153 7850 4219 7853
rect 3988 7848 4219 7850
rect 3988 7792 4158 7848
rect 4214 7792 4219 7848
rect 3988 7790 4219 7792
rect 3988 7788 3994 7790
rect 4153 7787 4219 7790
rect 4797 7850 4863 7853
rect 6453 7850 6519 7853
rect 4797 7848 6519 7850
rect 4797 7792 4802 7848
rect 4858 7792 6458 7848
rect 6514 7792 6519 7848
rect 4797 7790 6519 7792
rect 4797 7787 4863 7790
rect 6453 7787 6519 7790
rect 7465 7850 7531 7853
rect 8661 7850 8727 7853
rect 7465 7848 8727 7850
rect 7465 7792 7470 7848
rect 7526 7792 8666 7848
rect 8722 7792 8727 7848
rect 7465 7790 8727 7792
rect 7465 7787 7531 7790
rect 8661 7787 8727 7790
rect 9213 7850 9279 7853
rect 9622 7850 9628 7852
rect 9213 7848 9628 7850
rect 9213 7792 9218 7848
rect 9274 7792 9628 7848
rect 9213 7790 9628 7792
rect 9213 7787 9279 7790
rect 9622 7788 9628 7790
rect 9692 7788 9698 7852
rect 10409 7850 10475 7853
rect 10869 7850 10935 7853
rect 10409 7848 10935 7850
rect 10409 7792 10414 7848
rect 10470 7792 10874 7848
rect 10930 7792 10935 7848
rect 10409 7790 10935 7792
rect 10409 7787 10475 7790
rect 10869 7787 10935 7790
rect 11237 7848 11303 7853
rect 11237 7792 11242 7848
rect 11298 7792 11303 7848
rect 11237 7787 11303 7792
rect 12525 7850 12591 7853
rect 19885 7850 19951 7853
rect 12525 7848 19951 7850
rect 12525 7792 12530 7848
rect 12586 7792 19890 7848
rect 19946 7792 19951 7848
rect 12525 7790 19951 7792
rect 12525 7787 12591 7790
rect 19885 7787 19951 7790
rect -300 7714 160 7744
rect 1393 7714 1459 7717
rect -300 7712 1459 7714
rect -300 7656 1398 7712
rect 1454 7656 1459 7712
rect -300 7654 1459 7656
rect -300 7624 160 7654
rect 1393 7651 1459 7654
rect 2078 7652 2084 7716
rect 2148 7714 2154 7716
rect 3785 7714 3851 7717
rect 5165 7714 5231 7717
rect 2148 7654 3434 7714
rect 2148 7652 2154 7654
rect 1025 7578 1091 7581
rect 1158 7578 1164 7580
rect 1025 7576 1164 7578
rect 1025 7520 1030 7576
rect 1086 7520 1164 7576
rect 1025 7518 1164 7520
rect 1025 7515 1091 7518
rect 1158 7516 1164 7518
rect 1228 7516 1234 7580
rect 3374 7578 3434 7654
rect 3785 7712 5231 7714
rect 3785 7656 3790 7712
rect 3846 7656 5170 7712
rect 5226 7656 5231 7712
rect 3785 7654 5231 7656
rect 3785 7651 3851 7654
rect 5165 7651 5231 7654
rect 8661 7714 8727 7717
rect 9673 7714 9739 7717
rect 8661 7712 9739 7714
rect 8661 7656 8666 7712
rect 8722 7656 9678 7712
rect 9734 7656 9739 7712
rect 8661 7654 9739 7656
rect 11240 7714 11300 7787
rect 15009 7714 15075 7717
rect 11240 7712 15075 7714
rect 11240 7656 15014 7712
rect 15070 7656 15075 7712
rect 11240 7654 15075 7656
rect 8661 7651 8727 7654
rect 9673 7651 9739 7654
rect 15009 7651 15075 7654
rect 16205 7712 16271 7717
rect 16205 7656 16210 7712
rect 16266 7656 16271 7712
rect 16205 7651 16271 7656
rect 16389 7714 16455 7717
rect 18873 7714 18939 7717
rect 21840 7714 22300 7744
rect 16389 7712 18939 7714
rect 16389 7656 16394 7712
rect 16450 7656 18878 7712
rect 18934 7656 18939 7712
rect 16389 7654 18939 7656
rect 16389 7651 16455 7654
rect 18873 7651 18939 7654
rect 21176 7654 22300 7714
rect 5890 7648 6206 7649
rect 5890 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6206 7648
rect 5890 7583 6206 7584
rect 10835 7648 11151 7649
rect 10835 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11151 7648
rect 10835 7583 11151 7584
rect 15780 7648 16096 7649
rect 15780 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16096 7648
rect 15780 7583 16096 7584
rect 5390 7578 5396 7580
rect 3374 7518 5396 7578
rect 5390 7516 5396 7518
rect 5460 7516 5466 7580
rect 6453 7578 6519 7581
rect 9857 7578 9923 7581
rect 6453 7576 9923 7578
rect 6453 7520 6458 7576
rect 6514 7520 9862 7576
rect 9918 7520 9923 7576
rect 6453 7518 9923 7520
rect 6453 7515 6519 7518
rect 9857 7515 9923 7518
rect 12157 7578 12223 7581
rect 12750 7578 12756 7580
rect 12157 7576 12756 7578
rect 12157 7520 12162 7576
rect 12218 7520 12756 7576
rect 12157 7518 12756 7520
rect 12157 7515 12223 7518
rect 12750 7516 12756 7518
rect 12820 7516 12826 7580
rect 12934 7516 12940 7580
rect 13004 7578 13010 7580
rect 14641 7578 14707 7581
rect 13004 7576 14707 7578
rect 13004 7520 14646 7576
rect 14702 7520 14707 7576
rect 13004 7518 14707 7520
rect 16208 7578 16268 7651
rect 20725 7648 21041 7649
rect 20725 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21041 7648
rect 20725 7583 21041 7584
rect 16208 7518 17924 7578
rect 13004 7516 13010 7518
rect 14641 7515 14707 7518
rect -300 7442 160 7472
rect 2037 7442 2103 7445
rect -300 7440 2103 7442
rect -300 7384 2042 7440
rect 2098 7384 2103 7440
rect -300 7382 2103 7384
rect -300 7352 160 7382
rect 2037 7379 2103 7382
rect 2681 7442 2747 7445
rect 3182 7442 3188 7444
rect 2681 7440 3188 7442
rect 2681 7384 2686 7440
rect 2742 7384 3188 7440
rect 2681 7382 3188 7384
rect 2681 7379 2747 7382
rect 3182 7380 3188 7382
rect 3252 7380 3258 7444
rect 3877 7442 3943 7445
rect 13905 7442 13971 7445
rect 3877 7440 13971 7442
rect 3877 7384 3882 7440
rect 3938 7384 13910 7440
rect 13966 7384 13971 7440
rect 3877 7382 13971 7384
rect 3877 7379 3943 7382
rect 13905 7379 13971 7382
rect 14825 7442 14891 7445
rect 17677 7442 17743 7445
rect 14825 7440 17743 7442
rect 14825 7384 14830 7440
rect 14886 7384 17682 7440
rect 17738 7384 17743 7440
rect 14825 7382 17743 7384
rect 17864 7442 17924 7518
rect 21176 7442 21236 7654
rect 21840 7624 22300 7654
rect 17864 7382 21236 7442
rect 14825 7379 14891 7382
rect 17677 7379 17743 7382
rect 565 7306 631 7309
rect 1342 7306 1348 7308
rect 565 7304 1348 7306
rect 565 7248 570 7304
rect 626 7248 1348 7304
rect 565 7246 1348 7248
rect 565 7243 631 7246
rect 1342 7244 1348 7246
rect 1412 7244 1418 7308
rect 2681 7306 2747 7309
rect 2957 7306 3023 7309
rect 2681 7304 3023 7306
rect 2681 7248 2686 7304
rect 2742 7248 2962 7304
rect 3018 7248 3023 7304
rect 2681 7246 3023 7248
rect 2681 7243 2747 7246
rect 2957 7243 3023 7246
rect 3969 7306 4035 7309
rect 6913 7306 6979 7309
rect 11329 7306 11395 7309
rect 3969 7304 6979 7306
rect 3969 7248 3974 7304
rect 4030 7248 6918 7304
rect 6974 7248 6979 7304
rect 3969 7246 6979 7248
rect 3969 7243 4035 7246
rect 6913 7243 6979 7246
rect 8158 7304 11395 7306
rect 8158 7248 11334 7304
rect 11390 7248 11395 7304
rect 8158 7246 11395 7248
rect -300 7170 160 7200
rect 2957 7170 3023 7173
rect -300 7168 3023 7170
rect -300 7112 2962 7168
rect 3018 7112 3023 7168
rect -300 7110 3023 7112
rect -300 7080 160 7110
rect 2957 7107 3023 7110
rect 4153 7170 4219 7173
rect 7557 7170 7623 7173
rect 4153 7168 7623 7170
rect 4153 7112 4158 7168
rect 4214 7112 7562 7168
rect 7618 7112 7623 7168
rect 4153 7110 7623 7112
rect 4153 7107 4219 7110
rect 7557 7107 7623 7110
rect 3418 7104 3734 7105
rect 3418 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3734 7104
rect 3418 7039 3734 7040
rect 2221 7034 2287 7037
rect 3233 7034 3299 7037
rect 8158 7034 8218 7246
rect 11329 7243 11395 7246
rect 11513 7306 11579 7309
rect 12249 7306 12315 7309
rect 11513 7304 12315 7306
rect 11513 7248 11518 7304
rect 11574 7248 12254 7304
rect 12310 7248 12315 7304
rect 11513 7246 12315 7248
rect 11513 7243 11579 7246
rect 12249 7243 12315 7246
rect 12750 7244 12756 7308
rect 12820 7306 12826 7308
rect 16573 7306 16639 7309
rect 12820 7304 16639 7306
rect 12820 7248 16578 7304
rect 16634 7248 16639 7304
rect 12820 7246 16639 7248
rect 12820 7244 12826 7246
rect 16573 7243 16639 7246
rect 17125 7308 17191 7309
rect 17125 7304 17172 7308
rect 17236 7306 17242 7308
rect 17585 7306 17651 7309
rect 17718 7306 17724 7308
rect 17125 7248 17130 7304
rect 17125 7244 17172 7248
rect 17236 7246 17282 7306
rect 17585 7304 17724 7306
rect 17585 7248 17590 7304
rect 17646 7248 17724 7304
rect 17585 7246 17724 7248
rect 17236 7244 17242 7246
rect 17125 7243 17191 7244
rect 17585 7243 17651 7246
rect 17718 7244 17724 7246
rect 17788 7244 17794 7308
rect 18094 7246 18706 7306
rect 9673 7170 9739 7173
rect 10869 7170 10935 7173
rect 9673 7168 10935 7170
rect 9673 7112 9678 7168
rect 9734 7112 10874 7168
rect 10930 7112 10935 7168
rect 9673 7110 10935 7112
rect 9673 7107 9739 7110
rect 10869 7107 10935 7110
rect 11053 7170 11119 7173
rect 12709 7170 12775 7173
rect 11053 7168 12775 7170
rect 11053 7112 11058 7168
rect 11114 7112 12714 7168
rect 12770 7112 12775 7168
rect 11053 7110 12775 7112
rect 11053 7107 11119 7110
rect 12709 7107 12775 7110
rect 13905 7170 13971 7173
rect 18094 7170 18154 7246
rect 13905 7168 18154 7170
rect 13905 7112 13910 7168
rect 13966 7112 18154 7168
rect 13905 7110 18154 7112
rect 18646 7170 18706 7246
rect 21840 7170 22300 7200
rect 18646 7110 22300 7170
rect 13905 7107 13971 7110
rect 8363 7104 8679 7105
rect 8363 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8679 7104
rect 8363 7039 8679 7040
rect 13308 7104 13624 7105
rect 13308 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13624 7104
rect 13308 7039 13624 7040
rect 18253 7104 18569 7105
rect 18253 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18569 7104
rect 21840 7080 22300 7110
rect 18253 7039 18569 7040
rect 2221 7032 3299 7034
rect 2221 6976 2226 7032
rect 2282 6976 3238 7032
rect 3294 6976 3299 7032
rect 2221 6974 3299 6976
rect 2221 6971 2287 6974
rect 3233 6971 3299 6974
rect 5076 6974 8218 7034
rect 10501 7034 10567 7037
rect 11513 7034 11579 7037
rect 12617 7034 12683 7037
rect 12934 7034 12940 7036
rect 10501 7032 11162 7034
rect 10501 6976 10506 7032
rect 10562 6976 11162 7032
rect 10501 6974 11162 6976
rect -300 6898 160 6928
rect 3969 6898 4035 6901
rect -300 6896 4035 6898
rect -300 6840 3974 6896
rect 4030 6840 4035 6896
rect -300 6838 4035 6840
rect -300 6808 160 6838
rect 3969 6835 4035 6838
rect 2221 6762 2287 6765
rect 5076 6762 5136 6974
rect 10501 6971 10567 6974
rect 5257 6900 5323 6901
rect 5206 6836 5212 6900
rect 5276 6898 5323 6900
rect 6085 6898 6151 6901
rect 10961 6898 11027 6901
rect 5276 6896 5368 6898
rect 5318 6840 5368 6896
rect 5276 6838 5368 6840
rect 6085 6896 7298 6898
rect 6085 6840 6090 6896
rect 6146 6840 7298 6896
rect 6085 6838 7298 6840
rect 5276 6836 5323 6838
rect 5257 6835 5323 6836
rect 6085 6835 6151 6838
rect 2221 6760 5136 6762
rect 2221 6704 2226 6760
rect 2282 6704 5136 6760
rect 7238 6796 7298 6838
rect 7606 6896 11027 6898
rect 7606 6840 10966 6896
rect 11022 6840 11027 6896
rect 7606 6838 11027 6840
rect 11102 6898 11162 6974
rect 11513 7032 12683 7034
rect 11513 6976 11518 7032
rect 11574 6976 12622 7032
rect 12678 6976 12683 7032
rect 11513 6974 12683 6976
rect 11513 6971 11579 6974
rect 12617 6971 12683 6974
rect 12758 6974 12940 7034
rect 11697 6898 11763 6901
rect 12758 6898 12818 6974
rect 12934 6972 12940 6974
rect 13004 6972 13010 7036
rect 14181 7034 14247 7037
rect 16389 7034 16455 7037
rect 18045 7036 18111 7037
rect 18045 7034 18092 7036
rect 14181 7032 16455 7034
rect 14181 6976 14186 7032
rect 14242 6976 16394 7032
rect 16450 6976 16455 7032
rect 14181 6974 16455 6976
rect 18000 7032 18092 7034
rect 18000 6976 18050 7032
rect 18000 6974 18092 6976
rect 14181 6971 14247 6974
rect 16389 6971 16455 6974
rect 18045 6972 18092 6974
rect 18156 6972 18162 7036
rect 18045 6971 18111 6972
rect 11102 6838 11484 6898
rect 7606 6796 7666 6838
rect 10961 6835 11027 6838
rect 7238 6736 7666 6796
rect 2221 6702 5136 6704
rect 7560 6702 7666 6736
rect 7925 6762 7991 6765
rect 9673 6762 9739 6765
rect 11424 6762 11484 6838
rect 11697 6896 12818 6898
rect 11697 6840 11702 6896
rect 11758 6840 12818 6896
rect 11697 6838 12818 6840
rect 11697 6835 11763 6838
rect 12934 6836 12940 6900
rect 13004 6898 13010 6900
rect 13004 6838 19994 6898
rect 13004 6836 13010 6838
rect 12709 6762 12775 6765
rect 7925 6760 9739 6762
rect 7925 6704 7930 6760
rect 7986 6704 9678 6760
rect 9734 6704 9739 6760
rect 7925 6702 9739 6704
rect 2221 6699 2287 6702
rect 7925 6699 7991 6702
rect 9673 6699 9739 6702
rect 10504 6702 11346 6762
rect 11424 6760 12775 6762
rect 11424 6704 12714 6760
rect 12770 6704 12775 6760
rect 11424 6702 12775 6704
rect -300 6626 160 6656
rect 565 6626 631 6629
rect -300 6624 631 6626
rect -300 6568 570 6624
rect 626 6568 631 6624
rect -300 6566 631 6568
rect -300 6536 160 6566
rect 565 6563 631 6566
rect 4061 6626 4127 6629
rect 4705 6626 4771 6629
rect 4061 6624 4771 6626
rect 4061 6568 4066 6624
rect 4122 6568 4710 6624
rect 4766 6568 4771 6624
rect 4061 6566 4771 6568
rect 4061 6563 4127 6566
rect 4705 6563 4771 6566
rect 7097 6626 7163 6629
rect 7281 6626 7347 6629
rect 7097 6624 7347 6626
rect 7097 6568 7102 6624
rect 7158 6568 7286 6624
rect 7342 6568 7347 6624
rect 7097 6566 7347 6568
rect 7097 6563 7163 6566
rect 7281 6563 7347 6566
rect 8385 6626 8451 6629
rect 9990 6626 9996 6628
rect 8385 6624 9996 6626
rect 8385 6568 8390 6624
rect 8446 6568 9996 6624
rect 8385 6566 9996 6568
rect 8385 6563 8451 6566
rect 9990 6564 9996 6566
rect 10060 6564 10066 6628
rect 5890 6560 6206 6561
rect 5890 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6206 6560
rect 5890 6495 6206 6496
rect 4061 6492 4127 6493
rect 4061 6490 4108 6492
rect 4016 6488 4108 6490
rect 4016 6432 4066 6488
rect 4016 6430 4108 6432
rect 4061 6428 4108 6430
rect 4172 6428 4178 6492
rect 5625 6490 5691 6493
rect 4340 6488 5691 6490
rect 4340 6432 5630 6488
rect 5686 6432 5691 6488
rect 4340 6430 5691 6432
rect 4061 6427 4127 6428
rect -300 6354 160 6384
rect 1853 6354 1919 6357
rect 4340 6354 4400 6430
rect 5625 6427 5691 6430
rect 6453 6490 6519 6493
rect 7281 6490 7347 6493
rect 6453 6488 7068 6490
rect 6453 6432 6458 6488
rect 6514 6432 7068 6488
rect 6453 6430 7068 6432
rect 6453 6427 6519 6430
rect 4521 6356 4587 6357
rect -300 6352 1919 6354
rect -300 6296 1858 6352
rect 1914 6296 1919 6352
rect -300 6294 1919 6296
rect -300 6264 160 6294
rect 1853 6291 1919 6294
rect 2132 6294 4400 6354
rect 238 6156 244 6220
rect 308 6218 314 6220
rect 2132 6218 2192 6294
rect 4470 6292 4476 6356
rect 4540 6354 4587 6356
rect 4981 6354 5047 6357
rect 6862 6354 6868 6356
rect 4540 6352 4632 6354
rect 4582 6296 4632 6352
rect 4540 6294 4632 6296
rect 4981 6352 6868 6354
rect 4981 6296 4986 6352
rect 5042 6296 6868 6352
rect 4981 6294 6868 6296
rect 4540 6292 4587 6294
rect 4521 6291 4587 6292
rect 4981 6291 5047 6294
rect 6862 6292 6868 6294
rect 6932 6292 6938 6356
rect 7008 6354 7068 6430
rect 7281 6488 9690 6490
rect 7281 6432 7286 6488
rect 7342 6432 9690 6488
rect 7281 6430 9690 6432
rect 7281 6427 7347 6430
rect 9630 6356 9690 6430
rect 9990 6428 9996 6492
rect 10060 6490 10066 6492
rect 10504 6490 10564 6702
rect 11286 6626 11346 6702
rect 12709 6699 12775 6702
rect 12985 6762 13051 6765
rect 14825 6762 14891 6765
rect 12985 6760 14891 6762
rect 12985 6704 12990 6760
rect 13046 6704 14830 6760
rect 14886 6704 14891 6760
rect 12985 6702 14891 6704
rect 12985 6699 13051 6702
rect 14825 6699 14891 6702
rect 14958 6700 14964 6764
rect 15028 6762 15034 6764
rect 15285 6762 15351 6765
rect 16849 6762 16915 6765
rect 19701 6762 19767 6765
rect 15028 6760 15351 6762
rect 15028 6704 15290 6760
rect 15346 6704 15351 6760
rect 15028 6702 15351 6704
rect 15028 6700 15034 6702
rect 15285 6699 15351 6702
rect 15472 6702 16268 6762
rect 14089 6626 14155 6629
rect 11286 6624 14155 6626
rect 11286 6568 14094 6624
rect 14150 6568 14155 6624
rect 11286 6566 14155 6568
rect 14089 6563 14155 6566
rect 14222 6564 14228 6628
rect 14292 6626 14298 6628
rect 15472 6626 15532 6702
rect 14292 6566 15532 6626
rect 16208 6626 16268 6702
rect 16849 6760 19767 6762
rect 16849 6704 16854 6760
rect 16910 6704 19706 6760
rect 19762 6704 19767 6760
rect 16849 6702 19767 6704
rect 16849 6699 16915 6702
rect 19701 6699 19767 6702
rect 18505 6626 18571 6629
rect 16208 6624 18571 6626
rect 16208 6568 18510 6624
rect 18566 6568 18571 6624
rect 16208 6566 18571 6568
rect 14292 6564 14298 6566
rect 18505 6563 18571 6566
rect 10835 6560 11151 6561
rect 10835 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11151 6560
rect 10835 6495 11151 6496
rect 15780 6560 16096 6561
rect 15780 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16096 6560
rect 15780 6495 16096 6496
rect 12801 6490 12867 6493
rect 15285 6490 15351 6493
rect 15561 6492 15627 6493
rect 10060 6430 10564 6490
rect 11884 6430 12634 6490
rect 10060 6428 10066 6430
rect 7008 6294 9506 6354
rect 308 6158 2192 6218
rect 2313 6218 2379 6221
rect 6361 6218 6427 6221
rect 2313 6216 6427 6218
rect 2313 6160 2318 6216
rect 2374 6160 6366 6216
rect 6422 6160 6427 6216
rect 2313 6158 6427 6160
rect 308 6156 314 6158
rect 2313 6155 2379 6158
rect 6361 6155 6427 6158
rect 6545 6218 6611 6221
rect 7005 6218 7071 6221
rect 6545 6216 7071 6218
rect 6545 6160 6550 6216
rect 6606 6160 7010 6216
rect 7066 6160 7071 6216
rect 6545 6158 7071 6160
rect 6545 6155 6611 6158
rect 7005 6155 7071 6158
rect 7598 6156 7604 6220
rect 7668 6218 7674 6220
rect 7925 6218 7991 6221
rect 7668 6216 7991 6218
rect 7668 6160 7930 6216
rect 7986 6160 7991 6216
rect 7668 6158 7991 6160
rect 7668 6156 7674 6158
rect 7925 6155 7991 6158
rect 8569 6218 8635 6221
rect 9305 6218 9371 6221
rect 8569 6216 9371 6218
rect 8569 6160 8574 6216
rect 8630 6160 9310 6216
rect 9366 6160 9371 6216
rect 8569 6158 9371 6160
rect 8569 6155 8635 6158
rect 9305 6155 9371 6158
rect -300 6082 160 6112
rect 3141 6082 3207 6085
rect -300 6080 3207 6082
rect -300 6024 3146 6080
rect 3202 6024 3207 6080
rect -300 6022 3207 6024
rect -300 5992 160 6022
rect 3141 6019 3207 6022
rect 3877 6082 3943 6085
rect 4889 6082 4955 6085
rect 3877 6080 4955 6082
rect 3877 6024 3882 6080
rect 3938 6024 4894 6080
rect 4950 6024 4955 6080
rect 3877 6022 4955 6024
rect 3877 6019 3943 6022
rect 4889 6019 4955 6022
rect 5022 6020 5028 6084
rect 5092 6082 5098 6084
rect 7281 6082 7347 6085
rect 5092 6080 7347 6082
rect 5092 6024 7286 6080
rect 7342 6024 7347 6080
rect 5092 6022 7347 6024
rect 9446 6082 9506 6294
rect 9622 6292 9628 6356
rect 9692 6292 9698 6356
rect 9765 6354 9831 6357
rect 10501 6354 10567 6357
rect 9765 6352 10567 6354
rect 9765 6296 9770 6352
rect 9826 6296 10506 6352
rect 10562 6296 10567 6352
rect 9765 6294 10567 6296
rect 9765 6291 9831 6294
rect 10501 6291 10567 6294
rect 11145 6354 11211 6357
rect 11884 6354 11944 6430
rect 12341 6354 12407 6357
rect 11145 6352 11944 6354
rect 11145 6296 11150 6352
rect 11206 6296 11944 6352
rect 11145 6294 11944 6296
rect 12022 6352 12407 6354
rect 12022 6296 12346 6352
rect 12402 6296 12407 6352
rect 12022 6294 12407 6296
rect 12574 6354 12634 6430
rect 12801 6488 15351 6490
rect 12801 6432 12806 6488
rect 12862 6432 15290 6488
rect 15346 6432 15351 6488
rect 12801 6430 15351 6432
rect 12801 6427 12867 6430
rect 15285 6427 15351 6430
rect 15510 6428 15516 6492
rect 15580 6490 15627 6492
rect 16205 6490 16271 6493
rect 18229 6490 18295 6493
rect 15580 6488 15672 6490
rect 15622 6432 15672 6488
rect 15580 6430 15672 6432
rect 16205 6488 18295 6490
rect 16205 6432 16210 6488
rect 16266 6432 18234 6488
rect 18290 6432 18295 6488
rect 16205 6430 18295 6432
rect 15580 6428 15627 6430
rect 15561 6427 15627 6428
rect 16205 6427 16271 6430
rect 18229 6427 18295 6430
rect 18505 6490 18571 6493
rect 18873 6490 18939 6493
rect 18505 6488 18939 6490
rect 18505 6432 18510 6488
rect 18566 6432 18878 6488
rect 18934 6432 18939 6488
rect 18505 6430 18939 6432
rect 18505 6427 18571 6430
rect 18873 6427 18939 6430
rect 19517 6490 19583 6493
rect 19934 6490 19994 6838
rect 21840 6626 22300 6656
rect 21176 6566 22300 6626
rect 20725 6560 21041 6561
rect 20725 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21041 6560
rect 20725 6495 21041 6496
rect 19517 6488 19994 6490
rect 19517 6432 19522 6488
rect 19578 6432 19994 6488
rect 19517 6430 19994 6432
rect 19517 6427 19583 6430
rect 13077 6354 13143 6357
rect 12574 6352 13143 6354
rect 12574 6296 13082 6352
rect 13138 6296 13143 6352
rect 12574 6294 13143 6296
rect 11145 6291 11211 6294
rect 11053 6218 11119 6221
rect 11605 6218 11671 6221
rect 11053 6216 11671 6218
rect 11053 6160 11058 6216
rect 11114 6160 11610 6216
rect 11666 6160 11671 6216
rect 11053 6158 11671 6160
rect 11053 6155 11119 6158
rect 11605 6155 11671 6158
rect 11789 6218 11855 6221
rect 12022 6218 12082 6294
rect 12341 6291 12407 6294
rect 13077 6291 13143 6294
rect 13629 6354 13695 6357
rect 16757 6354 16823 6357
rect 13629 6352 16823 6354
rect 13629 6296 13634 6352
rect 13690 6296 16762 6352
rect 16818 6296 16823 6352
rect 13629 6294 16823 6296
rect 13629 6291 13695 6294
rect 16757 6291 16823 6294
rect 11789 6216 12082 6218
rect 11789 6160 11794 6216
rect 11850 6160 12082 6216
rect 11789 6158 12082 6160
rect 12341 6218 12407 6221
rect 15009 6218 15075 6221
rect 21176 6218 21236 6566
rect 21840 6536 22300 6566
rect 12341 6216 15075 6218
rect 12341 6160 12346 6216
rect 12402 6160 15014 6216
rect 15070 6160 15075 6216
rect 12341 6158 15075 6160
rect 11789 6155 11855 6158
rect 12341 6155 12407 6158
rect 15009 6155 15075 6158
rect 15150 6158 21236 6218
rect 11053 6082 11119 6085
rect 9446 6080 11119 6082
rect 9446 6024 11058 6080
rect 11114 6024 11119 6080
rect 9446 6022 11119 6024
rect 5092 6020 5098 6022
rect 7281 6019 7347 6022
rect 11053 6019 11119 6022
rect 11421 6082 11487 6085
rect 12893 6082 12959 6085
rect 11421 6080 12959 6082
rect 11421 6024 11426 6080
rect 11482 6024 12898 6080
rect 12954 6024 12959 6080
rect 11421 6022 12959 6024
rect 11421 6019 11487 6022
rect 12893 6019 12959 6022
rect 13905 6082 13971 6085
rect 15150 6082 15210 6158
rect 13905 6080 15210 6082
rect 13905 6024 13910 6080
rect 13966 6024 15210 6080
rect 13905 6022 15210 6024
rect 15285 6082 15351 6085
rect 17677 6082 17743 6085
rect 21840 6082 22300 6112
rect 15285 6080 17743 6082
rect 15285 6024 15290 6080
rect 15346 6024 17682 6080
rect 17738 6024 17743 6080
rect 15285 6022 17743 6024
rect 13905 6019 13971 6022
rect 15285 6019 15351 6022
rect 17677 6019 17743 6022
rect 19290 6022 22300 6082
rect 3418 6016 3734 6017
rect 3418 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3734 6016
rect 3418 5951 3734 5952
rect 8363 6016 8679 6017
rect 8363 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8679 6016
rect 8363 5951 8679 5952
rect 13308 6016 13624 6017
rect 13308 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13624 6016
rect 13308 5951 13624 5952
rect 18253 6016 18569 6017
rect 18253 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18569 6016
rect 18253 5951 18569 5952
rect 2865 5946 2931 5949
rect 2998 5946 3004 5948
rect 2865 5944 3004 5946
rect 2865 5888 2870 5944
rect 2926 5888 3004 5944
rect 2865 5886 3004 5888
rect 2865 5883 2931 5886
rect 2998 5884 3004 5886
rect 3068 5884 3074 5948
rect 6453 5946 6519 5949
rect 6678 5946 6684 5948
rect 6453 5944 6684 5946
rect 6453 5888 6458 5944
rect 6514 5888 6684 5944
rect 6453 5886 6684 5888
rect 6453 5883 6519 5886
rect 6678 5884 6684 5886
rect 6748 5884 6754 5948
rect 10409 5946 10475 5949
rect 9998 5944 10475 5946
rect 9998 5888 10414 5944
rect 10470 5888 10475 5944
rect 9998 5886 10475 5888
rect -300 5810 160 5840
rect 1393 5810 1459 5813
rect -300 5808 1459 5810
rect -300 5752 1398 5808
rect 1454 5752 1459 5808
rect -300 5750 1459 5752
rect -300 5720 160 5750
rect 1393 5747 1459 5750
rect 3049 5810 3115 5813
rect 6494 5810 6500 5812
rect 3049 5808 6500 5810
rect 3049 5752 3054 5808
rect 3110 5752 6500 5808
rect 3049 5750 6500 5752
rect 3049 5747 3115 5750
rect 6494 5748 6500 5750
rect 6564 5748 6570 5812
rect 6913 5810 6979 5813
rect 7782 5810 7788 5812
rect 6913 5808 7788 5810
rect 6913 5752 6918 5808
rect 6974 5752 7788 5808
rect 6913 5750 7788 5752
rect 6913 5747 6979 5750
rect 7782 5748 7788 5750
rect 7852 5748 7858 5812
rect 8661 5810 8727 5813
rect 9213 5812 9279 5813
rect 8886 5810 8892 5812
rect 8661 5808 8892 5810
rect 8661 5752 8666 5808
rect 8722 5752 8892 5808
rect 8661 5750 8892 5752
rect 8661 5747 8727 5750
rect 8886 5748 8892 5750
rect 8956 5748 8962 5812
rect 9213 5810 9260 5812
rect 9168 5808 9260 5810
rect 9168 5752 9218 5808
rect 9168 5750 9260 5752
rect 9213 5748 9260 5750
rect 9324 5748 9330 5812
rect 9213 5747 9279 5748
rect 1945 5674 2011 5677
rect 4153 5674 4219 5677
rect 1945 5672 4219 5674
rect 1945 5616 1950 5672
rect 2006 5616 4158 5672
rect 4214 5616 4219 5672
rect 1945 5614 4219 5616
rect 1945 5611 2011 5614
rect 4153 5611 4219 5614
rect 5533 5676 5599 5677
rect 5533 5672 5580 5676
rect 5644 5674 5650 5676
rect 9213 5674 9279 5677
rect 5644 5672 9279 5674
rect 5533 5616 5538 5672
rect 5644 5616 9218 5672
rect 9274 5616 9279 5672
rect 5533 5612 5580 5616
rect 5644 5614 9279 5616
rect 5644 5612 5650 5614
rect 5533 5611 5599 5612
rect 9213 5611 9279 5614
rect -300 5538 160 5568
rect 3049 5538 3115 5541
rect 6729 5540 6795 5541
rect 6678 5538 6684 5540
rect -300 5536 3115 5538
rect -300 5480 3054 5536
rect 3110 5480 3115 5536
rect -300 5478 3115 5480
rect 6638 5478 6684 5538
rect 6748 5536 6795 5540
rect 6790 5480 6795 5536
rect -300 5448 160 5478
rect 3049 5475 3115 5478
rect 6678 5476 6684 5478
rect 6748 5476 6795 5480
rect 6862 5476 6868 5540
rect 6932 5538 6938 5540
rect 9029 5538 9095 5541
rect 9765 5538 9831 5541
rect 6932 5478 8954 5538
rect 6932 5476 6938 5478
rect 6729 5475 6795 5476
rect 5890 5472 6206 5473
rect 5890 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6206 5472
rect 5890 5407 6206 5408
rect 2405 5402 2471 5405
rect 5349 5402 5415 5405
rect 2405 5400 5415 5402
rect 2405 5344 2410 5400
rect 2466 5344 5354 5400
rect 5410 5344 5415 5400
rect 2405 5342 5415 5344
rect 2405 5339 2471 5342
rect 5349 5339 5415 5342
rect 7414 5340 7420 5404
rect 7484 5402 7490 5404
rect 7649 5402 7715 5405
rect 7484 5400 7715 5402
rect 7484 5344 7654 5400
rect 7710 5344 7715 5400
rect 7484 5342 7715 5344
rect 8894 5402 8954 5478
rect 9029 5536 9831 5538
rect 9029 5480 9034 5536
rect 9090 5480 9770 5536
rect 9826 5480 9831 5536
rect 9029 5478 9831 5480
rect 9029 5475 9095 5478
rect 9765 5475 9831 5478
rect 9998 5402 10058 5886
rect 10409 5883 10475 5886
rect 10777 5946 10843 5949
rect 12198 5946 12204 5948
rect 10777 5944 12204 5946
rect 10777 5888 10782 5944
rect 10838 5888 12204 5944
rect 10777 5886 12204 5888
rect 10777 5883 10843 5886
rect 12198 5884 12204 5886
rect 12268 5884 12274 5948
rect 12341 5946 12407 5949
rect 13118 5946 13124 5948
rect 12341 5944 13124 5946
rect 12341 5888 12346 5944
rect 12402 5888 13124 5944
rect 12341 5886 13124 5888
rect 12341 5883 12407 5886
rect 13118 5884 13124 5886
rect 13188 5884 13194 5948
rect 13854 5884 13860 5948
rect 13924 5946 13930 5948
rect 13997 5946 14063 5949
rect 13924 5944 14063 5946
rect 13924 5888 14002 5944
rect 14058 5888 14063 5944
rect 13924 5886 14063 5888
rect 13924 5884 13930 5886
rect 13997 5883 14063 5886
rect 14181 5946 14247 5949
rect 14406 5946 14412 5948
rect 14181 5944 14412 5946
rect 14181 5888 14186 5944
rect 14242 5888 14412 5944
rect 14181 5886 14412 5888
rect 14181 5883 14247 5886
rect 14406 5884 14412 5886
rect 14476 5884 14482 5948
rect 14549 5946 14615 5949
rect 14549 5944 18154 5946
rect 14549 5888 14554 5944
rect 14610 5888 18154 5944
rect 14549 5886 18154 5888
rect 14549 5883 14615 5886
rect 10409 5810 10475 5813
rect 12014 5810 12020 5812
rect 10409 5808 12020 5810
rect 10409 5752 10414 5808
rect 10470 5752 12020 5808
rect 10409 5750 12020 5752
rect 10409 5747 10475 5750
rect 12014 5748 12020 5750
rect 12084 5748 12090 5812
rect 12709 5810 12775 5813
rect 14825 5810 14891 5813
rect 12709 5808 14891 5810
rect 12709 5752 12714 5808
rect 12770 5752 14830 5808
rect 14886 5752 14891 5808
rect 12709 5750 14891 5752
rect 12709 5747 12775 5750
rect 14825 5747 14891 5750
rect 15009 5810 15075 5813
rect 16665 5810 16731 5813
rect 15009 5808 16731 5810
rect 15009 5752 15014 5808
rect 15070 5752 16670 5808
rect 16726 5752 16731 5808
rect 15009 5750 16731 5752
rect 15009 5747 15075 5750
rect 16665 5747 16731 5750
rect 16849 5810 16915 5813
rect 17677 5810 17743 5813
rect 16849 5808 17743 5810
rect 16849 5752 16854 5808
rect 16910 5752 17682 5808
rect 17738 5752 17743 5808
rect 16849 5750 17743 5752
rect 18094 5810 18154 5886
rect 19290 5810 19350 6022
rect 21840 5992 22300 6022
rect 18094 5750 19350 5810
rect 16849 5747 16915 5750
rect 17677 5747 17743 5750
rect 11053 5674 11119 5677
rect 12525 5674 12591 5677
rect 11053 5672 12450 5674
rect 11053 5616 11058 5672
rect 11114 5616 12450 5672
rect 11053 5614 12450 5616
rect 11053 5611 11119 5614
rect 11513 5538 11579 5541
rect 11646 5538 11652 5540
rect 11513 5536 11652 5538
rect 11513 5480 11518 5536
rect 11574 5480 11652 5536
rect 11513 5478 11652 5480
rect 11513 5475 11579 5478
rect 11646 5476 11652 5478
rect 11716 5476 11722 5540
rect 12390 5538 12450 5614
rect 12525 5672 21236 5674
rect 12525 5616 12530 5672
rect 12586 5616 21236 5672
rect 12525 5614 21236 5616
rect 12525 5611 12591 5614
rect 16205 5538 16271 5541
rect 18137 5538 18203 5541
rect 12390 5478 15578 5538
rect 10835 5472 11151 5473
rect 10835 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11151 5472
rect 10835 5407 11151 5408
rect 8894 5342 10058 5402
rect 11697 5402 11763 5405
rect 12750 5402 12756 5404
rect 11697 5400 12756 5402
rect 11697 5344 11702 5400
rect 11758 5344 12756 5400
rect 11697 5342 12756 5344
rect 7484 5340 7490 5342
rect 7649 5339 7715 5342
rect 11697 5339 11763 5342
rect 12750 5340 12756 5342
rect 12820 5340 12826 5404
rect 12893 5402 12959 5405
rect 13537 5402 13603 5405
rect 12893 5400 13603 5402
rect 12893 5344 12898 5400
rect 12954 5344 13542 5400
rect 13598 5344 13603 5400
rect 12893 5342 13603 5344
rect 12893 5339 12959 5342
rect 13537 5339 13603 5342
rect -300 5266 160 5296
rect 1301 5266 1367 5269
rect -300 5264 1367 5266
rect -300 5208 1306 5264
rect 1362 5208 1367 5264
rect -300 5206 1367 5208
rect -300 5176 160 5206
rect 1301 5203 1367 5206
rect 2865 5266 2931 5269
rect 4429 5266 4495 5269
rect 7833 5266 7899 5269
rect 2865 5264 7899 5266
rect 2865 5208 2870 5264
rect 2926 5208 4434 5264
rect 4490 5208 7838 5264
rect 7894 5208 7899 5264
rect 2865 5206 7899 5208
rect 2865 5203 2931 5206
rect 4429 5203 4495 5206
rect 7833 5203 7899 5206
rect 7966 5204 7972 5268
rect 8036 5266 8042 5268
rect 9397 5266 9463 5269
rect 8036 5264 9463 5266
rect 8036 5208 9402 5264
rect 9458 5208 9463 5264
rect 8036 5206 9463 5208
rect 8036 5204 8042 5206
rect 9397 5203 9463 5206
rect 10542 5204 10548 5268
rect 10612 5266 10618 5268
rect 10777 5266 10843 5269
rect 14181 5266 14247 5269
rect 15142 5266 15148 5268
rect 10612 5264 10843 5266
rect 10612 5208 10782 5264
rect 10838 5208 10843 5264
rect 10612 5206 10843 5208
rect 10612 5204 10618 5206
rect 10777 5203 10843 5206
rect 12942 5264 14247 5266
rect 12942 5208 14186 5264
rect 14242 5208 14247 5264
rect 12942 5206 14247 5208
rect 5206 5068 5212 5132
rect 5276 5130 5282 5132
rect 9070 5130 9076 5132
rect 5276 5070 9076 5130
rect 5276 5068 5282 5070
rect 9070 5068 9076 5070
rect 9140 5068 9146 5132
rect 9305 5130 9371 5133
rect 11053 5130 11119 5133
rect 11329 5132 11395 5133
rect 11278 5130 11284 5132
rect 9305 5128 11119 5130
rect 9305 5072 9310 5128
rect 9366 5072 11058 5128
rect 11114 5072 11119 5128
rect 9305 5070 11119 5072
rect 11238 5070 11284 5130
rect 11348 5128 11395 5132
rect 11605 5132 11671 5133
rect 11605 5130 11652 5132
rect 11390 5072 11395 5128
rect 9305 5067 9371 5070
rect 11053 5067 11119 5070
rect 11278 5068 11284 5070
rect 11348 5068 11395 5072
rect 11560 5128 11652 5130
rect 11560 5072 11610 5128
rect 11560 5070 11652 5072
rect 11329 5067 11395 5068
rect 11605 5068 11652 5070
rect 11716 5068 11722 5132
rect 11881 5130 11947 5133
rect 12801 5130 12867 5133
rect 11881 5128 12867 5130
rect 11881 5072 11886 5128
rect 11942 5072 12806 5128
rect 12862 5072 12867 5128
rect 11881 5070 12867 5072
rect 11605 5067 11671 5068
rect 11881 5067 11947 5070
rect 12801 5067 12867 5070
rect -300 4994 160 5024
rect 4521 4994 4587 4997
rect 7649 4994 7715 4997
rect -300 4934 2100 4994
rect -300 4904 160 4934
rect 2040 4586 2100 4934
rect 4521 4992 7715 4994
rect 4521 4936 4526 4992
rect 4582 4936 7654 4992
rect 7710 4936 7715 4992
rect 4521 4934 7715 4936
rect 4521 4931 4587 4934
rect 7649 4931 7715 4934
rect 9765 4994 9831 4997
rect 10317 4994 10383 4997
rect 9765 4992 10383 4994
rect 9765 4936 9770 4992
rect 9826 4936 10322 4992
rect 10378 4936 10383 4992
rect 9765 4934 10383 4936
rect 9765 4931 9831 4934
rect 10317 4931 10383 4934
rect 10542 4932 10548 4996
rect 10612 4994 10618 4996
rect 10869 4994 10935 4997
rect 12942 4994 13002 5206
rect 14181 5203 14247 5206
rect 14368 5206 15148 5266
rect 13118 5068 13124 5132
rect 13188 5130 13194 5132
rect 14368 5130 14428 5206
rect 15142 5204 15148 5206
rect 15212 5204 15218 5268
rect 15377 5266 15443 5269
rect 15518 5266 15578 5478
rect 16205 5536 18203 5538
rect 16205 5480 16210 5536
rect 16266 5480 18142 5536
rect 18198 5480 18203 5536
rect 16205 5478 18203 5480
rect 16205 5475 16271 5478
rect 18137 5475 18203 5478
rect 18781 5538 18847 5541
rect 19374 5538 19380 5540
rect 18781 5536 19380 5538
rect 18781 5480 18786 5536
rect 18842 5480 19380 5536
rect 18781 5478 19380 5480
rect 18781 5475 18847 5478
rect 19374 5476 19380 5478
rect 19444 5476 19450 5540
rect 21176 5538 21236 5614
rect 21840 5538 22300 5568
rect 21176 5478 22300 5538
rect 15780 5472 16096 5473
rect 15780 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16096 5472
rect 15780 5407 16096 5408
rect 20725 5472 21041 5473
rect 20725 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21041 5472
rect 21840 5448 22300 5478
rect 20725 5407 21041 5408
rect 17033 5402 17099 5405
rect 17953 5402 18019 5405
rect 17033 5400 18019 5402
rect 17033 5344 17038 5400
rect 17094 5344 17958 5400
rect 18014 5344 18019 5400
rect 17033 5342 18019 5344
rect 17033 5339 17099 5342
rect 17953 5339 18019 5342
rect 15377 5264 15578 5266
rect 15377 5208 15382 5264
rect 15438 5208 15578 5264
rect 15377 5206 15578 5208
rect 15745 5266 15811 5269
rect 16481 5266 16547 5269
rect 15745 5264 16547 5266
rect 15745 5208 15750 5264
rect 15806 5208 16486 5264
rect 16542 5208 16547 5264
rect 15745 5206 16547 5208
rect 15377 5203 15443 5206
rect 15745 5203 15811 5206
rect 16481 5203 16547 5206
rect 16849 5266 16915 5269
rect 16849 5264 20730 5266
rect 16849 5208 16854 5264
rect 16910 5208 20730 5264
rect 16849 5206 20730 5208
rect 16849 5203 16915 5206
rect 13188 5070 14428 5130
rect 14549 5130 14615 5133
rect 14733 5130 14799 5133
rect 14549 5128 14799 5130
rect 14549 5072 14554 5128
rect 14610 5072 14738 5128
rect 14794 5072 14799 5128
rect 14549 5070 14799 5072
rect 13188 5068 13194 5070
rect 14549 5067 14615 5070
rect 14733 5067 14799 5070
rect 15193 5130 15259 5133
rect 19425 5130 19491 5133
rect 15193 5128 19491 5130
rect 15193 5072 15198 5128
rect 15254 5072 19430 5128
rect 19486 5072 19491 5128
rect 15193 5070 19491 5072
rect 15193 5067 15259 5070
rect 19425 5067 19491 5070
rect 10612 4992 10935 4994
rect 10612 4936 10874 4992
rect 10930 4936 10935 4992
rect 10612 4934 10935 4936
rect 10612 4932 10618 4934
rect 10869 4931 10935 4934
rect 11102 4934 13002 4994
rect 14181 4994 14247 4997
rect 14549 4994 14615 4997
rect 17033 4994 17099 4997
rect 14181 4992 14290 4994
rect 14181 4936 14186 4992
rect 14242 4936 14290 4992
rect 3418 4928 3734 4929
rect 3418 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3734 4928
rect 3418 4863 3734 4864
rect 8363 4928 8679 4929
rect 8363 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8679 4928
rect 8363 4863 8679 4864
rect 4981 4858 5047 4861
rect 7005 4860 7071 4861
rect 6862 4858 6868 4860
rect 4110 4798 4584 4858
rect 3601 4722 3667 4725
rect 3785 4722 3851 4725
rect 4110 4722 4170 4798
rect 3601 4720 4170 4722
rect 3601 4664 3606 4720
rect 3662 4664 3790 4720
rect 3846 4664 4170 4720
rect 3601 4662 4170 4664
rect 3601 4659 3667 4662
rect 3785 4659 3851 4662
rect 3969 4586 4035 4589
rect 2040 4584 4035 4586
rect 2040 4528 3974 4584
rect 4030 4528 4035 4584
rect 2040 4526 4035 4528
rect 4524 4586 4584 4798
rect 4981 4856 6868 4858
rect 4981 4800 4986 4856
rect 5042 4800 6868 4856
rect 4981 4798 6868 4800
rect 4981 4795 5047 4798
rect 6862 4796 6868 4798
rect 6932 4796 6938 4860
rect 7005 4856 7052 4860
rect 7116 4858 7122 4860
rect 7005 4800 7010 4856
rect 7005 4796 7052 4800
rect 7116 4798 7162 4858
rect 7116 4796 7122 4798
rect 7966 4796 7972 4860
rect 8036 4858 8042 4860
rect 8201 4858 8267 4861
rect 8036 4856 8267 4858
rect 8036 4800 8206 4856
rect 8262 4800 8267 4856
rect 8036 4798 8267 4800
rect 8036 4796 8042 4798
rect 7005 4795 7071 4796
rect 8201 4795 8267 4798
rect 9765 4858 9831 4861
rect 11102 4858 11162 4934
rect 14181 4931 14290 4936
rect 14549 4992 17099 4994
rect 14549 4936 14554 4992
rect 14610 4936 17038 4992
rect 17094 4936 17099 4992
rect 14549 4934 17099 4936
rect 20670 4994 20730 5206
rect 21840 4994 22300 5024
rect 20670 4934 22300 4994
rect 14549 4931 14615 4934
rect 17033 4931 17099 4934
rect 13308 4928 13624 4929
rect 13308 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13624 4928
rect 13308 4863 13624 4864
rect 11697 4860 11763 4861
rect 11646 4858 11652 4860
rect 9765 4856 11162 4858
rect 9765 4800 9770 4856
rect 9826 4800 11162 4856
rect 9765 4798 11162 4800
rect 11606 4798 11652 4858
rect 11716 4856 11763 4860
rect 11758 4800 11763 4856
rect 9765 4795 9831 4798
rect 11646 4796 11652 4798
rect 11716 4796 11763 4800
rect 11830 4796 11836 4860
rect 11900 4858 11906 4860
rect 12065 4858 12131 4861
rect 11900 4856 12131 4858
rect 11900 4800 12070 4856
rect 12126 4800 12131 4856
rect 11900 4798 12131 4800
rect 11900 4796 11906 4798
rect 11697 4795 11763 4796
rect 12065 4795 12131 4798
rect 12198 4796 12204 4860
rect 12268 4858 12274 4860
rect 12433 4858 12499 4861
rect 12268 4856 12499 4858
rect 12268 4800 12438 4856
rect 12494 4800 12499 4856
rect 12268 4798 12499 4800
rect 12268 4796 12274 4798
rect 12433 4795 12499 4798
rect 12709 4858 12775 4861
rect 13169 4858 13235 4861
rect 12709 4856 13235 4858
rect 12709 4800 12714 4856
rect 12770 4800 13174 4856
rect 13230 4800 13235 4856
rect 12709 4798 13235 4800
rect 12709 4795 12775 4798
rect 13169 4795 13235 4798
rect 4705 4722 4771 4725
rect 5441 4722 5507 4725
rect 4705 4720 5507 4722
rect 4705 4664 4710 4720
rect 4766 4664 5446 4720
rect 5502 4664 5507 4720
rect 4705 4662 5507 4664
rect 4705 4659 4771 4662
rect 5441 4659 5507 4662
rect 5574 4660 5580 4724
rect 5644 4722 5650 4724
rect 6862 4722 6868 4724
rect 5644 4662 6868 4722
rect 5644 4660 5650 4662
rect 6862 4660 6868 4662
rect 6932 4660 6938 4724
rect 10358 4660 10364 4724
rect 10428 4722 10434 4724
rect 10501 4722 10567 4725
rect 10428 4720 10567 4722
rect 10428 4664 10506 4720
rect 10562 4664 10567 4720
rect 10428 4662 10567 4664
rect 10428 4660 10434 4662
rect 10501 4659 10567 4662
rect 10869 4722 10935 4725
rect 12014 4722 12020 4724
rect 10869 4720 12020 4722
rect 10869 4664 10874 4720
rect 10930 4664 12020 4720
rect 10869 4662 12020 4664
rect 10869 4659 10935 4662
rect 12014 4660 12020 4662
rect 12084 4660 12090 4724
rect 12157 4722 12223 4725
rect 12341 4722 12407 4725
rect 12157 4720 12407 4722
rect 12157 4664 12162 4720
rect 12218 4664 12346 4720
rect 12402 4664 12407 4720
rect 12157 4662 12407 4664
rect 12157 4659 12223 4662
rect 12341 4659 12407 4662
rect 12566 4660 12572 4724
rect 12636 4722 12642 4724
rect 13169 4722 13235 4725
rect 14089 4722 14155 4725
rect 12636 4662 13002 4722
rect 12636 4660 12642 4662
rect 6729 4586 6795 4589
rect 4524 4584 6795 4586
rect 4524 4528 6734 4584
rect 6790 4528 6795 4584
rect 4524 4526 6795 4528
rect 3969 4523 4035 4526
rect 6729 4523 6795 4526
rect 6862 4524 6868 4588
rect 6932 4586 6938 4588
rect 10041 4586 10107 4589
rect 6932 4584 10107 4586
rect 6932 4528 10046 4584
rect 10102 4528 10107 4584
rect 6932 4526 10107 4528
rect 6932 4524 6938 4526
rect 10041 4523 10107 4526
rect 11053 4586 11119 4589
rect 11278 4586 11284 4588
rect 11053 4584 11284 4586
rect 11053 4528 11058 4584
rect 11114 4528 11284 4584
rect 11053 4526 11284 4528
rect 11053 4523 11119 4526
rect 11278 4524 11284 4526
rect 11348 4524 11354 4588
rect 11421 4584 11487 4589
rect 11421 4528 11426 4584
rect 11482 4528 11487 4584
rect 11421 4523 11487 4528
rect 11605 4586 11671 4589
rect 12198 4586 12204 4588
rect 11605 4584 12204 4586
rect 11605 4528 11610 4584
rect 11666 4528 12204 4584
rect 11605 4526 12204 4528
rect 11605 4523 11671 4526
rect 12198 4524 12204 4526
rect 12268 4524 12274 4588
rect 12942 4586 13002 4662
rect 13169 4720 14155 4722
rect 13169 4664 13174 4720
rect 13230 4664 14094 4720
rect 14150 4664 14155 4720
rect 13169 4662 14155 4664
rect 14230 4722 14290 4931
rect 18253 4928 18569 4929
rect 18253 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18569 4928
rect 21840 4904 22300 4934
rect 18253 4863 18569 4864
rect 14365 4858 14431 4861
rect 17493 4858 17559 4861
rect 14365 4856 17559 4858
rect 14365 4800 14370 4856
rect 14426 4800 17498 4856
rect 17554 4800 17559 4856
rect 14365 4798 17559 4800
rect 14365 4795 14431 4798
rect 17493 4795 17559 4798
rect 14230 4662 14474 4722
rect 13169 4659 13235 4662
rect 14089 4659 14155 4662
rect 14222 4586 14228 4588
rect 12942 4526 14228 4586
rect 14222 4524 14228 4526
rect 14292 4524 14298 4588
rect 3785 4450 3851 4453
rect 6729 4452 6795 4453
rect 4838 4450 4844 4452
rect 3785 4448 4844 4450
rect 3785 4392 3790 4448
rect 3846 4392 4844 4448
rect 3785 4390 4844 4392
rect 3785 4387 3851 4390
rect 4838 4388 4844 4390
rect 4908 4388 4914 4452
rect 6678 4388 6684 4452
rect 6748 4450 6795 4452
rect 6748 4448 6840 4450
rect 6790 4392 6840 4448
rect 6748 4390 6840 4392
rect 6748 4388 6795 4390
rect 7046 4388 7052 4452
rect 7116 4450 7122 4452
rect 7281 4450 7347 4453
rect 7116 4448 7347 4450
rect 7116 4392 7286 4448
rect 7342 4392 7347 4448
rect 7116 4390 7347 4392
rect 7116 4388 7122 4390
rect 6729 4387 6795 4388
rect 7281 4387 7347 4390
rect 5890 4384 6206 4385
rect 5890 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6206 4384
rect 5890 4319 6206 4320
rect 10835 4384 11151 4385
rect 10835 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11151 4384
rect 10835 4319 11151 4320
rect 4153 4314 4219 4317
rect 11424 4314 11484 4523
rect 11973 4450 12039 4453
rect 12433 4450 12499 4453
rect 11973 4448 12499 4450
rect 11973 4392 11978 4448
rect 12034 4392 12438 4448
rect 12494 4392 12499 4448
rect 11973 4390 12499 4392
rect 11973 4387 12039 4390
rect 12433 4387 12499 4390
rect 12750 4388 12756 4452
rect 12820 4450 12826 4452
rect 12893 4450 12959 4453
rect 12820 4448 12959 4450
rect 12820 4392 12898 4448
rect 12954 4392 12959 4448
rect 12820 4390 12959 4392
rect 12820 4388 12826 4390
rect 12893 4387 12959 4390
rect 13118 4388 13124 4452
rect 13188 4450 13194 4452
rect 14181 4450 14247 4453
rect 13188 4448 14247 4450
rect 13188 4392 14186 4448
rect 14242 4392 14247 4448
rect 13188 4390 14247 4392
rect 14414 4450 14474 4662
rect 15142 4660 15148 4724
rect 15212 4722 15218 4724
rect 16849 4722 16915 4725
rect 15212 4720 16915 4722
rect 15212 4664 16854 4720
rect 16910 4664 16915 4720
rect 15212 4662 16915 4664
rect 15212 4660 15218 4662
rect 16849 4659 16915 4662
rect 16982 4660 16988 4724
rect 17052 4722 17058 4724
rect 18229 4722 18295 4725
rect 17052 4720 18295 4722
rect 17052 4664 18234 4720
rect 18290 4664 18295 4720
rect 17052 4662 18295 4664
rect 17052 4660 17058 4662
rect 18229 4659 18295 4662
rect 14641 4586 14707 4589
rect 19885 4586 19951 4589
rect 14641 4584 19951 4586
rect 14641 4528 14646 4584
rect 14702 4528 19890 4584
rect 19946 4528 19951 4584
rect 14641 4526 19951 4528
rect 14641 4523 14707 4526
rect 19885 4523 19951 4526
rect 15653 4450 15719 4453
rect 14414 4448 15719 4450
rect 14414 4392 15658 4448
rect 15714 4392 15719 4448
rect 14414 4390 15719 4392
rect 13188 4388 13194 4390
rect 14181 4387 14247 4390
rect 15653 4387 15719 4390
rect 16297 4450 16363 4453
rect 19926 4450 19932 4452
rect 16297 4448 19932 4450
rect 16297 4392 16302 4448
rect 16358 4392 19932 4448
rect 16297 4390 19932 4392
rect 16297 4387 16363 4390
rect 19926 4388 19932 4390
rect 19996 4388 20002 4452
rect 21840 4450 22300 4480
rect 21636 4390 22300 4450
rect 15780 4384 16096 4385
rect 15780 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16096 4384
rect 15780 4319 16096 4320
rect 20725 4384 21041 4385
rect 20725 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21041 4384
rect 20725 4319 21041 4320
rect 11881 4314 11947 4317
rect 4153 4312 5780 4314
rect 4153 4256 4158 4312
rect 4214 4256 5780 4312
rect 4153 4254 5780 4256
rect 11424 4312 11947 4314
rect 11424 4256 11886 4312
rect 11942 4256 11947 4312
rect 11424 4254 11947 4256
rect 4153 4251 4219 4254
rect 1526 4116 1532 4180
rect 1596 4178 1602 4180
rect 5574 4178 5580 4180
rect 1596 4118 5580 4178
rect 1596 4116 1602 4118
rect 5574 4116 5580 4118
rect 5644 4116 5650 4180
rect 5720 4178 5780 4254
rect 11881 4251 11947 4254
rect 12249 4314 12315 4317
rect 12382 4314 12388 4316
rect 12249 4312 12388 4314
rect 12249 4256 12254 4312
rect 12310 4256 12388 4312
rect 12249 4254 12388 4256
rect 12249 4251 12315 4254
rect 12382 4252 12388 4254
rect 12452 4252 12458 4316
rect 12750 4252 12756 4316
rect 12820 4314 12826 4316
rect 15285 4314 15351 4317
rect 19241 4316 19307 4317
rect 12820 4312 15351 4314
rect 12820 4256 15290 4312
rect 15346 4256 15351 4312
rect 12820 4254 15351 4256
rect 12820 4252 12826 4254
rect 15285 4251 15351 4254
rect 19190 4252 19196 4316
rect 19260 4314 19307 4316
rect 21636 4314 21696 4390
rect 21840 4360 22300 4390
rect 19260 4312 19352 4314
rect 19302 4256 19352 4312
rect 19260 4254 19352 4256
rect 21590 4254 21696 4314
rect 19260 4252 19307 4254
rect 19241 4251 19307 4252
rect 13169 4178 13235 4181
rect 5720 4176 13235 4178
rect 5720 4120 13174 4176
rect 13230 4120 13235 4176
rect 5720 4118 13235 4120
rect 13169 4115 13235 4118
rect 13353 4178 13419 4181
rect 14774 4178 14780 4180
rect 13353 4176 14780 4178
rect 13353 4120 13358 4176
rect 13414 4120 14780 4176
rect 13353 4118 14780 4120
rect 13353 4115 13419 4118
rect 14774 4116 14780 4118
rect 14844 4116 14850 4180
rect 16481 4178 16547 4181
rect 21590 4178 21650 4254
rect 15196 4176 16547 4178
rect 15196 4120 16486 4176
rect 16542 4120 16547 4176
rect 15196 4118 16547 4120
rect 3182 3980 3188 4044
rect 3252 4042 3258 4044
rect 4061 4042 4127 4045
rect 7281 4042 7347 4045
rect 3252 3982 3986 4042
rect 3252 3980 3258 3982
rect 3926 3906 3986 3982
rect 4061 4040 7347 4042
rect 4061 3984 4066 4040
rect 4122 3984 7286 4040
rect 7342 3984 7347 4040
rect 4061 3982 7347 3984
rect 4061 3979 4127 3982
rect 7281 3979 7347 3982
rect 11145 4042 11211 4045
rect 12014 4042 12020 4044
rect 11145 4040 12020 4042
rect 11145 3984 11150 4040
rect 11206 3984 12020 4040
rect 11145 3982 12020 3984
rect 11145 3979 11211 3982
rect 12014 3980 12020 3982
rect 12084 4042 12090 4044
rect 12433 4042 12499 4045
rect 13261 4042 13327 4045
rect 12084 4040 12499 4042
rect 12084 3984 12438 4040
rect 12494 3984 12499 4040
rect 12084 3982 12499 3984
rect 12084 3980 12090 3982
rect 12433 3979 12499 3982
rect 12574 4040 13327 4042
rect 12574 3984 13266 4040
rect 13322 3984 13327 4040
rect 12574 3982 13327 3984
rect 4153 3906 4219 3909
rect 7833 3906 7899 3909
rect 9990 3906 9996 3908
rect 3926 3904 7899 3906
rect 3926 3848 4158 3904
rect 4214 3848 7838 3904
rect 7894 3848 7899 3904
rect 3926 3846 7899 3848
rect 4153 3843 4219 3846
rect 7833 3843 7899 3846
rect 9814 3846 9996 3906
rect 3418 3840 3734 3841
rect 3418 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3734 3840
rect 3418 3775 3734 3776
rect 8363 3840 8679 3841
rect 8363 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8679 3840
rect 8363 3775 8679 3776
rect 4245 3770 4311 3773
rect 4470 3770 4476 3772
rect 4245 3768 4476 3770
rect 4245 3712 4250 3768
rect 4306 3712 4476 3768
rect 4245 3710 4476 3712
rect 4245 3707 4311 3710
rect 4470 3708 4476 3710
rect 4540 3708 4546 3772
rect 9814 3637 9874 3846
rect 9990 3844 9996 3846
rect 10060 3844 10066 3908
rect 10225 3906 10291 3909
rect 11646 3906 11652 3908
rect 10225 3904 11652 3906
rect 10225 3848 10230 3904
rect 10286 3848 11652 3904
rect 10225 3846 11652 3848
rect 10225 3843 10291 3846
rect 11646 3844 11652 3846
rect 11716 3844 11722 3908
rect 11789 3906 11855 3909
rect 12574 3906 12634 3982
rect 13261 3979 13327 3982
rect 13445 4042 13511 4045
rect 15196 4042 15256 4118
rect 16481 4115 16547 4118
rect 16806 4118 21650 4178
rect 16806 4042 16866 4118
rect 13445 4040 15256 4042
rect 13445 3984 13450 4040
rect 13506 3984 15256 4040
rect 13445 3982 15256 3984
rect 15380 3982 16866 4042
rect 16941 4042 17007 4045
rect 17350 4042 17356 4044
rect 16941 4040 17356 4042
rect 16941 3984 16946 4040
rect 17002 3984 17356 4040
rect 16941 3982 17356 3984
rect 13445 3979 13511 3982
rect 11789 3904 12634 3906
rect 11789 3848 11794 3904
rect 11850 3848 12634 3904
rect 11789 3846 12634 3848
rect 12801 3906 12867 3909
rect 13010 3906 13076 3909
rect 12801 3904 13076 3906
rect 12801 3848 12806 3904
rect 12862 3848 13015 3904
rect 13071 3848 13076 3904
rect 12801 3846 13076 3848
rect 11789 3843 11855 3846
rect 12801 3843 12867 3846
rect 13010 3843 13076 3846
rect 13905 3906 13971 3909
rect 15380 3906 15440 3982
rect 16941 3979 17007 3982
rect 17350 3980 17356 3982
rect 17420 3980 17426 4044
rect 13905 3904 15440 3906
rect 13905 3848 13910 3904
rect 13966 3848 15440 3904
rect 13905 3846 15440 3848
rect 13905 3843 13971 3846
rect 15510 3844 15516 3908
rect 15580 3906 15586 3908
rect 15745 3906 15811 3909
rect 15580 3904 15811 3906
rect 15580 3848 15750 3904
rect 15806 3848 15811 3904
rect 15580 3846 15811 3848
rect 15580 3844 15586 3846
rect 15745 3843 15811 3846
rect 16481 3906 16547 3909
rect 17585 3906 17651 3909
rect 16481 3904 17651 3906
rect 16481 3848 16486 3904
rect 16542 3848 17590 3904
rect 17646 3848 17651 3904
rect 16481 3846 17651 3848
rect 16481 3843 16547 3846
rect 17585 3843 17651 3846
rect 18689 3906 18755 3909
rect 21840 3906 22300 3936
rect 18689 3904 22300 3906
rect 18689 3848 18694 3904
rect 18750 3848 22300 3904
rect 18689 3846 22300 3848
rect 18689 3843 18755 3846
rect 13308 3840 13624 3841
rect 13308 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13624 3840
rect 13308 3775 13624 3776
rect 18253 3840 18569 3841
rect 18253 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18569 3840
rect 21840 3816 22300 3846
rect 18253 3775 18569 3776
rect 10041 3770 10107 3773
rect 12566 3770 12572 3772
rect 10041 3768 12572 3770
rect 10041 3712 10046 3768
rect 10102 3712 12572 3768
rect 10041 3710 12572 3712
rect 10041 3707 10107 3710
rect 12566 3708 12572 3710
rect 12636 3708 12642 3772
rect 12893 3770 12959 3773
rect 13118 3770 13124 3772
rect 12893 3768 13124 3770
rect 12893 3712 12898 3768
rect 12954 3712 13124 3768
rect 12893 3710 13124 3712
rect 12893 3707 12959 3710
rect 13118 3708 13124 3710
rect 13188 3708 13194 3772
rect 13900 3708 13906 3772
rect 13970 3770 13976 3772
rect 14089 3770 14155 3773
rect 13970 3768 14155 3770
rect 13970 3712 14094 3768
rect 14150 3712 14155 3768
rect 13970 3710 14155 3712
rect 13970 3708 13976 3710
rect 14089 3707 14155 3710
rect 14222 3708 14228 3772
rect 14292 3770 14298 3772
rect 14590 3770 14596 3772
rect 14292 3710 14596 3770
rect 14292 3708 14298 3710
rect 14590 3708 14596 3710
rect 14660 3708 14666 3772
rect 14733 3770 14799 3773
rect 14958 3770 14964 3772
rect 14733 3768 14964 3770
rect 14733 3712 14738 3768
rect 14794 3712 14964 3768
rect 14733 3710 14964 3712
rect 14733 3707 14799 3710
rect 14958 3708 14964 3710
rect 15028 3708 15034 3772
rect 15142 3708 15148 3772
rect 15212 3770 15218 3772
rect 16757 3770 16823 3773
rect 15212 3768 16823 3770
rect 15212 3712 16762 3768
rect 16818 3712 16823 3768
rect 15212 3710 16823 3712
rect 15212 3708 15218 3710
rect 16757 3707 16823 3710
rect 17493 3772 17559 3773
rect 17493 3768 17540 3772
rect 17604 3770 17610 3772
rect 17493 3712 17498 3768
rect 17493 3708 17540 3712
rect 17604 3710 17650 3770
rect 17604 3708 17610 3710
rect 17493 3707 17559 3708
rect 2589 3634 2655 3637
rect 6545 3634 6611 3637
rect 2589 3632 6611 3634
rect 2589 3576 2594 3632
rect 2650 3576 6550 3632
rect 6606 3576 6611 3632
rect 2589 3574 6611 3576
rect 2589 3571 2655 3574
rect 6545 3571 6611 3574
rect 7598 3572 7604 3636
rect 7668 3634 7674 3636
rect 8385 3634 8451 3637
rect 7668 3632 8451 3634
rect 7668 3576 8390 3632
rect 8446 3576 8451 3632
rect 7668 3574 8451 3576
rect 9814 3632 9923 3637
rect 9814 3576 9862 3632
rect 9918 3576 9923 3632
rect 9814 3574 9923 3576
rect 7668 3572 7674 3574
rect 8385 3571 8451 3574
rect 9857 3571 9923 3574
rect 10501 3634 10567 3637
rect 11237 3634 11303 3637
rect 10501 3632 11303 3634
rect 10501 3576 10506 3632
rect 10562 3576 11242 3632
rect 11298 3576 11303 3632
rect 10501 3574 11303 3576
rect 10501 3571 10567 3574
rect 11237 3571 11303 3574
rect 11605 3634 11671 3637
rect 12433 3634 12499 3637
rect 11605 3632 12499 3634
rect 11605 3576 11610 3632
rect 11666 3576 12438 3632
rect 12494 3576 12499 3632
rect 11605 3574 12499 3576
rect 11605 3571 11671 3574
rect 12433 3571 12499 3574
rect 12566 3572 12572 3636
rect 12636 3634 12642 3636
rect 14958 3634 14964 3636
rect 12636 3574 14964 3634
rect 12636 3572 12642 3574
rect 14958 3572 14964 3574
rect 15028 3572 15034 3636
rect 15101 3634 15167 3637
rect 18229 3634 18295 3637
rect 15101 3632 18295 3634
rect 15101 3576 15106 3632
rect 15162 3576 18234 3632
rect 18290 3576 18295 3632
rect 15101 3574 18295 3576
rect 15101 3571 15167 3574
rect 18229 3571 18295 3574
rect 2405 3498 2471 3501
rect 6821 3498 6887 3501
rect 2405 3496 6887 3498
rect 2405 3440 2410 3496
rect 2466 3440 6826 3496
rect 6882 3440 6887 3496
rect 2405 3438 6887 3440
rect 2405 3435 2471 3438
rect 6821 3435 6887 3438
rect 9305 3498 9371 3501
rect 15837 3498 15903 3501
rect 9305 3496 15903 3498
rect 9305 3440 9310 3496
rect 9366 3440 15842 3496
rect 15898 3440 15903 3496
rect 9305 3438 15903 3440
rect 9305 3435 9371 3438
rect 15837 3435 15903 3438
rect 16021 3498 16087 3501
rect 18597 3498 18663 3501
rect 16021 3496 18663 3498
rect 16021 3440 16026 3496
rect 16082 3440 18602 3496
rect 18658 3440 18663 3496
rect 16021 3438 18663 3440
rect 16021 3435 16087 3438
rect 18597 3435 18663 3438
rect 6678 3300 6684 3364
rect 6748 3362 6754 3364
rect 7005 3362 7071 3365
rect 6748 3360 7071 3362
rect 6748 3304 7010 3360
rect 7066 3304 7071 3360
rect 6748 3302 7071 3304
rect 6748 3300 6754 3302
rect 7005 3299 7071 3302
rect 9029 3362 9095 3365
rect 9806 3362 9812 3364
rect 9029 3360 9812 3362
rect 9029 3304 9034 3360
rect 9090 3304 9812 3360
rect 9029 3302 9812 3304
rect 9029 3299 9095 3302
rect 9806 3300 9812 3302
rect 9876 3300 9882 3364
rect 10542 3300 10548 3364
rect 10612 3362 10618 3364
rect 10685 3362 10751 3365
rect 10612 3360 10751 3362
rect 10612 3304 10690 3360
rect 10746 3304 10751 3360
rect 10612 3302 10751 3304
rect 10612 3300 10618 3302
rect 10685 3299 10751 3302
rect 11278 3300 11284 3364
rect 11348 3362 11354 3364
rect 11513 3362 11579 3365
rect 12433 3364 12499 3365
rect 12382 3362 12388 3364
rect 11348 3360 11579 3362
rect 11348 3304 11518 3360
rect 11574 3304 11579 3360
rect 11348 3302 11579 3304
rect 12342 3302 12388 3362
rect 12452 3360 12499 3364
rect 12494 3304 12499 3360
rect 11348 3300 11354 3302
rect 11513 3299 11579 3302
rect 12382 3300 12388 3302
rect 12452 3300 12499 3304
rect 12433 3299 12499 3300
rect 12709 3362 12775 3365
rect 15101 3362 15167 3365
rect 15469 3362 15535 3365
rect 12709 3360 15167 3362
rect 12709 3304 12714 3360
rect 12770 3304 15106 3360
rect 15162 3304 15167 3360
rect 12709 3302 15167 3304
rect 12709 3299 12775 3302
rect 15101 3299 15167 3302
rect 15334 3360 15535 3362
rect 15334 3304 15474 3360
rect 15530 3304 15535 3360
rect 15334 3302 15535 3304
rect 5890 3296 6206 3297
rect 5890 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6206 3296
rect 5890 3231 6206 3232
rect 10835 3296 11151 3297
rect 10835 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11151 3296
rect 10835 3231 11151 3232
rect 6269 3228 6335 3229
rect 6269 3224 6316 3228
rect 6380 3226 6386 3228
rect 7189 3226 7255 3229
rect 6269 3168 6274 3224
rect 6269 3164 6316 3168
rect 6380 3166 6426 3226
rect 7054 3224 7255 3226
rect 7054 3168 7194 3224
rect 7250 3168 7255 3224
rect 7054 3166 7255 3168
rect 6380 3164 6386 3166
rect 6269 3163 6335 3164
rect 4981 3090 5047 3093
rect 5206 3090 5212 3092
rect 4981 3088 5212 3090
rect 4981 3032 4986 3088
rect 5042 3032 5212 3088
rect 4981 3030 5212 3032
rect 4981 3027 5047 3030
rect 5206 3028 5212 3030
rect 5276 3028 5282 3092
rect 5574 3028 5580 3092
rect 5644 3090 5650 3092
rect 6177 3090 6243 3093
rect 5644 3088 6243 3090
rect 5644 3032 6182 3088
rect 6238 3032 6243 3088
rect 5644 3030 6243 3032
rect 5644 3028 5650 3030
rect 6177 3027 6243 3030
rect 6913 3090 6979 3093
rect 7054 3090 7114 3166
rect 7189 3163 7255 3166
rect 7925 3226 7991 3229
rect 8150 3226 8156 3228
rect 7925 3224 8156 3226
rect 7925 3168 7930 3224
rect 7986 3168 8156 3224
rect 7925 3166 8156 3168
rect 7925 3163 7991 3166
rect 8150 3164 8156 3166
rect 8220 3164 8226 3228
rect 9213 3226 9279 3229
rect 10174 3226 10180 3228
rect 9213 3224 10180 3226
rect 9213 3168 9218 3224
rect 9274 3168 10180 3224
rect 9213 3166 10180 3168
rect 9213 3163 9279 3166
rect 10174 3164 10180 3166
rect 10244 3164 10250 3228
rect 11278 3164 11284 3228
rect 11348 3226 11354 3228
rect 11881 3226 11947 3229
rect 12985 3226 13051 3229
rect 11348 3166 11714 3226
rect 11348 3164 11354 3166
rect 9438 3090 9444 3092
rect 6913 3088 7114 3090
rect 6913 3032 6918 3088
rect 6974 3032 7114 3088
rect 6913 3030 7114 3032
rect 8158 3030 9444 3090
rect 6913 3027 6979 3030
rect 6729 2954 6795 2957
rect 7598 2954 7604 2956
rect 6729 2952 7604 2954
rect 6729 2896 6734 2952
rect 6790 2896 7604 2952
rect 6729 2894 7604 2896
rect 6729 2891 6795 2894
rect 7598 2892 7604 2894
rect 7668 2892 7674 2956
rect 3418 2752 3734 2753
rect 3418 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3734 2752
rect 3418 2687 3734 2688
rect 473 2684 539 2685
rect 422 2682 428 2684
rect 382 2622 428 2682
rect 492 2680 539 2684
rect 534 2624 539 2680
rect 422 2620 428 2622
rect 492 2620 539 2624
rect 606 2620 612 2684
rect 676 2682 682 2684
rect 1853 2682 1919 2685
rect 676 2680 1919 2682
rect 676 2624 1858 2680
rect 1914 2624 1919 2680
rect 676 2622 1919 2624
rect 676 2620 682 2622
rect 473 2619 539 2620
rect 1853 2619 1919 2622
rect 2497 2682 2563 2685
rect 4337 2684 4403 2685
rect 2630 2682 2636 2684
rect 2497 2680 2636 2682
rect 2497 2624 2502 2680
rect 2558 2624 2636 2680
rect 2497 2622 2636 2624
rect 2497 2619 2563 2622
rect 2630 2620 2636 2622
rect 2700 2620 2706 2684
rect 4286 2620 4292 2684
rect 4356 2682 4403 2684
rect 7281 2682 7347 2685
rect 8158 2682 8218 3030
rect 9438 3028 9444 3030
rect 9508 3028 9514 3092
rect 9990 3028 9996 3092
rect 10060 3028 10066 3092
rect 10777 3090 10843 3093
rect 11462 3090 11468 3092
rect 10777 3088 11468 3090
rect 10777 3032 10782 3088
rect 10838 3032 11468 3088
rect 10777 3030 11468 3032
rect 9305 2954 9371 2957
rect 9998 2954 10058 3028
rect 10777 3027 10843 3030
rect 11462 3028 11468 3030
rect 11532 3028 11538 3092
rect 11654 3090 11714 3166
rect 11881 3224 13051 3226
rect 11881 3168 11886 3224
rect 11942 3168 12990 3224
rect 13046 3168 13051 3224
rect 11881 3166 13051 3168
rect 11881 3163 11947 3166
rect 12985 3163 13051 3166
rect 13118 3164 13124 3228
rect 13188 3226 13194 3228
rect 14181 3226 14247 3229
rect 13188 3224 14247 3226
rect 13188 3168 14186 3224
rect 14242 3168 14247 3224
rect 13188 3166 14247 3168
rect 13188 3164 13194 3166
rect 14181 3163 14247 3166
rect 14365 3226 14431 3229
rect 14825 3226 14891 3229
rect 14365 3224 14891 3226
rect 14365 3168 14370 3224
rect 14426 3168 14830 3224
rect 14886 3168 14891 3224
rect 14365 3166 14891 3168
rect 14365 3163 14431 3166
rect 14825 3163 14891 3166
rect 15101 3226 15167 3229
rect 15334 3226 15394 3302
rect 15469 3299 15535 3302
rect 16389 3362 16455 3365
rect 16614 3362 16620 3364
rect 16389 3360 16620 3362
rect 16389 3304 16394 3360
rect 16450 3304 16620 3360
rect 16389 3302 16620 3304
rect 16389 3299 16455 3302
rect 16614 3300 16620 3302
rect 16684 3300 16690 3364
rect 16757 3362 16823 3365
rect 18597 3362 18663 3365
rect 16757 3360 18663 3362
rect 16757 3304 16762 3360
rect 16818 3304 18602 3360
rect 18658 3304 18663 3360
rect 16757 3302 18663 3304
rect 16757 3299 16823 3302
rect 18597 3299 18663 3302
rect 21265 3362 21331 3365
rect 21840 3362 22300 3392
rect 21265 3360 22300 3362
rect 21265 3304 21270 3360
rect 21326 3304 22300 3360
rect 21265 3302 22300 3304
rect 21265 3299 21331 3302
rect 15780 3296 16096 3297
rect 15780 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16096 3296
rect 15780 3231 16096 3232
rect 20725 3296 21041 3297
rect 20725 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21041 3296
rect 21840 3272 22300 3302
rect 20725 3231 21041 3232
rect 15101 3224 15394 3226
rect 15101 3168 15106 3224
rect 15162 3168 15394 3224
rect 15101 3166 15394 3168
rect 15469 3226 15535 3229
rect 15653 3226 15719 3229
rect 15469 3224 15719 3226
rect 15469 3168 15474 3224
rect 15530 3168 15658 3224
rect 15714 3168 15719 3224
rect 15469 3166 15719 3168
rect 15101 3163 15167 3166
rect 15469 3163 15535 3166
rect 15653 3163 15719 3166
rect 16481 3224 16547 3229
rect 16481 3168 16486 3224
rect 16542 3168 16547 3224
rect 16481 3163 16547 3168
rect 16665 3226 16731 3229
rect 18873 3226 18939 3229
rect 16665 3224 18939 3226
rect 16665 3168 16670 3224
rect 16726 3168 18878 3224
rect 18934 3168 18939 3224
rect 16665 3166 18939 3168
rect 16665 3163 16731 3166
rect 18873 3163 18939 3166
rect 11881 3090 11947 3093
rect 11654 3088 11947 3090
rect 11654 3032 11886 3088
rect 11942 3032 11947 3088
rect 11654 3030 11947 3032
rect 11881 3027 11947 3030
rect 12065 3090 12131 3093
rect 16297 3090 16363 3093
rect 12065 3088 16363 3090
rect 12065 3032 12070 3088
rect 12126 3032 16302 3088
rect 16358 3032 16363 3088
rect 12065 3030 16363 3032
rect 16484 3090 16544 3163
rect 16484 3030 21696 3090
rect 12065 3027 12131 3030
rect 16297 3027 16363 3030
rect 9305 2952 10058 2954
rect 9305 2896 9310 2952
rect 9366 2896 10058 2952
rect 9305 2894 10058 2896
rect 10409 2954 10475 2957
rect 11053 2954 11119 2957
rect 10409 2952 11119 2954
rect 10409 2896 10414 2952
rect 10470 2896 11058 2952
rect 11114 2896 11119 2952
rect 10409 2894 11119 2896
rect 9305 2891 9371 2894
rect 10409 2891 10475 2894
rect 11053 2891 11119 2894
rect 11697 2954 11763 2957
rect 12801 2954 12867 2957
rect 16573 2954 16639 2957
rect 19609 2954 19675 2957
rect 11697 2952 16639 2954
rect 11697 2896 11702 2952
rect 11758 2896 12806 2952
rect 12862 2896 16578 2952
rect 16634 2896 16639 2952
rect 11697 2894 16639 2896
rect 11697 2891 11763 2894
rect 12801 2891 12867 2894
rect 16573 2891 16639 2894
rect 17726 2952 19675 2954
rect 17726 2896 19614 2952
rect 19670 2896 19675 2952
rect 17726 2894 19675 2896
rect 9990 2756 9996 2820
rect 10060 2818 10066 2820
rect 10409 2818 10475 2821
rect 10060 2816 10475 2818
rect 10060 2760 10414 2816
rect 10470 2760 10475 2816
rect 10060 2758 10475 2760
rect 10060 2756 10066 2758
rect 10409 2755 10475 2758
rect 10685 2816 10751 2821
rect 10685 2760 10690 2816
rect 10746 2760 10751 2816
rect 10685 2755 10751 2760
rect 11145 2818 11211 2821
rect 12249 2820 12315 2821
rect 12014 2818 12020 2820
rect 11145 2816 12020 2818
rect 11145 2760 11150 2816
rect 11206 2760 12020 2816
rect 11145 2758 12020 2760
rect 11145 2755 11211 2758
rect 12014 2756 12020 2758
rect 12084 2756 12090 2820
rect 12198 2756 12204 2820
rect 12268 2818 12315 2820
rect 12433 2818 12499 2821
rect 13118 2818 13124 2820
rect 12268 2816 12360 2818
rect 12310 2760 12360 2816
rect 12268 2758 12360 2760
rect 12433 2816 13124 2818
rect 12433 2760 12438 2816
rect 12494 2760 13124 2816
rect 12433 2758 13124 2760
rect 12268 2756 12315 2758
rect 12249 2755 12315 2756
rect 12433 2755 12499 2758
rect 13118 2756 13124 2758
rect 13188 2756 13194 2820
rect 13721 2818 13787 2821
rect 14222 2818 14228 2820
rect 13721 2816 14228 2818
rect 13721 2760 13726 2816
rect 13782 2760 14228 2816
rect 13721 2758 14228 2760
rect 13721 2755 13787 2758
rect 14222 2756 14228 2758
rect 14292 2756 14298 2820
rect 14365 2818 14431 2821
rect 15377 2818 15443 2821
rect 17726 2818 17786 2894
rect 19609 2891 19675 2894
rect 14365 2816 15443 2818
rect 14365 2760 14370 2816
rect 14426 2760 15382 2816
rect 15438 2760 15443 2816
rect 14365 2758 15443 2760
rect 14365 2755 14431 2758
rect 15377 2755 15443 2758
rect 16070 2758 17786 2818
rect 8363 2752 8679 2753
rect 8363 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8679 2752
rect 8363 2687 8679 2688
rect 4356 2680 4448 2682
rect 4398 2624 4448 2680
rect 4356 2622 4448 2624
rect 7281 2680 8218 2682
rect 7281 2624 7286 2680
rect 7342 2624 8218 2680
rect 7281 2622 8218 2624
rect 4356 2620 4403 2622
rect 4337 2619 4403 2620
rect 7281 2619 7347 2622
rect 1710 2484 1716 2548
rect 1780 2546 1786 2548
rect 3785 2546 3851 2549
rect 10133 2546 10199 2549
rect 1780 2544 3851 2546
rect 1780 2488 3790 2544
rect 3846 2488 3851 2544
rect 1780 2486 3851 2488
rect 1780 2484 1786 2486
rect 3785 2483 3851 2486
rect 3926 2544 10199 2546
rect 3926 2488 10138 2544
rect 10194 2488 10199 2544
rect 3926 2486 10199 2488
rect 10688 2546 10748 2755
rect 13308 2752 13624 2753
rect 13308 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13624 2752
rect 13308 2687 13624 2688
rect 10869 2682 10935 2685
rect 13813 2684 13879 2685
rect 12750 2682 12756 2684
rect 10869 2680 12756 2682
rect 10869 2624 10874 2680
rect 10930 2624 12756 2680
rect 10869 2622 12756 2624
rect 10869 2619 10935 2622
rect 12750 2620 12756 2622
rect 12820 2620 12826 2684
rect 13813 2682 13860 2684
rect 13768 2680 13860 2682
rect 13768 2624 13818 2680
rect 13768 2622 13860 2624
rect 13813 2620 13860 2622
rect 13924 2620 13930 2684
rect 13997 2682 14063 2685
rect 16070 2682 16130 2758
rect 18638 2756 18644 2820
rect 18708 2818 18714 2820
rect 18873 2818 18939 2821
rect 19609 2820 19675 2821
rect 19558 2818 19564 2820
rect 18708 2816 18939 2818
rect 18708 2760 18878 2816
rect 18934 2760 18939 2816
rect 18708 2758 18939 2760
rect 19518 2758 19564 2818
rect 19628 2816 19675 2820
rect 19670 2760 19675 2816
rect 18708 2756 18714 2758
rect 18873 2755 18939 2758
rect 19558 2756 19564 2758
rect 19628 2756 19675 2760
rect 21636 2818 21696 3030
rect 21840 2818 22300 2848
rect 21636 2758 22300 2818
rect 19609 2755 19675 2756
rect 18253 2752 18569 2753
rect 18253 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18569 2752
rect 21840 2728 22300 2758
rect 18253 2687 18569 2688
rect 13997 2680 16130 2682
rect 13997 2624 14002 2680
rect 14058 2624 16130 2680
rect 13997 2622 16130 2624
rect 13813 2619 13879 2620
rect 13997 2619 14063 2622
rect 11789 2546 11855 2549
rect 12566 2546 12572 2548
rect 10688 2486 11346 2546
rect 790 2348 796 2412
rect 860 2410 866 2412
rect 3926 2410 3986 2486
rect 10133 2483 10199 2486
rect 860 2350 3986 2410
rect 4153 2410 4219 2413
rect 4470 2410 4476 2412
rect 4153 2408 4476 2410
rect 4153 2352 4158 2408
rect 4214 2352 4476 2408
rect 4153 2350 4476 2352
rect 860 2348 866 2350
rect 4153 2347 4219 2350
rect 4470 2348 4476 2350
rect 4540 2348 4546 2412
rect 4654 2348 4660 2412
rect 4724 2410 4730 2412
rect 5165 2410 5231 2413
rect 4724 2408 5231 2410
rect 4724 2352 5170 2408
rect 5226 2352 5231 2408
rect 4724 2350 5231 2352
rect 4724 2348 4730 2350
rect 5165 2347 5231 2350
rect 5574 2348 5580 2412
rect 5644 2410 5650 2412
rect 7005 2410 7071 2413
rect 7782 2410 7788 2412
rect 5644 2350 6378 2410
rect 5644 2348 5650 2350
rect 5890 2208 6206 2209
rect 5890 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6206 2208
rect 5890 2143 6206 2144
rect 6318 2138 6378 2350
rect 7005 2408 7788 2410
rect 7005 2352 7010 2408
rect 7066 2352 7788 2408
rect 7005 2350 7788 2352
rect 7005 2347 7071 2350
rect 7782 2348 7788 2350
rect 7852 2348 7858 2412
rect 9029 2410 9095 2413
rect 11145 2410 11211 2413
rect 9029 2408 11211 2410
rect 9029 2352 9034 2408
rect 9090 2352 11150 2408
rect 11206 2352 11211 2408
rect 9029 2350 11211 2352
rect 9029 2347 9095 2350
rect 11145 2347 11211 2350
rect 7465 2276 7531 2277
rect 7414 2212 7420 2276
rect 7484 2274 7531 2276
rect 9121 2274 9187 2277
rect 10358 2274 10364 2276
rect 7484 2272 7576 2274
rect 7526 2216 7576 2272
rect 7484 2214 7576 2216
rect 9078 2272 9187 2274
rect 9078 2216 9126 2272
rect 9182 2216 9187 2272
rect 7484 2212 7531 2214
rect 7465 2211 7531 2212
rect 9078 2211 9187 2216
rect 9262 2214 10364 2274
rect 9078 2138 9138 2211
rect 6318 2078 9138 2138
rect 841 2002 907 2005
rect 6085 2002 6151 2005
rect 841 2000 6151 2002
rect 841 1944 846 2000
rect 902 1944 6090 2000
rect 6146 1944 6151 2000
rect 841 1942 6151 1944
rect 841 1939 907 1942
rect 6085 1939 6151 1942
rect 6637 2002 6703 2005
rect 7230 2002 7236 2004
rect 6637 2000 7236 2002
rect 6637 1944 6642 2000
rect 6698 1944 7236 2000
rect 6637 1942 7236 1944
rect 6637 1939 6703 1942
rect 7230 1940 7236 1942
rect 7300 1940 7306 2004
rect 8477 2002 8543 2005
rect 9262 2002 9322 2214
rect 10358 2212 10364 2214
rect 10428 2212 10434 2276
rect 10835 2208 11151 2209
rect 10835 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11151 2208
rect 10835 2143 11151 2144
rect 11286 2138 11346 2486
rect 11789 2544 12572 2546
rect 11789 2488 11794 2544
rect 11850 2488 12572 2544
rect 11789 2486 12572 2488
rect 11789 2483 11855 2486
rect 12566 2484 12572 2486
rect 12636 2484 12642 2548
rect 12709 2546 12775 2549
rect 13721 2546 13787 2549
rect 12709 2544 13787 2546
rect 12709 2488 12714 2544
rect 12770 2488 13726 2544
rect 13782 2488 13787 2544
rect 12709 2486 13787 2488
rect 12709 2483 12775 2486
rect 13721 2483 13787 2486
rect 13997 2546 14063 2549
rect 16481 2546 16547 2549
rect 13997 2544 16547 2546
rect 13997 2488 14002 2544
rect 14058 2488 16486 2544
rect 16542 2488 16547 2544
rect 13997 2486 16547 2488
rect 13997 2483 14063 2486
rect 16481 2483 16547 2486
rect 12433 2410 12499 2413
rect 12750 2410 12756 2412
rect 12433 2408 12756 2410
rect 12433 2352 12438 2408
rect 12494 2352 12756 2408
rect 12433 2350 12756 2352
rect 12433 2347 12499 2350
rect 12750 2348 12756 2350
rect 12820 2348 12826 2412
rect 12985 2410 13051 2413
rect 16481 2410 16547 2413
rect 12985 2408 16547 2410
rect 12985 2352 12990 2408
rect 13046 2352 16486 2408
rect 16542 2352 16547 2408
rect 12985 2350 16547 2352
rect 12985 2347 13051 2350
rect 16481 2347 16547 2350
rect 16757 2410 16823 2413
rect 16982 2410 16988 2412
rect 16757 2408 16988 2410
rect 16757 2352 16762 2408
rect 16818 2352 16988 2408
rect 16757 2350 16988 2352
rect 16757 2347 16823 2350
rect 16982 2348 16988 2350
rect 17052 2348 17058 2412
rect 17953 2410 18019 2413
rect 19006 2410 19012 2412
rect 17953 2408 19012 2410
rect 17953 2352 17958 2408
rect 18014 2352 19012 2408
rect 17953 2350 19012 2352
rect 17953 2347 18019 2350
rect 19006 2348 19012 2350
rect 19076 2348 19082 2412
rect 11421 2274 11487 2277
rect 12801 2274 12867 2277
rect 12934 2274 12940 2276
rect 11421 2272 12940 2274
rect 11421 2216 11426 2272
rect 11482 2216 12806 2272
rect 12862 2216 12940 2272
rect 11421 2214 12940 2216
rect 11421 2211 11487 2214
rect 12801 2211 12867 2214
rect 12934 2212 12940 2214
rect 13004 2212 13010 2276
rect 13353 2274 13419 2277
rect 15326 2274 15332 2276
rect 13353 2272 15332 2274
rect 13353 2216 13358 2272
rect 13414 2216 15332 2272
rect 13353 2214 15332 2216
rect 13353 2211 13419 2214
rect 15326 2212 15332 2214
rect 15396 2212 15402 2276
rect 16205 2274 16271 2277
rect 16941 2274 17007 2277
rect 21840 2274 22300 2304
rect 16205 2272 17007 2274
rect 16205 2216 16210 2272
rect 16266 2216 16946 2272
rect 17002 2216 17007 2272
rect 16205 2214 17007 2216
rect 16205 2211 16271 2214
rect 16941 2211 17007 2214
rect 21222 2214 22300 2274
rect 15780 2208 16096 2209
rect 15780 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16096 2208
rect 15780 2143 16096 2144
rect 20725 2208 21041 2209
rect 20725 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21041 2208
rect 20725 2143 21041 2144
rect 12617 2138 12683 2141
rect 11286 2136 12683 2138
rect 11286 2080 12622 2136
rect 12678 2080 12683 2136
rect 11286 2078 12683 2080
rect 12617 2075 12683 2078
rect 12893 2138 12959 2141
rect 12893 2136 15716 2138
rect 12893 2080 12898 2136
rect 12954 2080 15716 2136
rect 12893 2078 15716 2080
rect 12893 2075 12959 2078
rect 8477 2000 9322 2002
rect 8477 1944 8482 2000
rect 8538 1944 9322 2000
rect 8477 1942 9322 1944
rect 8477 1939 8543 1942
rect 11830 1940 11836 2004
rect 11900 2002 11906 2004
rect 14549 2002 14615 2005
rect 11900 2000 14615 2002
rect 11900 1944 14554 2000
rect 14610 1944 14615 2000
rect 11900 1942 14615 1944
rect 11900 1940 11906 1942
rect 14549 1939 14615 1942
rect 14774 1940 14780 2004
rect 14844 2002 14850 2004
rect 14917 2002 14983 2005
rect 14844 2000 14983 2002
rect 14844 1944 14922 2000
rect 14978 1944 14983 2000
rect 14844 1942 14983 1944
rect 15656 2002 15716 2078
rect 16246 2076 16252 2140
rect 16316 2138 16322 2140
rect 17769 2138 17835 2141
rect 16316 2136 17835 2138
rect 16316 2080 17774 2136
rect 17830 2080 17835 2136
rect 16316 2078 17835 2080
rect 16316 2076 16322 2078
rect 17769 2075 17835 2078
rect 19742 2002 19748 2004
rect 15656 1942 19748 2002
rect 14844 1940 14850 1942
rect 14917 1939 14983 1942
rect 19742 1940 19748 1942
rect 19812 1940 19818 2004
rect 974 1804 980 1868
rect 1044 1866 1050 1868
rect 6821 1866 6887 1869
rect 1044 1864 6887 1866
rect 1044 1808 6826 1864
rect 6882 1808 6887 1864
rect 1044 1806 6887 1808
rect 1044 1804 1050 1806
rect 6821 1803 6887 1806
rect 7966 1804 7972 1868
rect 8036 1866 8042 1868
rect 9305 1866 9371 1869
rect 11789 1866 11855 1869
rect 8036 1806 8954 1866
rect 8036 1804 8042 1806
rect 6862 1668 6868 1732
rect 6932 1730 6938 1732
rect 8201 1730 8267 1733
rect 6932 1728 8267 1730
rect 6932 1672 8206 1728
rect 8262 1672 8267 1728
rect 6932 1670 8267 1672
rect 6932 1668 6938 1670
rect 8201 1667 8267 1670
rect 3418 1664 3734 1665
rect 3418 1600 3424 1664
rect 3488 1600 3504 1664
rect 3568 1600 3584 1664
rect 3648 1600 3664 1664
rect 3728 1600 3734 1664
rect 3418 1599 3734 1600
rect 8363 1664 8679 1665
rect 8363 1600 8369 1664
rect 8433 1600 8449 1664
rect 8513 1600 8529 1664
rect 8593 1600 8609 1664
rect 8673 1600 8679 1664
rect 8363 1599 8679 1600
rect 8109 1594 8175 1597
rect 4110 1592 8175 1594
rect 4110 1536 8114 1592
rect 8170 1536 8175 1592
rect 4110 1534 8175 1536
rect 8894 1594 8954 1806
rect 9305 1864 11855 1866
rect 9305 1808 9310 1864
rect 9366 1808 11794 1864
rect 11850 1808 11855 1864
rect 9305 1806 11855 1808
rect 9305 1803 9371 1806
rect 11789 1803 11855 1806
rect 11973 1866 12039 1869
rect 12934 1866 12940 1868
rect 11973 1864 12940 1866
rect 11973 1808 11978 1864
rect 12034 1808 12940 1864
rect 11973 1806 12940 1808
rect 11973 1803 12039 1806
rect 12934 1804 12940 1806
rect 13004 1804 13010 1868
rect 21222 1866 21282 2214
rect 21840 2184 22300 2214
rect 13172 1806 21282 1866
rect 9622 1668 9628 1732
rect 9692 1730 9698 1732
rect 12617 1730 12683 1733
rect 9692 1728 12683 1730
rect 9692 1672 12622 1728
rect 12678 1672 12683 1728
rect 9692 1670 12683 1672
rect 9692 1668 9698 1670
rect 12617 1667 12683 1670
rect 12801 1730 12867 1733
rect 13172 1730 13232 1806
rect 14038 1730 14044 1732
rect 12801 1728 13232 1730
rect 12801 1672 12806 1728
rect 12862 1672 13232 1728
rect 12801 1670 13232 1672
rect 13724 1670 14044 1730
rect 12801 1667 12867 1670
rect 13308 1664 13624 1665
rect 13308 1600 13314 1664
rect 13378 1600 13394 1664
rect 13458 1600 13474 1664
rect 13538 1600 13554 1664
rect 13618 1600 13624 1664
rect 13308 1599 13624 1600
rect 10869 1594 10935 1597
rect 8894 1592 10935 1594
rect 8894 1536 10874 1592
rect 10930 1536 10935 1592
rect 8894 1534 10935 1536
rect 1342 1396 1348 1460
rect 1412 1458 1418 1460
rect 4110 1458 4170 1534
rect 8109 1531 8175 1534
rect 10869 1531 10935 1534
rect 11010 1534 12404 1594
rect 9305 1460 9371 1461
rect 1412 1398 4170 1458
rect 1412 1396 1418 1398
rect 6494 1396 6500 1460
rect 6564 1458 6570 1460
rect 9254 1458 9260 1460
rect 6564 1398 8402 1458
rect 9214 1398 9260 1458
rect 9324 1456 9371 1460
rect 9366 1400 9371 1456
rect 6564 1396 6570 1398
rect 5533 1322 5599 1325
rect 8109 1322 8175 1325
rect 5533 1320 8175 1322
rect 5533 1264 5538 1320
rect 5594 1264 8114 1320
rect 8170 1264 8175 1320
rect 5533 1262 8175 1264
rect 8342 1322 8402 1398
rect 9254 1396 9260 1398
rect 9324 1396 9371 1400
rect 9305 1395 9371 1396
rect 11010 1322 11070 1534
rect 11789 1410 11855 1413
rect 11789 1408 11898 1410
rect 11789 1352 11794 1408
rect 11850 1352 11898 1408
rect 12198 1396 12204 1460
rect 12268 1396 12274 1460
rect 12344 1458 12404 1534
rect 13724 1458 13784 1670
rect 14038 1668 14044 1670
rect 14108 1668 14114 1732
rect 14958 1668 14964 1732
rect 15028 1730 15034 1732
rect 17309 1730 17375 1733
rect 21840 1730 22300 1760
rect 15028 1728 17375 1730
rect 15028 1672 17314 1728
rect 17370 1672 17375 1728
rect 15028 1670 17375 1672
rect 15028 1668 15034 1670
rect 17309 1667 17375 1670
rect 19290 1670 22300 1730
rect 18253 1664 18569 1665
rect 18253 1600 18259 1664
rect 18323 1600 18339 1664
rect 18403 1600 18419 1664
rect 18483 1600 18499 1664
rect 18563 1600 18569 1664
rect 18253 1599 18569 1600
rect 14181 1594 14247 1597
rect 12344 1398 13784 1458
rect 13908 1592 14247 1594
rect 13908 1536 14186 1592
rect 14242 1536 14247 1592
rect 13908 1534 14247 1536
rect 11789 1347 11898 1352
rect 8342 1262 11070 1322
rect 5533 1259 5599 1262
rect 8109 1259 8175 1262
rect 2262 1124 2268 1188
rect 2332 1186 2338 1188
rect 5349 1186 5415 1189
rect 2332 1184 5415 1186
rect 2332 1128 5354 1184
rect 5410 1128 5415 1184
rect 2332 1126 5415 1128
rect 2332 1124 2338 1126
rect 5349 1123 5415 1126
rect 7598 1124 7604 1188
rect 7668 1186 7674 1188
rect 8201 1186 8267 1189
rect 10041 1186 10107 1189
rect 10225 1186 10291 1189
rect 7668 1184 8267 1186
rect 7668 1128 8206 1184
rect 8262 1128 8267 1184
rect 7668 1126 8267 1128
rect 7668 1124 7674 1126
rect 8201 1123 8267 1126
rect 9998 1184 10107 1186
rect 9998 1128 10046 1184
rect 10102 1128 10107 1184
rect 9998 1123 10107 1128
rect 10182 1184 10291 1186
rect 10182 1128 10230 1184
rect 10286 1128 10291 1184
rect 10182 1123 10291 1128
rect 11838 1186 11898 1347
rect 12206 1322 12266 1396
rect 13353 1322 13419 1325
rect 12206 1320 13419 1322
rect 12206 1264 13358 1320
rect 13414 1264 13419 1320
rect 12206 1262 13419 1264
rect 13353 1259 13419 1262
rect 13537 1322 13603 1325
rect 13908 1322 13968 1534
rect 14181 1531 14247 1534
rect 14406 1532 14412 1596
rect 14476 1594 14482 1596
rect 16941 1594 17007 1597
rect 14476 1592 17007 1594
rect 14476 1536 16946 1592
rect 17002 1536 17007 1592
rect 14476 1534 17007 1536
rect 14476 1532 14482 1534
rect 16941 1531 17007 1534
rect 15929 1458 15995 1461
rect 19290 1458 19350 1670
rect 21840 1640 22300 1670
rect 13537 1320 13968 1322
rect 13537 1264 13542 1320
rect 13598 1264 13968 1320
rect 13537 1262 13968 1264
rect 14046 1456 15995 1458
rect 14046 1400 15934 1456
rect 15990 1400 15995 1456
rect 14046 1398 15995 1400
rect 13537 1259 13603 1262
rect 12525 1186 12591 1189
rect 11838 1184 12591 1186
rect 11838 1128 12530 1184
rect 12586 1128 12591 1184
rect 11838 1126 12591 1128
rect 12525 1123 12591 1126
rect 12750 1124 12756 1188
rect 12820 1186 12826 1188
rect 14046 1186 14106 1398
rect 15929 1395 15995 1398
rect 16116 1398 19350 1458
rect 14222 1260 14228 1324
rect 14292 1260 14298 1324
rect 14733 1322 14799 1325
rect 16116 1322 16176 1398
rect 14733 1320 16176 1322
rect 14733 1264 14738 1320
rect 14794 1264 16176 1320
rect 14733 1262 16176 1264
rect 16297 1322 16363 1325
rect 16430 1322 16436 1324
rect 16297 1320 16436 1322
rect 16297 1264 16302 1320
rect 16358 1264 16436 1320
rect 16297 1262 16436 1264
rect 12820 1126 14106 1186
rect 14230 1186 14290 1260
rect 14733 1259 14799 1262
rect 16297 1259 16363 1262
rect 16430 1260 16436 1262
rect 16500 1260 16506 1324
rect 18045 1322 18111 1325
rect 20110 1322 20116 1324
rect 18045 1320 20116 1322
rect 18045 1264 18050 1320
rect 18106 1264 20116 1320
rect 18045 1262 20116 1264
rect 18045 1259 18111 1262
rect 20110 1260 20116 1262
rect 20180 1260 20186 1324
rect 15326 1186 15332 1188
rect 14230 1126 15332 1186
rect 12820 1124 12826 1126
rect 15326 1124 15332 1126
rect 15396 1124 15402 1188
rect 16297 1186 16363 1189
rect 17902 1186 17908 1188
rect 16297 1184 17908 1186
rect 16297 1128 16302 1184
rect 16358 1128 17908 1184
rect 16297 1126 17908 1128
rect 16297 1123 16363 1126
rect 17902 1124 17908 1126
rect 17972 1124 17978 1188
rect 21173 1186 21239 1189
rect 21840 1186 22300 1216
rect 21173 1184 22300 1186
rect 21173 1128 21178 1184
rect 21234 1128 22300 1184
rect 21173 1126 22300 1128
rect 21173 1123 21239 1126
rect 5890 1120 6206 1121
rect 5890 1056 5896 1120
rect 5960 1056 5976 1120
rect 6040 1056 6056 1120
rect 6120 1056 6136 1120
rect 6200 1056 6206 1120
rect 5890 1055 6206 1056
rect 9998 1053 10058 1123
rect 10182 1053 10242 1123
rect 10835 1120 11151 1121
rect 10835 1056 10841 1120
rect 10905 1056 10921 1120
rect 10985 1056 11001 1120
rect 11065 1056 11081 1120
rect 11145 1056 11151 1120
rect 10835 1055 11151 1056
rect 15780 1120 16096 1121
rect 15780 1056 15786 1120
rect 15850 1056 15866 1120
rect 15930 1056 15946 1120
rect 16010 1056 16026 1120
rect 16090 1056 16096 1120
rect 15780 1055 16096 1056
rect 20725 1120 21041 1121
rect 20725 1056 20731 1120
rect 20795 1056 20811 1120
rect 20875 1056 20891 1120
rect 20955 1056 20971 1120
rect 21035 1056 21041 1120
rect 21840 1096 22300 1126
rect 20725 1055 21041 1056
rect 9998 1048 10107 1053
rect 9998 992 10046 1048
rect 10102 992 10107 1048
rect 9998 990 10107 992
rect 10182 1048 10291 1053
rect 10182 992 10230 1048
rect 10286 992 10291 1048
rect 10182 990 10291 992
rect 10041 987 10107 990
rect 10225 987 10291 990
rect 12065 1050 12131 1053
rect 15510 1050 15516 1052
rect 12065 1048 15516 1050
rect 12065 992 12070 1048
rect 12126 992 15516 1048
rect 12065 990 15516 992
rect 12065 987 12131 990
rect 15510 988 15516 990
rect 15580 988 15586 1052
rect 16205 1050 16271 1053
rect 18965 1050 19031 1053
rect 16205 1048 19031 1050
rect 16205 992 16210 1048
rect 16266 992 18970 1048
rect 19026 992 19031 1048
rect 16205 990 19031 992
rect 16205 987 16271 990
rect 18965 987 19031 990
rect 9806 852 9812 916
rect 9876 914 9882 916
rect 10041 914 10107 917
rect 9876 912 10107 914
rect 9876 856 10046 912
rect 10102 856 10107 912
rect 9876 854 10107 856
rect 9876 852 9882 854
rect 10041 851 10107 854
rect 10174 852 10180 916
rect 10244 914 10250 916
rect 11145 914 11211 917
rect 10244 912 11211 914
rect 10244 856 11150 912
rect 11206 856 11211 912
rect 10244 854 11211 856
rect 10244 852 10250 854
rect 11145 851 11211 854
rect 11278 852 11284 916
rect 11348 914 11354 916
rect 18413 914 18479 917
rect 11348 912 18479 914
rect 11348 856 18418 912
rect 18474 856 18479 912
rect 11348 854 18479 856
rect 11348 852 11354 854
rect 18413 851 18479 854
rect 381 778 447 781
rect 7557 778 7623 781
rect 381 776 7623 778
rect 381 720 386 776
rect 442 720 7562 776
rect 7618 720 7623 776
rect 381 718 7623 720
rect 381 715 447 718
rect 7557 715 7623 718
rect 9990 716 9996 780
rect 10060 778 10066 780
rect 10225 778 10291 781
rect 10060 776 10291 778
rect 10060 720 10230 776
rect 10286 720 10291 776
rect 10060 718 10291 720
rect 10060 716 10066 718
rect 10225 715 10291 718
rect 10542 716 10548 780
rect 10612 778 10618 780
rect 11513 778 11579 781
rect 10612 776 11579 778
rect 10612 720 11518 776
rect 11574 720 11579 776
rect 10612 718 11579 720
rect 10612 716 10618 718
rect 11513 715 11579 718
rect 12014 716 12020 780
rect 12084 778 12090 780
rect 13353 778 13419 781
rect 12084 776 13419 778
rect 12084 720 13358 776
rect 13414 720 13419 776
rect 12084 718 13419 720
rect 12084 716 12090 718
rect 13353 715 13419 718
rect 13537 778 13603 781
rect 16757 778 16823 781
rect 19057 778 19123 781
rect 13537 776 16823 778
rect 13537 720 13542 776
rect 13598 720 16762 776
rect 16818 720 16823 776
rect 13537 718 16823 720
rect 13537 715 13603 718
rect 16757 715 16823 718
rect 16944 776 19123 778
rect 16944 720 19062 776
rect 19118 720 19123 776
rect 16944 718 19123 720
rect 3877 642 3943 645
rect 12893 642 12959 645
rect 3877 640 12959 642
rect 3877 584 3882 640
rect 3938 584 12898 640
rect 12954 584 12959 640
rect 3877 582 12959 584
rect 3877 579 3943 582
rect 12893 579 12959 582
rect 13261 642 13327 645
rect 15694 642 15700 644
rect 13261 640 15700 642
rect 13261 584 13266 640
rect 13322 584 15700 640
rect 13261 582 15700 584
rect 13261 579 13327 582
rect 15694 580 15700 582
rect 15764 580 15770 644
rect 16944 642 17004 718
rect 19057 715 19123 718
rect 15840 582 17004 642
rect 17585 642 17651 645
rect 21840 642 22300 672
rect 17585 640 22300 642
rect 17585 584 17590 640
rect 17646 584 22300 640
rect 17585 582 22300 584
rect 12566 444 12572 508
rect 12636 506 12642 508
rect 12636 446 14336 506
rect 12636 444 12642 446
rect 11646 308 11652 372
rect 11716 370 11722 372
rect 14084 370 14090 372
rect 11716 310 14090 370
rect 11716 308 11722 310
rect 14084 308 14090 310
rect 14154 308 14160 372
rect 14276 370 14336 446
rect 14406 444 14412 508
rect 14476 506 14482 508
rect 15840 506 15900 582
rect 17585 579 17651 582
rect 21840 552 22300 582
rect 14476 446 15900 506
rect 14476 444 14482 446
rect 16062 444 16068 508
rect 16132 506 16138 508
rect 18137 506 18203 509
rect 16132 504 18203 506
rect 16132 448 18142 504
rect 18198 448 18203 504
rect 16132 446 18203 448
rect 16132 444 16138 446
rect 18137 443 18203 446
rect 14641 370 14707 373
rect 14276 368 14707 370
rect 14276 312 14646 368
rect 14702 312 14707 368
rect 14276 310 14707 312
rect 14641 307 14707 310
rect 14774 308 14780 372
rect 14844 370 14850 372
rect 15285 370 15351 373
rect 14844 368 15351 370
rect 14844 312 15290 368
rect 15346 312 15351 368
rect 14844 310 15351 312
rect 14844 308 14850 310
rect 15285 307 15351 310
rect 15745 370 15811 373
rect 18781 370 18847 373
rect 15745 368 18847 370
rect 15745 312 15750 368
rect 15806 312 18786 368
rect 18842 312 18847 368
rect 15745 310 18847 312
rect 15745 307 15811 310
rect 18781 307 18847 310
rect 12382 172 12388 236
rect 12452 234 12458 236
rect 18505 234 18571 237
rect 12452 232 18571 234
rect 12452 176 18510 232
rect 18566 176 18571 232
rect 12452 174 18571 176
rect 12452 172 12458 174
rect 18505 171 18571 174
rect 6678 36 6684 100
rect 6748 98 6754 100
rect 7465 98 7531 101
rect 6748 96 7531 98
rect 6748 40 7470 96
rect 7526 40 7531 96
rect 6748 38 7531 40
rect 6748 36 6754 38
rect 7465 35 7531 38
rect 8150 36 8156 100
rect 8220 98 8226 100
rect 8569 98 8635 101
rect 8220 96 8635 98
rect 8220 40 8574 96
rect 8630 40 8635 96
rect 8220 38 8635 40
rect 8220 36 8226 38
rect 8569 35 8635 38
rect 12934 36 12940 100
rect 13004 98 13010 100
rect 17951 98 18017 101
rect 13004 96 18017 98
rect 13004 40 17956 96
rect 18012 40 18017 96
rect 13004 38 18017 40
rect 13004 36 13010 38
rect 17951 35 18017 38
<< via3 >>
rect 14596 44508 14660 44572
rect 16620 43692 16684 43756
rect 5896 43548 5960 43552
rect 5896 43492 5900 43548
rect 5900 43492 5956 43548
rect 5956 43492 5960 43548
rect 5896 43488 5960 43492
rect 5976 43548 6040 43552
rect 5976 43492 5980 43548
rect 5980 43492 6036 43548
rect 6036 43492 6040 43548
rect 5976 43488 6040 43492
rect 6056 43548 6120 43552
rect 6056 43492 6060 43548
rect 6060 43492 6116 43548
rect 6116 43492 6120 43548
rect 6056 43488 6120 43492
rect 6136 43548 6200 43552
rect 6136 43492 6140 43548
rect 6140 43492 6196 43548
rect 6196 43492 6200 43548
rect 6136 43488 6200 43492
rect 10841 43548 10905 43552
rect 10841 43492 10845 43548
rect 10845 43492 10901 43548
rect 10901 43492 10905 43548
rect 10841 43488 10905 43492
rect 10921 43548 10985 43552
rect 10921 43492 10925 43548
rect 10925 43492 10981 43548
rect 10981 43492 10985 43548
rect 10921 43488 10985 43492
rect 11001 43548 11065 43552
rect 11001 43492 11005 43548
rect 11005 43492 11061 43548
rect 11061 43492 11065 43548
rect 11001 43488 11065 43492
rect 11081 43548 11145 43552
rect 11081 43492 11085 43548
rect 11085 43492 11141 43548
rect 11141 43492 11145 43548
rect 11081 43488 11145 43492
rect 15786 43548 15850 43552
rect 15786 43492 15790 43548
rect 15790 43492 15846 43548
rect 15846 43492 15850 43548
rect 15786 43488 15850 43492
rect 15866 43548 15930 43552
rect 15866 43492 15870 43548
rect 15870 43492 15926 43548
rect 15926 43492 15930 43548
rect 15866 43488 15930 43492
rect 15946 43548 16010 43552
rect 15946 43492 15950 43548
rect 15950 43492 16006 43548
rect 16006 43492 16010 43548
rect 15946 43488 16010 43492
rect 16026 43548 16090 43552
rect 16026 43492 16030 43548
rect 16030 43492 16086 43548
rect 16086 43492 16090 43548
rect 16026 43488 16090 43492
rect 20731 43548 20795 43552
rect 20731 43492 20735 43548
rect 20735 43492 20791 43548
rect 20791 43492 20795 43548
rect 20731 43488 20795 43492
rect 20811 43548 20875 43552
rect 20811 43492 20815 43548
rect 20815 43492 20871 43548
rect 20871 43492 20875 43548
rect 20811 43488 20875 43492
rect 20891 43548 20955 43552
rect 20891 43492 20895 43548
rect 20895 43492 20951 43548
rect 20951 43492 20955 43548
rect 20891 43488 20955 43492
rect 20971 43548 21035 43552
rect 20971 43492 20975 43548
rect 20975 43492 21031 43548
rect 21031 43492 21035 43548
rect 20971 43488 21035 43492
rect 5028 43148 5092 43212
rect 16252 43148 16316 43212
rect 5580 43012 5644 43076
rect 3424 43004 3488 43008
rect 3424 42948 3428 43004
rect 3428 42948 3484 43004
rect 3484 42948 3488 43004
rect 3424 42944 3488 42948
rect 3504 43004 3568 43008
rect 3504 42948 3508 43004
rect 3508 42948 3564 43004
rect 3564 42948 3568 43004
rect 3504 42944 3568 42948
rect 3584 43004 3648 43008
rect 3584 42948 3588 43004
rect 3588 42948 3644 43004
rect 3644 42948 3648 43004
rect 3584 42944 3648 42948
rect 3664 43004 3728 43008
rect 3664 42948 3668 43004
rect 3668 42948 3724 43004
rect 3724 42948 3728 43004
rect 3664 42944 3728 42948
rect 8369 43004 8433 43008
rect 8369 42948 8373 43004
rect 8373 42948 8429 43004
rect 8429 42948 8433 43004
rect 8369 42944 8433 42948
rect 8449 43004 8513 43008
rect 8449 42948 8453 43004
rect 8453 42948 8509 43004
rect 8509 42948 8513 43004
rect 8449 42944 8513 42948
rect 8529 43004 8593 43008
rect 8529 42948 8533 43004
rect 8533 42948 8589 43004
rect 8589 42948 8593 43004
rect 8529 42944 8593 42948
rect 8609 43004 8673 43008
rect 8609 42948 8613 43004
rect 8613 42948 8669 43004
rect 8669 42948 8673 43004
rect 8609 42944 8673 42948
rect 13314 43004 13378 43008
rect 13314 42948 13318 43004
rect 13318 42948 13374 43004
rect 13374 42948 13378 43004
rect 13314 42944 13378 42948
rect 13394 43004 13458 43008
rect 13394 42948 13398 43004
rect 13398 42948 13454 43004
rect 13454 42948 13458 43004
rect 13394 42944 13458 42948
rect 13474 43004 13538 43008
rect 13474 42948 13478 43004
rect 13478 42948 13534 43004
rect 13534 42948 13538 43004
rect 13474 42944 13538 42948
rect 13554 43004 13618 43008
rect 13554 42948 13558 43004
rect 13558 42948 13614 43004
rect 13614 42948 13618 43004
rect 13554 42944 13618 42948
rect 18259 43004 18323 43008
rect 18259 42948 18263 43004
rect 18263 42948 18319 43004
rect 18319 42948 18323 43004
rect 18259 42944 18323 42948
rect 18339 43004 18403 43008
rect 18339 42948 18343 43004
rect 18343 42948 18399 43004
rect 18399 42948 18403 43004
rect 18339 42944 18403 42948
rect 18419 43004 18483 43008
rect 18419 42948 18423 43004
rect 18423 42948 18479 43004
rect 18479 42948 18483 43004
rect 18419 42944 18483 42948
rect 18499 43004 18563 43008
rect 18499 42948 18503 43004
rect 18503 42948 18559 43004
rect 18559 42948 18563 43004
rect 18499 42944 18563 42948
rect 10548 42876 10612 42940
rect 15516 42604 15580 42668
rect 5896 42460 5960 42464
rect 5896 42404 5900 42460
rect 5900 42404 5956 42460
rect 5956 42404 5960 42460
rect 5896 42400 5960 42404
rect 5976 42460 6040 42464
rect 5976 42404 5980 42460
rect 5980 42404 6036 42460
rect 6036 42404 6040 42460
rect 5976 42400 6040 42404
rect 6056 42460 6120 42464
rect 6056 42404 6060 42460
rect 6060 42404 6116 42460
rect 6116 42404 6120 42460
rect 6056 42400 6120 42404
rect 6136 42460 6200 42464
rect 6136 42404 6140 42460
rect 6140 42404 6196 42460
rect 6196 42404 6200 42460
rect 6136 42400 6200 42404
rect 10841 42460 10905 42464
rect 10841 42404 10845 42460
rect 10845 42404 10901 42460
rect 10901 42404 10905 42460
rect 10841 42400 10905 42404
rect 10921 42460 10985 42464
rect 10921 42404 10925 42460
rect 10925 42404 10981 42460
rect 10981 42404 10985 42460
rect 10921 42400 10985 42404
rect 11001 42460 11065 42464
rect 11001 42404 11005 42460
rect 11005 42404 11061 42460
rect 11061 42404 11065 42460
rect 11001 42400 11065 42404
rect 11081 42460 11145 42464
rect 11081 42404 11085 42460
rect 11085 42404 11141 42460
rect 11141 42404 11145 42460
rect 11081 42400 11145 42404
rect 15786 42460 15850 42464
rect 15786 42404 15790 42460
rect 15790 42404 15846 42460
rect 15846 42404 15850 42460
rect 15786 42400 15850 42404
rect 15866 42460 15930 42464
rect 15866 42404 15870 42460
rect 15870 42404 15926 42460
rect 15926 42404 15930 42460
rect 15866 42400 15930 42404
rect 15946 42460 16010 42464
rect 15946 42404 15950 42460
rect 15950 42404 16006 42460
rect 16006 42404 16010 42460
rect 15946 42400 16010 42404
rect 16026 42460 16090 42464
rect 16026 42404 16030 42460
rect 16030 42404 16086 42460
rect 16086 42404 16090 42460
rect 16026 42400 16090 42404
rect 20731 42460 20795 42464
rect 20731 42404 20735 42460
rect 20735 42404 20791 42460
rect 20791 42404 20795 42460
rect 20731 42400 20795 42404
rect 20811 42460 20875 42464
rect 20811 42404 20815 42460
rect 20815 42404 20871 42460
rect 20871 42404 20875 42460
rect 20811 42400 20875 42404
rect 20891 42460 20955 42464
rect 20891 42404 20895 42460
rect 20895 42404 20951 42460
rect 20951 42404 20955 42460
rect 20891 42400 20955 42404
rect 20971 42460 21035 42464
rect 20971 42404 20975 42460
rect 20975 42404 21031 42460
rect 21031 42404 21035 42460
rect 20971 42400 21035 42404
rect 7420 42196 7484 42260
rect 5396 42060 5460 42124
rect 9444 42060 9508 42124
rect 12940 42060 13004 42124
rect 18092 42060 18156 42124
rect 3424 41916 3488 41920
rect 3424 41860 3428 41916
rect 3428 41860 3484 41916
rect 3484 41860 3488 41916
rect 3424 41856 3488 41860
rect 3504 41916 3568 41920
rect 3504 41860 3508 41916
rect 3508 41860 3564 41916
rect 3564 41860 3568 41916
rect 3504 41856 3568 41860
rect 3584 41916 3648 41920
rect 3584 41860 3588 41916
rect 3588 41860 3644 41916
rect 3644 41860 3648 41916
rect 3584 41856 3648 41860
rect 3664 41916 3728 41920
rect 3664 41860 3668 41916
rect 3668 41860 3724 41916
rect 3724 41860 3728 41916
rect 3664 41856 3728 41860
rect 8369 41916 8433 41920
rect 8369 41860 8373 41916
rect 8373 41860 8429 41916
rect 8429 41860 8433 41916
rect 8369 41856 8433 41860
rect 8449 41916 8513 41920
rect 8449 41860 8453 41916
rect 8453 41860 8509 41916
rect 8509 41860 8513 41916
rect 8449 41856 8513 41860
rect 8529 41916 8593 41920
rect 8529 41860 8533 41916
rect 8533 41860 8589 41916
rect 8589 41860 8593 41916
rect 8529 41856 8593 41860
rect 8609 41916 8673 41920
rect 8609 41860 8613 41916
rect 8613 41860 8669 41916
rect 8669 41860 8673 41916
rect 8609 41856 8673 41860
rect 13314 41916 13378 41920
rect 13314 41860 13318 41916
rect 13318 41860 13374 41916
rect 13374 41860 13378 41916
rect 13314 41856 13378 41860
rect 13394 41916 13458 41920
rect 13394 41860 13398 41916
rect 13398 41860 13454 41916
rect 13454 41860 13458 41916
rect 13394 41856 13458 41860
rect 13474 41916 13538 41920
rect 13474 41860 13478 41916
rect 13478 41860 13534 41916
rect 13534 41860 13538 41916
rect 13474 41856 13538 41860
rect 13554 41916 13618 41920
rect 13554 41860 13558 41916
rect 13558 41860 13614 41916
rect 13614 41860 13618 41916
rect 13554 41856 13618 41860
rect 18259 41916 18323 41920
rect 18259 41860 18263 41916
rect 18263 41860 18319 41916
rect 18319 41860 18323 41916
rect 18259 41856 18323 41860
rect 18339 41916 18403 41920
rect 18339 41860 18343 41916
rect 18343 41860 18399 41916
rect 18399 41860 18403 41916
rect 18339 41856 18403 41860
rect 18419 41916 18483 41920
rect 18419 41860 18423 41916
rect 18423 41860 18479 41916
rect 18479 41860 18483 41916
rect 18419 41856 18483 41860
rect 18499 41916 18563 41920
rect 18499 41860 18503 41916
rect 18503 41860 18559 41916
rect 18559 41860 18563 41916
rect 18499 41856 18563 41860
rect 15332 41788 15396 41852
rect 1164 41652 1228 41716
rect 6500 41652 6564 41716
rect 13124 41712 13188 41716
rect 13124 41656 13174 41712
rect 13174 41656 13188 41712
rect 13124 41652 13188 41656
rect 2084 41380 2148 41444
rect 3924 41516 3988 41580
rect 9260 41516 9324 41580
rect 11652 41516 11716 41580
rect 15516 41380 15580 41444
rect 5896 41372 5960 41376
rect 5896 41316 5900 41372
rect 5900 41316 5956 41372
rect 5956 41316 5960 41372
rect 5896 41312 5960 41316
rect 5976 41372 6040 41376
rect 5976 41316 5980 41372
rect 5980 41316 6036 41372
rect 6036 41316 6040 41372
rect 5976 41312 6040 41316
rect 6056 41372 6120 41376
rect 6056 41316 6060 41372
rect 6060 41316 6116 41372
rect 6116 41316 6120 41372
rect 6056 41312 6120 41316
rect 6136 41372 6200 41376
rect 6136 41316 6140 41372
rect 6140 41316 6196 41372
rect 6196 41316 6200 41372
rect 6136 41312 6200 41316
rect 10841 41372 10905 41376
rect 10841 41316 10845 41372
rect 10845 41316 10901 41372
rect 10901 41316 10905 41372
rect 10841 41312 10905 41316
rect 10921 41372 10985 41376
rect 10921 41316 10925 41372
rect 10925 41316 10981 41372
rect 10981 41316 10985 41372
rect 10921 41312 10985 41316
rect 11001 41372 11065 41376
rect 11001 41316 11005 41372
rect 11005 41316 11061 41372
rect 11061 41316 11065 41372
rect 11001 41312 11065 41316
rect 11081 41372 11145 41376
rect 11081 41316 11085 41372
rect 11085 41316 11141 41372
rect 11141 41316 11145 41372
rect 11081 41312 11145 41316
rect 15786 41372 15850 41376
rect 15786 41316 15790 41372
rect 15790 41316 15846 41372
rect 15846 41316 15850 41372
rect 15786 41312 15850 41316
rect 15866 41372 15930 41376
rect 15866 41316 15870 41372
rect 15870 41316 15926 41372
rect 15926 41316 15930 41372
rect 15866 41312 15930 41316
rect 15946 41372 16010 41376
rect 15946 41316 15950 41372
rect 15950 41316 16006 41372
rect 16006 41316 16010 41372
rect 15946 41312 16010 41316
rect 16026 41372 16090 41376
rect 16026 41316 16030 41372
rect 16030 41316 16086 41372
rect 16086 41316 16090 41372
rect 16026 41312 16090 41316
rect 20731 41372 20795 41376
rect 20731 41316 20735 41372
rect 20735 41316 20791 41372
rect 20791 41316 20795 41372
rect 20731 41312 20795 41316
rect 20811 41372 20875 41376
rect 20811 41316 20815 41372
rect 20815 41316 20871 41372
rect 20871 41316 20875 41372
rect 20811 41312 20875 41316
rect 20891 41372 20955 41376
rect 20891 41316 20895 41372
rect 20895 41316 20951 41372
rect 20951 41316 20955 41372
rect 20891 41312 20955 41316
rect 20971 41372 21035 41376
rect 20971 41316 20975 41372
rect 20975 41316 21031 41372
rect 21031 41316 21035 41372
rect 20971 41312 21035 41316
rect 16436 41244 16500 41308
rect 14596 41168 14660 41172
rect 14596 41112 14610 41168
rect 14610 41112 14660 41168
rect 14596 41108 14660 41112
rect 14964 41108 15028 41172
rect 3188 40972 3252 41036
rect 18092 40836 18156 40900
rect 3424 40828 3488 40832
rect 3424 40772 3428 40828
rect 3428 40772 3484 40828
rect 3484 40772 3488 40828
rect 3424 40768 3488 40772
rect 3504 40828 3568 40832
rect 3504 40772 3508 40828
rect 3508 40772 3564 40828
rect 3564 40772 3568 40828
rect 3504 40768 3568 40772
rect 3584 40828 3648 40832
rect 3584 40772 3588 40828
rect 3588 40772 3644 40828
rect 3644 40772 3648 40828
rect 3584 40768 3648 40772
rect 3664 40828 3728 40832
rect 3664 40772 3668 40828
rect 3668 40772 3724 40828
rect 3724 40772 3728 40828
rect 3664 40768 3728 40772
rect 8369 40828 8433 40832
rect 8369 40772 8373 40828
rect 8373 40772 8429 40828
rect 8429 40772 8433 40828
rect 8369 40768 8433 40772
rect 8449 40828 8513 40832
rect 8449 40772 8453 40828
rect 8453 40772 8509 40828
rect 8509 40772 8513 40828
rect 8449 40768 8513 40772
rect 8529 40828 8593 40832
rect 8529 40772 8533 40828
rect 8533 40772 8589 40828
rect 8589 40772 8593 40828
rect 8529 40768 8593 40772
rect 8609 40828 8673 40832
rect 8609 40772 8613 40828
rect 8613 40772 8669 40828
rect 8669 40772 8673 40828
rect 8609 40768 8673 40772
rect 13314 40828 13378 40832
rect 13314 40772 13318 40828
rect 13318 40772 13374 40828
rect 13374 40772 13378 40828
rect 13314 40768 13378 40772
rect 13394 40828 13458 40832
rect 13394 40772 13398 40828
rect 13398 40772 13454 40828
rect 13454 40772 13458 40828
rect 13394 40768 13458 40772
rect 13474 40828 13538 40832
rect 13474 40772 13478 40828
rect 13478 40772 13534 40828
rect 13534 40772 13538 40828
rect 13474 40768 13538 40772
rect 13554 40828 13618 40832
rect 13554 40772 13558 40828
rect 13558 40772 13614 40828
rect 13614 40772 13618 40828
rect 13554 40768 13618 40772
rect 18259 40828 18323 40832
rect 18259 40772 18263 40828
rect 18263 40772 18319 40828
rect 18319 40772 18323 40828
rect 18259 40768 18323 40772
rect 18339 40828 18403 40832
rect 18339 40772 18343 40828
rect 18343 40772 18399 40828
rect 18399 40772 18403 40828
rect 18339 40768 18403 40772
rect 18419 40828 18483 40832
rect 18419 40772 18423 40828
rect 18423 40772 18479 40828
rect 18479 40772 18483 40828
rect 18419 40768 18483 40772
rect 18499 40828 18563 40832
rect 18499 40772 18503 40828
rect 18503 40772 18559 40828
rect 18559 40772 18563 40828
rect 18499 40768 18563 40772
rect 16620 40700 16684 40764
rect 12204 40564 12268 40628
rect 1716 40428 1780 40492
rect 15332 40292 15396 40356
rect 5896 40284 5960 40288
rect 5896 40228 5900 40284
rect 5900 40228 5956 40284
rect 5956 40228 5960 40284
rect 5896 40224 5960 40228
rect 5976 40284 6040 40288
rect 5976 40228 5980 40284
rect 5980 40228 6036 40284
rect 6036 40228 6040 40284
rect 5976 40224 6040 40228
rect 6056 40284 6120 40288
rect 6056 40228 6060 40284
rect 6060 40228 6116 40284
rect 6116 40228 6120 40284
rect 6056 40224 6120 40228
rect 6136 40284 6200 40288
rect 6136 40228 6140 40284
rect 6140 40228 6196 40284
rect 6196 40228 6200 40284
rect 6136 40224 6200 40228
rect 10841 40284 10905 40288
rect 10841 40228 10845 40284
rect 10845 40228 10901 40284
rect 10901 40228 10905 40284
rect 10841 40224 10905 40228
rect 10921 40284 10985 40288
rect 10921 40228 10925 40284
rect 10925 40228 10981 40284
rect 10981 40228 10985 40284
rect 10921 40224 10985 40228
rect 11001 40284 11065 40288
rect 11001 40228 11005 40284
rect 11005 40228 11061 40284
rect 11061 40228 11065 40284
rect 11001 40224 11065 40228
rect 11081 40284 11145 40288
rect 11081 40228 11085 40284
rect 11085 40228 11141 40284
rect 11141 40228 11145 40284
rect 11081 40224 11145 40228
rect 15786 40284 15850 40288
rect 15786 40228 15790 40284
rect 15790 40228 15846 40284
rect 15846 40228 15850 40284
rect 15786 40224 15850 40228
rect 15866 40284 15930 40288
rect 15866 40228 15870 40284
rect 15870 40228 15926 40284
rect 15926 40228 15930 40284
rect 15866 40224 15930 40228
rect 15946 40284 16010 40288
rect 15946 40228 15950 40284
rect 15950 40228 16006 40284
rect 16006 40228 16010 40284
rect 15946 40224 16010 40228
rect 16026 40284 16090 40288
rect 16026 40228 16030 40284
rect 16030 40228 16086 40284
rect 16086 40228 16090 40284
rect 16026 40224 16090 40228
rect 20731 40284 20795 40288
rect 20731 40228 20735 40284
rect 20735 40228 20791 40284
rect 20791 40228 20795 40284
rect 20731 40224 20795 40228
rect 20811 40284 20875 40288
rect 20811 40228 20815 40284
rect 20815 40228 20871 40284
rect 20871 40228 20875 40284
rect 20811 40224 20875 40228
rect 20891 40284 20955 40288
rect 20891 40228 20895 40284
rect 20895 40228 20951 40284
rect 20951 40228 20955 40284
rect 20891 40224 20955 40228
rect 20971 40284 21035 40288
rect 20971 40228 20975 40284
rect 20975 40228 21031 40284
rect 21031 40228 21035 40284
rect 20971 40224 21035 40228
rect 7972 40080 8036 40084
rect 7972 40024 7986 40080
rect 7986 40024 8036 40080
rect 7972 40020 8036 40024
rect 12756 40020 12820 40084
rect 16988 40080 17052 40084
rect 16988 40024 17002 40080
rect 17002 40024 17052 40080
rect 16988 40020 17052 40024
rect 17908 40020 17972 40084
rect 18644 40080 18708 40084
rect 18644 40024 18658 40080
rect 18658 40024 18708 40080
rect 18644 40020 18708 40024
rect 17540 39748 17604 39812
rect 3424 39740 3488 39744
rect 3424 39684 3428 39740
rect 3428 39684 3484 39740
rect 3484 39684 3488 39740
rect 3424 39680 3488 39684
rect 3504 39740 3568 39744
rect 3504 39684 3508 39740
rect 3508 39684 3564 39740
rect 3564 39684 3568 39740
rect 3504 39680 3568 39684
rect 3584 39740 3648 39744
rect 3584 39684 3588 39740
rect 3588 39684 3644 39740
rect 3644 39684 3648 39740
rect 3584 39680 3648 39684
rect 3664 39740 3728 39744
rect 3664 39684 3668 39740
rect 3668 39684 3724 39740
rect 3724 39684 3728 39740
rect 3664 39680 3728 39684
rect 8369 39740 8433 39744
rect 8369 39684 8373 39740
rect 8373 39684 8429 39740
rect 8429 39684 8433 39740
rect 8369 39680 8433 39684
rect 8449 39740 8513 39744
rect 8449 39684 8453 39740
rect 8453 39684 8509 39740
rect 8509 39684 8513 39740
rect 8449 39680 8513 39684
rect 8529 39740 8593 39744
rect 8529 39684 8533 39740
rect 8533 39684 8589 39740
rect 8589 39684 8593 39740
rect 8529 39680 8593 39684
rect 8609 39740 8673 39744
rect 8609 39684 8613 39740
rect 8613 39684 8669 39740
rect 8669 39684 8673 39740
rect 8609 39680 8673 39684
rect 13314 39740 13378 39744
rect 13314 39684 13318 39740
rect 13318 39684 13374 39740
rect 13374 39684 13378 39740
rect 13314 39680 13378 39684
rect 13394 39740 13458 39744
rect 13394 39684 13398 39740
rect 13398 39684 13454 39740
rect 13454 39684 13458 39740
rect 13394 39680 13458 39684
rect 13474 39740 13538 39744
rect 13474 39684 13478 39740
rect 13478 39684 13534 39740
rect 13534 39684 13538 39740
rect 13474 39680 13538 39684
rect 13554 39740 13618 39744
rect 13554 39684 13558 39740
rect 13558 39684 13614 39740
rect 13614 39684 13618 39740
rect 13554 39680 13618 39684
rect 18259 39740 18323 39744
rect 18259 39684 18263 39740
rect 18263 39684 18319 39740
rect 18319 39684 18323 39740
rect 18259 39680 18323 39684
rect 18339 39740 18403 39744
rect 18339 39684 18343 39740
rect 18343 39684 18399 39740
rect 18399 39684 18403 39740
rect 18339 39680 18403 39684
rect 18419 39740 18483 39744
rect 18419 39684 18423 39740
rect 18423 39684 18479 39740
rect 18479 39684 18483 39740
rect 18419 39680 18483 39684
rect 18499 39740 18563 39744
rect 18499 39684 18503 39740
rect 18503 39684 18559 39740
rect 18559 39684 18563 39740
rect 18499 39680 18563 39684
rect 9996 39612 10060 39676
rect 16252 39264 16316 39268
rect 16252 39208 16266 39264
rect 16266 39208 16316 39264
rect 16252 39204 16316 39208
rect 18644 39264 18708 39268
rect 18644 39208 18658 39264
rect 18658 39208 18708 39264
rect 18644 39204 18708 39208
rect 5896 39196 5960 39200
rect 5896 39140 5900 39196
rect 5900 39140 5956 39196
rect 5956 39140 5960 39196
rect 5896 39136 5960 39140
rect 5976 39196 6040 39200
rect 5976 39140 5980 39196
rect 5980 39140 6036 39196
rect 6036 39140 6040 39196
rect 5976 39136 6040 39140
rect 6056 39196 6120 39200
rect 6056 39140 6060 39196
rect 6060 39140 6116 39196
rect 6116 39140 6120 39196
rect 6056 39136 6120 39140
rect 6136 39196 6200 39200
rect 6136 39140 6140 39196
rect 6140 39140 6196 39196
rect 6196 39140 6200 39196
rect 6136 39136 6200 39140
rect 10841 39196 10905 39200
rect 10841 39140 10845 39196
rect 10845 39140 10901 39196
rect 10901 39140 10905 39196
rect 10841 39136 10905 39140
rect 10921 39196 10985 39200
rect 10921 39140 10925 39196
rect 10925 39140 10981 39196
rect 10981 39140 10985 39196
rect 10921 39136 10985 39140
rect 11001 39196 11065 39200
rect 11001 39140 11005 39196
rect 11005 39140 11061 39196
rect 11061 39140 11065 39196
rect 11001 39136 11065 39140
rect 11081 39196 11145 39200
rect 11081 39140 11085 39196
rect 11085 39140 11141 39196
rect 11141 39140 11145 39196
rect 11081 39136 11145 39140
rect 15786 39196 15850 39200
rect 15786 39140 15790 39196
rect 15790 39140 15846 39196
rect 15846 39140 15850 39196
rect 15786 39136 15850 39140
rect 15866 39196 15930 39200
rect 15866 39140 15870 39196
rect 15870 39140 15926 39196
rect 15926 39140 15930 39196
rect 15866 39136 15930 39140
rect 15946 39196 16010 39200
rect 15946 39140 15950 39196
rect 15950 39140 16006 39196
rect 16006 39140 16010 39196
rect 15946 39136 16010 39140
rect 16026 39196 16090 39200
rect 16026 39140 16030 39196
rect 16030 39140 16086 39196
rect 16086 39140 16090 39196
rect 16026 39136 16090 39140
rect 20731 39196 20795 39200
rect 20731 39140 20735 39196
rect 20735 39140 20791 39196
rect 20791 39140 20795 39196
rect 20731 39136 20795 39140
rect 20811 39196 20875 39200
rect 20811 39140 20815 39196
rect 20815 39140 20871 39196
rect 20871 39140 20875 39196
rect 20811 39136 20875 39140
rect 20891 39196 20955 39200
rect 20891 39140 20895 39196
rect 20895 39140 20951 39196
rect 20951 39140 20955 39196
rect 20891 39136 20955 39140
rect 20971 39196 21035 39200
rect 20971 39140 20975 39196
rect 20975 39140 21031 39196
rect 21031 39140 21035 39196
rect 20971 39136 21035 39140
rect 5028 39068 5092 39132
rect 13860 39068 13924 39132
rect 980 38796 1044 38860
rect 3424 38652 3488 38656
rect 3424 38596 3428 38652
rect 3428 38596 3484 38652
rect 3484 38596 3488 38652
rect 3424 38592 3488 38596
rect 3504 38652 3568 38656
rect 3504 38596 3508 38652
rect 3508 38596 3564 38652
rect 3564 38596 3568 38652
rect 3504 38592 3568 38596
rect 3584 38652 3648 38656
rect 3584 38596 3588 38652
rect 3588 38596 3644 38652
rect 3644 38596 3648 38652
rect 3584 38592 3648 38596
rect 3664 38652 3728 38656
rect 3664 38596 3668 38652
rect 3668 38596 3724 38652
rect 3724 38596 3728 38652
rect 3664 38592 3728 38596
rect 8369 38652 8433 38656
rect 8369 38596 8373 38652
rect 8373 38596 8429 38652
rect 8429 38596 8433 38652
rect 8369 38592 8433 38596
rect 8449 38652 8513 38656
rect 8449 38596 8453 38652
rect 8453 38596 8509 38652
rect 8509 38596 8513 38652
rect 8449 38592 8513 38596
rect 8529 38652 8593 38656
rect 8529 38596 8533 38652
rect 8533 38596 8589 38652
rect 8589 38596 8593 38652
rect 8529 38592 8593 38596
rect 8609 38652 8673 38656
rect 8609 38596 8613 38652
rect 8613 38596 8669 38652
rect 8669 38596 8673 38652
rect 8609 38592 8673 38596
rect 13314 38652 13378 38656
rect 13314 38596 13318 38652
rect 13318 38596 13374 38652
rect 13374 38596 13378 38652
rect 13314 38592 13378 38596
rect 13394 38652 13458 38656
rect 13394 38596 13398 38652
rect 13398 38596 13454 38652
rect 13454 38596 13458 38652
rect 13394 38592 13458 38596
rect 13474 38652 13538 38656
rect 13474 38596 13478 38652
rect 13478 38596 13534 38652
rect 13534 38596 13538 38652
rect 13474 38592 13538 38596
rect 13554 38652 13618 38656
rect 13554 38596 13558 38652
rect 13558 38596 13614 38652
rect 13614 38596 13618 38652
rect 13554 38592 13618 38596
rect 17172 38720 17236 38724
rect 17172 38664 17186 38720
rect 17186 38664 17236 38720
rect 17172 38660 17236 38664
rect 18259 38652 18323 38656
rect 18259 38596 18263 38652
rect 18263 38596 18319 38652
rect 18319 38596 18323 38652
rect 18259 38592 18323 38596
rect 18339 38652 18403 38656
rect 18339 38596 18343 38652
rect 18343 38596 18399 38652
rect 18399 38596 18403 38652
rect 18339 38592 18403 38596
rect 18419 38652 18483 38656
rect 18419 38596 18423 38652
rect 18423 38596 18479 38652
rect 18479 38596 18483 38652
rect 18419 38592 18483 38596
rect 18499 38652 18563 38656
rect 18499 38596 18503 38652
rect 18503 38596 18559 38652
rect 18559 38596 18563 38652
rect 18499 38592 18563 38596
rect 12572 38116 12636 38180
rect 5896 38108 5960 38112
rect 5896 38052 5900 38108
rect 5900 38052 5956 38108
rect 5956 38052 5960 38108
rect 5896 38048 5960 38052
rect 5976 38108 6040 38112
rect 5976 38052 5980 38108
rect 5980 38052 6036 38108
rect 6036 38052 6040 38108
rect 5976 38048 6040 38052
rect 6056 38108 6120 38112
rect 6056 38052 6060 38108
rect 6060 38052 6116 38108
rect 6116 38052 6120 38108
rect 6056 38048 6120 38052
rect 6136 38108 6200 38112
rect 6136 38052 6140 38108
rect 6140 38052 6196 38108
rect 6196 38052 6200 38108
rect 6136 38048 6200 38052
rect 10841 38108 10905 38112
rect 10841 38052 10845 38108
rect 10845 38052 10901 38108
rect 10901 38052 10905 38108
rect 10841 38048 10905 38052
rect 10921 38108 10985 38112
rect 10921 38052 10925 38108
rect 10925 38052 10981 38108
rect 10981 38052 10985 38108
rect 10921 38048 10985 38052
rect 11001 38108 11065 38112
rect 11001 38052 11005 38108
rect 11005 38052 11061 38108
rect 11061 38052 11065 38108
rect 11001 38048 11065 38052
rect 11081 38108 11145 38112
rect 11081 38052 11085 38108
rect 11085 38052 11141 38108
rect 11141 38052 11145 38108
rect 11081 38048 11145 38052
rect 15786 38108 15850 38112
rect 15786 38052 15790 38108
rect 15790 38052 15846 38108
rect 15846 38052 15850 38108
rect 15786 38048 15850 38052
rect 15866 38108 15930 38112
rect 15866 38052 15870 38108
rect 15870 38052 15926 38108
rect 15926 38052 15930 38108
rect 15866 38048 15930 38052
rect 15946 38108 16010 38112
rect 15946 38052 15950 38108
rect 15950 38052 16006 38108
rect 16006 38052 16010 38108
rect 15946 38048 16010 38052
rect 16026 38108 16090 38112
rect 16026 38052 16030 38108
rect 16030 38052 16086 38108
rect 16086 38052 16090 38108
rect 16026 38048 16090 38052
rect 20731 38108 20795 38112
rect 20731 38052 20735 38108
rect 20735 38052 20791 38108
rect 20791 38052 20795 38108
rect 20731 38048 20795 38052
rect 20811 38108 20875 38112
rect 20811 38052 20815 38108
rect 20815 38052 20871 38108
rect 20871 38052 20875 38108
rect 20811 38048 20875 38052
rect 20891 38108 20955 38112
rect 20891 38052 20895 38108
rect 20895 38052 20951 38108
rect 20951 38052 20955 38108
rect 20891 38048 20955 38052
rect 20971 38108 21035 38112
rect 20971 38052 20975 38108
rect 20975 38052 21031 38108
rect 21031 38052 21035 38108
rect 20971 38048 21035 38052
rect 16436 37844 16500 37908
rect 19012 37844 19076 37908
rect 3424 37564 3488 37568
rect 3424 37508 3428 37564
rect 3428 37508 3484 37564
rect 3484 37508 3488 37564
rect 3424 37504 3488 37508
rect 3504 37564 3568 37568
rect 3504 37508 3508 37564
rect 3508 37508 3564 37564
rect 3564 37508 3568 37564
rect 3504 37504 3568 37508
rect 3584 37564 3648 37568
rect 3584 37508 3588 37564
rect 3588 37508 3644 37564
rect 3644 37508 3648 37564
rect 3584 37504 3648 37508
rect 3664 37564 3728 37568
rect 3664 37508 3668 37564
rect 3668 37508 3724 37564
rect 3724 37508 3728 37564
rect 3664 37504 3728 37508
rect 8369 37564 8433 37568
rect 8369 37508 8373 37564
rect 8373 37508 8429 37564
rect 8429 37508 8433 37564
rect 8369 37504 8433 37508
rect 8449 37564 8513 37568
rect 8449 37508 8453 37564
rect 8453 37508 8509 37564
rect 8509 37508 8513 37564
rect 8449 37504 8513 37508
rect 8529 37564 8593 37568
rect 8529 37508 8533 37564
rect 8533 37508 8589 37564
rect 8589 37508 8593 37564
rect 8529 37504 8593 37508
rect 8609 37564 8673 37568
rect 8609 37508 8613 37564
rect 8613 37508 8669 37564
rect 8669 37508 8673 37564
rect 8609 37504 8673 37508
rect 13314 37564 13378 37568
rect 13314 37508 13318 37564
rect 13318 37508 13374 37564
rect 13374 37508 13378 37564
rect 13314 37504 13378 37508
rect 13394 37564 13458 37568
rect 13394 37508 13398 37564
rect 13398 37508 13454 37564
rect 13454 37508 13458 37564
rect 13394 37504 13458 37508
rect 13474 37564 13538 37568
rect 13474 37508 13478 37564
rect 13478 37508 13534 37564
rect 13534 37508 13538 37564
rect 13474 37504 13538 37508
rect 13554 37564 13618 37568
rect 13554 37508 13558 37564
rect 13558 37508 13614 37564
rect 13614 37508 13618 37564
rect 13554 37504 13618 37508
rect 18259 37564 18323 37568
rect 18259 37508 18263 37564
rect 18263 37508 18319 37564
rect 18319 37508 18323 37564
rect 18259 37504 18323 37508
rect 18339 37564 18403 37568
rect 18339 37508 18343 37564
rect 18343 37508 18399 37564
rect 18399 37508 18403 37564
rect 18339 37504 18403 37508
rect 18419 37564 18483 37568
rect 18419 37508 18423 37564
rect 18423 37508 18479 37564
rect 18479 37508 18483 37564
rect 18419 37504 18483 37508
rect 18499 37564 18563 37568
rect 18499 37508 18503 37564
rect 18503 37508 18559 37564
rect 18559 37508 18563 37564
rect 18499 37504 18563 37508
rect 16804 37436 16868 37500
rect 6868 37300 6932 37364
rect 13124 37300 13188 37364
rect 19932 37300 19996 37364
rect 12204 37028 12268 37092
rect 5896 37020 5960 37024
rect 5896 36964 5900 37020
rect 5900 36964 5956 37020
rect 5956 36964 5960 37020
rect 5896 36960 5960 36964
rect 5976 37020 6040 37024
rect 5976 36964 5980 37020
rect 5980 36964 6036 37020
rect 6036 36964 6040 37020
rect 5976 36960 6040 36964
rect 6056 37020 6120 37024
rect 6056 36964 6060 37020
rect 6060 36964 6116 37020
rect 6116 36964 6120 37020
rect 6056 36960 6120 36964
rect 6136 37020 6200 37024
rect 6136 36964 6140 37020
rect 6140 36964 6196 37020
rect 6196 36964 6200 37020
rect 6136 36960 6200 36964
rect 10841 37020 10905 37024
rect 10841 36964 10845 37020
rect 10845 36964 10901 37020
rect 10901 36964 10905 37020
rect 10841 36960 10905 36964
rect 10921 37020 10985 37024
rect 10921 36964 10925 37020
rect 10925 36964 10981 37020
rect 10981 36964 10985 37020
rect 10921 36960 10985 36964
rect 11001 37020 11065 37024
rect 11001 36964 11005 37020
rect 11005 36964 11061 37020
rect 11061 36964 11065 37020
rect 11001 36960 11065 36964
rect 11081 37020 11145 37024
rect 11081 36964 11085 37020
rect 11085 36964 11141 37020
rect 11141 36964 11145 37020
rect 11081 36960 11145 36964
rect 15786 37020 15850 37024
rect 15786 36964 15790 37020
rect 15790 36964 15846 37020
rect 15846 36964 15850 37020
rect 15786 36960 15850 36964
rect 15866 37020 15930 37024
rect 15866 36964 15870 37020
rect 15870 36964 15926 37020
rect 15926 36964 15930 37020
rect 15866 36960 15930 36964
rect 15946 37020 16010 37024
rect 15946 36964 15950 37020
rect 15950 36964 16006 37020
rect 16006 36964 16010 37020
rect 15946 36960 16010 36964
rect 16026 37020 16090 37024
rect 16026 36964 16030 37020
rect 16030 36964 16086 37020
rect 16086 36964 16090 37020
rect 16026 36960 16090 36964
rect 20731 37020 20795 37024
rect 20731 36964 20735 37020
rect 20735 36964 20791 37020
rect 20791 36964 20795 37020
rect 20731 36960 20795 36964
rect 20811 37020 20875 37024
rect 20811 36964 20815 37020
rect 20815 36964 20871 37020
rect 20871 36964 20875 37020
rect 20811 36960 20875 36964
rect 20891 37020 20955 37024
rect 20891 36964 20895 37020
rect 20895 36964 20951 37020
rect 20951 36964 20955 37020
rect 20891 36960 20955 36964
rect 20971 37020 21035 37024
rect 20971 36964 20975 37020
rect 20975 36964 21031 37020
rect 21031 36964 21035 37020
rect 20971 36960 21035 36964
rect 18092 36892 18156 36956
rect 5396 36620 5460 36684
rect 10548 36756 10612 36820
rect 3424 36476 3488 36480
rect 3424 36420 3428 36476
rect 3428 36420 3484 36476
rect 3484 36420 3488 36476
rect 3424 36416 3488 36420
rect 3504 36476 3568 36480
rect 3504 36420 3508 36476
rect 3508 36420 3564 36476
rect 3564 36420 3568 36476
rect 3504 36416 3568 36420
rect 3584 36476 3648 36480
rect 3584 36420 3588 36476
rect 3588 36420 3644 36476
rect 3644 36420 3648 36476
rect 3584 36416 3648 36420
rect 3664 36476 3728 36480
rect 3664 36420 3668 36476
rect 3668 36420 3724 36476
rect 3724 36420 3728 36476
rect 3664 36416 3728 36420
rect 8369 36476 8433 36480
rect 8369 36420 8373 36476
rect 8373 36420 8429 36476
rect 8429 36420 8433 36476
rect 8369 36416 8433 36420
rect 8449 36476 8513 36480
rect 8449 36420 8453 36476
rect 8453 36420 8509 36476
rect 8509 36420 8513 36476
rect 8449 36416 8513 36420
rect 8529 36476 8593 36480
rect 8529 36420 8533 36476
rect 8533 36420 8589 36476
rect 8589 36420 8593 36476
rect 8529 36416 8593 36420
rect 8609 36476 8673 36480
rect 8609 36420 8613 36476
rect 8613 36420 8669 36476
rect 8669 36420 8673 36476
rect 8609 36416 8673 36420
rect 13314 36476 13378 36480
rect 13314 36420 13318 36476
rect 13318 36420 13374 36476
rect 13374 36420 13378 36476
rect 13314 36416 13378 36420
rect 13394 36476 13458 36480
rect 13394 36420 13398 36476
rect 13398 36420 13454 36476
rect 13454 36420 13458 36476
rect 13394 36416 13458 36420
rect 13474 36476 13538 36480
rect 13474 36420 13478 36476
rect 13478 36420 13534 36476
rect 13534 36420 13538 36476
rect 13474 36416 13538 36420
rect 13554 36476 13618 36480
rect 13554 36420 13558 36476
rect 13558 36420 13614 36476
rect 13614 36420 13618 36476
rect 13554 36416 13618 36420
rect 18259 36476 18323 36480
rect 18259 36420 18263 36476
rect 18263 36420 18319 36476
rect 18319 36420 18323 36476
rect 18259 36416 18323 36420
rect 18339 36476 18403 36480
rect 18339 36420 18343 36476
rect 18343 36420 18399 36476
rect 18399 36420 18403 36476
rect 18339 36416 18403 36420
rect 18419 36476 18483 36480
rect 18419 36420 18423 36476
rect 18423 36420 18479 36476
rect 18479 36420 18483 36476
rect 18419 36416 18483 36420
rect 18499 36476 18563 36480
rect 18499 36420 18503 36476
rect 18503 36420 18559 36476
rect 18559 36420 18563 36476
rect 18499 36416 18563 36420
rect 8156 36212 8220 36276
rect 4476 35940 4540 36004
rect 18644 36408 18708 36412
rect 18644 36352 18694 36408
rect 18694 36352 18708 36408
rect 18644 36348 18708 36352
rect 19012 36212 19076 36276
rect 18828 36076 18892 36140
rect 5896 35932 5960 35936
rect 5896 35876 5900 35932
rect 5900 35876 5956 35932
rect 5956 35876 5960 35932
rect 5896 35872 5960 35876
rect 5976 35932 6040 35936
rect 5976 35876 5980 35932
rect 5980 35876 6036 35932
rect 6036 35876 6040 35932
rect 5976 35872 6040 35876
rect 6056 35932 6120 35936
rect 6056 35876 6060 35932
rect 6060 35876 6116 35932
rect 6116 35876 6120 35932
rect 6056 35872 6120 35876
rect 6136 35932 6200 35936
rect 6136 35876 6140 35932
rect 6140 35876 6196 35932
rect 6196 35876 6200 35932
rect 6136 35872 6200 35876
rect 10841 35932 10905 35936
rect 10841 35876 10845 35932
rect 10845 35876 10901 35932
rect 10901 35876 10905 35932
rect 10841 35872 10905 35876
rect 10921 35932 10985 35936
rect 10921 35876 10925 35932
rect 10925 35876 10981 35932
rect 10981 35876 10985 35932
rect 10921 35872 10985 35876
rect 11001 35932 11065 35936
rect 11001 35876 11005 35932
rect 11005 35876 11061 35932
rect 11061 35876 11065 35932
rect 11001 35872 11065 35876
rect 11081 35932 11145 35936
rect 11081 35876 11085 35932
rect 11085 35876 11141 35932
rect 11141 35876 11145 35932
rect 11081 35872 11145 35876
rect 15786 35932 15850 35936
rect 15786 35876 15790 35932
rect 15790 35876 15846 35932
rect 15846 35876 15850 35932
rect 15786 35872 15850 35876
rect 15866 35932 15930 35936
rect 15866 35876 15870 35932
rect 15870 35876 15926 35932
rect 15926 35876 15930 35932
rect 15866 35872 15930 35876
rect 15946 35932 16010 35936
rect 15946 35876 15950 35932
rect 15950 35876 16006 35932
rect 16006 35876 16010 35932
rect 15946 35872 16010 35876
rect 16026 35932 16090 35936
rect 16026 35876 16030 35932
rect 16030 35876 16086 35932
rect 16086 35876 16090 35932
rect 16026 35872 16090 35876
rect 20731 35932 20795 35936
rect 20731 35876 20735 35932
rect 20735 35876 20791 35932
rect 20791 35876 20795 35932
rect 20731 35872 20795 35876
rect 20811 35932 20875 35936
rect 20811 35876 20815 35932
rect 20815 35876 20871 35932
rect 20871 35876 20875 35932
rect 20811 35872 20875 35876
rect 20891 35932 20955 35936
rect 20891 35876 20895 35932
rect 20895 35876 20951 35932
rect 20951 35876 20955 35932
rect 20891 35872 20955 35876
rect 20971 35932 21035 35936
rect 20971 35876 20975 35932
rect 20975 35876 21031 35932
rect 21031 35876 21035 35932
rect 20971 35872 21035 35876
rect 9076 35804 9140 35868
rect 8892 35668 8956 35732
rect 14412 35804 14476 35868
rect 19196 35804 19260 35868
rect 11468 35532 11532 35596
rect 3424 35388 3488 35392
rect 3424 35332 3428 35388
rect 3428 35332 3484 35388
rect 3484 35332 3488 35388
rect 3424 35328 3488 35332
rect 3504 35388 3568 35392
rect 3504 35332 3508 35388
rect 3508 35332 3564 35388
rect 3564 35332 3568 35388
rect 3504 35328 3568 35332
rect 3584 35388 3648 35392
rect 3584 35332 3588 35388
rect 3588 35332 3644 35388
rect 3644 35332 3648 35388
rect 3584 35328 3648 35332
rect 3664 35388 3728 35392
rect 3664 35332 3668 35388
rect 3668 35332 3724 35388
rect 3724 35332 3728 35388
rect 3664 35328 3728 35332
rect 8369 35388 8433 35392
rect 8369 35332 8373 35388
rect 8373 35332 8429 35388
rect 8429 35332 8433 35388
rect 8369 35328 8433 35332
rect 8449 35388 8513 35392
rect 8449 35332 8453 35388
rect 8453 35332 8509 35388
rect 8509 35332 8513 35388
rect 8449 35328 8513 35332
rect 8529 35388 8593 35392
rect 8529 35332 8533 35388
rect 8533 35332 8589 35388
rect 8589 35332 8593 35388
rect 8529 35328 8593 35332
rect 8609 35388 8673 35392
rect 8609 35332 8613 35388
rect 8613 35332 8669 35388
rect 8669 35332 8673 35388
rect 8609 35328 8673 35332
rect 13314 35388 13378 35392
rect 13314 35332 13318 35388
rect 13318 35332 13374 35388
rect 13374 35332 13378 35388
rect 13314 35328 13378 35332
rect 13394 35388 13458 35392
rect 13394 35332 13398 35388
rect 13398 35332 13454 35388
rect 13454 35332 13458 35388
rect 13394 35328 13458 35332
rect 13474 35388 13538 35392
rect 13474 35332 13478 35388
rect 13478 35332 13534 35388
rect 13534 35332 13538 35388
rect 13474 35328 13538 35332
rect 13554 35388 13618 35392
rect 13554 35332 13558 35388
rect 13558 35332 13614 35388
rect 13614 35332 13618 35388
rect 13554 35328 13618 35332
rect 18259 35388 18323 35392
rect 18259 35332 18263 35388
rect 18263 35332 18319 35388
rect 18319 35332 18323 35388
rect 18259 35328 18323 35332
rect 18339 35388 18403 35392
rect 18339 35332 18343 35388
rect 18343 35332 18399 35388
rect 18399 35332 18403 35388
rect 18339 35328 18403 35332
rect 18419 35388 18483 35392
rect 18419 35332 18423 35388
rect 18423 35332 18479 35388
rect 18479 35332 18483 35388
rect 18419 35328 18483 35332
rect 18499 35388 18563 35392
rect 18499 35332 18503 35388
rect 18503 35332 18559 35388
rect 18559 35332 18563 35388
rect 18499 35328 18563 35332
rect 796 35260 860 35324
rect 11284 35260 11348 35324
rect 14044 35260 14108 35324
rect 7788 35124 7852 35188
rect 14596 35184 14660 35188
rect 14596 35128 14610 35184
rect 14610 35128 14660 35184
rect 14596 35124 14660 35128
rect 5896 34844 5960 34848
rect 5896 34788 5900 34844
rect 5900 34788 5956 34844
rect 5956 34788 5960 34844
rect 5896 34784 5960 34788
rect 5976 34844 6040 34848
rect 5976 34788 5980 34844
rect 5980 34788 6036 34844
rect 6036 34788 6040 34844
rect 5976 34784 6040 34788
rect 6056 34844 6120 34848
rect 6056 34788 6060 34844
rect 6060 34788 6116 34844
rect 6116 34788 6120 34844
rect 6056 34784 6120 34788
rect 6136 34844 6200 34848
rect 6136 34788 6140 34844
rect 6140 34788 6196 34844
rect 6196 34788 6200 34844
rect 6136 34784 6200 34788
rect 10180 34640 10244 34644
rect 10180 34584 10194 34640
rect 10194 34584 10244 34640
rect 10180 34580 10244 34584
rect 6500 34444 6564 34508
rect 10364 34444 10428 34508
rect 10841 34844 10905 34848
rect 10841 34788 10845 34844
rect 10845 34788 10901 34844
rect 10901 34788 10905 34844
rect 10841 34784 10905 34788
rect 10921 34844 10985 34848
rect 10921 34788 10925 34844
rect 10925 34788 10981 34844
rect 10981 34788 10985 34844
rect 10921 34784 10985 34788
rect 11001 34844 11065 34848
rect 11001 34788 11005 34844
rect 11005 34788 11061 34844
rect 11061 34788 11065 34844
rect 11001 34784 11065 34788
rect 11081 34844 11145 34848
rect 11081 34788 11085 34844
rect 11085 34788 11141 34844
rect 11141 34788 11145 34844
rect 11081 34784 11145 34788
rect 15786 34844 15850 34848
rect 15786 34788 15790 34844
rect 15790 34788 15846 34844
rect 15846 34788 15850 34844
rect 15786 34784 15850 34788
rect 15866 34844 15930 34848
rect 15866 34788 15870 34844
rect 15870 34788 15926 34844
rect 15926 34788 15930 34844
rect 15866 34784 15930 34788
rect 15946 34844 16010 34848
rect 15946 34788 15950 34844
rect 15950 34788 16006 34844
rect 16006 34788 16010 34844
rect 15946 34784 16010 34788
rect 16026 34844 16090 34848
rect 16026 34788 16030 34844
rect 16030 34788 16086 34844
rect 16086 34788 16090 34844
rect 16026 34784 16090 34788
rect 20731 34844 20795 34848
rect 20731 34788 20735 34844
rect 20735 34788 20791 34844
rect 20791 34788 20795 34844
rect 20731 34784 20795 34788
rect 20811 34844 20875 34848
rect 20811 34788 20815 34844
rect 20815 34788 20871 34844
rect 20871 34788 20875 34844
rect 20811 34784 20875 34788
rect 20891 34844 20955 34848
rect 20891 34788 20895 34844
rect 20895 34788 20951 34844
rect 20951 34788 20955 34844
rect 20891 34784 20955 34788
rect 20971 34844 21035 34848
rect 20971 34788 20975 34844
rect 20975 34788 21031 34844
rect 21031 34788 21035 34844
rect 20971 34784 21035 34788
rect 11652 34716 11716 34780
rect 15148 34716 15212 34780
rect 15516 34776 15580 34780
rect 15516 34720 15530 34776
rect 15530 34720 15580 34776
rect 15516 34716 15580 34720
rect 11652 34640 11716 34644
rect 11652 34584 11666 34640
rect 11666 34584 11716 34640
rect 11652 34580 11716 34584
rect 12020 34580 12084 34644
rect 12204 34444 12268 34508
rect 4844 34308 4908 34372
rect 7420 34308 7484 34372
rect 3424 34300 3488 34304
rect 3424 34244 3428 34300
rect 3428 34244 3484 34300
rect 3484 34244 3488 34300
rect 3424 34240 3488 34244
rect 3504 34300 3568 34304
rect 3504 34244 3508 34300
rect 3508 34244 3564 34300
rect 3564 34244 3568 34300
rect 3504 34240 3568 34244
rect 3584 34300 3648 34304
rect 3584 34244 3588 34300
rect 3588 34244 3644 34300
rect 3644 34244 3648 34300
rect 3584 34240 3648 34244
rect 3664 34300 3728 34304
rect 3664 34244 3668 34300
rect 3668 34244 3724 34300
rect 3724 34244 3728 34300
rect 3664 34240 3728 34244
rect 8369 34300 8433 34304
rect 8369 34244 8373 34300
rect 8373 34244 8429 34300
rect 8429 34244 8433 34300
rect 8369 34240 8433 34244
rect 8449 34300 8513 34304
rect 8449 34244 8453 34300
rect 8453 34244 8509 34300
rect 8509 34244 8513 34300
rect 8449 34240 8513 34244
rect 8529 34300 8593 34304
rect 8529 34244 8533 34300
rect 8533 34244 8589 34300
rect 8589 34244 8593 34300
rect 8529 34240 8593 34244
rect 8609 34300 8673 34304
rect 8609 34244 8613 34300
rect 8613 34244 8669 34300
rect 8669 34244 8673 34300
rect 8609 34240 8673 34244
rect 13314 34300 13378 34304
rect 13314 34244 13318 34300
rect 13318 34244 13374 34300
rect 13374 34244 13378 34300
rect 13314 34240 13378 34244
rect 13394 34300 13458 34304
rect 13394 34244 13398 34300
rect 13398 34244 13454 34300
rect 13454 34244 13458 34300
rect 13394 34240 13458 34244
rect 13474 34300 13538 34304
rect 13474 34244 13478 34300
rect 13478 34244 13534 34300
rect 13534 34244 13538 34300
rect 13474 34240 13538 34244
rect 13554 34300 13618 34304
rect 13554 34244 13558 34300
rect 13558 34244 13614 34300
rect 13614 34244 13618 34300
rect 13554 34240 13618 34244
rect 18259 34300 18323 34304
rect 18259 34244 18263 34300
rect 18263 34244 18319 34300
rect 18319 34244 18323 34300
rect 18259 34240 18323 34244
rect 18339 34300 18403 34304
rect 18339 34244 18343 34300
rect 18343 34244 18399 34300
rect 18399 34244 18403 34300
rect 18339 34240 18403 34244
rect 18419 34300 18483 34304
rect 18419 34244 18423 34300
rect 18423 34244 18479 34300
rect 18479 34244 18483 34300
rect 18419 34240 18483 34244
rect 18499 34300 18563 34304
rect 18499 34244 18503 34300
rect 18503 34244 18559 34300
rect 18559 34244 18563 34300
rect 18499 34240 18563 34244
rect 4108 34172 4172 34236
rect 7420 34172 7484 34236
rect 7604 34172 7668 34236
rect 17356 34172 17420 34236
rect 19380 34096 19444 34100
rect 19380 34040 19430 34096
rect 19430 34040 19444 34096
rect 19380 34036 19444 34040
rect 3004 33900 3068 33964
rect 6500 33900 6564 33964
rect 16620 33900 16684 33964
rect 6316 33764 6380 33828
rect 19748 33764 19812 33828
rect 5896 33756 5960 33760
rect 5896 33700 5900 33756
rect 5900 33700 5956 33756
rect 5956 33700 5960 33756
rect 5896 33696 5960 33700
rect 5976 33756 6040 33760
rect 5976 33700 5980 33756
rect 5980 33700 6036 33756
rect 6036 33700 6040 33756
rect 5976 33696 6040 33700
rect 6056 33756 6120 33760
rect 6056 33700 6060 33756
rect 6060 33700 6116 33756
rect 6116 33700 6120 33756
rect 6056 33696 6120 33700
rect 6136 33756 6200 33760
rect 6136 33700 6140 33756
rect 6140 33700 6196 33756
rect 6196 33700 6200 33756
rect 6136 33696 6200 33700
rect 10841 33756 10905 33760
rect 10841 33700 10845 33756
rect 10845 33700 10901 33756
rect 10901 33700 10905 33756
rect 10841 33696 10905 33700
rect 10921 33756 10985 33760
rect 10921 33700 10925 33756
rect 10925 33700 10981 33756
rect 10981 33700 10985 33756
rect 10921 33696 10985 33700
rect 11001 33756 11065 33760
rect 11001 33700 11005 33756
rect 11005 33700 11061 33756
rect 11061 33700 11065 33756
rect 11001 33696 11065 33700
rect 11081 33756 11145 33760
rect 11081 33700 11085 33756
rect 11085 33700 11141 33756
rect 11141 33700 11145 33756
rect 11081 33696 11145 33700
rect 15786 33756 15850 33760
rect 15786 33700 15790 33756
rect 15790 33700 15846 33756
rect 15846 33700 15850 33756
rect 15786 33696 15850 33700
rect 15866 33756 15930 33760
rect 15866 33700 15870 33756
rect 15870 33700 15926 33756
rect 15926 33700 15930 33756
rect 15866 33696 15930 33700
rect 15946 33756 16010 33760
rect 15946 33700 15950 33756
rect 15950 33700 16006 33756
rect 16006 33700 16010 33756
rect 15946 33696 16010 33700
rect 16026 33756 16090 33760
rect 16026 33700 16030 33756
rect 16030 33700 16086 33756
rect 16086 33700 16090 33756
rect 16026 33696 16090 33700
rect 20731 33756 20795 33760
rect 20731 33700 20735 33756
rect 20735 33700 20791 33756
rect 20791 33700 20795 33756
rect 20731 33696 20795 33700
rect 20811 33756 20875 33760
rect 20811 33700 20815 33756
rect 20815 33700 20871 33756
rect 20871 33700 20875 33756
rect 20811 33696 20875 33700
rect 20891 33756 20955 33760
rect 20891 33700 20895 33756
rect 20895 33700 20951 33756
rect 20951 33700 20955 33756
rect 20891 33696 20955 33700
rect 20971 33756 21035 33760
rect 20971 33700 20975 33756
rect 20975 33700 21031 33756
rect 21031 33700 21035 33756
rect 20971 33696 21035 33700
rect 4476 33492 4540 33556
rect 428 33356 492 33420
rect 4292 33356 4356 33420
rect 3424 33212 3488 33216
rect 3424 33156 3428 33212
rect 3428 33156 3484 33212
rect 3484 33156 3488 33212
rect 3424 33152 3488 33156
rect 3504 33212 3568 33216
rect 3504 33156 3508 33212
rect 3508 33156 3564 33212
rect 3564 33156 3568 33212
rect 3504 33152 3568 33156
rect 3584 33212 3648 33216
rect 3584 33156 3588 33212
rect 3588 33156 3644 33212
rect 3644 33156 3648 33212
rect 3584 33152 3648 33156
rect 3664 33212 3728 33216
rect 3664 33156 3668 33212
rect 3668 33156 3724 33212
rect 3724 33156 3728 33212
rect 3664 33152 3728 33156
rect 18828 33220 18892 33284
rect 8369 33212 8433 33216
rect 8369 33156 8373 33212
rect 8373 33156 8429 33212
rect 8429 33156 8433 33212
rect 8369 33152 8433 33156
rect 8449 33212 8513 33216
rect 8449 33156 8453 33212
rect 8453 33156 8509 33212
rect 8509 33156 8513 33212
rect 8449 33152 8513 33156
rect 8529 33212 8593 33216
rect 8529 33156 8533 33212
rect 8533 33156 8589 33212
rect 8589 33156 8593 33212
rect 8529 33152 8593 33156
rect 8609 33212 8673 33216
rect 8609 33156 8613 33212
rect 8613 33156 8669 33212
rect 8669 33156 8673 33212
rect 8609 33152 8673 33156
rect 13314 33212 13378 33216
rect 13314 33156 13318 33212
rect 13318 33156 13374 33212
rect 13374 33156 13378 33212
rect 13314 33152 13378 33156
rect 13394 33212 13458 33216
rect 13394 33156 13398 33212
rect 13398 33156 13454 33212
rect 13454 33156 13458 33212
rect 13394 33152 13458 33156
rect 13474 33212 13538 33216
rect 13474 33156 13478 33212
rect 13478 33156 13534 33212
rect 13534 33156 13538 33212
rect 13474 33152 13538 33156
rect 13554 33212 13618 33216
rect 13554 33156 13558 33212
rect 13558 33156 13614 33212
rect 13614 33156 13618 33212
rect 13554 33152 13618 33156
rect 18259 33212 18323 33216
rect 18259 33156 18263 33212
rect 18263 33156 18319 33212
rect 18319 33156 18323 33212
rect 18259 33152 18323 33156
rect 18339 33212 18403 33216
rect 18339 33156 18343 33212
rect 18343 33156 18399 33212
rect 18399 33156 18403 33212
rect 18339 33152 18403 33156
rect 18419 33212 18483 33216
rect 18419 33156 18423 33212
rect 18423 33156 18479 33212
rect 18479 33156 18483 33212
rect 18419 33152 18483 33156
rect 18499 33212 18563 33216
rect 18499 33156 18503 33212
rect 18503 33156 18559 33212
rect 18559 33156 18563 33212
rect 18499 33152 18563 33156
rect 18828 32948 18892 33012
rect 19380 33280 19444 33284
rect 19380 33224 19394 33280
rect 19394 33224 19444 33280
rect 19380 33220 19444 33224
rect 19748 33280 19812 33284
rect 19748 33224 19762 33280
rect 19762 33224 19812 33280
rect 19748 33220 19812 33224
rect 19380 32948 19444 33012
rect 2452 32812 2516 32876
rect 6316 32812 6380 32876
rect 8892 32812 8956 32876
rect 5896 32668 5960 32672
rect 5896 32612 5900 32668
rect 5900 32612 5956 32668
rect 5956 32612 5960 32668
rect 5896 32608 5960 32612
rect 5976 32668 6040 32672
rect 5976 32612 5980 32668
rect 5980 32612 6036 32668
rect 6036 32612 6040 32668
rect 5976 32608 6040 32612
rect 6056 32668 6120 32672
rect 6056 32612 6060 32668
rect 6060 32612 6116 32668
rect 6116 32612 6120 32668
rect 6056 32608 6120 32612
rect 6136 32668 6200 32672
rect 6136 32612 6140 32668
rect 6140 32612 6196 32668
rect 6196 32612 6200 32668
rect 6136 32608 6200 32612
rect 10841 32668 10905 32672
rect 10841 32612 10845 32668
rect 10845 32612 10901 32668
rect 10901 32612 10905 32668
rect 10841 32608 10905 32612
rect 10921 32668 10985 32672
rect 10921 32612 10925 32668
rect 10925 32612 10981 32668
rect 10981 32612 10985 32668
rect 10921 32608 10985 32612
rect 11001 32668 11065 32672
rect 11001 32612 11005 32668
rect 11005 32612 11061 32668
rect 11061 32612 11065 32668
rect 11001 32608 11065 32612
rect 11081 32668 11145 32672
rect 11081 32612 11085 32668
rect 11085 32612 11141 32668
rect 11141 32612 11145 32668
rect 11081 32608 11145 32612
rect 15786 32668 15850 32672
rect 15786 32612 15790 32668
rect 15790 32612 15846 32668
rect 15846 32612 15850 32668
rect 15786 32608 15850 32612
rect 15866 32668 15930 32672
rect 15866 32612 15870 32668
rect 15870 32612 15926 32668
rect 15926 32612 15930 32668
rect 15866 32608 15930 32612
rect 15946 32668 16010 32672
rect 15946 32612 15950 32668
rect 15950 32612 16006 32668
rect 16006 32612 16010 32668
rect 15946 32608 16010 32612
rect 16026 32668 16090 32672
rect 16026 32612 16030 32668
rect 16030 32612 16086 32668
rect 16086 32612 16090 32668
rect 16026 32608 16090 32612
rect 20731 32668 20795 32672
rect 20731 32612 20735 32668
rect 20735 32612 20791 32668
rect 20791 32612 20795 32668
rect 20731 32608 20795 32612
rect 20811 32668 20875 32672
rect 20811 32612 20815 32668
rect 20815 32612 20871 32668
rect 20871 32612 20875 32668
rect 20811 32608 20875 32612
rect 20891 32668 20955 32672
rect 20891 32612 20895 32668
rect 20895 32612 20951 32668
rect 20951 32612 20955 32668
rect 20891 32608 20955 32612
rect 20971 32668 21035 32672
rect 20971 32612 20975 32668
rect 20975 32612 21031 32668
rect 21031 32612 21035 32668
rect 20971 32608 21035 32612
rect 13124 32600 13188 32604
rect 13124 32544 13138 32600
rect 13138 32544 13188 32600
rect 13124 32540 13188 32544
rect 17724 32540 17788 32604
rect 4660 32132 4724 32196
rect 3424 32124 3488 32128
rect 3424 32068 3428 32124
rect 3428 32068 3484 32124
rect 3484 32068 3488 32124
rect 3424 32064 3488 32068
rect 3504 32124 3568 32128
rect 3504 32068 3508 32124
rect 3508 32068 3564 32124
rect 3564 32068 3568 32124
rect 3504 32064 3568 32068
rect 3584 32124 3648 32128
rect 3584 32068 3588 32124
rect 3588 32068 3644 32124
rect 3644 32068 3648 32124
rect 3584 32064 3648 32068
rect 3664 32124 3728 32128
rect 3664 32068 3668 32124
rect 3668 32068 3724 32124
rect 3724 32068 3728 32124
rect 3664 32064 3728 32068
rect 8369 32124 8433 32128
rect 8369 32068 8373 32124
rect 8373 32068 8429 32124
rect 8429 32068 8433 32124
rect 8369 32064 8433 32068
rect 8449 32124 8513 32128
rect 8449 32068 8453 32124
rect 8453 32068 8509 32124
rect 8509 32068 8513 32124
rect 8449 32064 8513 32068
rect 8529 32124 8593 32128
rect 8529 32068 8533 32124
rect 8533 32068 8589 32124
rect 8589 32068 8593 32124
rect 8529 32064 8593 32068
rect 8609 32124 8673 32128
rect 8609 32068 8613 32124
rect 8613 32068 8669 32124
rect 8669 32068 8673 32124
rect 8609 32064 8673 32068
rect 13314 32124 13378 32128
rect 13314 32068 13318 32124
rect 13318 32068 13374 32124
rect 13374 32068 13378 32124
rect 13314 32064 13378 32068
rect 13394 32124 13458 32128
rect 13394 32068 13398 32124
rect 13398 32068 13454 32124
rect 13454 32068 13458 32124
rect 13394 32064 13458 32068
rect 13474 32124 13538 32128
rect 13474 32068 13478 32124
rect 13478 32068 13534 32124
rect 13534 32068 13538 32124
rect 13474 32064 13538 32068
rect 13554 32124 13618 32128
rect 13554 32068 13558 32124
rect 13558 32068 13614 32124
rect 13614 32068 13618 32124
rect 13554 32064 13618 32068
rect 18259 32124 18323 32128
rect 18259 32068 18263 32124
rect 18263 32068 18319 32124
rect 18319 32068 18323 32124
rect 18259 32064 18323 32068
rect 18339 32124 18403 32128
rect 18339 32068 18343 32124
rect 18343 32068 18399 32124
rect 18399 32068 18403 32124
rect 18339 32064 18403 32068
rect 18419 32124 18483 32128
rect 18419 32068 18423 32124
rect 18423 32068 18479 32124
rect 18479 32068 18483 32124
rect 18419 32064 18483 32068
rect 18499 32124 18563 32128
rect 18499 32068 18503 32124
rect 18503 32068 18559 32124
rect 18559 32068 18563 32124
rect 18499 32064 18563 32068
rect 5028 31860 5092 31924
rect 6868 31588 6932 31652
rect 7236 31588 7300 31652
rect 9812 31588 9876 31652
rect 5896 31580 5960 31584
rect 5896 31524 5900 31580
rect 5900 31524 5956 31580
rect 5956 31524 5960 31580
rect 5896 31520 5960 31524
rect 5976 31580 6040 31584
rect 5976 31524 5980 31580
rect 5980 31524 6036 31580
rect 6036 31524 6040 31580
rect 5976 31520 6040 31524
rect 6056 31580 6120 31584
rect 6056 31524 6060 31580
rect 6060 31524 6116 31580
rect 6116 31524 6120 31580
rect 6056 31520 6120 31524
rect 6136 31580 6200 31584
rect 6136 31524 6140 31580
rect 6140 31524 6196 31580
rect 6196 31524 6200 31580
rect 6136 31520 6200 31524
rect 10841 31580 10905 31584
rect 10841 31524 10845 31580
rect 10845 31524 10901 31580
rect 10901 31524 10905 31580
rect 10841 31520 10905 31524
rect 10921 31580 10985 31584
rect 10921 31524 10925 31580
rect 10925 31524 10981 31580
rect 10981 31524 10985 31580
rect 10921 31520 10985 31524
rect 11001 31580 11065 31584
rect 11001 31524 11005 31580
rect 11005 31524 11061 31580
rect 11061 31524 11065 31580
rect 11001 31520 11065 31524
rect 11081 31580 11145 31584
rect 11081 31524 11085 31580
rect 11085 31524 11141 31580
rect 11141 31524 11145 31580
rect 11081 31520 11145 31524
rect 15786 31580 15850 31584
rect 15786 31524 15790 31580
rect 15790 31524 15846 31580
rect 15846 31524 15850 31580
rect 15786 31520 15850 31524
rect 15866 31580 15930 31584
rect 15866 31524 15870 31580
rect 15870 31524 15926 31580
rect 15926 31524 15930 31580
rect 15866 31520 15930 31524
rect 15946 31580 16010 31584
rect 15946 31524 15950 31580
rect 15950 31524 16006 31580
rect 16006 31524 16010 31580
rect 15946 31520 16010 31524
rect 16026 31580 16090 31584
rect 16026 31524 16030 31580
rect 16030 31524 16086 31580
rect 16086 31524 16090 31580
rect 16026 31520 16090 31524
rect 20731 31580 20795 31584
rect 20731 31524 20735 31580
rect 20735 31524 20791 31580
rect 20791 31524 20795 31580
rect 20731 31520 20795 31524
rect 20811 31580 20875 31584
rect 20811 31524 20815 31580
rect 20815 31524 20871 31580
rect 20871 31524 20875 31580
rect 20811 31520 20875 31524
rect 20891 31580 20955 31584
rect 20891 31524 20895 31580
rect 20895 31524 20951 31580
rect 20951 31524 20955 31580
rect 20891 31520 20955 31524
rect 20971 31580 21035 31584
rect 20971 31524 20975 31580
rect 20975 31524 21031 31580
rect 21031 31524 21035 31580
rect 20971 31520 21035 31524
rect 16436 31452 16500 31516
rect 19748 31452 19812 31516
rect 2268 31316 2332 31380
rect 16436 31316 16500 31380
rect 18092 31316 18156 31380
rect 7420 31180 7484 31244
rect 11284 31180 11348 31244
rect 4660 31044 4724 31108
rect 5212 31044 5276 31108
rect 5396 31044 5460 31108
rect 19932 31180 19996 31244
rect 3424 31036 3488 31040
rect 3424 30980 3428 31036
rect 3428 30980 3484 31036
rect 3484 30980 3488 31036
rect 3424 30976 3488 30980
rect 3504 31036 3568 31040
rect 3504 30980 3508 31036
rect 3508 30980 3564 31036
rect 3564 30980 3568 31036
rect 3504 30976 3568 30980
rect 3584 31036 3648 31040
rect 3584 30980 3588 31036
rect 3588 30980 3644 31036
rect 3644 30980 3648 31036
rect 3584 30976 3648 30980
rect 3664 31036 3728 31040
rect 3664 30980 3668 31036
rect 3668 30980 3724 31036
rect 3724 30980 3728 31036
rect 3664 30976 3728 30980
rect 8369 31036 8433 31040
rect 8369 30980 8373 31036
rect 8373 30980 8429 31036
rect 8429 30980 8433 31036
rect 8369 30976 8433 30980
rect 8449 31036 8513 31040
rect 8449 30980 8453 31036
rect 8453 30980 8509 31036
rect 8509 30980 8513 31036
rect 8449 30976 8513 30980
rect 8529 31036 8593 31040
rect 8529 30980 8533 31036
rect 8533 30980 8589 31036
rect 8589 30980 8593 31036
rect 8529 30976 8593 30980
rect 8609 31036 8673 31040
rect 8609 30980 8613 31036
rect 8613 30980 8669 31036
rect 8669 30980 8673 31036
rect 8609 30976 8673 30980
rect 5212 30772 5276 30836
rect 8156 30696 8220 30700
rect 8156 30640 8206 30696
rect 8206 30640 8220 30696
rect 8156 30636 8220 30640
rect 5896 30492 5960 30496
rect 5896 30436 5900 30492
rect 5900 30436 5956 30492
rect 5956 30436 5960 30492
rect 5896 30432 5960 30436
rect 5976 30492 6040 30496
rect 5976 30436 5980 30492
rect 5980 30436 6036 30492
rect 6036 30436 6040 30492
rect 5976 30432 6040 30436
rect 6056 30492 6120 30496
rect 6056 30436 6060 30492
rect 6060 30436 6116 30492
rect 6116 30436 6120 30492
rect 6056 30432 6120 30436
rect 6136 30492 6200 30496
rect 6136 30436 6140 30492
rect 6140 30436 6196 30492
rect 6196 30436 6200 30492
rect 6136 30432 6200 30436
rect 16804 31044 16868 31108
rect 13314 31036 13378 31040
rect 13314 30980 13318 31036
rect 13318 30980 13374 31036
rect 13374 30980 13378 31036
rect 13314 30976 13378 30980
rect 13394 31036 13458 31040
rect 13394 30980 13398 31036
rect 13398 30980 13454 31036
rect 13454 30980 13458 31036
rect 13394 30976 13458 30980
rect 13474 31036 13538 31040
rect 13474 30980 13478 31036
rect 13478 30980 13534 31036
rect 13534 30980 13538 31036
rect 13474 30976 13538 30980
rect 13554 31036 13618 31040
rect 13554 30980 13558 31036
rect 13558 30980 13614 31036
rect 13614 30980 13618 31036
rect 13554 30976 13618 30980
rect 18259 31036 18323 31040
rect 18259 30980 18263 31036
rect 18263 30980 18319 31036
rect 18319 30980 18323 31036
rect 18259 30976 18323 30980
rect 18339 31036 18403 31040
rect 18339 30980 18343 31036
rect 18343 30980 18399 31036
rect 18399 30980 18403 31036
rect 18339 30976 18403 30980
rect 18419 31036 18483 31040
rect 18419 30980 18423 31036
rect 18423 30980 18479 31036
rect 18479 30980 18483 31036
rect 18419 30976 18483 30980
rect 18499 31036 18563 31040
rect 18499 30980 18503 31036
rect 18503 30980 18559 31036
rect 18559 30980 18563 31036
rect 18499 30976 18563 30980
rect 14044 30500 14108 30564
rect 10841 30492 10905 30496
rect 10841 30436 10845 30492
rect 10845 30436 10901 30492
rect 10901 30436 10905 30492
rect 10841 30432 10905 30436
rect 10921 30492 10985 30496
rect 10921 30436 10925 30492
rect 10925 30436 10981 30492
rect 10981 30436 10985 30492
rect 10921 30432 10985 30436
rect 11001 30492 11065 30496
rect 11001 30436 11005 30492
rect 11005 30436 11061 30492
rect 11061 30436 11065 30492
rect 11001 30432 11065 30436
rect 11081 30492 11145 30496
rect 11081 30436 11085 30492
rect 11085 30436 11141 30492
rect 11141 30436 11145 30492
rect 11081 30432 11145 30436
rect 16620 30636 16684 30700
rect 15786 30492 15850 30496
rect 15786 30436 15790 30492
rect 15790 30436 15846 30492
rect 15846 30436 15850 30492
rect 15786 30432 15850 30436
rect 15866 30492 15930 30496
rect 15866 30436 15870 30492
rect 15870 30436 15926 30492
rect 15926 30436 15930 30492
rect 15866 30432 15930 30436
rect 15946 30492 16010 30496
rect 15946 30436 15950 30492
rect 15950 30436 16006 30492
rect 16006 30436 16010 30492
rect 15946 30432 16010 30436
rect 16026 30492 16090 30496
rect 16026 30436 16030 30492
rect 16030 30436 16086 30492
rect 16086 30436 16090 30492
rect 16026 30432 16090 30436
rect 19012 30500 19076 30564
rect 20731 30492 20795 30496
rect 20731 30436 20735 30492
rect 20735 30436 20791 30492
rect 20791 30436 20795 30492
rect 20731 30432 20795 30436
rect 20811 30492 20875 30496
rect 20811 30436 20815 30492
rect 20815 30436 20871 30492
rect 20871 30436 20875 30492
rect 20811 30432 20875 30436
rect 20891 30492 20955 30496
rect 20891 30436 20895 30492
rect 20895 30436 20951 30492
rect 20951 30436 20955 30492
rect 20891 30432 20955 30436
rect 20971 30492 21035 30496
rect 20971 30436 20975 30492
rect 20975 30436 21031 30492
rect 21031 30436 21035 30492
rect 20971 30432 21035 30436
rect 17356 30364 17420 30428
rect 19012 30364 19076 30428
rect 980 30152 1044 30156
rect 980 30096 1030 30152
rect 1030 30096 1044 30152
rect 980 30092 1044 30096
rect 2084 30092 2148 30156
rect 16804 30092 16868 30156
rect 3924 30016 3988 30020
rect 3924 29960 3974 30016
rect 3974 29960 3988 30016
rect 3924 29956 3988 29960
rect 3424 29948 3488 29952
rect 3424 29892 3428 29948
rect 3428 29892 3484 29948
rect 3484 29892 3488 29948
rect 3424 29888 3488 29892
rect 3504 29948 3568 29952
rect 3504 29892 3508 29948
rect 3508 29892 3564 29948
rect 3564 29892 3568 29948
rect 3504 29888 3568 29892
rect 3584 29948 3648 29952
rect 3584 29892 3588 29948
rect 3588 29892 3644 29948
rect 3644 29892 3648 29948
rect 3584 29888 3648 29892
rect 3664 29948 3728 29952
rect 3664 29892 3668 29948
rect 3668 29892 3724 29948
rect 3724 29892 3728 29948
rect 3664 29888 3728 29892
rect 8369 29948 8433 29952
rect 8369 29892 8373 29948
rect 8373 29892 8429 29948
rect 8429 29892 8433 29948
rect 8369 29888 8433 29892
rect 8449 29948 8513 29952
rect 8449 29892 8453 29948
rect 8453 29892 8509 29948
rect 8509 29892 8513 29948
rect 8449 29888 8513 29892
rect 8529 29948 8593 29952
rect 8529 29892 8533 29948
rect 8533 29892 8589 29948
rect 8589 29892 8593 29948
rect 8529 29888 8593 29892
rect 8609 29948 8673 29952
rect 8609 29892 8613 29948
rect 8613 29892 8669 29948
rect 8669 29892 8673 29948
rect 8609 29888 8673 29892
rect 13314 29948 13378 29952
rect 13314 29892 13318 29948
rect 13318 29892 13374 29948
rect 13374 29892 13378 29948
rect 13314 29888 13378 29892
rect 13394 29948 13458 29952
rect 13394 29892 13398 29948
rect 13398 29892 13454 29948
rect 13454 29892 13458 29948
rect 13394 29888 13458 29892
rect 13474 29948 13538 29952
rect 13474 29892 13478 29948
rect 13478 29892 13534 29948
rect 13534 29892 13538 29948
rect 13474 29888 13538 29892
rect 13554 29948 13618 29952
rect 13554 29892 13558 29948
rect 13558 29892 13614 29948
rect 13614 29892 13618 29948
rect 13554 29888 13618 29892
rect 18259 29948 18323 29952
rect 18259 29892 18263 29948
rect 18263 29892 18319 29948
rect 18319 29892 18323 29948
rect 18259 29888 18323 29892
rect 18339 29948 18403 29952
rect 18339 29892 18343 29948
rect 18343 29892 18399 29948
rect 18399 29892 18403 29948
rect 18339 29888 18403 29892
rect 18419 29948 18483 29952
rect 18419 29892 18423 29948
rect 18423 29892 18479 29948
rect 18479 29892 18483 29948
rect 18419 29888 18483 29892
rect 18499 29948 18563 29952
rect 18499 29892 18503 29948
rect 18503 29892 18559 29948
rect 18559 29892 18563 29948
rect 18499 29888 18563 29892
rect 4292 29820 4356 29884
rect 7420 29820 7484 29884
rect 5212 29684 5276 29748
rect 14228 29684 14292 29748
rect 7788 29412 7852 29476
rect 5896 29404 5960 29408
rect 5896 29348 5900 29404
rect 5900 29348 5956 29404
rect 5956 29348 5960 29404
rect 5896 29344 5960 29348
rect 5976 29404 6040 29408
rect 5976 29348 5980 29404
rect 5980 29348 6036 29404
rect 6036 29348 6040 29404
rect 5976 29344 6040 29348
rect 6056 29404 6120 29408
rect 6056 29348 6060 29404
rect 6060 29348 6116 29404
rect 6116 29348 6120 29404
rect 6056 29344 6120 29348
rect 6136 29404 6200 29408
rect 6136 29348 6140 29404
rect 6140 29348 6196 29404
rect 6196 29348 6200 29404
rect 6136 29344 6200 29348
rect 10841 29404 10905 29408
rect 10841 29348 10845 29404
rect 10845 29348 10901 29404
rect 10901 29348 10905 29404
rect 10841 29344 10905 29348
rect 10921 29404 10985 29408
rect 10921 29348 10925 29404
rect 10925 29348 10981 29404
rect 10981 29348 10985 29404
rect 10921 29344 10985 29348
rect 11001 29404 11065 29408
rect 11001 29348 11005 29404
rect 11005 29348 11061 29404
rect 11061 29348 11065 29404
rect 11001 29344 11065 29348
rect 11081 29404 11145 29408
rect 11081 29348 11085 29404
rect 11085 29348 11141 29404
rect 11141 29348 11145 29404
rect 11081 29344 11145 29348
rect 3004 29276 3068 29340
rect 4660 29276 4724 29340
rect 5028 29276 5092 29340
rect 19380 29548 19444 29612
rect 15786 29404 15850 29408
rect 15786 29348 15790 29404
rect 15790 29348 15846 29404
rect 15846 29348 15850 29404
rect 15786 29344 15850 29348
rect 15866 29404 15930 29408
rect 15866 29348 15870 29404
rect 15870 29348 15926 29404
rect 15926 29348 15930 29404
rect 15866 29344 15930 29348
rect 15946 29404 16010 29408
rect 15946 29348 15950 29404
rect 15950 29348 16006 29404
rect 16006 29348 16010 29404
rect 15946 29344 16010 29348
rect 16026 29404 16090 29408
rect 16026 29348 16030 29404
rect 16030 29348 16086 29404
rect 16086 29348 16090 29404
rect 16026 29344 16090 29348
rect 20731 29404 20795 29408
rect 20731 29348 20735 29404
rect 20735 29348 20791 29404
rect 20791 29348 20795 29404
rect 20731 29344 20795 29348
rect 20811 29404 20875 29408
rect 20811 29348 20815 29404
rect 20815 29348 20871 29404
rect 20871 29348 20875 29404
rect 20811 29344 20875 29348
rect 20891 29404 20955 29408
rect 20891 29348 20895 29404
rect 20895 29348 20951 29404
rect 20951 29348 20955 29404
rect 20891 29344 20955 29348
rect 20971 29404 21035 29408
rect 20971 29348 20975 29404
rect 20975 29348 21031 29404
rect 21031 29348 21035 29404
rect 20971 29344 21035 29348
rect 1164 29004 1228 29068
rect 1532 29004 1596 29068
rect 9444 29140 9508 29204
rect 13124 29276 13188 29340
rect 14228 29140 14292 29204
rect 16436 29140 16500 29204
rect 18644 29140 18708 29204
rect 1900 28868 1964 28932
rect 9260 29004 9324 29068
rect 9444 29064 9508 29068
rect 9444 29008 9458 29064
rect 9458 29008 9508 29064
rect 9444 29004 9508 29008
rect 10548 29004 10612 29068
rect 14412 29004 14476 29068
rect 15148 29064 15212 29068
rect 15148 29008 15198 29064
rect 15198 29008 15212 29064
rect 15148 29004 15212 29008
rect 16988 29004 17052 29068
rect 17724 29004 17788 29068
rect 12756 28928 12820 28932
rect 12756 28872 12770 28928
rect 12770 28872 12820 28928
rect 12756 28868 12820 28872
rect 12940 28868 13004 28932
rect 3424 28860 3488 28864
rect 3424 28804 3428 28860
rect 3428 28804 3484 28860
rect 3484 28804 3488 28860
rect 3424 28800 3488 28804
rect 3504 28860 3568 28864
rect 3504 28804 3508 28860
rect 3508 28804 3564 28860
rect 3564 28804 3568 28860
rect 3504 28800 3568 28804
rect 3584 28860 3648 28864
rect 3584 28804 3588 28860
rect 3588 28804 3644 28860
rect 3644 28804 3648 28860
rect 3584 28800 3648 28804
rect 3664 28860 3728 28864
rect 3664 28804 3668 28860
rect 3668 28804 3724 28860
rect 3724 28804 3728 28860
rect 3664 28800 3728 28804
rect 8369 28860 8433 28864
rect 8369 28804 8373 28860
rect 8373 28804 8429 28860
rect 8429 28804 8433 28860
rect 8369 28800 8433 28804
rect 8449 28860 8513 28864
rect 8449 28804 8453 28860
rect 8453 28804 8509 28860
rect 8509 28804 8513 28860
rect 8449 28800 8513 28804
rect 8529 28860 8593 28864
rect 8529 28804 8533 28860
rect 8533 28804 8589 28860
rect 8589 28804 8593 28860
rect 8529 28800 8593 28804
rect 8609 28860 8673 28864
rect 8609 28804 8613 28860
rect 8613 28804 8669 28860
rect 8669 28804 8673 28860
rect 8609 28800 8673 28804
rect 13314 28860 13378 28864
rect 13314 28804 13318 28860
rect 13318 28804 13374 28860
rect 13374 28804 13378 28860
rect 13314 28800 13378 28804
rect 13394 28860 13458 28864
rect 13394 28804 13398 28860
rect 13398 28804 13454 28860
rect 13454 28804 13458 28860
rect 13394 28800 13458 28804
rect 13474 28860 13538 28864
rect 13474 28804 13478 28860
rect 13478 28804 13534 28860
rect 13534 28804 13538 28860
rect 13474 28800 13538 28804
rect 13554 28860 13618 28864
rect 13554 28804 13558 28860
rect 13558 28804 13614 28860
rect 13614 28804 13618 28860
rect 13554 28800 13618 28804
rect 18259 28860 18323 28864
rect 18259 28804 18263 28860
rect 18263 28804 18319 28860
rect 18319 28804 18323 28860
rect 18259 28800 18323 28804
rect 18339 28860 18403 28864
rect 18339 28804 18343 28860
rect 18343 28804 18399 28860
rect 18399 28804 18403 28860
rect 18339 28800 18403 28804
rect 18419 28860 18483 28864
rect 18419 28804 18423 28860
rect 18423 28804 18479 28860
rect 18479 28804 18483 28860
rect 18419 28800 18483 28804
rect 18499 28860 18563 28864
rect 18499 28804 18503 28860
rect 18503 28804 18559 28860
rect 18559 28804 18563 28860
rect 18499 28800 18563 28804
rect 7420 28732 7484 28796
rect 2268 28596 2332 28660
rect 14044 28596 14108 28660
rect 5896 28316 5960 28320
rect 5896 28260 5900 28316
rect 5900 28260 5956 28316
rect 5956 28260 5960 28316
rect 5896 28256 5960 28260
rect 5976 28316 6040 28320
rect 5976 28260 5980 28316
rect 5980 28260 6036 28316
rect 6036 28260 6040 28316
rect 5976 28256 6040 28260
rect 6056 28316 6120 28320
rect 6056 28260 6060 28316
rect 6060 28260 6116 28316
rect 6116 28260 6120 28316
rect 6056 28256 6120 28260
rect 6136 28316 6200 28320
rect 6136 28260 6140 28316
rect 6140 28260 6196 28316
rect 6196 28260 6200 28316
rect 6136 28256 6200 28260
rect 10841 28316 10905 28320
rect 10841 28260 10845 28316
rect 10845 28260 10901 28316
rect 10901 28260 10905 28316
rect 10841 28256 10905 28260
rect 10921 28316 10985 28320
rect 10921 28260 10925 28316
rect 10925 28260 10981 28316
rect 10981 28260 10985 28316
rect 10921 28256 10985 28260
rect 11001 28316 11065 28320
rect 11001 28260 11005 28316
rect 11005 28260 11061 28316
rect 11061 28260 11065 28316
rect 11001 28256 11065 28260
rect 11081 28316 11145 28320
rect 11081 28260 11085 28316
rect 11085 28260 11141 28316
rect 11141 28260 11145 28316
rect 11081 28256 11145 28260
rect 2084 28188 2148 28252
rect 2820 28188 2884 28252
rect 12756 28460 12820 28524
rect 5028 28052 5092 28116
rect 2636 27916 2700 27980
rect 15786 28316 15850 28320
rect 15786 28260 15790 28316
rect 15790 28260 15846 28316
rect 15846 28260 15850 28316
rect 15786 28256 15850 28260
rect 15866 28316 15930 28320
rect 15866 28260 15870 28316
rect 15870 28260 15926 28316
rect 15926 28260 15930 28316
rect 15866 28256 15930 28260
rect 15946 28316 16010 28320
rect 15946 28260 15950 28316
rect 15950 28260 16006 28316
rect 16006 28260 16010 28316
rect 15946 28256 16010 28260
rect 16026 28316 16090 28320
rect 16026 28260 16030 28316
rect 16030 28260 16086 28316
rect 16086 28260 16090 28316
rect 16026 28256 16090 28260
rect 20731 28316 20795 28320
rect 20731 28260 20735 28316
rect 20735 28260 20791 28316
rect 20791 28260 20795 28316
rect 20731 28256 20795 28260
rect 20811 28316 20875 28320
rect 20811 28260 20815 28316
rect 20815 28260 20871 28316
rect 20871 28260 20875 28316
rect 20811 28256 20875 28260
rect 20891 28316 20955 28320
rect 20891 28260 20895 28316
rect 20895 28260 20951 28316
rect 20951 28260 20955 28316
rect 20891 28256 20955 28260
rect 20971 28316 21035 28320
rect 20971 28260 20975 28316
rect 20975 28260 21031 28316
rect 21031 28260 21035 28316
rect 20971 28256 21035 28260
rect 15148 28188 15212 28252
rect 19380 28188 19444 28252
rect 2268 27780 2332 27844
rect 2452 27780 2516 27844
rect 3424 27772 3488 27776
rect 3424 27716 3428 27772
rect 3428 27716 3484 27772
rect 3484 27716 3488 27772
rect 3424 27712 3488 27716
rect 3504 27772 3568 27776
rect 3504 27716 3508 27772
rect 3508 27716 3564 27772
rect 3564 27716 3568 27772
rect 3504 27712 3568 27716
rect 3584 27772 3648 27776
rect 3584 27716 3588 27772
rect 3588 27716 3644 27772
rect 3644 27716 3648 27772
rect 3584 27712 3648 27716
rect 3664 27772 3728 27776
rect 3664 27716 3668 27772
rect 3668 27716 3724 27772
rect 3724 27716 3728 27772
rect 3664 27712 3728 27716
rect 8369 27772 8433 27776
rect 8369 27716 8373 27772
rect 8373 27716 8429 27772
rect 8429 27716 8433 27772
rect 8369 27712 8433 27716
rect 8449 27772 8513 27776
rect 8449 27716 8453 27772
rect 8453 27716 8509 27772
rect 8509 27716 8513 27772
rect 8449 27712 8513 27716
rect 8529 27772 8593 27776
rect 8529 27716 8533 27772
rect 8533 27716 8589 27772
rect 8589 27716 8593 27772
rect 8529 27712 8593 27716
rect 8609 27772 8673 27776
rect 8609 27716 8613 27772
rect 8613 27716 8669 27772
rect 8669 27716 8673 27772
rect 8609 27712 8673 27716
rect 13314 27772 13378 27776
rect 13314 27716 13318 27772
rect 13318 27716 13374 27772
rect 13374 27716 13378 27772
rect 13314 27712 13378 27716
rect 13394 27772 13458 27776
rect 13394 27716 13398 27772
rect 13398 27716 13454 27772
rect 13454 27716 13458 27772
rect 13394 27712 13458 27716
rect 13474 27772 13538 27776
rect 13474 27716 13478 27772
rect 13478 27716 13534 27772
rect 13534 27716 13538 27772
rect 13474 27712 13538 27716
rect 13554 27772 13618 27776
rect 13554 27716 13558 27772
rect 13558 27716 13614 27772
rect 13614 27716 13618 27772
rect 13554 27712 13618 27716
rect 18259 27772 18323 27776
rect 18259 27716 18263 27772
rect 18263 27716 18319 27772
rect 18319 27716 18323 27772
rect 18259 27712 18323 27716
rect 18339 27772 18403 27776
rect 18339 27716 18343 27772
rect 18343 27716 18399 27772
rect 18399 27716 18403 27772
rect 18339 27712 18403 27716
rect 18419 27772 18483 27776
rect 18419 27716 18423 27772
rect 18423 27716 18479 27772
rect 18479 27716 18483 27772
rect 18419 27712 18483 27716
rect 18499 27772 18563 27776
rect 18499 27716 18503 27772
rect 18503 27716 18559 27772
rect 18559 27716 18563 27772
rect 18499 27712 18563 27716
rect 3004 27644 3068 27708
rect 3924 27704 3988 27708
rect 3924 27648 3974 27704
rect 3974 27648 3988 27704
rect 3924 27644 3988 27648
rect 14964 27644 15028 27708
rect 4108 27508 4172 27572
rect 19196 27644 19260 27708
rect 1348 27372 1412 27436
rect 4292 27236 4356 27300
rect 5896 27228 5960 27232
rect 5896 27172 5900 27228
rect 5900 27172 5956 27228
rect 5956 27172 5960 27228
rect 5896 27168 5960 27172
rect 5976 27228 6040 27232
rect 5976 27172 5980 27228
rect 5980 27172 6036 27228
rect 6036 27172 6040 27228
rect 5976 27168 6040 27172
rect 6056 27228 6120 27232
rect 6056 27172 6060 27228
rect 6060 27172 6116 27228
rect 6116 27172 6120 27228
rect 6056 27168 6120 27172
rect 6136 27228 6200 27232
rect 6136 27172 6140 27228
rect 6140 27172 6196 27228
rect 6196 27172 6200 27228
rect 6136 27168 6200 27172
rect 10841 27228 10905 27232
rect 10841 27172 10845 27228
rect 10845 27172 10901 27228
rect 10901 27172 10905 27228
rect 10841 27168 10905 27172
rect 10921 27228 10985 27232
rect 10921 27172 10925 27228
rect 10925 27172 10981 27228
rect 10981 27172 10985 27228
rect 10921 27168 10985 27172
rect 11001 27228 11065 27232
rect 11001 27172 11005 27228
rect 11005 27172 11061 27228
rect 11061 27172 11065 27228
rect 11001 27168 11065 27172
rect 11081 27228 11145 27232
rect 11081 27172 11085 27228
rect 11085 27172 11141 27228
rect 11141 27172 11145 27228
rect 11081 27168 11145 27172
rect 15786 27228 15850 27232
rect 15786 27172 15790 27228
rect 15790 27172 15846 27228
rect 15846 27172 15850 27228
rect 15786 27168 15850 27172
rect 15866 27228 15930 27232
rect 15866 27172 15870 27228
rect 15870 27172 15926 27228
rect 15926 27172 15930 27228
rect 15866 27168 15930 27172
rect 15946 27228 16010 27232
rect 15946 27172 15950 27228
rect 15950 27172 16006 27228
rect 16006 27172 16010 27228
rect 15946 27168 16010 27172
rect 16026 27228 16090 27232
rect 16026 27172 16030 27228
rect 16030 27172 16086 27228
rect 16086 27172 16090 27228
rect 16026 27168 16090 27172
rect 20731 27228 20795 27232
rect 20731 27172 20735 27228
rect 20735 27172 20791 27228
rect 20791 27172 20795 27228
rect 20731 27168 20795 27172
rect 20811 27228 20875 27232
rect 20811 27172 20815 27228
rect 20815 27172 20871 27228
rect 20871 27172 20875 27228
rect 20811 27168 20875 27172
rect 20891 27228 20955 27232
rect 20891 27172 20895 27228
rect 20895 27172 20951 27228
rect 20951 27172 20955 27228
rect 20891 27168 20955 27172
rect 20971 27228 21035 27232
rect 20971 27172 20975 27228
rect 20975 27172 21031 27228
rect 21031 27172 21035 27228
rect 20971 27168 21035 27172
rect 1716 27100 1780 27164
rect 9628 27100 9692 27164
rect 8156 27024 8220 27028
rect 8156 26968 8206 27024
rect 8206 26968 8220 27024
rect 8156 26964 8220 26968
rect 9812 26964 9876 27028
rect 12388 27024 12452 27028
rect 12388 26968 12402 27024
rect 12402 26968 12452 27024
rect 12388 26964 12452 26968
rect 17724 26964 17788 27028
rect 3424 26684 3488 26688
rect 3424 26628 3428 26684
rect 3428 26628 3484 26684
rect 3484 26628 3488 26684
rect 3424 26624 3488 26628
rect 3504 26684 3568 26688
rect 3504 26628 3508 26684
rect 3508 26628 3564 26684
rect 3564 26628 3568 26684
rect 3504 26624 3568 26628
rect 3584 26684 3648 26688
rect 3584 26628 3588 26684
rect 3588 26628 3644 26684
rect 3644 26628 3648 26684
rect 3584 26624 3648 26628
rect 3664 26684 3728 26688
rect 3664 26628 3668 26684
rect 3668 26628 3724 26684
rect 3724 26628 3728 26684
rect 3664 26624 3728 26628
rect 8369 26684 8433 26688
rect 8369 26628 8373 26684
rect 8373 26628 8429 26684
rect 8429 26628 8433 26684
rect 8369 26624 8433 26628
rect 8449 26684 8513 26688
rect 8449 26628 8453 26684
rect 8453 26628 8509 26684
rect 8509 26628 8513 26684
rect 8449 26624 8513 26628
rect 8529 26684 8593 26688
rect 8529 26628 8533 26684
rect 8533 26628 8589 26684
rect 8589 26628 8593 26684
rect 8529 26624 8593 26628
rect 8609 26684 8673 26688
rect 8609 26628 8613 26684
rect 8613 26628 8669 26684
rect 8669 26628 8673 26684
rect 8609 26624 8673 26628
rect 13314 26684 13378 26688
rect 13314 26628 13318 26684
rect 13318 26628 13374 26684
rect 13374 26628 13378 26684
rect 13314 26624 13378 26628
rect 13394 26684 13458 26688
rect 13394 26628 13398 26684
rect 13398 26628 13454 26684
rect 13454 26628 13458 26684
rect 13394 26624 13458 26628
rect 13474 26684 13538 26688
rect 13474 26628 13478 26684
rect 13478 26628 13534 26684
rect 13534 26628 13538 26684
rect 13474 26624 13538 26628
rect 13554 26684 13618 26688
rect 13554 26628 13558 26684
rect 13558 26628 13614 26684
rect 13614 26628 13618 26684
rect 13554 26624 13618 26628
rect 18259 26684 18323 26688
rect 18259 26628 18263 26684
rect 18263 26628 18319 26684
rect 18319 26628 18323 26684
rect 18259 26624 18323 26628
rect 18339 26684 18403 26688
rect 18339 26628 18343 26684
rect 18343 26628 18399 26684
rect 18399 26628 18403 26684
rect 18339 26624 18403 26628
rect 18419 26684 18483 26688
rect 18419 26628 18423 26684
rect 18423 26628 18479 26684
rect 18479 26628 18483 26684
rect 18419 26624 18483 26628
rect 18499 26684 18563 26688
rect 18499 26628 18503 26684
rect 18503 26628 18559 26684
rect 18559 26628 18563 26684
rect 18499 26624 18563 26628
rect 9812 26556 9876 26620
rect 13124 26556 13188 26620
rect 16620 26556 16684 26620
rect 4108 26284 4172 26348
rect 6868 26148 6932 26212
rect 11652 26148 11716 26212
rect 5896 26140 5960 26144
rect 5896 26084 5900 26140
rect 5900 26084 5956 26140
rect 5956 26084 5960 26140
rect 5896 26080 5960 26084
rect 5976 26140 6040 26144
rect 5976 26084 5980 26140
rect 5980 26084 6036 26140
rect 6036 26084 6040 26140
rect 5976 26080 6040 26084
rect 6056 26140 6120 26144
rect 6056 26084 6060 26140
rect 6060 26084 6116 26140
rect 6116 26084 6120 26140
rect 6056 26080 6120 26084
rect 6136 26140 6200 26144
rect 6136 26084 6140 26140
rect 6140 26084 6196 26140
rect 6196 26084 6200 26140
rect 6136 26080 6200 26084
rect 10841 26140 10905 26144
rect 10841 26084 10845 26140
rect 10845 26084 10901 26140
rect 10901 26084 10905 26140
rect 10841 26080 10905 26084
rect 10921 26140 10985 26144
rect 10921 26084 10925 26140
rect 10925 26084 10981 26140
rect 10981 26084 10985 26140
rect 10921 26080 10985 26084
rect 11001 26140 11065 26144
rect 11001 26084 11005 26140
rect 11005 26084 11061 26140
rect 11061 26084 11065 26140
rect 11001 26080 11065 26084
rect 11081 26140 11145 26144
rect 11081 26084 11085 26140
rect 11085 26084 11141 26140
rect 11141 26084 11145 26140
rect 11081 26080 11145 26084
rect 5396 25876 5460 25940
rect 3004 25740 3068 25804
rect 2452 25604 2516 25668
rect 6500 25740 6564 25804
rect 15786 26140 15850 26144
rect 15786 26084 15790 26140
rect 15790 26084 15846 26140
rect 15846 26084 15850 26140
rect 15786 26080 15850 26084
rect 15866 26140 15930 26144
rect 15866 26084 15870 26140
rect 15870 26084 15926 26140
rect 15926 26084 15930 26140
rect 15866 26080 15930 26084
rect 15946 26140 16010 26144
rect 15946 26084 15950 26140
rect 15950 26084 16006 26140
rect 16006 26084 16010 26140
rect 15946 26080 16010 26084
rect 16026 26140 16090 26144
rect 16026 26084 16030 26140
rect 16030 26084 16086 26140
rect 16086 26084 16090 26140
rect 16026 26080 16090 26084
rect 20731 26140 20795 26144
rect 20731 26084 20735 26140
rect 20735 26084 20791 26140
rect 20791 26084 20795 26140
rect 20731 26080 20795 26084
rect 20811 26140 20875 26144
rect 20811 26084 20815 26140
rect 20815 26084 20871 26140
rect 20871 26084 20875 26140
rect 20811 26080 20875 26084
rect 20891 26140 20955 26144
rect 20891 26084 20895 26140
rect 20895 26084 20951 26140
rect 20951 26084 20955 26140
rect 20891 26080 20955 26084
rect 20971 26140 21035 26144
rect 20971 26084 20975 26140
rect 20975 26084 21031 26140
rect 21031 26084 21035 26140
rect 20971 26080 21035 26084
rect 3424 25596 3488 25600
rect 3424 25540 3428 25596
rect 3428 25540 3484 25596
rect 3484 25540 3488 25596
rect 3424 25536 3488 25540
rect 3504 25596 3568 25600
rect 3504 25540 3508 25596
rect 3508 25540 3564 25596
rect 3564 25540 3568 25596
rect 3504 25536 3568 25540
rect 3584 25596 3648 25600
rect 3584 25540 3588 25596
rect 3588 25540 3644 25596
rect 3644 25540 3648 25596
rect 3584 25536 3648 25540
rect 3664 25596 3728 25600
rect 3664 25540 3668 25596
rect 3668 25540 3724 25596
rect 3724 25540 3728 25596
rect 3664 25536 3728 25540
rect 8369 25596 8433 25600
rect 8369 25540 8373 25596
rect 8373 25540 8429 25596
rect 8429 25540 8433 25596
rect 8369 25536 8433 25540
rect 8449 25596 8513 25600
rect 8449 25540 8453 25596
rect 8453 25540 8509 25596
rect 8509 25540 8513 25596
rect 8449 25536 8513 25540
rect 8529 25596 8593 25600
rect 8529 25540 8533 25596
rect 8533 25540 8589 25596
rect 8589 25540 8593 25596
rect 8529 25536 8593 25540
rect 8609 25596 8673 25600
rect 8609 25540 8613 25596
rect 8613 25540 8669 25596
rect 8669 25540 8673 25596
rect 8609 25536 8673 25540
rect 13314 25596 13378 25600
rect 13314 25540 13318 25596
rect 13318 25540 13374 25596
rect 13374 25540 13378 25596
rect 13314 25536 13378 25540
rect 13394 25596 13458 25600
rect 13394 25540 13398 25596
rect 13398 25540 13454 25596
rect 13454 25540 13458 25596
rect 13394 25536 13458 25540
rect 13474 25596 13538 25600
rect 13474 25540 13478 25596
rect 13478 25540 13534 25596
rect 13534 25540 13538 25596
rect 13474 25536 13538 25540
rect 13554 25596 13618 25600
rect 13554 25540 13558 25596
rect 13558 25540 13614 25596
rect 13614 25540 13618 25596
rect 13554 25536 13618 25540
rect 796 25468 860 25532
rect 2820 25392 2884 25396
rect 5028 25468 5092 25532
rect 9260 25468 9324 25532
rect 9628 25468 9692 25532
rect 2820 25336 2870 25392
rect 2870 25336 2884 25392
rect 2820 25332 2884 25336
rect 12940 25060 13004 25124
rect 15516 25120 15580 25124
rect 15516 25064 15566 25120
rect 15566 25064 15580 25120
rect 15516 25060 15580 25064
rect 5896 25052 5960 25056
rect 5896 24996 5900 25052
rect 5900 24996 5956 25052
rect 5956 24996 5960 25052
rect 5896 24992 5960 24996
rect 5976 25052 6040 25056
rect 5976 24996 5980 25052
rect 5980 24996 6036 25052
rect 6036 24996 6040 25052
rect 5976 24992 6040 24996
rect 6056 25052 6120 25056
rect 6056 24996 6060 25052
rect 6060 24996 6116 25052
rect 6116 24996 6120 25052
rect 6056 24992 6120 24996
rect 6136 25052 6200 25056
rect 6136 24996 6140 25052
rect 6140 24996 6196 25052
rect 6196 24996 6200 25052
rect 6136 24992 6200 24996
rect 8892 24924 8956 24988
rect 10841 25052 10905 25056
rect 10841 24996 10845 25052
rect 10845 24996 10901 25052
rect 10901 24996 10905 25052
rect 10841 24992 10905 24996
rect 10921 25052 10985 25056
rect 10921 24996 10925 25052
rect 10925 24996 10981 25052
rect 10981 24996 10985 25052
rect 10921 24992 10985 24996
rect 11001 25052 11065 25056
rect 11001 24996 11005 25052
rect 11005 24996 11061 25052
rect 11061 24996 11065 25052
rect 11001 24992 11065 24996
rect 11081 25052 11145 25056
rect 11081 24996 11085 25052
rect 11085 24996 11141 25052
rect 11141 24996 11145 25052
rect 11081 24992 11145 24996
rect 15786 25052 15850 25056
rect 15786 24996 15790 25052
rect 15790 24996 15846 25052
rect 15846 24996 15850 25052
rect 15786 24992 15850 24996
rect 15866 25052 15930 25056
rect 15866 24996 15870 25052
rect 15870 24996 15926 25052
rect 15926 24996 15930 25052
rect 15866 24992 15930 24996
rect 15946 25052 16010 25056
rect 15946 24996 15950 25052
rect 15950 24996 16006 25052
rect 16006 24996 16010 25052
rect 15946 24992 16010 24996
rect 16026 25052 16090 25056
rect 16026 24996 16030 25052
rect 16030 24996 16086 25052
rect 16086 24996 16090 25052
rect 16026 24992 16090 24996
rect 11284 24924 11348 24988
rect 6684 24848 6748 24852
rect 6684 24792 6734 24848
rect 6734 24792 6748 24848
rect 6684 24788 6748 24792
rect 18259 25596 18323 25600
rect 18259 25540 18263 25596
rect 18263 25540 18319 25596
rect 18319 25540 18323 25596
rect 18259 25536 18323 25540
rect 18339 25596 18403 25600
rect 18339 25540 18343 25596
rect 18343 25540 18399 25596
rect 18399 25540 18403 25596
rect 18339 25536 18403 25540
rect 18419 25596 18483 25600
rect 18419 25540 18423 25596
rect 18423 25540 18479 25596
rect 18479 25540 18483 25596
rect 18419 25536 18483 25540
rect 18499 25596 18563 25600
rect 18499 25540 18503 25596
rect 18503 25540 18559 25596
rect 18559 25540 18563 25596
rect 18499 25536 18563 25540
rect 19564 25060 19628 25124
rect 20731 25052 20795 25056
rect 20731 24996 20735 25052
rect 20735 24996 20791 25052
rect 20791 24996 20795 25052
rect 20731 24992 20795 24996
rect 20811 25052 20875 25056
rect 20811 24996 20815 25052
rect 20815 24996 20871 25052
rect 20871 24996 20875 25052
rect 20811 24992 20875 24996
rect 20891 25052 20955 25056
rect 20891 24996 20895 25052
rect 20895 24996 20951 25052
rect 20951 24996 20955 25052
rect 20891 24992 20955 24996
rect 20971 25052 21035 25056
rect 20971 24996 20975 25052
rect 20975 24996 21031 25052
rect 21031 24996 21035 25052
rect 20971 24992 21035 24996
rect 19196 24788 19260 24852
rect 6316 24516 6380 24580
rect 9628 24516 9692 24580
rect 3424 24508 3488 24512
rect 3424 24452 3428 24508
rect 3428 24452 3484 24508
rect 3484 24452 3488 24508
rect 3424 24448 3488 24452
rect 3504 24508 3568 24512
rect 3504 24452 3508 24508
rect 3508 24452 3564 24508
rect 3564 24452 3568 24508
rect 3504 24448 3568 24452
rect 3584 24508 3648 24512
rect 3584 24452 3588 24508
rect 3588 24452 3644 24508
rect 3644 24452 3648 24508
rect 3584 24448 3648 24452
rect 3664 24508 3728 24512
rect 3664 24452 3668 24508
rect 3668 24452 3724 24508
rect 3724 24452 3728 24508
rect 3664 24448 3728 24452
rect 8369 24508 8433 24512
rect 8369 24452 8373 24508
rect 8373 24452 8429 24508
rect 8429 24452 8433 24508
rect 8369 24448 8433 24452
rect 8449 24508 8513 24512
rect 8449 24452 8453 24508
rect 8453 24452 8509 24508
rect 8509 24452 8513 24508
rect 8449 24448 8513 24452
rect 8529 24508 8593 24512
rect 8529 24452 8533 24508
rect 8533 24452 8589 24508
rect 8589 24452 8593 24508
rect 8529 24448 8593 24452
rect 8609 24508 8673 24512
rect 8609 24452 8613 24508
rect 8613 24452 8669 24508
rect 8669 24452 8673 24508
rect 8609 24448 8673 24452
rect 13314 24508 13378 24512
rect 13314 24452 13318 24508
rect 13318 24452 13374 24508
rect 13374 24452 13378 24508
rect 13314 24448 13378 24452
rect 13394 24508 13458 24512
rect 13394 24452 13398 24508
rect 13398 24452 13454 24508
rect 13454 24452 13458 24508
rect 13394 24448 13458 24452
rect 13474 24508 13538 24512
rect 13474 24452 13478 24508
rect 13478 24452 13534 24508
rect 13534 24452 13538 24508
rect 13474 24448 13538 24452
rect 13554 24508 13618 24512
rect 13554 24452 13558 24508
rect 13558 24452 13614 24508
rect 13614 24452 13618 24508
rect 13554 24448 13618 24452
rect 18259 24508 18323 24512
rect 18259 24452 18263 24508
rect 18263 24452 18319 24508
rect 18319 24452 18323 24508
rect 18259 24448 18323 24452
rect 18339 24508 18403 24512
rect 18339 24452 18343 24508
rect 18343 24452 18399 24508
rect 18399 24452 18403 24508
rect 18339 24448 18403 24452
rect 18419 24508 18483 24512
rect 18419 24452 18423 24508
rect 18423 24452 18479 24508
rect 18479 24452 18483 24508
rect 18419 24448 18483 24452
rect 18499 24508 18563 24512
rect 18499 24452 18503 24508
rect 18503 24452 18559 24508
rect 18559 24452 18563 24508
rect 18499 24448 18563 24452
rect 4108 24244 4172 24308
rect 4660 24304 4724 24308
rect 4660 24248 4674 24304
rect 4674 24248 4724 24304
rect 4660 24244 4724 24248
rect 6316 24244 6380 24308
rect 1716 24108 1780 24172
rect 2636 24108 2700 24172
rect 16620 24108 16684 24172
rect 12572 23972 12636 24036
rect 5896 23964 5960 23968
rect 5896 23908 5900 23964
rect 5900 23908 5956 23964
rect 5956 23908 5960 23964
rect 5896 23904 5960 23908
rect 5976 23964 6040 23968
rect 5976 23908 5980 23964
rect 5980 23908 6036 23964
rect 6036 23908 6040 23964
rect 5976 23904 6040 23908
rect 6056 23964 6120 23968
rect 6056 23908 6060 23964
rect 6060 23908 6116 23964
rect 6116 23908 6120 23964
rect 6056 23904 6120 23908
rect 6136 23964 6200 23968
rect 6136 23908 6140 23964
rect 6140 23908 6196 23964
rect 6196 23908 6200 23964
rect 6136 23904 6200 23908
rect 10841 23964 10905 23968
rect 10841 23908 10845 23964
rect 10845 23908 10901 23964
rect 10901 23908 10905 23964
rect 10841 23904 10905 23908
rect 10921 23964 10985 23968
rect 10921 23908 10925 23964
rect 10925 23908 10981 23964
rect 10981 23908 10985 23964
rect 10921 23904 10985 23908
rect 11001 23964 11065 23968
rect 11001 23908 11005 23964
rect 11005 23908 11061 23964
rect 11061 23908 11065 23964
rect 11001 23904 11065 23908
rect 11081 23964 11145 23968
rect 11081 23908 11085 23964
rect 11085 23908 11141 23964
rect 11141 23908 11145 23964
rect 11081 23904 11145 23908
rect 15786 23964 15850 23968
rect 15786 23908 15790 23964
rect 15790 23908 15846 23964
rect 15846 23908 15850 23964
rect 15786 23904 15850 23908
rect 15866 23964 15930 23968
rect 15866 23908 15870 23964
rect 15870 23908 15926 23964
rect 15926 23908 15930 23964
rect 15866 23904 15930 23908
rect 15946 23964 16010 23968
rect 15946 23908 15950 23964
rect 15950 23908 16006 23964
rect 16006 23908 16010 23964
rect 15946 23904 16010 23908
rect 16026 23964 16090 23968
rect 16026 23908 16030 23964
rect 16030 23908 16086 23964
rect 16086 23908 16090 23964
rect 16026 23904 16090 23908
rect 20731 23964 20795 23968
rect 20731 23908 20735 23964
rect 20735 23908 20791 23964
rect 20791 23908 20795 23964
rect 20731 23904 20795 23908
rect 20811 23964 20875 23968
rect 20811 23908 20815 23964
rect 20815 23908 20871 23964
rect 20871 23908 20875 23964
rect 20811 23904 20875 23908
rect 20891 23964 20955 23968
rect 20891 23908 20895 23964
rect 20895 23908 20951 23964
rect 20951 23908 20955 23964
rect 20891 23904 20955 23908
rect 20971 23964 21035 23968
rect 20971 23908 20975 23964
rect 20975 23908 21031 23964
rect 21031 23908 21035 23964
rect 20971 23904 21035 23908
rect 1164 23836 1228 23900
rect 5028 23836 5092 23900
rect 5212 23896 5276 23900
rect 5212 23840 5226 23896
rect 5226 23840 5276 23896
rect 5212 23836 5276 23840
rect 7420 23836 7484 23900
rect 9628 23836 9692 23900
rect 4844 23564 4908 23628
rect 5212 23564 5276 23628
rect 9812 23700 9876 23764
rect 9260 23624 9324 23628
rect 9260 23568 9274 23624
rect 9274 23568 9324 23624
rect 1900 23428 1964 23492
rect 7052 23428 7116 23492
rect 3424 23420 3488 23424
rect 3424 23364 3428 23420
rect 3428 23364 3484 23420
rect 3484 23364 3488 23420
rect 3424 23360 3488 23364
rect 3504 23420 3568 23424
rect 3504 23364 3508 23420
rect 3508 23364 3564 23420
rect 3564 23364 3568 23420
rect 3504 23360 3568 23364
rect 3584 23420 3648 23424
rect 3584 23364 3588 23420
rect 3588 23364 3644 23420
rect 3644 23364 3648 23420
rect 3584 23360 3648 23364
rect 3664 23420 3728 23424
rect 3664 23364 3668 23420
rect 3668 23364 3724 23420
rect 3724 23364 3728 23420
rect 3664 23360 3728 23364
rect 4660 23292 4724 23356
rect 8369 23420 8433 23424
rect 8369 23364 8373 23420
rect 8373 23364 8429 23420
rect 8429 23364 8433 23420
rect 8369 23360 8433 23364
rect 8449 23420 8513 23424
rect 8449 23364 8453 23420
rect 8453 23364 8509 23420
rect 8509 23364 8513 23420
rect 8449 23360 8513 23364
rect 8529 23420 8593 23424
rect 8529 23364 8533 23420
rect 8533 23364 8589 23420
rect 8589 23364 8593 23420
rect 8529 23360 8593 23364
rect 8609 23420 8673 23424
rect 8609 23364 8613 23420
rect 8613 23364 8669 23420
rect 8669 23364 8673 23420
rect 8609 23360 8673 23364
rect 9260 23564 9324 23568
rect 9812 23564 9876 23628
rect 12756 23836 12820 23900
rect 12572 23700 12636 23764
rect 14596 23564 14660 23628
rect 17540 23564 17604 23628
rect 9628 23428 9692 23492
rect 16252 23428 16316 23492
rect 17356 23428 17420 23492
rect 13314 23420 13378 23424
rect 13314 23364 13318 23420
rect 13318 23364 13374 23420
rect 13374 23364 13378 23420
rect 13314 23360 13378 23364
rect 13394 23420 13458 23424
rect 13394 23364 13398 23420
rect 13398 23364 13454 23420
rect 13454 23364 13458 23420
rect 13394 23360 13458 23364
rect 13474 23420 13538 23424
rect 13474 23364 13478 23420
rect 13478 23364 13534 23420
rect 13534 23364 13538 23420
rect 13474 23360 13538 23364
rect 13554 23420 13618 23424
rect 13554 23364 13558 23420
rect 13558 23364 13614 23420
rect 13614 23364 13618 23420
rect 13554 23360 13618 23364
rect 18259 23420 18323 23424
rect 18259 23364 18263 23420
rect 18263 23364 18319 23420
rect 18319 23364 18323 23420
rect 18259 23360 18323 23364
rect 18339 23420 18403 23424
rect 18339 23364 18343 23420
rect 18343 23364 18399 23420
rect 18399 23364 18403 23420
rect 18339 23360 18403 23364
rect 18419 23420 18483 23424
rect 18419 23364 18423 23420
rect 18423 23364 18479 23420
rect 18479 23364 18483 23420
rect 18419 23360 18483 23364
rect 18499 23420 18563 23424
rect 18499 23364 18503 23420
rect 18503 23364 18559 23420
rect 18559 23364 18563 23420
rect 18499 23360 18563 23364
rect 3188 23020 3252 23084
rect 4844 23020 4908 23084
rect 9260 23020 9324 23084
rect 12020 23080 12084 23084
rect 12020 23024 12070 23080
rect 12070 23024 12084 23080
rect 12020 23020 12084 23024
rect 10180 22884 10244 22948
rect 5896 22876 5960 22880
rect 5896 22820 5900 22876
rect 5900 22820 5956 22876
rect 5956 22820 5960 22876
rect 5896 22816 5960 22820
rect 5976 22876 6040 22880
rect 5976 22820 5980 22876
rect 5980 22820 6036 22876
rect 6036 22820 6040 22876
rect 5976 22816 6040 22820
rect 6056 22876 6120 22880
rect 6056 22820 6060 22876
rect 6060 22820 6116 22876
rect 6116 22820 6120 22876
rect 6056 22816 6120 22820
rect 6136 22876 6200 22880
rect 6136 22820 6140 22876
rect 6140 22820 6196 22876
rect 6196 22820 6200 22876
rect 6136 22816 6200 22820
rect 10841 22876 10905 22880
rect 10841 22820 10845 22876
rect 10845 22820 10901 22876
rect 10901 22820 10905 22876
rect 10841 22816 10905 22820
rect 10921 22876 10985 22880
rect 10921 22820 10925 22876
rect 10925 22820 10981 22876
rect 10981 22820 10985 22876
rect 10921 22816 10985 22820
rect 11001 22876 11065 22880
rect 11001 22820 11005 22876
rect 11005 22820 11061 22876
rect 11061 22820 11065 22876
rect 11001 22816 11065 22820
rect 11081 22876 11145 22880
rect 11081 22820 11085 22876
rect 11085 22820 11141 22876
rect 11141 22820 11145 22876
rect 11081 22816 11145 22820
rect 15786 22876 15850 22880
rect 15786 22820 15790 22876
rect 15790 22820 15846 22876
rect 15846 22820 15850 22876
rect 15786 22816 15850 22820
rect 15866 22876 15930 22880
rect 15866 22820 15870 22876
rect 15870 22820 15926 22876
rect 15926 22820 15930 22876
rect 15866 22816 15930 22820
rect 15946 22876 16010 22880
rect 15946 22820 15950 22876
rect 15950 22820 16006 22876
rect 16006 22820 16010 22876
rect 15946 22816 16010 22820
rect 16026 22876 16090 22880
rect 16026 22820 16030 22876
rect 16030 22820 16086 22876
rect 16086 22820 16090 22876
rect 16026 22816 16090 22820
rect 20731 22876 20795 22880
rect 20731 22820 20735 22876
rect 20735 22820 20791 22876
rect 20791 22820 20795 22876
rect 20731 22816 20795 22820
rect 20811 22876 20875 22880
rect 20811 22820 20815 22876
rect 20815 22820 20871 22876
rect 20871 22820 20875 22876
rect 20811 22816 20875 22820
rect 20891 22876 20955 22880
rect 20891 22820 20895 22876
rect 20895 22820 20951 22876
rect 20951 22820 20955 22876
rect 20891 22816 20955 22820
rect 20971 22876 21035 22880
rect 20971 22820 20975 22876
rect 20975 22820 21031 22876
rect 21031 22820 21035 22876
rect 20971 22816 21035 22820
rect 2820 22748 2884 22812
rect 5580 22748 5644 22812
rect 7236 22748 7300 22812
rect 9076 22748 9140 22812
rect 10548 22808 10612 22812
rect 10548 22752 10598 22808
rect 10598 22752 10612 22808
rect 10548 22748 10612 22752
rect 9996 22612 10060 22676
rect 12204 22612 12268 22676
rect 14596 22672 14660 22676
rect 14596 22616 14646 22672
rect 14646 22616 14660 22672
rect 14596 22612 14660 22616
rect 14780 22612 14844 22676
rect 19932 22612 19996 22676
rect 18092 22476 18156 22540
rect 19748 22536 19812 22540
rect 19748 22480 19762 22536
rect 19762 22480 19812 22536
rect 19748 22476 19812 22480
rect 15516 22340 15580 22404
rect 16252 22340 16316 22404
rect 19380 22340 19444 22404
rect 3424 22332 3488 22336
rect 3424 22276 3428 22332
rect 3428 22276 3484 22332
rect 3484 22276 3488 22332
rect 3424 22272 3488 22276
rect 3504 22332 3568 22336
rect 3504 22276 3508 22332
rect 3508 22276 3564 22332
rect 3564 22276 3568 22332
rect 3504 22272 3568 22276
rect 3584 22332 3648 22336
rect 3584 22276 3588 22332
rect 3588 22276 3644 22332
rect 3644 22276 3648 22332
rect 3584 22272 3648 22276
rect 3664 22332 3728 22336
rect 3664 22276 3668 22332
rect 3668 22276 3724 22332
rect 3724 22276 3728 22332
rect 3664 22272 3728 22276
rect 8369 22332 8433 22336
rect 8369 22276 8373 22332
rect 8373 22276 8429 22332
rect 8429 22276 8433 22332
rect 8369 22272 8433 22276
rect 8449 22332 8513 22336
rect 8449 22276 8453 22332
rect 8453 22276 8509 22332
rect 8509 22276 8513 22332
rect 8449 22272 8513 22276
rect 8529 22332 8593 22336
rect 8529 22276 8533 22332
rect 8533 22276 8589 22332
rect 8589 22276 8593 22332
rect 8529 22272 8593 22276
rect 8609 22332 8673 22336
rect 8609 22276 8613 22332
rect 8613 22276 8669 22332
rect 8669 22276 8673 22332
rect 8609 22272 8673 22276
rect 13314 22332 13378 22336
rect 13314 22276 13318 22332
rect 13318 22276 13374 22332
rect 13374 22276 13378 22332
rect 13314 22272 13378 22276
rect 13394 22332 13458 22336
rect 13394 22276 13398 22332
rect 13398 22276 13454 22332
rect 13454 22276 13458 22332
rect 13394 22272 13458 22276
rect 13474 22332 13538 22336
rect 13474 22276 13478 22332
rect 13478 22276 13534 22332
rect 13534 22276 13538 22332
rect 13474 22272 13538 22276
rect 13554 22332 13618 22336
rect 13554 22276 13558 22332
rect 13558 22276 13614 22332
rect 13614 22276 13618 22332
rect 13554 22272 13618 22276
rect 18259 22332 18323 22336
rect 18259 22276 18263 22332
rect 18263 22276 18319 22332
rect 18319 22276 18323 22332
rect 18259 22272 18323 22276
rect 18339 22332 18403 22336
rect 18339 22276 18343 22332
rect 18343 22276 18399 22332
rect 18399 22276 18403 22332
rect 18339 22272 18403 22276
rect 18419 22332 18483 22336
rect 18419 22276 18423 22332
rect 18423 22276 18479 22332
rect 18479 22276 18483 22332
rect 18419 22272 18483 22276
rect 18499 22332 18563 22336
rect 18499 22276 18503 22332
rect 18503 22276 18559 22332
rect 18559 22276 18563 22332
rect 18499 22272 18563 22276
rect 4292 22204 4356 22268
rect 7420 22264 7484 22268
rect 7420 22208 7470 22264
rect 7470 22208 7484 22264
rect 7420 22204 7484 22208
rect 10548 22264 10612 22268
rect 10548 22208 10562 22264
rect 10562 22208 10612 22264
rect 10548 22204 10612 22208
rect 4108 22068 4172 22132
rect 15332 22068 15396 22132
rect 1900 21932 1964 21996
rect 11836 21932 11900 21996
rect 5896 21788 5960 21792
rect 5896 21732 5900 21788
rect 5900 21732 5956 21788
rect 5956 21732 5960 21788
rect 5896 21728 5960 21732
rect 5976 21788 6040 21792
rect 5976 21732 5980 21788
rect 5980 21732 6036 21788
rect 6036 21732 6040 21788
rect 5976 21728 6040 21732
rect 6056 21788 6120 21792
rect 6056 21732 6060 21788
rect 6060 21732 6116 21788
rect 6116 21732 6120 21788
rect 6056 21728 6120 21732
rect 6136 21788 6200 21792
rect 6136 21732 6140 21788
rect 6140 21732 6196 21788
rect 6196 21732 6200 21788
rect 6136 21728 6200 21732
rect 10841 21788 10905 21792
rect 10841 21732 10845 21788
rect 10845 21732 10901 21788
rect 10901 21732 10905 21788
rect 10841 21728 10905 21732
rect 10921 21788 10985 21792
rect 10921 21732 10925 21788
rect 10925 21732 10981 21788
rect 10981 21732 10985 21788
rect 10921 21728 10985 21732
rect 11001 21788 11065 21792
rect 11001 21732 11005 21788
rect 11005 21732 11061 21788
rect 11061 21732 11065 21788
rect 11001 21728 11065 21732
rect 11081 21788 11145 21792
rect 11081 21732 11085 21788
rect 11085 21732 11141 21788
rect 11141 21732 11145 21788
rect 11081 21728 11145 21732
rect 15786 21788 15850 21792
rect 15786 21732 15790 21788
rect 15790 21732 15846 21788
rect 15846 21732 15850 21788
rect 15786 21728 15850 21732
rect 15866 21788 15930 21792
rect 15866 21732 15870 21788
rect 15870 21732 15926 21788
rect 15926 21732 15930 21788
rect 15866 21728 15930 21732
rect 15946 21788 16010 21792
rect 15946 21732 15950 21788
rect 15950 21732 16006 21788
rect 16006 21732 16010 21788
rect 15946 21728 16010 21732
rect 16026 21788 16090 21792
rect 16026 21732 16030 21788
rect 16030 21732 16086 21788
rect 16086 21732 16090 21788
rect 16026 21728 16090 21732
rect 20731 21788 20795 21792
rect 20731 21732 20735 21788
rect 20735 21732 20791 21788
rect 20791 21732 20795 21788
rect 20731 21728 20795 21732
rect 20811 21788 20875 21792
rect 20811 21732 20815 21788
rect 20815 21732 20871 21788
rect 20871 21732 20875 21788
rect 20811 21728 20875 21732
rect 20891 21788 20955 21792
rect 20891 21732 20895 21788
rect 20895 21732 20951 21788
rect 20951 21732 20955 21788
rect 20891 21728 20955 21732
rect 20971 21788 21035 21792
rect 20971 21732 20975 21788
rect 20975 21732 21031 21788
rect 21031 21732 21035 21788
rect 20971 21728 21035 21732
rect 3004 21660 3068 21724
rect 5580 21660 5644 21724
rect 6684 21660 6748 21724
rect 14228 21524 14292 21588
rect 796 21388 860 21452
rect 3424 21244 3488 21248
rect 3424 21188 3428 21244
rect 3428 21188 3484 21244
rect 3484 21188 3488 21244
rect 3424 21184 3488 21188
rect 3504 21244 3568 21248
rect 3504 21188 3508 21244
rect 3508 21188 3564 21244
rect 3564 21188 3568 21244
rect 3504 21184 3568 21188
rect 3584 21244 3648 21248
rect 3584 21188 3588 21244
rect 3588 21188 3644 21244
rect 3644 21188 3648 21244
rect 3584 21184 3648 21188
rect 3664 21244 3728 21248
rect 3664 21188 3668 21244
rect 3668 21188 3724 21244
rect 3724 21188 3728 21244
rect 3664 21184 3728 21188
rect 8369 21244 8433 21248
rect 8369 21188 8373 21244
rect 8373 21188 8429 21244
rect 8429 21188 8433 21244
rect 8369 21184 8433 21188
rect 8449 21244 8513 21248
rect 8449 21188 8453 21244
rect 8453 21188 8509 21244
rect 8509 21188 8513 21244
rect 8449 21184 8513 21188
rect 8529 21244 8593 21248
rect 8529 21188 8533 21244
rect 8533 21188 8589 21244
rect 8589 21188 8593 21244
rect 8529 21184 8593 21188
rect 8609 21244 8673 21248
rect 8609 21188 8613 21244
rect 8613 21188 8669 21244
rect 8669 21188 8673 21244
rect 8609 21184 8673 21188
rect 13314 21244 13378 21248
rect 13314 21188 13318 21244
rect 13318 21188 13374 21244
rect 13374 21188 13378 21244
rect 13314 21184 13378 21188
rect 13394 21244 13458 21248
rect 13394 21188 13398 21244
rect 13398 21188 13454 21244
rect 13454 21188 13458 21244
rect 13394 21184 13458 21188
rect 13474 21244 13538 21248
rect 13474 21188 13478 21244
rect 13478 21188 13534 21244
rect 13534 21188 13538 21244
rect 13474 21184 13538 21188
rect 13554 21244 13618 21248
rect 13554 21188 13558 21244
rect 13558 21188 13614 21244
rect 13614 21188 13618 21244
rect 13554 21184 13618 21188
rect 2084 21116 2148 21180
rect 5396 21116 5460 21180
rect 12388 20980 12452 21044
rect 18259 21244 18323 21248
rect 18259 21188 18263 21244
rect 18263 21188 18319 21244
rect 18319 21188 18323 21244
rect 18259 21184 18323 21188
rect 18339 21244 18403 21248
rect 18339 21188 18343 21244
rect 18343 21188 18399 21244
rect 18399 21188 18403 21244
rect 18339 21184 18403 21188
rect 18419 21244 18483 21248
rect 18419 21188 18423 21244
rect 18423 21188 18479 21244
rect 18479 21188 18483 21244
rect 18419 21184 18483 21188
rect 18499 21244 18563 21248
rect 18499 21188 18503 21244
rect 18503 21188 18559 21244
rect 18559 21188 18563 21244
rect 18499 21184 18563 21188
rect 15516 21116 15580 21180
rect 16436 21116 16500 21180
rect 6868 20844 6932 20908
rect 7788 20844 7852 20908
rect 13124 20844 13188 20908
rect 19012 20844 19076 20908
rect 4844 20708 4908 20772
rect 6500 20708 6564 20772
rect 6868 20708 6932 20772
rect 7972 20708 8036 20772
rect 14964 20708 15028 20772
rect 16436 20768 16500 20772
rect 16436 20712 16486 20768
rect 16486 20712 16500 20768
rect 16436 20708 16500 20712
rect 5896 20700 5960 20704
rect 5896 20644 5900 20700
rect 5900 20644 5956 20700
rect 5956 20644 5960 20700
rect 5896 20640 5960 20644
rect 5976 20700 6040 20704
rect 5976 20644 5980 20700
rect 5980 20644 6036 20700
rect 6036 20644 6040 20700
rect 5976 20640 6040 20644
rect 6056 20700 6120 20704
rect 6056 20644 6060 20700
rect 6060 20644 6116 20700
rect 6116 20644 6120 20700
rect 6056 20640 6120 20644
rect 6136 20700 6200 20704
rect 6136 20644 6140 20700
rect 6140 20644 6196 20700
rect 6196 20644 6200 20700
rect 6136 20640 6200 20644
rect 10841 20700 10905 20704
rect 10841 20644 10845 20700
rect 10845 20644 10901 20700
rect 10901 20644 10905 20700
rect 10841 20640 10905 20644
rect 10921 20700 10985 20704
rect 10921 20644 10925 20700
rect 10925 20644 10981 20700
rect 10981 20644 10985 20700
rect 10921 20640 10985 20644
rect 11001 20700 11065 20704
rect 11001 20644 11005 20700
rect 11005 20644 11061 20700
rect 11061 20644 11065 20700
rect 11001 20640 11065 20644
rect 11081 20700 11145 20704
rect 11081 20644 11085 20700
rect 11085 20644 11141 20700
rect 11141 20644 11145 20700
rect 11081 20640 11145 20644
rect 15786 20700 15850 20704
rect 15786 20644 15790 20700
rect 15790 20644 15846 20700
rect 15846 20644 15850 20700
rect 15786 20640 15850 20644
rect 15866 20700 15930 20704
rect 15866 20644 15870 20700
rect 15870 20644 15926 20700
rect 15926 20644 15930 20700
rect 15866 20640 15930 20644
rect 15946 20700 16010 20704
rect 15946 20644 15950 20700
rect 15950 20644 16006 20700
rect 16006 20644 16010 20700
rect 15946 20640 16010 20644
rect 16026 20700 16090 20704
rect 16026 20644 16030 20700
rect 16030 20644 16086 20700
rect 16086 20644 16090 20700
rect 16026 20640 16090 20644
rect 20731 20700 20795 20704
rect 20731 20644 20735 20700
rect 20735 20644 20791 20700
rect 20791 20644 20795 20700
rect 20731 20640 20795 20644
rect 20811 20700 20875 20704
rect 20811 20644 20815 20700
rect 20815 20644 20871 20700
rect 20871 20644 20875 20700
rect 20811 20640 20875 20644
rect 20891 20700 20955 20704
rect 20891 20644 20895 20700
rect 20895 20644 20951 20700
rect 20951 20644 20955 20700
rect 20891 20640 20955 20644
rect 20971 20700 21035 20704
rect 20971 20644 20975 20700
rect 20975 20644 21031 20700
rect 21031 20644 21035 20700
rect 20971 20640 21035 20644
rect 18092 20572 18156 20636
rect 5212 20436 5276 20500
rect 5580 20436 5644 20500
rect 12756 20436 12820 20500
rect 14780 20436 14844 20500
rect 8156 20300 8220 20364
rect 3188 20224 3252 20228
rect 3188 20168 3238 20224
rect 3238 20168 3252 20224
rect 3188 20164 3252 20168
rect 10548 20164 10612 20228
rect 14044 20224 14108 20228
rect 14044 20168 14058 20224
rect 14058 20168 14108 20224
rect 14044 20164 14108 20168
rect 3424 20156 3488 20160
rect 3424 20100 3428 20156
rect 3428 20100 3484 20156
rect 3484 20100 3488 20156
rect 3424 20096 3488 20100
rect 3504 20156 3568 20160
rect 3504 20100 3508 20156
rect 3508 20100 3564 20156
rect 3564 20100 3568 20156
rect 3504 20096 3568 20100
rect 3584 20156 3648 20160
rect 3584 20100 3588 20156
rect 3588 20100 3644 20156
rect 3644 20100 3648 20156
rect 3584 20096 3648 20100
rect 3664 20156 3728 20160
rect 3664 20100 3668 20156
rect 3668 20100 3724 20156
rect 3724 20100 3728 20156
rect 3664 20096 3728 20100
rect 8369 20156 8433 20160
rect 8369 20100 8373 20156
rect 8373 20100 8429 20156
rect 8429 20100 8433 20156
rect 8369 20096 8433 20100
rect 8449 20156 8513 20160
rect 8449 20100 8453 20156
rect 8453 20100 8509 20156
rect 8509 20100 8513 20156
rect 8449 20096 8513 20100
rect 8529 20156 8593 20160
rect 8529 20100 8533 20156
rect 8533 20100 8589 20156
rect 8589 20100 8593 20156
rect 8529 20096 8593 20100
rect 8609 20156 8673 20160
rect 8609 20100 8613 20156
rect 8613 20100 8669 20156
rect 8669 20100 8673 20156
rect 8609 20096 8673 20100
rect 13314 20156 13378 20160
rect 13314 20100 13318 20156
rect 13318 20100 13374 20156
rect 13374 20100 13378 20156
rect 13314 20096 13378 20100
rect 13394 20156 13458 20160
rect 13394 20100 13398 20156
rect 13398 20100 13454 20156
rect 13454 20100 13458 20156
rect 13394 20096 13458 20100
rect 13474 20156 13538 20160
rect 13474 20100 13478 20156
rect 13478 20100 13534 20156
rect 13534 20100 13538 20156
rect 13474 20096 13538 20100
rect 13554 20156 13618 20160
rect 13554 20100 13558 20156
rect 13558 20100 13614 20156
rect 13614 20100 13618 20156
rect 13554 20096 13618 20100
rect 18259 20156 18323 20160
rect 18259 20100 18263 20156
rect 18263 20100 18319 20156
rect 18319 20100 18323 20156
rect 18259 20096 18323 20100
rect 18339 20156 18403 20160
rect 18339 20100 18343 20156
rect 18343 20100 18399 20156
rect 18399 20100 18403 20156
rect 18339 20096 18403 20100
rect 18419 20156 18483 20160
rect 18419 20100 18423 20156
rect 18423 20100 18479 20156
rect 18479 20100 18483 20156
rect 18419 20096 18483 20100
rect 18499 20156 18563 20160
rect 18499 20100 18503 20156
rect 18503 20100 18559 20156
rect 18559 20100 18563 20156
rect 18499 20096 18563 20100
rect 2820 20028 2884 20092
rect 5396 20028 5460 20092
rect 12020 19892 12084 19956
rect 13860 19892 13924 19956
rect 17724 19756 17788 19820
rect 8156 19620 8220 19684
rect 5896 19612 5960 19616
rect 5896 19556 5900 19612
rect 5900 19556 5956 19612
rect 5956 19556 5960 19612
rect 5896 19552 5960 19556
rect 5976 19612 6040 19616
rect 5976 19556 5980 19612
rect 5980 19556 6036 19612
rect 6036 19556 6040 19612
rect 5976 19552 6040 19556
rect 6056 19612 6120 19616
rect 6056 19556 6060 19612
rect 6060 19556 6116 19612
rect 6116 19556 6120 19612
rect 6056 19552 6120 19556
rect 6136 19612 6200 19616
rect 6136 19556 6140 19612
rect 6140 19556 6196 19612
rect 6196 19556 6200 19612
rect 6136 19552 6200 19556
rect 10841 19612 10905 19616
rect 10841 19556 10845 19612
rect 10845 19556 10901 19612
rect 10901 19556 10905 19612
rect 10841 19552 10905 19556
rect 10921 19612 10985 19616
rect 10921 19556 10925 19612
rect 10925 19556 10981 19612
rect 10981 19556 10985 19612
rect 10921 19552 10985 19556
rect 11001 19612 11065 19616
rect 11001 19556 11005 19612
rect 11005 19556 11061 19612
rect 11061 19556 11065 19612
rect 11001 19552 11065 19556
rect 11081 19612 11145 19616
rect 11081 19556 11085 19612
rect 11085 19556 11141 19612
rect 11141 19556 11145 19612
rect 11081 19552 11145 19556
rect 15786 19612 15850 19616
rect 15786 19556 15790 19612
rect 15790 19556 15846 19612
rect 15846 19556 15850 19612
rect 15786 19552 15850 19556
rect 15866 19612 15930 19616
rect 15866 19556 15870 19612
rect 15870 19556 15926 19612
rect 15926 19556 15930 19612
rect 15866 19552 15930 19556
rect 15946 19612 16010 19616
rect 15946 19556 15950 19612
rect 15950 19556 16006 19612
rect 16006 19556 16010 19612
rect 15946 19552 16010 19556
rect 16026 19612 16090 19616
rect 16026 19556 16030 19612
rect 16030 19556 16086 19612
rect 16086 19556 16090 19612
rect 16026 19552 16090 19556
rect 20731 19612 20795 19616
rect 20731 19556 20735 19612
rect 20735 19556 20791 19612
rect 20791 19556 20795 19612
rect 20731 19552 20795 19556
rect 20811 19612 20875 19616
rect 20811 19556 20815 19612
rect 20815 19556 20871 19612
rect 20871 19556 20875 19612
rect 20811 19552 20875 19556
rect 20891 19612 20955 19616
rect 20891 19556 20895 19612
rect 20895 19556 20951 19612
rect 20951 19556 20955 19612
rect 20891 19552 20955 19556
rect 20971 19612 21035 19616
rect 20971 19556 20975 19612
rect 20975 19556 21031 19612
rect 21031 19556 21035 19612
rect 20971 19552 21035 19556
rect 3188 19348 3252 19412
rect 3924 19484 3988 19548
rect 9260 19348 9324 19412
rect 10364 19484 10428 19548
rect 11652 19484 11716 19548
rect 11284 19348 11348 19412
rect 10548 19212 10612 19276
rect 3424 19068 3488 19072
rect 3424 19012 3428 19068
rect 3428 19012 3484 19068
rect 3484 19012 3488 19068
rect 3424 19008 3488 19012
rect 3504 19068 3568 19072
rect 3504 19012 3508 19068
rect 3508 19012 3564 19068
rect 3564 19012 3568 19068
rect 3504 19008 3568 19012
rect 3584 19068 3648 19072
rect 3584 19012 3588 19068
rect 3588 19012 3644 19068
rect 3644 19012 3648 19068
rect 3584 19008 3648 19012
rect 3664 19068 3728 19072
rect 3664 19012 3668 19068
rect 3668 19012 3724 19068
rect 3724 19012 3728 19068
rect 3664 19008 3728 19012
rect 8369 19068 8433 19072
rect 8369 19012 8373 19068
rect 8373 19012 8429 19068
rect 8429 19012 8433 19068
rect 8369 19008 8433 19012
rect 8449 19068 8513 19072
rect 8449 19012 8453 19068
rect 8453 19012 8509 19068
rect 8509 19012 8513 19068
rect 8449 19008 8513 19012
rect 8529 19068 8593 19072
rect 8529 19012 8533 19068
rect 8533 19012 8589 19068
rect 8589 19012 8593 19068
rect 8529 19008 8593 19012
rect 8609 19068 8673 19072
rect 8609 19012 8613 19068
rect 8613 19012 8669 19068
rect 8669 19012 8673 19068
rect 8609 19008 8673 19012
rect 13314 19068 13378 19072
rect 13314 19012 13318 19068
rect 13318 19012 13374 19068
rect 13374 19012 13378 19068
rect 13314 19008 13378 19012
rect 13394 19068 13458 19072
rect 13394 19012 13398 19068
rect 13398 19012 13454 19068
rect 13454 19012 13458 19068
rect 13394 19008 13458 19012
rect 13474 19068 13538 19072
rect 13474 19012 13478 19068
rect 13478 19012 13534 19068
rect 13534 19012 13538 19068
rect 13474 19008 13538 19012
rect 13554 19068 13618 19072
rect 13554 19012 13558 19068
rect 13558 19012 13614 19068
rect 13614 19012 13618 19068
rect 13554 19008 13618 19012
rect 18259 19068 18323 19072
rect 18259 19012 18263 19068
rect 18263 19012 18319 19068
rect 18319 19012 18323 19068
rect 18259 19008 18323 19012
rect 18339 19068 18403 19072
rect 18339 19012 18343 19068
rect 18343 19012 18399 19068
rect 18399 19012 18403 19068
rect 18339 19008 18403 19012
rect 18419 19068 18483 19072
rect 18419 19012 18423 19068
rect 18423 19012 18479 19068
rect 18479 19012 18483 19068
rect 18419 19008 18483 19012
rect 18499 19068 18563 19072
rect 18499 19012 18503 19068
rect 18503 19012 18559 19068
rect 18559 19012 18563 19068
rect 18499 19008 18563 19012
rect 12388 19000 12452 19004
rect 12388 18944 12402 19000
rect 12402 18944 12452 19000
rect 12388 18940 12452 18944
rect 6684 18804 6748 18868
rect 7420 18804 7484 18868
rect 7972 18804 8036 18868
rect 9260 18804 9324 18868
rect 14596 18804 14660 18868
rect 11836 18668 11900 18732
rect 5896 18524 5960 18528
rect 5896 18468 5900 18524
rect 5900 18468 5956 18524
rect 5956 18468 5960 18524
rect 5896 18464 5960 18468
rect 5976 18524 6040 18528
rect 5976 18468 5980 18524
rect 5980 18468 6036 18524
rect 6036 18468 6040 18524
rect 5976 18464 6040 18468
rect 6056 18524 6120 18528
rect 6056 18468 6060 18524
rect 6060 18468 6116 18524
rect 6116 18468 6120 18524
rect 6056 18464 6120 18468
rect 6136 18524 6200 18528
rect 6136 18468 6140 18524
rect 6140 18468 6196 18524
rect 6196 18468 6200 18524
rect 6136 18464 6200 18468
rect 10841 18524 10905 18528
rect 10841 18468 10845 18524
rect 10845 18468 10901 18524
rect 10901 18468 10905 18524
rect 10841 18464 10905 18468
rect 10921 18524 10985 18528
rect 10921 18468 10925 18524
rect 10925 18468 10981 18524
rect 10981 18468 10985 18524
rect 10921 18464 10985 18468
rect 11001 18524 11065 18528
rect 11001 18468 11005 18524
rect 11005 18468 11061 18524
rect 11061 18468 11065 18524
rect 11001 18464 11065 18468
rect 11081 18524 11145 18528
rect 11081 18468 11085 18524
rect 11085 18468 11141 18524
rect 11141 18468 11145 18524
rect 11081 18464 11145 18468
rect 15786 18524 15850 18528
rect 15786 18468 15790 18524
rect 15790 18468 15846 18524
rect 15846 18468 15850 18524
rect 15786 18464 15850 18468
rect 15866 18524 15930 18528
rect 15866 18468 15870 18524
rect 15870 18468 15926 18524
rect 15926 18468 15930 18524
rect 15866 18464 15930 18468
rect 15946 18524 16010 18528
rect 15946 18468 15950 18524
rect 15950 18468 16006 18524
rect 16006 18468 16010 18524
rect 15946 18464 16010 18468
rect 16026 18524 16090 18528
rect 16026 18468 16030 18524
rect 16030 18468 16086 18524
rect 16086 18468 16090 18524
rect 16026 18464 16090 18468
rect 20731 18524 20795 18528
rect 20731 18468 20735 18524
rect 20735 18468 20791 18524
rect 20791 18468 20795 18524
rect 20731 18464 20795 18468
rect 20811 18524 20875 18528
rect 20811 18468 20815 18524
rect 20815 18468 20871 18524
rect 20871 18468 20875 18524
rect 20811 18464 20875 18468
rect 20891 18524 20955 18528
rect 20891 18468 20895 18524
rect 20895 18468 20951 18524
rect 20951 18468 20955 18524
rect 20891 18464 20955 18468
rect 20971 18524 21035 18528
rect 20971 18468 20975 18524
rect 20975 18468 21031 18524
rect 21031 18468 21035 18524
rect 20971 18464 21035 18468
rect 2452 18396 2516 18460
rect 2636 18396 2700 18460
rect 3004 18456 3068 18460
rect 3004 18400 3054 18456
rect 3054 18400 3068 18456
rect 3004 18396 3068 18400
rect 5580 18396 5644 18460
rect 14412 18396 14476 18460
rect 2268 18260 2332 18324
rect 796 18184 860 18188
rect 796 18128 810 18184
rect 810 18128 860 18184
rect 796 18124 860 18128
rect 6316 18260 6380 18324
rect 19196 18260 19260 18324
rect 6684 18124 6748 18188
rect 9628 18124 9692 18188
rect 13124 18124 13188 18188
rect 20116 18124 20180 18188
rect 3424 17980 3488 17984
rect 3424 17924 3428 17980
rect 3428 17924 3484 17980
rect 3484 17924 3488 17980
rect 3424 17920 3488 17924
rect 3504 17980 3568 17984
rect 3504 17924 3508 17980
rect 3508 17924 3564 17980
rect 3564 17924 3568 17980
rect 3504 17920 3568 17924
rect 3584 17980 3648 17984
rect 3584 17924 3588 17980
rect 3588 17924 3644 17980
rect 3644 17924 3648 17980
rect 3584 17920 3648 17924
rect 3664 17980 3728 17984
rect 3664 17924 3668 17980
rect 3668 17924 3724 17980
rect 3724 17924 3728 17980
rect 3664 17920 3728 17924
rect 8369 17980 8433 17984
rect 8369 17924 8373 17980
rect 8373 17924 8429 17980
rect 8429 17924 8433 17980
rect 8369 17920 8433 17924
rect 8449 17980 8513 17984
rect 8449 17924 8453 17980
rect 8453 17924 8509 17980
rect 8509 17924 8513 17980
rect 8449 17920 8513 17924
rect 8529 17980 8593 17984
rect 8529 17924 8533 17980
rect 8533 17924 8589 17980
rect 8589 17924 8593 17980
rect 8529 17920 8593 17924
rect 8609 17980 8673 17984
rect 8609 17924 8613 17980
rect 8613 17924 8669 17980
rect 8669 17924 8673 17980
rect 8609 17920 8673 17924
rect 4108 17852 4172 17916
rect 13314 17980 13378 17984
rect 13314 17924 13318 17980
rect 13318 17924 13374 17980
rect 13374 17924 13378 17980
rect 13314 17920 13378 17924
rect 13394 17980 13458 17984
rect 13394 17924 13398 17980
rect 13398 17924 13454 17980
rect 13454 17924 13458 17980
rect 13394 17920 13458 17924
rect 13474 17980 13538 17984
rect 13474 17924 13478 17980
rect 13478 17924 13534 17980
rect 13534 17924 13538 17980
rect 13474 17920 13538 17924
rect 13554 17980 13618 17984
rect 13554 17924 13558 17980
rect 13558 17924 13614 17980
rect 13614 17924 13618 17980
rect 13554 17920 13618 17924
rect 18259 17980 18323 17984
rect 18259 17924 18263 17980
rect 18263 17924 18319 17980
rect 18319 17924 18323 17980
rect 18259 17920 18323 17924
rect 18339 17980 18403 17984
rect 18339 17924 18343 17980
rect 18343 17924 18399 17980
rect 18399 17924 18403 17980
rect 18339 17920 18403 17924
rect 18419 17980 18483 17984
rect 18419 17924 18423 17980
rect 18423 17924 18479 17980
rect 18479 17924 18483 17980
rect 18419 17920 18483 17924
rect 18499 17980 18563 17984
rect 18499 17924 18503 17980
rect 18503 17924 18559 17980
rect 18559 17924 18563 17980
rect 18499 17920 18563 17924
rect 1900 17580 1964 17644
rect 14228 17716 14292 17780
rect 9812 17580 9876 17644
rect 4660 17444 4724 17508
rect 5896 17436 5960 17440
rect 5896 17380 5900 17436
rect 5900 17380 5956 17436
rect 5956 17380 5960 17436
rect 5896 17376 5960 17380
rect 5976 17436 6040 17440
rect 5976 17380 5980 17436
rect 5980 17380 6036 17436
rect 6036 17380 6040 17436
rect 5976 17376 6040 17380
rect 6056 17436 6120 17440
rect 6056 17380 6060 17436
rect 6060 17380 6116 17436
rect 6116 17380 6120 17436
rect 6056 17376 6120 17380
rect 6136 17436 6200 17440
rect 6136 17380 6140 17436
rect 6140 17380 6196 17436
rect 6196 17380 6200 17436
rect 6136 17376 6200 17380
rect 10180 17172 10244 17236
rect 10841 17436 10905 17440
rect 10841 17380 10845 17436
rect 10845 17380 10901 17436
rect 10901 17380 10905 17436
rect 10841 17376 10905 17380
rect 10921 17436 10985 17440
rect 10921 17380 10925 17436
rect 10925 17380 10981 17436
rect 10981 17380 10985 17436
rect 10921 17376 10985 17380
rect 11001 17436 11065 17440
rect 11001 17380 11005 17436
rect 11005 17380 11061 17436
rect 11061 17380 11065 17436
rect 11001 17376 11065 17380
rect 11081 17436 11145 17440
rect 11081 17380 11085 17436
rect 11085 17380 11141 17436
rect 11141 17380 11145 17436
rect 11081 17376 11145 17380
rect 15786 17436 15850 17440
rect 15786 17380 15790 17436
rect 15790 17380 15846 17436
rect 15846 17380 15850 17436
rect 15786 17376 15850 17380
rect 15866 17436 15930 17440
rect 15866 17380 15870 17436
rect 15870 17380 15926 17436
rect 15926 17380 15930 17436
rect 15866 17376 15930 17380
rect 15946 17436 16010 17440
rect 15946 17380 15950 17436
rect 15950 17380 16006 17436
rect 16006 17380 16010 17436
rect 15946 17376 16010 17380
rect 16026 17436 16090 17440
rect 16026 17380 16030 17436
rect 16030 17380 16086 17436
rect 16086 17380 16090 17436
rect 16026 17376 16090 17380
rect 20731 17436 20795 17440
rect 20731 17380 20735 17436
rect 20735 17380 20791 17436
rect 20791 17380 20795 17436
rect 20731 17376 20795 17380
rect 20811 17436 20875 17440
rect 20811 17380 20815 17436
rect 20815 17380 20871 17436
rect 20871 17380 20875 17436
rect 20811 17376 20875 17380
rect 20891 17436 20955 17440
rect 20891 17380 20895 17436
rect 20895 17380 20951 17436
rect 20951 17380 20955 17436
rect 20891 17376 20955 17380
rect 20971 17436 21035 17440
rect 20971 17380 20975 17436
rect 20975 17380 21031 17436
rect 21031 17380 21035 17436
rect 20971 17376 21035 17380
rect 11284 17308 11348 17372
rect 9812 17036 9876 17100
rect 11836 17096 11900 17100
rect 11836 17040 11850 17096
rect 11850 17040 11900 17096
rect 11836 17036 11900 17040
rect 5028 16900 5092 16964
rect 3424 16892 3488 16896
rect 3424 16836 3428 16892
rect 3428 16836 3484 16892
rect 3484 16836 3488 16892
rect 3424 16832 3488 16836
rect 3504 16892 3568 16896
rect 3504 16836 3508 16892
rect 3508 16836 3564 16892
rect 3564 16836 3568 16892
rect 3504 16832 3568 16836
rect 3584 16892 3648 16896
rect 3584 16836 3588 16892
rect 3588 16836 3644 16892
rect 3644 16836 3648 16892
rect 3584 16832 3648 16836
rect 3664 16892 3728 16896
rect 3664 16836 3668 16892
rect 3668 16836 3724 16892
rect 3724 16836 3728 16892
rect 3664 16832 3728 16836
rect 8369 16892 8433 16896
rect 8369 16836 8373 16892
rect 8373 16836 8429 16892
rect 8429 16836 8433 16892
rect 8369 16832 8433 16836
rect 8449 16892 8513 16896
rect 8449 16836 8453 16892
rect 8453 16836 8509 16892
rect 8509 16836 8513 16892
rect 8449 16832 8513 16836
rect 8529 16892 8593 16896
rect 8529 16836 8533 16892
rect 8533 16836 8589 16892
rect 8589 16836 8593 16892
rect 8529 16832 8593 16836
rect 8609 16892 8673 16896
rect 8609 16836 8613 16892
rect 8613 16836 8669 16892
rect 8669 16836 8673 16892
rect 8609 16832 8673 16836
rect 13314 16892 13378 16896
rect 13314 16836 13318 16892
rect 13318 16836 13374 16892
rect 13374 16836 13378 16892
rect 13314 16832 13378 16836
rect 13394 16892 13458 16896
rect 13394 16836 13398 16892
rect 13398 16836 13454 16892
rect 13454 16836 13458 16892
rect 13394 16832 13458 16836
rect 13474 16892 13538 16896
rect 13474 16836 13478 16892
rect 13478 16836 13534 16892
rect 13534 16836 13538 16892
rect 13474 16832 13538 16836
rect 13554 16892 13618 16896
rect 13554 16836 13558 16892
rect 13558 16836 13614 16892
rect 13614 16836 13618 16892
rect 13554 16832 13618 16836
rect 18259 16892 18323 16896
rect 18259 16836 18263 16892
rect 18263 16836 18319 16892
rect 18319 16836 18323 16892
rect 18259 16832 18323 16836
rect 18339 16892 18403 16896
rect 18339 16836 18343 16892
rect 18343 16836 18399 16892
rect 18399 16836 18403 16892
rect 18339 16832 18403 16836
rect 18419 16892 18483 16896
rect 18419 16836 18423 16892
rect 18423 16836 18479 16892
rect 18479 16836 18483 16892
rect 18419 16832 18483 16836
rect 18499 16892 18563 16896
rect 18499 16836 18503 16892
rect 18503 16836 18559 16892
rect 18559 16836 18563 16892
rect 18499 16832 18563 16836
rect 9628 16764 9692 16828
rect 14044 16764 14108 16828
rect 19748 16628 19812 16692
rect 2084 16492 2148 16556
rect 4108 16356 4172 16420
rect 6500 16356 6564 16420
rect 17356 16492 17420 16556
rect 18092 16552 18156 16556
rect 18092 16496 18106 16552
rect 18106 16496 18156 16552
rect 18092 16492 18156 16496
rect 19380 16356 19444 16420
rect 5896 16348 5960 16352
rect 5896 16292 5900 16348
rect 5900 16292 5956 16348
rect 5956 16292 5960 16348
rect 5896 16288 5960 16292
rect 5976 16348 6040 16352
rect 5976 16292 5980 16348
rect 5980 16292 6036 16348
rect 6036 16292 6040 16348
rect 5976 16288 6040 16292
rect 6056 16348 6120 16352
rect 6056 16292 6060 16348
rect 6060 16292 6116 16348
rect 6116 16292 6120 16348
rect 6056 16288 6120 16292
rect 6136 16348 6200 16352
rect 6136 16292 6140 16348
rect 6140 16292 6196 16348
rect 6196 16292 6200 16348
rect 6136 16288 6200 16292
rect 10841 16348 10905 16352
rect 10841 16292 10845 16348
rect 10845 16292 10901 16348
rect 10901 16292 10905 16348
rect 10841 16288 10905 16292
rect 10921 16348 10985 16352
rect 10921 16292 10925 16348
rect 10925 16292 10981 16348
rect 10981 16292 10985 16348
rect 10921 16288 10985 16292
rect 11001 16348 11065 16352
rect 11001 16292 11005 16348
rect 11005 16292 11061 16348
rect 11061 16292 11065 16348
rect 11001 16288 11065 16292
rect 11081 16348 11145 16352
rect 11081 16292 11085 16348
rect 11085 16292 11141 16348
rect 11141 16292 11145 16348
rect 11081 16288 11145 16292
rect 15786 16348 15850 16352
rect 15786 16292 15790 16348
rect 15790 16292 15846 16348
rect 15846 16292 15850 16348
rect 15786 16288 15850 16292
rect 15866 16348 15930 16352
rect 15866 16292 15870 16348
rect 15870 16292 15926 16348
rect 15926 16292 15930 16348
rect 15866 16288 15930 16292
rect 15946 16348 16010 16352
rect 15946 16292 15950 16348
rect 15950 16292 16006 16348
rect 16006 16292 16010 16348
rect 15946 16288 16010 16292
rect 16026 16348 16090 16352
rect 16026 16292 16030 16348
rect 16030 16292 16086 16348
rect 16086 16292 16090 16348
rect 16026 16288 16090 16292
rect 20731 16348 20795 16352
rect 20731 16292 20735 16348
rect 20735 16292 20791 16348
rect 20791 16292 20795 16348
rect 20731 16288 20795 16292
rect 20811 16348 20875 16352
rect 20811 16292 20815 16348
rect 20815 16292 20871 16348
rect 20871 16292 20875 16348
rect 20811 16288 20875 16292
rect 20891 16348 20955 16352
rect 20891 16292 20895 16348
rect 20895 16292 20951 16348
rect 20951 16292 20955 16348
rect 20891 16288 20955 16292
rect 20971 16348 21035 16352
rect 20971 16292 20975 16348
rect 20975 16292 21031 16348
rect 21031 16292 21035 16348
rect 20971 16288 21035 16292
rect 3924 16220 3988 16284
rect 3188 16084 3252 16148
rect 6316 16084 6380 16148
rect 7604 16084 7668 16148
rect 11652 16220 11716 16284
rect 15516 16220 15580 16284
rect 15516 16084 15580 16148
rect 1716 16008 1780 16012
rect 1716 15952 1766 16008
rect 1766 15952 1780 16008
rect 1716 15948 1780 15952
rect 17908 15948 17972 16012
rect 11836 15812 11900 15876
rect 3424 15804 3488 15808
rect 3424 15748 3428 15804
rect 3428 15748 3484 15804
rect 3484 15748 3488 15804
rect 3424 15744 3488 15748
rect 3504 15804 3568 15808
rect 3504 15748 3508 15804
rect 3508 15748 3564 15804
rect 3564 15748 3568 15804
rect 3504 15744 3568 15748
rect 3584 15804 3648 15808
rect 3584 15748 3588 15804
rect 3588 15748 3644 15804
rect 3644 15748 3648 15804
rect 3584 15744 3648 15748
rect 3664 15804 3728 15808
rect 3664 15748 3668 15804
rect 3668 15748 3724 15804
rect 3724 15748 3728 15804
rect 3664 15744 3728 15748
rect 8369 15804 8433 15808
rect 8369 15748 8373 15804
rect 8373 15748 8429 15804
rect 8429 15748 8433 15804
rect 8369 15744 8433 15748
rect 8449 15804 8513 15808
rect 8449 15748 8453 15804
rect 8453 15748 8509 15804
rect 8509 15748 8513 15804
rect 8449 15744 8513 15748
rect 8529 15804 8593 15808
rect 8529 15748 8533 15804
rect 8533 15748 8589 15804
rect 8589 15748 8593 15804
rect 8529 15744 8593 15748
rect 8609 15804 8673 15808
rect 8609 15748 8613 15804
rect 8613 15748 8669 15804
rect 8669 15748 8673 15804
rect 8609 15744 8673 15748
rect 4844 15540 4908 15604
rect 5580 15540 5644 15604
rect 6868 15540 6932 15604
rect 12940 15812 13004 15876
rect 13314 15804 13378 15808
rect 13314 15748 13318 15804
rect 13318 15748 13374 15804
rect 13374 15748 13378 15804
rect 13314 15744 13378 15748
rect 13394 15804 13458 15808
rect 13394 15748 13398 15804
rect 13398 15748 13454 15804
rect 13454 15748 13458 15804
rect 13394 15744 13458 15748
rect 13474 15804 13538 15808
rect 13474 15748 13478 15804
rect 13478 15748 13534 15804
rect 13534 15748 13538 15804
rect 13474 15744 13538 15748
rect 13554 15804 13618 15808
rect 13554 15748 13558 15804
rect 13558 15748 13614 15804
rect 13614 15748 13618 15804
rect 13554 15744 13618 15748
rect 18259 15804 18323 15808
rect 18259 15748 18263 15804
rect 18263 15748 18319 15804
rect 18319 15748 18323 15804
rect 18259 15744 18323 15748
rect 18339 15804 18403 15808
rect 18339 15748 18343 15804
rect 18343 15748 18399 15804
rect 18399 15748 18403 15804
rect 18339 15744 18403 15748
rect 18419 15804 18483 15808
rect 18419 15748 18423 15804
rect 18423 15748 18479 15804
rect 18479 15748 18483 15804
rect 18419 15744 18483 15748
rect 18499 15804 18563 15808
rect 18499 15748 18503 15804
rect 18503 15748 18559 15804
rect 18559 15748 18563 15804
rect 18499 15744 18563 15748
rect 14964 15540 15028 15604
rect 244 15404 308 15468
rect 5580 15328 5644 15332
rect 16804 15404 16868 15468
rect 5580 15272 5594 15328
rect 5594 15272 5644 15328
rect 5580 15268 5644 15272
rect 5896 15260 5960 15264
rect 5896 15204 5900 15260
rect 5900 15204 5956 15260
rect 5956 15204 5960 15260
rect 5896 15200 5960 15204
rect 5976 15260 6040 15264
rect 5976 15204 5980 15260
rect 5980 15204 6036 15260
rect 6036 15204 6040 15260
rect 5976 15200 6040 15204
rect 6056 15260 6120 15264
rect 6056 15204 6060 15260
rect 6060 15204 6116 15260
rect 6116 15204 6120 15260
rect 6056 15200 6120 15204
rect 6136 15260 6200 15264
rect 6136 15204 6140 15260
rect 6140 15204 6196 15260
rect 6196 15204 6200 15260
rect 6136 15200 6200 15204
rect 796 15132 860 15196
rect 6868 15132 6932 15196
rect 10364 15268 10428 15332
rect 10841 15260 10905 15264
rect 10841 15204 10845 15260
rect 10845 15204 10901 15260
rect 10901 15204 10905 15260
rect 10841 15200 10905 15204
rect 10921 15260 10985 15264
rect 10921 15204 10925 15260
rect 10925 15204 10981 15260
rect 10981 15204 10985 15260
rect 10921 15200 10985 15204
rect 11001 15260 11065 15264
rect 11001 15204 11005 15260
rect 11005 15204 11061 15260
rect 11061 15204 11065 15260
rect 11001 15200 11065 15204
rect 11081 15260 11145 15264
rect 11081 15204 11085 15260
rect 11085 15204 11141 15260
rect 11141 15204 11145 15260
rect 11081 15200 11145 15204
rect 15786 15260 15850 15264
rect 15786 15204 15790 15260
rect 15790 15204 15846 15260
rect 15846 15204 15850 15260
rect 15786 15200 15850 15204
rect 15866 15260 15930 15264
rect 15866 15204 15870 15260
rect 15870 15204 15926 15260
rect 15926 15204 15930 15260
rect 15866 15200 15930 15204
rect 15946 15260 16010 15264
rect 15946 15204 15950 15260
rect 15950 15204 16006 15260
rect 16006 15204 16010 15260
rect 15946 15200 16010 15204
rect 16026 15260 16090 15264
rect 16026 15204 16030 15260
rect 16030 15204 16086 15260
rect 16086 15204 16090 15260
rect 16026 15200 16090 15204
rect 20731 15260 20795 15264
rect 20731 15204 20735 15260
rect 20735 15204 20791 15260
rect 20791 15204 20795 15260
rect 20731 15200 20795 15204
rect 20811 15260 20875 15264
rect 20811 15204 20815 15260
rect 20815 15204 20871 15260
rect 20871 15204 20875 15260
rect 20811 15200 20875 15204
rect 20891 15260 20955 15264
rect 20891 15204 20895 15260
rect 20895 15204 20951 15260
rect 20951 15204 20955 15260
rect 20891 15200 20955 15204
rect 20971 15260 21035 15264
rect 20971 15204 20975 15260
rect 20975 15204 21031 15260
rect 21031 15204 21035 15260
rect 20971 15200 21035 15204
rect 18828 15132 18892 15196
rect 12204 15056 12268 15060
rect 12204 15000 12218 15056
rect 12218 15000 12268 15056
rect 12204 14996 12268 15000
rect 13860 14996 13924 15060
rect 16988 14996 17052 15060
rect 17356 14996 17420 15060
rect 18644 14996 18708 15060
rect 1900 14860 1964 14924
rect 5396 14724 5460 14788
rect 18644 14860 18708 14924
rect 3424 14716 3488 14720
rect 3424 14660 3428 14716
rect 3428 14660 3484 14716
rect 3484 14660 3488 14716
rect 3424 14656 3488 14660
rect 3504 14716 3568 14720
rect 3504 14660 3508 14716
rect 3508 14660 3564 14716
rect 3564 14660 3568 14716
rect 3504 14656 3568 14660
rect 3584 14716 3648 14720
rect 3584 14660 3588 14716
rect 3588 14660 3644 14716
rect 3644 14660 3648 14716
rect 3584 14656 3648 14660
rect 3664 14716 3728 14720
rect 3664 14660 3668 14716
rect 3668 14660 3724 14716
rect 3724 14660 3728 14716
rect 3664 14656 3728 14660
rect 8369 14716 8433 14720
rect 8369 14660 8373 14716
rect 8373 14660 8429 14716
rect 8429 14660 8433 14716
rect 8369 14656 8433 14660
rect 8449 14716 8513 14720
rect 8449 14660 8453 14716
rect 8453 14660 8509 14716
rect 8509 14660 8513 14716
rect 8449 14656 8513 14660
rect 8529 14716 8593 14720
rect 8529 14660 8533 14716
rect 8533 14660 8589 14716
rect 8589 14660 8593 14716
rect 8529 14656 8593 14660
rect 8609 14716 8673 14720
rect 8609 14660 8613 14716
rect 8613 14660 8669 14716
rect 8669 14660 8673 14716
rect 8609 14656 8673 14660
rect 2636 14648 2700 14652
rect 2636 14592 2686 14648
rect 2686 14592 2700 14648
rect 2636 14588 2700 14592
rect 3004 14588 3068 14652
rect 5212 14588 5276 14652
rect 13314 14716 13378 14720
rect 13314 14660 13318 14716
rect 13318 14660 13374 14716
rect 13374 14660 13378 14716
rect 13314 14656 13378 14660
rect 13394 14716 13458 14720
rect 13394 14660 13398 14716
rect 13398 14660 13454 14716
rect 13454 14660 13458 14716
rect 13394 14656 13458 14660
rect 13474 14716 13538 14720
rect 13474 14660 13478 14716
rect 13478 14660 13534 14716
rect 13534 14660 13538 14716
rect 13474 14656 13538 14660
rect 13554 14716 13618 14720
rect 13554 14660 13558 14716
rect 13558 14660 13614 14716
rect 13614 14660 13618 14716
rect 13554 14656 13618 14660
rect 612 14512 676 14516
rect 612 14456 626 14512
rect 626 14456 676 14512
rect 612 14452 676 14456
rect 1164 14452 1228 14516
rect 4292 14452 4356 14516
rect 14228 14588 14292 14652
rect 18259 14716 18323 14720
rect 18259 14660 18263 14716
rect 18263 14660 18319 14716
rect 18319 14660 18323 14716
rect 18259 14656 18323 14660
rect 18339 14716 18403 14720
rect 18339 14660 18343 14716
rect 18343 14660 18399 14716
rect 18399 14660 18403 14716
rect 18339 14656 18403 14660
rect 18419 14716 18483 14720
rect 18419 14660 18423 14716
rect 18423 14660 18479 14716
rect 18479 14660 18483 14716
rect 18419 14656 18483 14660
rect 18499 14716 18563 14720
rect 18499 14660 18503 14716
rect 18503 14660 18559 14716
rect 18559 14660 18563 14716
rect 18499 14656 18563 14660
rect 17540 14588 17604 14652
rect 15148 14452 15212 14516
rect 19196 14452 19260 14516
rect 9628 14316 9692 14380
rect 14412 14316 14476 14380
rect 15148 14376 15212 14380
rect 15148 14320 15162 14376
rect 15162 14320 15212 14376
rect 15148 14316 15212 14320
rect 1348 14180 1412 14244
rect 4108 14180 4172 14244
rect 13124 14180 13188 14244
rect 5896 14172 5960 14176
rect 5896 14116 5900 14172
rect 5900 14116 5956 14172
rect 5956 14116 5960 14172
rect 5896 14112 5960 14116
rect 5976 14172 6040 14176
rect 5976 14116 5980 14172
rect 5980 14116 6036 14172
rect 6036 14116 6040 14172
rect 5976 14112 6040 14116
rect 6056 14172 6120 14176
rect 6056 14116 6060 14172
rect 6060 14116 6116 14172
rect 6116 14116 6120 14172
rect 6056 14112 6120 14116
rect 6136 14172 6200 14176
rect 6136 14116 6140 14172
rect 6140 14116 6196 14172
rect 6196 14116 6200 14172
rect 6136 14112 6200 14116
rect 10841 14172 10905 14176
rect 10841 14116 10845 14172
rect 10845 14116 10901 14172
rect 10901 14116 10905 14172
rect 10841 14112 10905 14116
rect 10921 14172 10985 14176
rect 10921 14116 10925 14172
rect 10925 14116 10981 14172
rect 10981 14116 10985 14172
rect 10921 14112 10985 14116
rect 11001 14172 11065 14176
rect 11001 14116 11005 14172
rect 11005 14116 11061 14172
rect 11061 14116 11065 14172
rect 11001 14112 11065 14116
rect 11081 14172 11145 14176
rect 11081 14116 11085 14172
rect 11085 14116 11141 14172
rect 11141 14116 11145 14172
rect 11081 14112 11145 14116
rect 15786 14172 15850 14176
rect 15786 14116 15790 14172
rect 15790 14116 15846 14172
rect 15846 14116 15850 14172
rect 15786 14112 15850 14116
rect 15866 14172 15930 14176
rect 15866 14116 15870 14172
rect 15870 14116 15926 14172
rect 15926 14116 15930 14172
rect 15866 14112 15930 14116
rect 15946 14172 16010 14176
rect 15946 14116 15950 14172
rect 15950 14116 16006 14172
rect 16006 14116 16010 14172
rect 15946 14112 16010 14116
rect 16026 14172 16090 14176
rect 16026 14116 16030 14172
rect 16030 14116 16086 14172
rect 16086 14116 16090 14172
rect 16026 14112 16090 14116
rect 20731 14172 20795 14176
rect 20731 14116 20735 14172
rect 20735 14116 20791 14172
rect 20791 14116 20795 14172
rect 20731 14112 20795 14116
rect 20811 14172 20875 14176
rect 20811 14116 20815 14172
rect 20815 14116 20871 14172
rect 20871 14116 20875 14172
rect 20811 14112 20875 14116
rect 20891 14172 20955 14176
rect 20891 14116 20895 14172
rect 20895 14116 20951 14172
rect 20951 14116 20955 14172
rect 20891 14112 20955 14116
rect 20971 14172 21035 14176
rect 20971 14116 20975 14172
rect 20975 14116 21031 14172
rect 21031 14116 21035 14172
rect 20971 14112 21035 14116
rect 6316 14104 6380 14108
rect 6316 14048 6366 14104
rect 6366 14048 6380 14104
rect 6316 14044 6380 14048
rect 7420 14044 7484 14108
rect 14780 14044 14844 14108
rect 15332 13908 15396 13972
rect 20116 13908 20180 13972
rect 4108 13636 4172 13700
rect 7420 13636 7484 13700
rect 14780 13772 14844 13836
rect 3424 13628 3488 13632
rect 3424 13572 3428 13628
rect 3428 13572 3484 13628
rect 3484 13572 3488 13628
rect 3424 13568 3488 13572
rect 3504 13628 3568 13632
rect 3504 13572 3508 13628
rect 3508 13572 3564 13628
rect 3564 13572 3568 13628
rect 3504 13568 3568 13572
rect 3584 13628 3648 13632
rect 3584 13572 3588 13628
rect 3588 13572 3644 13628
rect 3644 13572 3648 13628
rect 3584 13568 3648 13572
rect 3664 13628 3728 13632
rect 3664 13572 3668 13628
rect 3668 13572 3724 13628
rect 3724 13572 3728 13628
rect 3664 13568 3728 13572
rect 8369 13628 8433 13632
rect 8369 13572 8373 13628
rect 8373 13572 8429 13628
rect 8429 13572 8433 13628
rect 8369 13568 8433 13572
rect 8449 13628 8513 13632
rect 8449 13572 8453 13628
rect 8453 13572 8509 13628
rect 8509 13572 8513 13628
rect 8449 13568 8513 13572
rect 8529 13628 8593 13632
rect 8529 13572 8533 13628
rect 8533 13572 8589 13628
rect 8589 13572 8593 13628
rect 8529 13568 8593 13572
rect 8609 13628 8673 13632
rect 8609 13572 8613 13628
rect 8613 13572 8669 13628
rect 8669 13572 8673 13628
rect 8609 13568 8673 13572
rect 13314 13628 13378 13632
rect 13314 13572 13318 13628
rect 13318 13572 13374 13628
rect 13374 13572 13378 13628
rect 13314 13568 13378 13572
rect 13394 13628 13458 13632
rect 13394 13572 13398 13628
rect 13398 13572 13454 13628
rect 13454 13572 13458 13628
rect 13394 13568 13458 13572
rect 13474 13628 13538 13632
rect 13474 13572 13478 13628
rect 13478 13572 13534 13628
rect 13534 13572 13538 13628
rect 13474 13568 13538 13572
rect 13554 13628 13618 13632
rect 13554 13572 13558 13628
rect 13558 13572 13614 13628
rect 13614 13572 13618 13628
rect 13554 13568 13618 13572
rect 18259 13628 18323 13632
rect 18259 13572 18263 13628
rect 18263 13572 18319 13628
rect 18319 13572 18323 13628
rect 18259 13568 18323 13572
rect 18339 13628 18403 13632
rect 18339 13572 18343 13628
rect 18343 13572 18399 13628
rect 18399 13572 18403 13628
rect 18339 13568 18403 13572
rect 18419 13628 18483 13632
rect 18419 13572 18423 13628
rect 18423 13572 18479 13628
rect 18479 13572 18483 13628
rect 18419 13568 18483 13572
rect 18499 13628 18563 13632
rect 18499 13572 18503 13628
rect 18503 13572 18559 13628
rect 18559 13572 18563 13628
rect 18499 13568 18563 13572
rect 9996 13500 10060 13564
rect 5580 13364 5644 13428
rect 11468 13364 11532 13428
rect 12572 13364 12636 13428
rect 16436 13500 16500 13564
rect 17724 13500 17788 13564
rect 14596 13364 14660 13428
rect 16620 13364 16684 13428
rect 2636 13228 2700 13292
rect 4108 13228 4172 13292
rect 5028 13288 5092 13292
rect 5028 13232 5042 13288
rect 5042 13232 5092 13288
rect 5028 13228 5092 13232
rect 16252 13228 16316 13292
rect 10364 13152 10428 13156
rect 10364 13096 10414 13152
rect 10414 13096 10428 13152
rect 10364 13092 10428 13096
rect 14412 13092 14476 13156
rect 15148 13152 15212 13156
rect 15148 13096 15162 13152
rect 15162 13096 15212 13152
rect 15148 13092 15212 13096
rect 15516 13092 15580 13156
rect 5896 13084 5960 13088
rect 5896 13028 5900 13084
rect 5900 13028 5956 13084
rect 5956 13028 5960 13084
rect 5896 13024 5960 13028
rect 5976 13084 6040 13088
rect 5976 13028 5980 13084
rect 5980 13028 6036 13084
rect 6036 13028 6040 13084
rect 5976 13024 6040 13028
rect 6056 13084 6120 13088
rect 6056 13028 6060 13084
rect 6060 13028 6116 13084
rect 6116 13028 6120 13084
rect 6056 13024 6120 13028
rect 6136 13084 6200 13088
rect 6136 13028 6140 13084
rect 6140 13028 6196 13084
rect 6196 13028 6200 13084
rect 6136 13024 6200 13028
rect 10841 13084 10905 13088
rect 10841 13028 10845 13084
rect 10845 13028 10901 13084
rect 10901 13028 10905 13084
rect 10841 13024 10905 13028
rect 10921 13084 10985 13088
rect 10921 13028 10925 13084
rect 10925 13028 10981 13084
rect 10981 13028 10985 13084
rect 10921 13024 10985 13028
rect 11001 13084 11065 13088
rect 11001 13028 11005 13084
rect 11005 13028 11061 13084
rect 11061 13028 11065 13084
rect 11001 13024 11065 13028
rect 11081 13084 11145 13088
rect 11081 13028 11085 13084
rect 11085 13028 11141 13084
rect 11141 13028 11145 13084
rect 11081 13024 11145 13028
rect 4844 12956 4908 13020
rect 15786 13084 15850 13088
rect 15786 13028 15790 13084
rect 15790 13028 15846 13084
rect 15846 13028 15850 13084
rect 15786 13024 15850 13028
rect 15866 13084 15930 13088
rect 15866 13028 15870 13084
rect 15870 13028 15926 13084
rect 15926 13028 15930 13084
rect 15866 13024 15930 13028
rect 15946 13084 16010 13088
rect 15946 13028 15950 13084
rect 15950 13028 16006 13084
rect 16006 13028 16010 13084
rect 15946 13024 16010 13028
rect 16026 13084 16090 13088
rect 16026 13028 16030 13084
rect 16030 13028 16086 13084
rect 16086 13028 16090 13084
rect 16026 13024 16090 13028
rect 20731 13084 20795 13088
rect 20731 13028 20735 13084
rect 20735 13028 20791 13084
rect 20791 13028 20795 13084
rect 20731 13024 20795 13028
rect 20811 13084 20875 13088
rect 20811 13028 20815 13084
rect 20815 13028 20871 13084
rect 20871 13028 20875 13084
rect 20811 13024 20875 13028
rect 20891 13084 20955 13088
rect 20891 13028 20895 13084
rect 20895 13028 20951 13084
rect 20951 13028 20955 13084
rect 20891 13024 20955 13028
rect 20971 13084 21035 13088
rect 20971 13028 20975 13084
rect 20975 13028 21031 13084
rect 21031 13028 21035 13084
rect 20971 13024 21035 13028
rect 2268 12684 2332 12748
rect 5396 12548 5460 12612
rect 3424 12540 3488 12544
rect 3424 12484 3428 12540
rect 3428 12484 3484 12540
rect 3484 12484 3488 12540
rect 3424 12480 3488 12484
rect 3504 12540 3568 12544
rect 3504 12484 3508 12540
rect 3508 12484 3564 12540
rect 3564 12484 3568 12540
rect 3504 12480 3568 12484
rect 3584 12540 3648 12544
rect 3584 12484 3588 12540
rect 3588 12484 3644 12540
rect 3644 12484 3648 12540
rect 3584 12480 3648 12484
rect 3664 12540 3728 12544
rect 3664 12484 3668 12540
rect 3668 12484 3724 12540
rect 3724 12484 3728 12540
rect 3664 12480 3728 12484
rect 8369 12540 8433 12544
rect 8369 12484 8373 12540
rect 8373 12484 8429 12540
rect 8429 12484 8433 12540
rect 8369 12480 8433 12484
rect 8449 12540 8513 12544
rect 8449 12484 8453 12540
rect 8453 12484 8509 12540
rect 8509 12484 8513 12540
rect 8449 12480 8513 12484
rect 8529 12540 8593 12544
rect 8529 12484 8533 12540
rect 8533 12484 8589 12540
rect 8589 12484 8593 12540
rect 8529 12480 8593 12484
rect 8609 12540 8673 12544
rect 8609 12484 8613 12540
rect 8613 12484 8669 12540
rect 8669 12484 8673 12540
rect 8609 12480 8673 12484
rect 5718 12412 5782 12476
rect 5580 12276 5644 12340
rect 16804 12684 16868 12748
rect 13314 12540 13378 12544
rect 13314 12484 13318 12540
rect 13318 12484 13374 12540
rect 13374 12484 13378 12540
rect 13314 12480 13378 12484
rect 13394 12540 13458 12544
rect 13394 12484 13398 12540
rect 13398 12484 13454 12540
rect 13454 12484 13458 12540
rect 13394 12480 13458 12484
rect 13474 12540 13538 12544
rect 13474 12484 13478 12540
rect 13478 12484 13534 12540
rect 13534 12484 13538 12540
rect 13474 12480 13538 12484
rect 13554 12540 13618 12544
rect 13554 12484 13558 12540
rect 13558 12484 13614 12540
rect 13614 12484 13618 12540
rect 13554 12480 13618 12484
rect 16252 12472 16316 12476
rect 20300 12684 20364 12748
rect 18259 12540 18323 12544
rect 18259 12484 18263 12540
rect 18263 12484 18319 12540
rect 18319 12484 18323 12540
rect 18259 12480 18323 12484
rect 18339 12540 18403 12544
rect 18339 12484 18343 12540
rect 18343 12484 18399 12540
rect 18399 12484 18403 12540
rect 18339 12480 18403 12484
rect 18419 12540 18483 12544
rect 18419 12484 18423 12540
rect 18423 12484 18479 12540
rect 18479 12484 18483 12540
rect 18419 12480 18483 12484
rect 18499 12540 18563 12544
rect 18499 12484 18503 12540
rect 18503 12484 18559 12540
rect 18559 12484 18563 12540
rect 18499 12480 18563 12484
rect 16252 12416 16302 12472
rect 16302 12416 16316 12472
rect 16252 12412 16316 12416
rect 17540 12276 17604 12340
rect 4844 12004 4908 12068
rect 7604 12004 7668 12068
rect 11468 12004 11532 12068
rect 13860 12004 13924 12068
rect 14412 12004 14476 12068
rect 19564 12004 19628 12068
rect 5896 11996 5960 12000
rect 5896 11940 5900 11996
rect 5900 11940 5956 11996
rect 5956 11940 5960 11996
rect 5896 11936 5960 11940
rect 5976 11996 6040 12000
rect 5976 11940 5980 11996
rect 5980 11940 6036 11996
rect 6036 11940 6040 11996
rect 5976 11936 6040 11940
rect 6056 11996 6120 12000
rect 6056 11940 6060 11996
rect 6060 11940 6116 11996
rect 6116 11940 6120 11996
rect 6056 11936 6120 11940
rect 6136 11996 6200 12000
rect 6136 11940 6140 11996
rect 6140 11940 6196 11996
rect 6196 11940 6200 11996
rect 6136 11936 6200 11940
rect 10841 11996 10905 12000
rect 10841 11940 10845 11996
rect 10845 11940 10901 11996
rect 10901 11940 10905 11996
rect 10841 11936 10905 11940
rect 10921 11996 10985 12000
rect 10921 11940 10925 11996
rect 10925 11940 10981 11996
rect 10981 11940 10985 11996
rect 10921 11936 10985 11940
rect 11001 11996 11065 12000
rect 11001 11940 11005 11996
rect 11005 11940 11061 11996
rect 11061 11940 11065 11996
rect 11001 11936 11065 11940
rect 11081 11996 11145 12000
rect 11081 11940 11085 11996
rect 11085 11940 11141 11996
rect 11141 11940 11145 11996
rect 11081 11936 11145 11940
rect 15786 11996 15850 12000
rect 15786 11940 15790 11996
rect 15790 11940 15846 11996
rect 15846 11940 15850 11996
rect 15786 11936 15850 11940
rect 15866 11996 15930 12000
rect 15866 11940 15870 11996
rect 15870 11940 15926 11996
rect 15926 11940 15930 11996
rect 15866 11936 15930 11940
rect 15946 11996 16010 12000
rect 15946 11940 15950 11996
rect 15950 11940 16006 11996
rect 16006 11940 16010 11996
rect 15946 11936 16010 11940
rect 16026 11996 16090 12000
rect 16026 11940 16030 11996
rect 16030 11940 16086 11996
rect 16086 11940 16090 11996
rect 16026 11936 16090 11940
rect 20731 11996 20795 12000
rect 20731 11940 20735 11996
rect 20735 11940 20791 11996
rect 20791 11940 20795 11996
rect 20731 11936 20795 11940
rect 20811 11996 20875 12000
rect 20811 11940 20815 11996
rect 20815 11940 20871 11996
rect 20871 11940 20875 11996
rect 20811 11936 20875 11940
rect 20891 11996 20955 12000
rect 20891 11940 20895 11996
rect 20895 11940 20951 11996
rect 20951 11940 20955 11996
rect 20891 11936 20955 11940
rect 20971 11996 21035 12000
rect 20971 11940 20975 11996
rect 20975 11940 21031 11996
rect 21031 11940 21035 11996
rect 20971 11936 21035 11940
rect 2452 11732 2516 11796
rect 5396 11732 5460 11796
rect 6868 11792 6932 11796
rect 6868 11736 6882 11792
rect 6882 11736 6932 11792
rect 6868 11732 6932 11736
rect 14228 11868 14292 11932
rect 17172 11868 17236 11932
rect 7420 11596 7484 11660
rect 4292 11460 4356 11524
rect 14964 11732 15028 11796
rect 15332 11792 15396 11796
rect 15332 11736 15382 11792
rect 15382 11736 15396 11792
rect 15332 11732 15396 11736
rect 15516 11732 15580 11796
rect 3424 11452 3488 11456
rect 3424 11396 3428 11452
rect 3428 11396 3484 11452
rect 3484 11396 3488 11452
rect 3424 11392 3488 11396
rect 3504 11452 3568 11456
rect 3504 11396 3508 11452
rect 3508 11396 3564 11452
rect 3564 11396 3568 11452
rect 3504 11392 3568 11396
rect 3584 11452 3648 11456
rect 3584 11396 3588 11452
rect 3588 11396 3644 11452
rect 3644 11396 3648 11452
rect 3584 11392 3648 11396
rect 3664 11452 3728 11456
rect 3664 11396 3668 11452
rect 3668 11396 3724 11452
rect 3724 11396 3728 11452
rect 3664 11392 3728 11396
rect 16252 11460 16316 11524
rect 16620 11460 16684 11524
rect 8369 11452 8433 11456
rect 8369 11396 8373 11452
rect 8373 11396 8429 11452
rect 8429 11396 8433 11452
rect 8369 11392 8433 11396
rect 8449 11452 8513 11456
rect 8449 11396 8453 11452
rect 8453 11396 8509 11452
rect 8509 11396 8513 11452
rect 8449 11392 8513 11396
rect 8529 11452 8593 11456
rect 8529 11396 8533 11452
rect 8533 11396 8589 11452
rect 8589 11396 8593 11452
rect 8529 11392 8593 11396
rect 8609 11452 8673 11456
rect 8609 11396 8613 11452
rect 8613 11396 8669 11452
rect 8669 11396 8673 11452
rect 8609 11392 8673 11396
rect 13314 11452 13378 11456
rect 13314 11396 13318 11452
rect 13318 11396 13374 11452
rect 13374 11396 13378 11452
rect 13314 11392 13378 11396
rect 13394 11452 13458 11456
rect 13394 11396 13398 11452
rect 13398 11396 13454 11452
rect 13454 11396 13458 11452
rect 13394 11392 13458 11396
rect 13474 11452 13538 11456
rect 13474 11396 13478 11452
rect 13478 11396 13534 11452
rect 13534 11396 13538 11452
rect 13474 11392 13538 11396
rect 13554 11452 13618 11456
rect 13554 11396 13558 11452
rect 13558 11396 13614 11452
rect 13614 11396 13618 11452
rect 13554 11392 13618 11396
rect 18259 11452 18323 11456
rect 18259 11396 18263 11452
rect 18263 11396 18319 11452
rect 18319 11396 18323 11452
rect 18259 11392 18323 11396
rect 18339 11452 18403 11456
rect 18339 11396 18343 11452
rect 18343 11396 18399 11452
rect 18399 11396 18403 11452
rect 18339 11392 18403 11396
rect 18419 11452 18483 11456
rect 18419 11396 18423 11452
rect 18423 11396 18479 11452
rect 18479 11396 18483 11452
rect 18419 11392 18483 11396
rect 18499 11452 18563 11456
rect 18499 11396 18503 11452
rect 18503 11396 18559 11452
rect 18559 11396 18563 11452
rect 18499 11392 18563 11396
rect 8754 11324 8818 11388
rect 2268 11052 2332 11116
rect 2452 11112 2516 11116
rect 2452 11056 2502 11112
rect 2502 11056 2516 11112
rect 2452 11052 2516 11056
rect 4844 11112 4908 11116
rect 4844 11056 4858 11112
rect 4858 11056 4908 11112
rect 4844 11052 4908 11056
rect 1532 10916 1596 10980
rect 4292 10916 4356 10980
rect 4844 10976 4908 10980
rect 4844 10920 4894 10976
rect 4894 10920 4908 10976
rect 4844 10916 4908 10920
rect 12020 11188 12084 11252
rect 6868 11052 6932 11116
rect 5896 10908 5960 10912
rect 5896 10852 5900 10908
rect 5900 10852 5956 10908
rect 5956 10852 5960 10908
rect 5896 10848 5960 10852
rect 5976 10908 6040 10912
rect 5976 10852 5980 10908
rect 5980 10852 6036 10908
rect 6036 10852 6040 10908
rect 5976 10848 6040 10852
rect 6056 10908 6120 10912
rect 6056 10852 6060 10908
rect 6060 10852 6116 10908
rect 6116 10852 6120 10908
rect 6056 10848 6120 10852
rect 6136 10908 6200 10912
rect 6136 10852 6140 10908
rect 6140 10852 6196 10908
rect 6196 10852 6200 10908
rect 6136 10848 6200 10852
rect 10841 10908 10905 10912
rect 10841 10852 10845 10908
rect 10845 10852 10901 10908
rect 10901 10852 10905 10908
rect 10841 10848 10905 10852
rect 10921 10908 10985 10912
rect 10921 10852 10925 10908
rect 10925 10852 10981 10908
rect 10981 10852 10985 10908
rect 10921 10848 10985 10852
rect 11001 10908 11065 10912
rect 11001 10852 11005 10908
rect 11005 10852 11061 10908
rect 11061 10852 11065 10908
rect 11001 10848 11065 10852
rect 11081 10908 11145 10912
rect 11081 10852 11085 10908
rect 11085 10852 11141 10908
rect 11141 10852 11145 10908
rect 11081 10848 11145 10852
rect 18828 10976 18892 10980
rect 18828 10920 18842 10976
rect 18842 10920 18892 10976
rect 18828 10916 18892 10920
rect 15786 10908 15850 10912
rect 15786 10852 15790 10908
rect 15790 10852 15846 10908
rect 15846 10852 15850 10908
rect 15786 10848 15850 10852
rect 15866 10908 15930 10912
rect 15866 10852 15870 10908
rect 15870 10852 15926 10908
rect 15926 10852 15930 10908
rect 15866 10848 15930 10852
rect 15946 10908 16010 10912
rect 15946 10852 15950 10908
rect 15950 10852 16006 10908
rect 16006 10852 16010 10908
rect 15946 10848 16010 10852
rect 16026 10908 16090 10912
rect 16026 10852 16030 10908
rect 16030 10852 16086 10908
rect 16086 10852 16090 10908
rect 16026 10848 16090 10852
rect 20731 10908 20795 10912
rect 20731 10852 20735 10908
rect 20735 10852 20791 10908
rect 20791 10852 20795 10908
rect 20731 10848 20795 10852
rect 20811 10908 20875 10912
rect 20811 10852 20815 10908
rect 20815 10852 20871 10908
rect 20871 10852 20875 10908
rect 20811 10848 20875 10852
rect 20891 10908 20955 10912
rect 20891 10852 20895 10908
rect 20895 10852 20951 10908
rect 20951 10852 20955 10908
rect 20891 10848 20955 10852
rect 20971 10908 21035 10912
rect 20971 10852 20975 10908
rect 20975 10852 21031 10908
rect 21031 10852 21035 10908
rect 20971 10848 21035 10852
rect 11652 10840 11716 10844
rect 11652 10784 11666 10840
rect 11666 10784 11716 10840
rect 11652 10780 11716 10784
rect 13860 10780 13924 10844
rect 2268 10644 2332 10708
rect 3004 10644 3068 10708
rect 3924 10704 3988 10708
rect 3924 10648 3974 10704
rect 3974 10648 3988 10704
rect 3924 10644 3988 10648
rect 5028 10644 5092 10708
rect 11468 10644 11532 10708
rect 17540 10644 17604 10708
rect 3004 10508 3068 10572
rect 11836 10508 11900 10572
rect 14044 10508 14108 10572
rect 14412 10508 14476 10572
rect 15516 10508 15580 10572
rect 5580 10432 5644 10436
rect 5580 10376 5594 10432
rect 5594 10376 5644 10432
rect 5580 10372 5644 10376
rect 7972 10432 8036 10436
rect 7972 10376 8022 10432
rect 8022 10376 8036 10432
rect 7972 10372 8036 10376
rect 8892 10372 8956 10436
rect 3424 10364 3488 10368
rect 3424 10308 3428 10364
rect 3428 10308 3484 10364
rect 3484 10308 3488 10364
rect 3424 10304 3488 10308
rect 3504 10364 3568 10368
rect 3504 10308 3508 10364
rect 3508 10308 3564 10364
rect 3564 10308 3568 10364
rect 3504 10304 3568 10308
rect 3584 10364 3648 10368
rect 3584 10308 3588 10364
rect 3588 10308 3644 10364
rect 3644 10308 3648 10364
rect 3584 10304 3648 10308
rect 3664 10364 3728 10368
rect 3664 10308 3668 10364
rect 3668 10308 3724 10364
rect 3724 10308 3728 10364
rect 3664 10304 3728 10308
rect 8369 10364 8433 10368
rect 8369 10308 8373 10364
rect 8373 10308 8429 10364
rect 8429 10308 8433 10364
rect 8369 10304 8433 10308
rect 8449 10364 8513 10368
rect 8449 10308 8453 10364
rect 8453 10308 8509 10364
rect 8509 10308 8513 10364
rect 8449 10304 8513 10308
rect 8529 10364 8593 10368
rect 8529 10308 8533 10364
rect 8533 10308 8589 10364
rect 8589 10308 8593 10364
rect 8529 10304 8593 10308
rect 8609 10364 8673 10368
rect 8609 10308 8613 10364
rect 8613 10308 8669 10364
rect 8669 10308 8673 10364
rect 8609 10304 8673 10308
rect 2636 10296 2700 10300
rect 2636 10240 2650 10296
rect 2650 10240 2700 10296
rect 2636 10236 2700 10240
rect 4108 10236 4172 10300
rect 5396 10236 5460 10300
rect 1900 9964 1964 10028
rect 7972 9964 8036 10028
rect 8892 10236 8956 10300
rect 9076 10236 9140 10300
rect 9444 10372 9508 10436
rect 10686 10372 10750 10436
rect 11468 10372 11532 10436
rect 13314 10364 13378 10368
rect 13314 10308 13318 10364
rect 13318 10308 13374 10364
rect 13374 10308 13378 10364
rect 13314 10304 13378 10308
rect 13394 10364 13458 10368
rect 13394 10308 13398 10364
rect 13398 10308 13454 10364
rect 13454 10308 13458 10364
rect 13394 10304 13458 10308
rect 13474 10364 13538 10368
rect 13474 10308 13478 10364
rect 13478 10308 13534 10364
rect 13534 10308 13538 10364
rect 13474 10304 13538 10308
rect 13554 10364 13618 10368
rect 13554 10308 13558 10364
rect 13558 10308 13614 10364
rect 13614 10308 13618 10364
rect 13554 10304 13618 10308
rect 9444 10236 9508 10300
rect 12756 10236 12820 10300
rect 14412 10160 14476 10164
rect 14412 10104 14462 10160
rect 14462 10104 14476 10160
rect 14412 10100 14476 10104
rect 17172 10100 17236 10164
rect 18259 10364 18323 10368
rect 18259 10308 18263 10364
rect 18263 10308 18319 10364
rect 18319 10308 18323 10364
rect 18259 10304 18323 10308
rect 18339 10364 18403 10368
rect 18339 10308 18343 10364
rect 18343 10308 18399 10364
rect 18399 10308 18403 10364
rect 18339 10304 18403 10308
rect 18419 10364 18483 10368
rect 18419 10308 18423 10364
rect 18423 10308 18479 10364
rect 18479 10308 18483 10364
rect 18419 10304 18483 10308
rect 18499 10364 18563 10368
rect 18499 10308 18503 10364
rect 18503 10308 18559 10364
rect 18559 10308 18563 10364
rect 18499 10304 18563 10308
rect 18828 10100 18892 10164
rect 17908 10024 17972 10028
rect 17908 9968 17922 10024
rect 17922 9968 17972 10024
rect 17908 9964 17972 9968
rect 18092 9964 18156 10028
rect 5896 9820 5960 9824
rect 5896 9764 5900 9820
rect 5900 9764 5956 9820
rect 5956 9764 5960 9820
rect 5896 9760 5960 9764
rect 5976 9820 6040 9824
rect 5976 9764 5980 9820
rect 5980 9764 6036 9820
rect 6036 9764 6040 9820
rect 5976 9760 6040 9764
rect 6056 9820 6120 9824
rect 6056 9764 6060 9820
rect 6060 9764 6116 9820
rect 6116 9764 6120 9820
rect 6056 9760 6120 9764
rect 6136 9820 6200 9824
rect 6136 9764 6140 9820
rect 6140 9764 6196 9820
rect 6196 9764 6200 9820
rect 6136 9760 6200 9764
rect 12756 9888 12820 9892
rect 12756 9832 12806 9888
rect 12806 9832 12820 9888
rect 12756 9828 12820 9832
rect 10841 9820 10905 9824
rect 10841 9764 10845 9820
rect 10845 9764 10901 9820
rect 10901 9764 10905 9820
rect 10841 9760 10905 9764
rect 10921 9820 10985 9824
rect 10921 9764 10925 9820
rect 10925 9764 10981 9820
rect 10981 9764 10985 9820
rect 10921 9760 10985 9764
rect 11001 9820 11065 9824
rect 11001 9764 11005 9820
rect 11005 9764 11061 9820
rect 11061 9764 11065 9820
rect 11001 9760 11065 9764
rect 11081 9820 11145 9824
rect 11081 9764 11085 9820
rect 11085 9764 11141 9820
rect 11141 9764 11145 9820
rect 11081 9760 11145 9764
rect 15786 9820 15850 9824
rect 15786 9764 15790 9820
rect 15790 9764 15846 9820
rect 15846 9764 15850 9820
rect 15786 9760 15850 9764
rect 15866 9820 15930 9824
rect 15866 9764 15870 9820
rect 15870 9764 15926 9820
rect 15926 9764 15930 9820
rect 15866 9760 15930 9764
rect 15946 9820 16010 9824
rect 15946 9764 15950 9820
rect 15950 9764 16006 9820
rect 16006 9764 16010 9820
rect 15946 9760 16010 9764
rect 16026 9820 16090 9824
rect 16026 9764 16030 9820
rect 16030 9764 16086 9820
rect 16086 9764 16090 9820
rect 16026 9760 16090 9764
rect 20731 9820 20795 9824
rect 20731 9764 20735 9820
rect 20735 9764 20791 9820
rect 20791 9764 20795 9820
rect 20731 9760 20795 9764
rect 20811 9820 20875 9824
rect 20811 9764 20815 9820
rect 20815 9764 20871 9820
rect 20871 9764 20875 9820
rect 20811 9760 20875 9764
rect 20891 9820 20955 9824
rect 20891 9764 20895 9820
rect 20895 9764 20951 9820
rect 20951 9764 20955 9820
rect 20891 9760 20955 9764
rect 20971 9820 21035 9824
rect 20971 9764 20975 9820
rect 20975 9764 21031 9820
rect 21031 9764 21035 9820
rect 20971 9760 21035 9764
rect 8156 9752 8220 9756
rect 8156 9696 8170 9752
rect 8170 9696 8220 9752
rect 8156 9692 8220 9696
rect 11652 9692 11716 9756
rect 2636 9556 2700 9620
rect 1348 9420 1412 9484
rect 4476 9556 4540 9620
rect 3188 9420 3252 9484
rect 2820 9284 2884 9348
rect 5028 9480 5092 9484
rect 5028 9424 5078 9480
rect 5078 9424 5092 9480
rect 5028 9420 5092 9424
rect 7788 9420 7852 9484
rect 5028 9284 5092 9348
rect 15148 9420 15212 9484
rect 10364 9284 10428 9348
rect 12940 9284 13004 9348
rect 3424 9276 3488 9280
rect 3424 9220 3428 9276
rect 3428 9220 3484 9276
rect 3484 9220 3488 9276
rect 3424 9216 3488 9220
rect 3504 9276 3568 9280
rect 3504 9220 3508 9276
rect 3508 9220 3564 9276
rect 3564 9220 3568 9276
rect 3504 9216 3568 9220
rect 3584 9276 3648 9280
rect 3584 9220 3588 9276
rect 3588 9220 3644 9276
rect 3644 9220 3648 9276
rect 3584 9216 3648 9220
rect 3664 9276 3728 9280
rect 3664 9220 3668 9276
rect 3668 9220 3724 9276
rect 3724 9220 3728 9276
rect 3664 9216 3728 9220
rect 8369 9276 8433 9280
rect 8369 9220 8373 9276
rect 8373 9220 8429 9276
rect 8429 9220 8433 9276
rect 8369 9216 8433 9220
rect 8449 9276 8513 9280
rect 8449 9220 8453 9276
rect 8453 9220 8509 9276
rect 8509 9220 8513 9276
rect 8449 9216 8513 9220
rect 8529 9276 8593 9280
rect 8529 9220 8533 9276
rect 8533 9220 8589 9276
rect 8589 9220 8593 9276
rect 8529 9216 8593 9220
rect 8609 9276 8673 9280
rect 8609 9220 8613 9276
rect 8613 9220 8669 9276
rect 8669 9220 8673 9276
rect 8609 9216 8673 9220
rect 8156 9208 8220 9212
rect 8156 9152 8206 9208
rect 8206 9152 8220 9208
rect 8156 9148 8220 9152
rect 8892 9148 8956 9212
rect 12204 9148 12268 9212
rect 1900 9012 1964 9076
rect 2268 9012 2332 9076
rect 4108 9012 4172 9076
rect 1716 8876 1780 8940
rect 2268 8876 2332 8940
rect 2636 8876 2700 8940
rect 5396 9012 5460 9076
rect 9812 9012 9876 9076
rect 10364 9012 10428 9076
rect 16804 9284 16868 9348
rect 18092 9284 18156 9348
rect 19380 9344 19444 9348
rect 19380 9288 19394 9344
rect 19394 9288 19444 9344
rect 19380 9284 19444 9288
rect 13314 9276 13378 9280
rect 13314 9220 13318 9276
rect 13318 9220 13374 9276
rect 13374 9220 13378 9276
rect 13314 9216 13378 9220
rect 13394 9276 13458 9280
rect 13394 9220 13398 9276
rect 13398 9220 13454 9276
rect 13454 9220 13458 9276
rect 13394 9216 13458 9220
rect 13474 9276 13538 9280
rect 13474 9220 13478 9276
rect 13478 9220 13534 9276
rect 13534 9220 13538 9276
rect 13474 9216 13538 9220
rect 13554 9276 13618 9280
rect 13554 9220 13558 9276
rect 13558 9220 13614 9276
rect 13614 9220 13618 9276
rect 13554 9216 13618 9220
rect 18259 9276 18323 9280
rect 18259 9220 18263 9276
rect 18263 9220 18319 9276
rect 18319 9220 18323 9276
rect 18259 9216 18323 9220
rect 18339 9276 18403 9280
rect 18339 9220 18343 9276
rect 18343 9220 18399 9276
rect 18399 9220 18403 9276
rect 18339 9216 18403 9220
rect 18419 9276 18483 9280
rect 18419 9220 18423 9276
rect 18423 9220 18479 9276
rect 18479 9220 18483 9276
rect 18419 9216 18483 9220
rect 18499 9276 18563 9280
rect 18499 9220 18503 9276
rect 18503 9220 18559 9276
rect 18559 9220 18563 9276
rect 18499 9216 18563 9220
rect 14964 9208 15028 9212
rect 14964 9152 14978 9208
rect 14978 9152 15028 9208
rect 14964 9148 15028 9152
rect 18828 9148 18892 9212
rect 20300 9148 20364 9212
rect 4476 8876 4540 8940
rect 19932 9012 19996 9076
rect 7788 8740 7852 8804
rect 10364 8740 10428 8804
rect 10548 8740 10612 8804
rect 5896 8732 5960 8736
rect 5896 8676 5900 8732
rect 5900 8676 5956 8732
rect 5956 8676 5960 8732
rect 5896 8672 5960 8676
rect 5976 8732 6040 8736
rect 5976 8676 5980 8732
rect 5980 8676 6036 8732
rect 6036 8676 6040 8732
rect 5976 8672 6040 8676
rect 6056 8732 6120 8736
rect 6056 8676 6060 8732
rect 6060 8676 6116 8732
rect 6116 8676 6120 8732
rect 6056 8672 6120 8676
rect 6136 8732 6200 8736
rect 6136 8676 6140 8732
rect 6140 8676 6196 8732
rect 6196 8676 6200 8732
rect 6136 8672 6200 8676
rect 12388 8740 12452 8804
rect 13860 8740 13924 8804
rect 16988 8876 17052 8940
rect 10841 8732 10905 8736
rect 10841 8676 10845 8732
rect 10845 8676 10901 8732
rect 10901 8676 10905 8732
rect 10841 8672 10905 8676
rect 10921 8732 10985 8736
rect 10921 8676 10925 8732
rect 10925 8676 10981 8732
rect 10981 8676 10985 8732
rect 10921 8672 10985 8676
rect 11001 8732 11065 8736
rect 11001 8676 11005 8732
rect 11005 8676 11061 8732
rect 11061 8676 11065 8732
rect 11001 8672 11065 8676
rect 11081 8732 11145 8736
rect 11081 8676 11085 8732
rect 11085 8676 11141 8732
rect 11141 8676 11145 8732
rect 11081 8672 11145 8676
rect 15786 8732 15850 8736
rect 15786 8676 15790 8732
rect 15790 8676 15846 8732
rect 15846 8676 15850 8732
rect 15786 8672 15850 8676
rect 15866 8732 15930 8736
rect 15866 8676 15870 8732
rect 15870 8676 15926 8732
rect 15926 8676 15930 8732
rect 15866 8672 15930 8676
rect 15946 8732 16010 8736
rect 15946 8676 15950 8732
rect 15950 8676 16006 8732
rect 16006 8676 16010 8732
rect 15946 8672 16010 8676
rect 16026 8732 16090 8736
rect 16026 8676 16030 8732
rect 16030 8676 16086 8732
rect 16086 8676 16090 8732
rect 16026 8672 16090 8676
rect 20731 8732 20795 8736
rect 20731 8676 20735 8732
rect 20735 8676 20791 8732
rect 20791 8676 20795 8732
rect 20731 8672 20795 8676
rect 20811 8732 20875 8736
rect 20811 8676 20815 8732
rect 20815 8676 20871 8732
rect 20871 8676 20875 8732
rect 20811 8672 20875 8676
rect 20891 8732 20955 8736
rect 20891 8676 20895 8732
rect 20895 8676 20951 8732
rect 20951 8676 20955 8732
rect 20891 8672 20955 8676
rect 20971 8732 21035 8736
rect 20971 8676 20975 8732
rect 20975 8676 21031 8732
rect 21031 8676 21035 8732
rect 20971 8672 21035 8676
rect 3004 8468 3068 8532
rect 3188 8468 3252 8532
rect 2452 8392 2516 8396
rect 2452 8336 2466 8392
rect 2466 8336 2516 8392
rect 2452 8332 2516 8336
rect 5396 8196 5460 8260
rect 6500 8196 6564 8260
rect 3424 8188 3488 8192
rect 3424 8132 3428 8188
rect 3428 8132 3484 8188
rect 3484 8132 3488 8188
rect 3424 8128 3488 8132
rect 3504 8188 3568 8192
rect 3504 8132 3508 8188
rect 3508 8132 3564 8188
rect 3564 8132 3568 8188
rect 3504 8128 3568 8132
rect 3584 8188 3648 8192
rect 3584 8132 3588 8188
rect 3588 8132 3644 8188
rect 3644 8132 3648 8188
rect 3584 8128 3648 8132
rect 3664 8188 3728 8192
rect 3664 8132 3668 8188
rect 3668 8132 3724 8188
rect 3724 8132 3728 8188
rect 3664 8128 3728 8132
rect 8369 8188 8433 8192
rect 8369 8132 8373 8188
rect 8373 8132 8429 8188
rect 8429 8132 8433 8188
rect 8369 8128 8433 8132
rect 8449 8188 8513 8192
rect 8449 8132 8453 8188
rect 8453 8132 8509 8188
rect 8509 8132 8513 8188
rect 8449 8128 8513 8132
rect 8529 8188 8593 8192
rect 8529 8132 8533 8188
rect 8533 8132 8589 8188
rect 8589 8132 8593 8188
rect 8529 8128 8593 8132
rect 8609 8188 8673 8192
rect 8609 8132 8613 8188
rect 8613 8132 8669 8188
rect 8669 8132 8673 8188
rect 8609 8128 8673 8132
rect 1716 8060 1780 8124
rect 4108 8120 4172 8124
rect 4108 8064 4122 8120
rect 4122 8064 4172 8120
rect 4108 8060 4172 8064
rect 13314 8188 13378 8192
rect 13314 8132 13318 8188
rect 13318 8132 13374 8188
rect 13374 8132 13378 8188
rect 13314 8128 13378 8132
rect 13394 8188 13458 8192
rect 13394 8132 13398 8188
rect 13398 8132 13454 8188
rect 13454 8132 13458 8188
rect 13394 8128 13458 8132
rect 13474 8188 13538 8192
rect 13474 8132 13478 8188
rect 13478 8132 13534 8188
rect 13534 8132 13538 8188
rect 13474 8128 13538 8132
rect 13554 8188 13618 8192
rect 13554 8132 13558 8188
rect 13558 8132 13614 8188
rect 13614 8132 13618 8188
rect 13554 8128 13618 8132
rect 18259 8188 18323 8192
rect 18259 8132 18263 8188
rect 18263 8132 18319 8188
rect 18319 8132 18323 8188
rect 18259 8128 18323 8132
rect 18339 8188 18403 8192
rect 18339 8132 18343 8188
rect 18343 8132 18399 8188
rect 18399 8132 18403 8188
rect 18339 8128 18403 8132
rect 18419 8188 18483 8192
rect 18419 8132 18423 8188
rect 18423 8132 18479 8188
rect 18479 8132 18483 8188
rect 18419 8128 18483 8132
rect 18499 8188 18563 8192
rect 18499 8132 18503 8188
rect 18503 8132 18559 8188
rect 18559 8132 18563 8188
rect 18499 8128 18563 8132
rect 10548 8060 10612 8124
rect 16804 8060 16868 8124
rect 10548 7924 10612 7988
rect 13860 7924 13924 7988
rect 19564 8060 19628 8124
rect 1348 7848 1412 7852
rect 1348 7792 1398 7848
rect 1398 7792 1412 7848
rect 1348 7788 1412 7792
rect 1900 7848 1964 7852
rect 1900 7792 1914 7848
rect 1914 7792 1964 7848
rect 1900 7788 1964 7792
rect 2820 7788 2884 7852
rect 3924 7788 3988 7852
rect 9628 7788 9692 7852
rect 2084 7652 2148 7716
rect 1164 7516 1228 7580
rect 5896 7644 5960 7648
rect 5896 7588 5900 7644
rect 5900 7588 5956 7644
rect 5956 7588 5960 7644
rect 5896 7584 5960 7588
rect 5976 7644 6040 7648
rect 5976 7588 5980 7644
rect 5980 7588 6036 7644
rect 6036 7588 6040 7644
rect 5976 7584 6040 7588
rect 6056 7644 6120 7648
rect 6056 7588 6060 7644
rect 6060 7588 6116 7644
rect 6116 7588 6120 7644
rect 6056 7584 6120 7588
rect 6136 7644 6200 7648
rect 6136 7588 6140 7644
rect 6140 7588 6196 7644
rect 6196 7588 6200 7644
rect 6136 7584 6200 7588
rect 10841 7644 10905 7648
rect 10841 7588 10845 7644
rect 10845 7588 10901 7644
rect 10901 7588 10905 7644
rect 10841 7584 10905 7588
rect 10921 7644 10985 7648
rect 10921 7588 10925 7644
rect 10925 7588 10981 7644
rect 10981 7588 10985 7644
rect 10921 7584 10985 7588
rect 11001 7644 11065 7648
rect 11001 7588 11005 7644
rect 11005 7588 11061 7644
rect 11061 7588 11065 7644
rect 11001 7584 11065 7588
rect 11081 7644 11145 7648
rect 11081 7588 11085 7644
rect 11085 7588 11141 7644
rect 11141 7588 11145 7644
rect 11081 7584 11145 7588
rect 15786 7644 15850 7648
rect 15786 7588 15790 7644
rect 15790 7588 15846 7644
rect 15846 7588 15850 7644
rect 15786 7584 15850 7588
rect 15866 7644 15930 7648
rect 15866 7588 15870 7644
rect 15870 7588 15926 7644
rect 15926 7588 15930 7644
rect 15866 7584 15930 7588
rect 15946 7644 16010 7648
rect 15946 7588 15950 7644
rect 15950 7588 16006 7644
rect 16006 7588 16010 7644
rect 15946 7584 16010 7588
rect 16026 7644 16090 7648
rect 16026 7588 16030 7644
rect 16030 7588 16086 7644
rect 16086 7588 16090 7644
rect 16026 7584 16090 7588
rect 5396 7516 5460 7580
rect 12756 7516 12820 7580
rect 12940 7516 13004 7580
rect 20731 7644 20795 7648
rect 20731 7588 20735 7644
rect 20735 7588 20791 7644
rect 20791 7588 20795 7644
rect 20731 7584 20795 7588
rect 20811 7644 20875 7648
rect 20811 7588 20815 7644
rect 20815 7588 20871 7644
rect 20871 7588 20875 7644
rect 20811 7584 20875 7588
rect 20891 7644 20955 7648
rect 20891 7588 20895 7644
rect 20895 7588 20951 7644
rect 20951 7588 20955 7644
rect 20891 7584 20955 7588
rect 20971 7644 21035 7648
rect 20971 7588 20975 7644
rect 20975 7588 21031 7644
rect 21031 7588 21035 7644
rect 20971 7584 21035 7588
rect 3188 7380 3252 7444
rect 1348 7244 1412 7308
rect 3424 7100 3488 7104
rect 3424 7044 3428 7100
rect 3428 7044 3484 7100
rect 3484 7044 3488 7100
rect 3424 7040 3488 7044
rect 3504 7100 3568 7104
rect 3504 7044 3508 7100
rect 3508 7044 3564 7100
rect 3564 7044 3568 7100
rect 3504 7040 3568 7044
rect 3584 7100 3648 7104
rect 3584 7044 3588 7100
rect 3588 7044 3644 7100
rect 3644 7044 3648 7100
rect 3584 7040 3648 7044
rect 3664 7100 3728 7104
rect 3664 7044 3668 7100
rect 3668 7044 3724 7100
rect 3724 7044 3728 7100
rect 3664 7040 3728 7044
rect 12756 7244 12820 7308
rect 17172 7304 17236 7308
rect 17172 7248 17186 7304
rect 17186 7248 17236 7304
rect 17172 7244 17236 7248
rect 17724 7244 17788 7308
rect 8369 7100 8433 7104
rect 8369 7044 8373 7100
rect 8373 7044 8429 7100
rect 8429 7044 8433 7100
rect 8369 7040 8433 7044
rect 8449 7100 8513 7104
rect 8449 7044 8453 7100
rect 8453 7044 8509 7100
rect 8509 7044 8513 7100
rect 8449 7040 8513 7044
rect 8529 7100 8593 7104
rect 8529 7044 8533 7100
rect 8533 7044 8589 7100
rect 8589 7044 8593 7100
rect 8529 7040 8593 7044
rect 8609 7100 8673 7104
rect 8609 7044 8613 7100
rect 8613 7044 8669 7100
rect 8669 7044 8673 7100
rect 8609 7040 8673 7044
rect 13314 7100 13378 7104
rect 13314 7044 13318 7100
rect 13318 7044 13374 7100
rect 13374 7044 13378 7100
rect 13314 7040 13378 7044
rect 13394 7100 13458 7104
rect 13394 7044 13398 7100
rect 13398 7044 13454 7100
rect 13454 7044 13458 7100
rect 13394 7040 13458 7044
rect 13474 7100 13538 7104
rect 13474 7044 13478 7100
rect 13478 7044 13534 7100
rect 13534 7044 13538 7100
rect 13474 7040 13538 7044
rect 13554 7100 13618 7104
rect 13554 7044 13558 7100
rect 13558 7044 13614 7100
rect 13614 7044 13618 7100
rect 13554 7040 13618 7044
rect 18259 7100 18323 7104
rect 18259 7044 18263 7100
rect 18263 7044 18319 7100
rect 18319 7044 18323 7100
rect 18259 7040 18323 7044
rect 18339 7100 18403 7104
rect 18339 7044 18343 7100
rect 18343 7044 18399 7100
rect 18399 7044 18403 7100
rect 18339 7040 18403 7044
rect 18419 7100 18483 7104
rect 18419 7044 18423 7100
rect 18423 7044 18479 7100
rect 18479 7044 18483 7100
rect 18419 7040 18483 7044
rect 18499 7100 18563 7104
rect 18499 7044 18503 7100
rect 18503 7044 18559 7100
rect 18559 7044 18563 7100
rect 18499 7040 18563 7044
rect 5212 6896 5276 6900
rect 5212 6840 5262 6896
rect 5262 6840 5276 6896
rect 5212 6836 5276 6840
rect 12940 6972 13004 7036
rect 18092 7032 18156 7036
rect 18092 6976 18106 7032
rect 18106 6976 18156 7032
rect 18092 6972 18156 6976
rect 12940 6836 13004 6900
rect 9996 6564 10060 6628
rect 5896 6556 5960 6560
rect 5896 6500 5900 6556
rect 5900 6500 5956 6556
rect 5956 6500 5960 6556
rect 5896 6496 5960 6500
rect 5976 6556 6040 6560
rect 5976 6500 5980 6556
rect 5980 6500 6036 6556
rect 6036 6500 6040 6556
rect 5976 6496 6040 6500
rect 6056 6556 6120 6560
rect 6056 6500 6060 6556
rect 6060 6500 6116 6556
rect 6116 6500 6120 6556
rect 6056 6496 6120 6500
rect 6136 6556 6200 6560
rect 6136 6500 6140 6556
rect 6140 6500 6196 6556
rect 6196 6500 6200 6556
rect 6136 6496 6200 6500
rect 4108 6488 4172 6492
rect 4108 6432 4122 6488
rect 4122 6432 4172 6488
rect 4108 6428 4172 6432
rect 244 6156 308 6220
rect 4476 6352 4540 6356
rect 4476 6296 4526 6352
rect 4526 6296 4540 6352
rect 4476 6292 4540 6296
rect 6868 6292 6932 6356
rect 9996 6428 10060 6492
rect 14964 6700 15028 6764
rect 14228 6564 14292 6628
rect 10841 6556 10905 6560
rect 10841 6500 10845 6556
rect 10845 6500 10901 6556
rect 10901 6500 10905 6556
rect 10841 6496 10905 6500
rect 10921 6556 10985 6560
rect 10921 6500 10925 6556
rect 10925 6500 10981 6556
rect 10981 6500 10985 6556
rect 10921 6496 10985 6500
rect 11001 6556 11065 6560
rect 11001 6500 11005 6556
rect 11005 6500 11061 6556
rect 11061 6500 11065 6556
rect 11001 6496 11065 6500
rect 11081 6556 11145 6560
rect 11081 6500 11085 6556
rect 11085 6500 11141 6556
rect 11141 6500 11145 6556
rect 11081 6496 11145 6500
rect 15786 6556 15850 6560
rect 15786 6500 15790 6556
rect 15790 6500 15846 6556
rect 15846 6500 15850 6556
rect 15786 6496 15850 6500
rect 15866 6556 15930 6560
rect 15866 6500 15870 6556
rect 15870 6500 15926 6556
rect 15926 6500 15930 6556
rect 15866 6496 15930 6500
rect 15946 6556 16010 6560
rect 15946 6500 15950 6556
rect 15950 6500 16006 6556
rect 16006 6500 16010 6556
rect 15946 6496 16010 6500
rect 16026 6556 16090 6560
rect 16026 6500 16030 6556
rect 16030 6500 16086 6556
rect 16086 6500 16090 6556
rect 16026 6496 16090 6500
rect 7604 6156 7668 6220
rect 5028 6020 5092 6084
rect 9628 6292 9692 6356
rect 15516 6488 15580 6492
rect 15516 6432 15566 6488
rect 15566 6432 15580 6488
rect 15516 6428 15580 6432
rect 20731 6556 20795 6560
rect 20731 6500 20735 6556
rect 20735 6500 20791 6556
rect 20791 6500 20795 6556
rect 20731 6496 20795 6500
rect 20811 6556 20875 6560
rect 20811 6500 20815 6556
rect 20815 6500 20871 6556
rect 20871 6500 20875 6556
rect 20811 6496 20875 6500
rect 20891 6556 20955 6560
rect 20891 6500 20895 6556
rect 20895 6500 20951 6556
rect 20951 6500 20955 6556
rect 20891 6496 20955 6500
rect 20971 6556 21035 6560
rect 20971 6500 20975 6556
rect 20975 6500 21031 6556
rect 21031 6500 21035 6556
rect 20971 6496 21035 6500
rect 3424 6012 3488 6016
rect 3424 5956 3428 6012
rect 3428 5956 3484 6012
rect 3484 5956 3488 6012
rect 3424 5952 3488 5956
rect 3504 6012 3568 6016
rect 3504 5956 3508 6012
rect 3508 5956 3564 6012
rect 3564 5956 3568 6012
rect 3504 5952 3568 5956
rect 3584 6012 3648 6016
rect 3584 5956 3588 6012
rect 3588 5956 3644 6012
rect 3644 5956 3648 6012
rect 3584 5952 3648 5956
rect 3664 6012 3728 6016
rect 3664 5956 3668 6012
rect 3668 5956 3724 6012
rect 3724 5956 3728 6012
rect 3664 5952 3728 5956
rect 8369 6012 8433 6016
rect 8369 5956 8373 6012
rect 8373 5956 8429 6012
rect 8429 5956 8433 6012
rect 8369 5952 8433 5956
rect 8449 6012 8513 6016
rect 8449 5956 8453 6012
rect 8453 5956 8509 6012
rect 8509 5956 8513 6012
rect 8449 5952 8513 5956
rect 8529 6012 8593 6016
rect 8529 5956 8533 6012
rect 8533 5956 8589 6012
rect 8589 5956 8593 6012
rect 8529 5952 8593 5956
rect 8609 6012 8673 6016
rect 8609 5956 8613 6012
rect 8613 5956 8669 6012
rect 8669 5956 8673 6012
rect 8609 5952 8673 5956
rect 13314 6012 13378 6016
rect 13314 5956 13318 6012
rect 13318 5956 13374 6012
rect 13374 5956 13378 6012
rect 13314 5952 13378 5956
rect 13394 6012 13458 6016
rect 13394 5956 13398 6012
rect 13398 5956 13454 6012
rect 13454 5956 13458 6012
rect 13394 5952 13458 5956
rect 13474 6012 13538 6016
rect 13474 5956 13478 6012
rect 13478 5956 13534 6012
rect 13534 5956 13538 6012
rect 13474 5952 13538 5956
rect 13554 6012 13618 6016
rect 13554 5956 13558 6012
rect 13558 5956 13614 6012
rect 13614 5956 13618 6012
rect 13554 5952 13618 5956
rect 18259 6012 18323 6016
rect 18259 5956 18263 6012
rect 18263 5956 18319 6012
rect 18319 5956 18323 6012
rect 18259 5952 18323 5956
rect 18339 6012 18403 6016
rect 18339 5956 18343 6012
rect 18343 5956 18399 6012
rect 18399 5956 18403 6012
rect 18339 5952 18403 5956
rect 18419 6012 18483 6016
rect 18419 5956 18423 6012
rect 18423 5956 18479 6012
rect 18479 5956 18483 6012
rect 18419 5952 18483 5956
rect 18499 6012 18563 6016
rect 18499 5956 18503 6012
rect 18503 5956 18559 6012
rect 18559 5956 18563 6012
rect 18499 5952 18563 5956
rect 3004 5884 3068 5948
rect 6684 5884 6748 5948
rect 6500 5748 6564 5812
rect 7788 5748 7852 5812
rect 8892 5748 8956 5812
rect 9260 5808 9324 5812
rect 9260 5752 9274 5808
rect 9274 5752 9324 5808
rect 9260 5748 9324 5752
rect 5580 5672 5644 5676
rect 5580 5616 5594 5672
rect 5594 5616 5644 5672
rect 5580 5612 5644 5616
rect 6684 5536 6748 5540
rect 6684 5480 6734 5536
rect 6734 5480 6748 5536
rect 6684 5476 6748 5480
rect 6868 5476 6932 5540
rect 5896 5468 5960 5472
rect 5896 5412 5900 5468
rect 5900 5412 5956 5468
rect 5956 5412 5960 5468
rect 5896 5408 5960 5412
rect 5976 5468 6040 5472
rect 5976 5412 5980 5468
rect 5980 5412 6036 5468
rect 6036 5412 6040 5468
rect 5976 5408 6040 5412
rect 6056 5468 6120 5472
rect 6056 5412 6060 5468
rect 6060 5412 6116 5468
rect 6116 5412 6120 5468
rect 6056 5408 6120 5412
rect 6136 5468 6200 5472
rect 6136 5412 6140 5468
rect 6140 5412 6196 5468
rect 6196 5412 6200 5468
rect 6136 5408 6200 5412
rect 7420 5340 7484 5404
rect 12204 5884 12268 5948
rect 13124 5884 13188 5948
rect 13860 5884 13924 5948
rect 14412 5884 14476 5948
rect 12020 5748 12084 5812
rect 11652 5476 11716 5540
rect 10841 5468 10905 5472
rect 10841 5412 10845 5468
rect 10845 5412 10901 5468
rect 10901 5412 10905 5468
rect 10841 5408 10905 5412
rect 10921 5468 10985 5472
rect 10921 5412 10925 5468
rect 10925 5412 10981 5468
rect 10981 5412 10985 5468
rect 10921 5408 10985 5412
rect 11001 5468 11065 5472
rect 11001 5412 11005 5468
rect 11005 5412 11061 5468
rect 11061 5412 11065 5468
rect 11001 5408 11065 5412
rect 11081 5468 11145 5472
rect 11081 5412 11085 5468
rect 11085 5412 11141 5468
rect 11141 5412 11145 5468
rect 11081 5408 11145 5412
rect 12756 5340 12820 5404
rect 7972 5204 8036 5268
rect 10548 5204 10612 5268
rect 5212 5068 5276 5132
rect 9076 5068 9140 5132
rect 11284 5128 11348 5132
rect 11284 5072 11334 5128
rect 11334 5072 11348 5128
rect 11284 5068 11348 5072
rect 11652 5128 11716 5132
rect 11652 5072 11666 5128
rect 11666 5072 11716 5128
rect 11652 5068 11716 5072
rect 10548 4932 10612 4996
rect 13124 5068 13188 5132
rect 15148 5204 15212 5268
rect 19380 5476 19444 5540
rect 15786 5468 15850 5472
rect 15786 5412 15790 5468
rect 15790 5412 15846 5468
rect 15846 5412 15850 5468
rect 15786 5408 15850 5412
rect 15866 5468 15930 5472
rect 15866 5412 15870 5468
rect 15870 5412 15926 5468
rect 15926 5412 15930 5468
rect 15866 5408 15930 5412
rect 15946 5468 16010 5472
rect 15946 5412 15950 5468
rect 15950 5412 16006 5468
rect 16006 5412 16010 5468
rect 15946 5408 16010 5412
rect 16026 5468 16090 5472
rect 16026 5412 16030 5468
rect 16030 5412 16086 5468
rect 16086 5412 16090 5468
rect 16026 5408 16090 5412
rect 20731 5468 20795 5472
rect 20731 5412 20735 5468
rect 20735 5412 20791 5468
rect 20791 5412 20795 5468
rect 20731 5408 20795 5412
rect 20811 5468 20875 5472
rect 20811 5412 20815 5468
rect 20815 5412 20871 5468
rect 20871 5412 20875 5468
rect 20811 5408 20875 5412
rect 20891 5468 20955 5472
rect 20891 5412 20895 5468
rect 20895 5412 20951 5468
rect 20951 5412 20955 5468
rect 20891 5408 20955 5412
rect 20971 5468 21035 5472
rect 20971 5412 20975 5468
rect 20975 5412 21031 5468
rect 21031 5412 21035 5468
rect 20971 5408 21035 5412
rect 3424 4924 3488 4928
rect 3424 4868 3428 4924
rect 3428 4868 3484 4924
rect 3484 4868 3488 4924
rect 3424 4864 3488 4868
rect 3504 4924 3568 4928
rect 3504 4868 3508 4924
rect 3508 4868 3564 4924
rect 3564 4868 3568 4924
rect 3504 4864 3568 4868
rect 3584 4924 3648 4928
rect 3584 4868 3588 4924
rect 3588 4868 3644 4924
rect 3644 4868 3648 4924
rect 3584 4864 3648 4868
rect 3664 4924 3728 4928
rect 3664 4868 3668 4924
rect 3668 4868 3724 4924
rect 3724 4868 3728 4924
rect 3664 4864 3728 4868
rect 8369 4924 8433 4928
rect 8369 4868 8373 4924
rect 8373 4868 8429 4924
rect 8429 4868 8433 4924
rect 8369 4864 8433 4868
rect 8449 4924 8513 4928
rect 8449 4868 8453 4924
rect 8453 4868 8509 4924
rect 8509 4868 8513 4924
rect 8449 4864 8513 4868
rect 8529 4924 8593 4928
rect 8529 4868 8533 4924
rect 8533 4868 8589 4924
rect 8589 4868 8593 4924
rect 8529 4864 8593 4868
rect 8609 4924 8673 4928
rect 8609 4868 8613 4924
rect 8613 4868 8669 4924
rect 8669 4868 8673 4924
rect 8609 4864 8673 4868
rect 6868 4796 6932 4860
rect 7052 4856 7116 4860
rect 7052 4800 7066 4856
rect 7066 4800 7116 4856
rect 7052 4796 7116 4800
rect 7972 4796 8036 4860
rect 13314 4924 13378 4928
rect 13314 4868 13318 4924
rect 13318 4868 13374 4924
rect 13374 4868 13378 4924
rect 13314 4864 13378 4868
rect 13394 4924 13458 4928
rect 13394 4868 13398 4924
rect 13398 4868 13454 4924
rect 13454 4868 13458 4924
rect 13394 4864 13458 4868
rect 13474 4924 13538 4928
rect 13474 4868 13478 4924
rect 13478 4868 13534 4924
rect 13534 4868 13538 4924
rect 13474 4864 13538 4868
rect 13554 4924 13618 4928
rect 13554 4868 13558 4924
rect 13558 4868 13614 4924
rect 13614 4868 13618 4924
rect 13554 4864 13618 4868
rect 11652 4856 11716 4860
rect 11652 4800 11702 4856
rect 11702 4800 11716 4856
rect 11652 4796 11716 4800
rect 11836 4796 11900 4860
rect 12204 4796 12268 4860
rect 5580 4660 5644 4724
rect 6868 4660 6932 4724
rect 10364 4660 10428 4724
rect 12020 4660 12084 4724
rect 12572 4660 12636 4724
rect 6868 4524 6932 4588
rect 11284 4524 11348 4588
rect 12204 4524 12268 4588
rect 18259 4924 18323 4928
rect 18259 4868 18263 4924
rect 18263 4868 18319 4924
rect 18319 4868 18323 4924
rect 18259 4864 18323 4868
rect 18339 4924 18403 4928
rect 18339 4868 18343 4924
rect 18343 4868 18399 4924
rect 18399 4868 18403 4924
rect 18339 4864 18403 4868
rect 18419 4924 18483 4928
rect 18419 4868 18423 4924
rect 18423 4868 18479 4924
rect 18479 4868 18483 4924
rect 18419 4864 18483 4868
rect 18499 4924 18563 4928
rect 18499 4868 18503 4924
rect 18503 4868 18559 4924
rect 18559 4868 18563 4924
rect 18499 4864 18563 4868
rect 14228 4524 14292 4588
rect 4844 4388 4908 4452
rect 6684 4448 6748 4452
rect 6684 4392 6734 4448
rect 6734 4392 6748 4448
rect 6684 4388 6748 4392
rect 7052 4388 7116 4452
rect 5896 4380 5960 4384
rect 5896 4324 5900 4380
rect 5900 4324 5956 4380
rect 5956 4324 5960 4380
rect 5896 4320 5960 4324
rect 5976 4380 6040 4384
rect 5976 4324 5980 4380
rect 5980 4324 6036 4380
rect 6036 4324 6040 4380
rect 5976 4320 6040 4324
rect 6056 4380 6120 4384
rect 6056 4324 6060 4380
rect 6060 4324 6116 4380
rect 6116 4324 6120 4380
rect 6056 4320 6120 4324
rect 6136 4380 6200 4384
rect 6136 4324 6140 4380
rect 6140 4324 6196 4380
rect 6196 4324 6200 4380
rect 6136 4320 6200 4324
rect 10841 4380 10905 4384
rect 10841 4324 10845 4380
rect 10845 4324 10901 4380
rect 10901 4324 10905 4380
rect 10841 4320 10905 4324
rect 10921 4380 10985 4384
rect 10921 4324 10925 4380
rect 10925 4324 10981 4380
rect 10981 4324 10985 4380
rect 10921 4320 10985 4324
rect 11001 4380 11065 4384
rect 11001 4324 11005 4380
rect 11005 4324 11061 4380
rect 11061 4324 11065 4380
rect 11001 4320 11065 4324
rect 11081 4380 11145 4384
rect 11081 4324 11085 4380
rect 11085 4324 11141 4380
rect 11141 4324 11145 4380
rect 11081 4320 11145 4324
rect 12756 4388 12820 4452
rect 13124 4388 13188 4452
rect 15148 4660 15212 4724
rect 16988 4660 17052 4724
rect 19932 4388 19996 4452
rect 15786 4380 15850 4384
rect 15786 4324 15790 4380
rect 15790 4324 15846 4380
rect 15846 4324 15850 4380
rect 15786 4320 15850 4324
rect 15866 4380 15930 4384
rect 15866 4324 15870 4380
rect 15870 4324 15926 4380
rect 15926 4324 15930 4380
rect 15866 4320 15930 4324
rect 15946 4380 16010 4384
rect 15946 4324 15950 4380
rect 15950 4324 16006 4380
rect 16006 4324 16010 4380
rect 15946 4320 16010 4324
rect 16026 4380 16090 4384
rect 16026 4324 16030 4380
rect 16030 4324 16086 4380
rect 16086 4324 16090 4380
rect 16026 4320 16090 4324
rect 20731 4380 20795 4384
rect 20731 4324 20735 4380
rect 20735 4324 20791 4380
rect 20791 4324 20795 4380
rect 20731 4320 20795 4324
rect 20811 4380 20875 4384
rect 20811 4324 20815 4380
rect 20815 4324 20871 4380
rect 20871 4324 20875 4380
rect 20811 4320 20875 4324
rect 20891 4380 20955 4384
rect 20891 4324 20895 4380
rect 20895 4324 20951 4380
rect 20951 4324 20955 4380
rect 20891 4320 20955 4324
rect 20971 4380 21035 4384
rect 20971 4324 20975 4380
rect 20975 4324 21031 4380
rect 21031 4324 21035 4380
rect 20971 4320 21035 4324
rect 1532 4116 1596 4180
rect 5580 4116 5644 4180
rect 12388 4252 12452 4316
rect 12756 4252 12820 4316
rect 19196 4312 19260 4316
rect 19196 4256 19246 4312
rect 19246 4256 19260 4312
rect 19196 4252 19260 4256
rect 14780 4116 14844 4180
rect 3188 3980 3252 4044
rect 12020 3980 12084 4044
rect 3424 3836 3488 3840
rect 3424 3780 3428 3836
rect 3428 3780 3484 3836
rect 3484 3780 3488 3836
rect 3424 3776 3488 3780
rect 3504 3836 3568 3840
rect 3504 3780 3508 3836
rect 3508 3780 3564 3836
rect 3564 3780 3568 3836
rect 3504 3776 3568 3780
rect 3584 3836 3648 3840
rect 3584 3780 3588 3836
rect 3588 3780 3644 3836
rect 3644 3780 3648 3836
rect 3584 3776 3648 3780
rect 3664 3836 3728 3840
rect 3664 3780 3668 3836
rect 3668 3780 3724 3836
rect 3724 3780 3728 3836
rect 3664 3776 3728 3780
rect 8369 3836 8433 3840
rect 8369 3780 8373 3836
rect 8373 3780 8429 3836
rect 8429 3780 8433 3836
rect 8369 3776 8433 3780
rect 8449 3836 8513 3840
rect 8449 3780 8453 3836
rect 8453 3780 8509 3836
rect 8509 3780 8513 3836
rect 8449 3776 8513 3780
rect 8529 3836 8593 3840
rect 8529 3780 8533 3836
rect 8533 3780 8589 3836
rect 8589 3780 8593 3836
rect 8529 3776 8593 3780
rect 8609 3836 8673 3840
rect 8609 3780 8613 3836
rect 8613 3780 8669 3836
rect 8669 3780 8673 3836
rect 8609 3776 8673 3780
rect 4476 3708 4540 3772
rect 9996 3844 10060 3908
rect 11652 3844 11716 3908
rect 17356 3980 17420 4044
rect 15516 3844 15580 3908
rect 13314 3836 13378 3840
rect 13314 3780 13318 3836
rect 13318 3780 13374 3836
rect 13374 3780 13378 3836
rect 13314 3776 13378 3780
rect 13394 3836 13458 3840
rect 13394 3780 13398 3836
rect 13398 3780 13454 3836
rect 13454 3780 13458 3836
rect 13394 3776 13458 3780
rect 13474 3836 13538 3840
rect 13474 3780 13478 3836
rect 13478 3780 13534 3836
rect 13534 3780 13538 3836
rect 13474 3776 13538 3780
rect 13554 3836 13618 3840
rect 13554 3780 13558 3836
rect 13558 3780 13614 3836
rect 13614 3780 13618 3836
rect 13554 3776 13618 3780
rect 18259 3836 18323 3840
rect 18259 3780 18263 3836
rect 18263 3780 18319 3836
rect 18319 3780 18323 3836
rect 18259 3776 18323 3780
rect 18339 3836 18403 3840
rect 18339 3780 18343 3836
rect 18343 3780 18399 3836
rect 18399 3780 18403 3836
rect 18339 3776 18403 3780
rect 18419 3836 18483 3840
rect 18419 3780 18423 3836
rect 18423 3780 18479 3836
rect 18479 3780 18483 3836
rect 18419 3776 18483 3780
rect 18499 3836 18563 3840
rect 18499 3780 18503 3836
rect 18503 3780 18559 3836
rect 18559 3780 18563 3836
rect 18499 3776 18563 3780
rect 12572 3708 12636 3772
rect 13124 3708 13188 3772
rect 13906 3708 13970 3772
rect 14228 3708 14292 3772
rect 14596 3708 14660 3772
rect 14964 3708 15028 3772
rect 15148 3708 15212 3772
rect 17540 3768 17604 3772
rect 17540 3712 17554 3768
rect 17554 3712 17604 3768
rect 17540 3708 17604 3712
rect 7604 3572 7668 3636
rect 12572 3572 12636 3636
rect 14964 3572 15028 3636
rect 6684 3300 6748 3364
rect 9812 3300 9876 3364
rect 10548 3300 10612 3364
rect 11284 3300 11348 3364
rect 12388 3360 12452 3364
rect 12388 3304 12438 3360
rect 12438 3304 12452 3360
rect 12388 3300 12452 3304
rect 5896 3292 5960 3296
rect 5896 3236 5900 3292
rect 5900 3236 5956 3292
rect 5956 3236 5960 3292
rect 5896 3232 5960 3236
rect 5976 3292 6040 3296
rect 5976 3236 5980 3292
rect 5980 3236 6036 3292
rect 6036 3236 6040 3292
rect 5976 3232 6040 3236
rect 6056 3292 6120 3296
rect 6056 3236 6060 3292
rect 6060 3236 6116 3292
rect 6116 3236 6120 3292
rect 6056 3232 6120 3236
rect 6136 3292 6200 3296
rect 6136 3236 6140 3292
rect 6140 3236 6196 3292
rect 6196 3236 6200 3292
rect 6136 3232 6200 3236
rect 10841 3292 10905 3296
rect 10841 3236 10845 3292
rect 10845 3236 10901 3292
rect 10901 3236 10905 3292
rect 10841 3232 10905 3236
rect 10921 3292 10985 3296
rect 10921 3236 10925 3292
rect 10925 3236 10981 3292
rect 10981 3236 10985 3292
rect 10921 3232 10985 3236
rect 11001 3292 11065 3296
rect 11001 3236 11005 3292
rect 11005 3236 11061 3292
rect 11061 3236 11065 3292
rect 11001 3232 11065 3236
rect 11081 3292 11145 3296
rect 11081 3236 11085 3292
rect 11085 3236 11141 3292
rect 11141 3236 11145 3292
rect 11081 3232 11145 3236
rect 6316 3224 6380 3228
rect 6316 3168 6330 3224
rect 6330 3168 6380 3224
rect 6316 3164 6380 3168
rect 5212 3028 5276 3092
rect 5580 3028 5644 3092
rect 8156 3164 8220 3228
rect 10180 3164 10244 3228
rect 11284 3164 11348 3228
rect 7604 2892 7668 2956
rect 3424 2748 3488 2752
rect 3424 2692 3428 2748
rect 3428 2692 3484 2748
rect 3484 2692 3488 2748
rect 3424 2688 3488 2692
rect 3504 2748 3568 2752
rect 3504 2692 3508 2748
rect 3508 2692 3564 2748
rect 3564 2692 3568 2748
rect 3504 2688 3568 2692
rect 3584 2748 3648 2752
rect 3584 2692 3588 2748
rect 3588 2692 3644 2748
rect 3644 2692 3648 2748
rect 3584 2688 3648 2692
rect 3664 2748 3728 2752
rect 3664 2692 3668 2748
rect 3668 2692 3724 2748
rect 3724 2692 3728 2748
rect 3664 2688 3728 2692
rect 428 2680 492 2684
rect 428 2624 478 2680
rect 478 2624 492 2680
rect 428 2620 492 2624
rect 612 2620 676 2684
rect 2636 2620 2700 2684
rect 4292 2680 4356 2684
rect 9444 3028 9508 3092
rect 9996 3028 10060 3092
rect 11468 3028 11532 3092
rect 13124 3164 13188 3228
rect 16620 3300 16684 3364
rect 15786 3292 15850 3296
rect 15786 3236 15790 3292
rect 15790 3236 15846 3292
rect 15846 3236 15850 3292
rect 15786 3232 15850 3236
rect 15866 3292 15930 3296
rect 15866 3236 15870 3292
rect 15870 3236 15926 3292
rect 15926 3236 15930 3292
rect 15866 3232 15930 3236
rect 15946 3292 16010 3296
rect 15946 3236 15950 3292
rect 15950 3236 16006 3292
rect 16006 3236 16010 3292
rect 15946 3232 16010 3236
rect 16026 3292 16090 3296
rect 16026 3236 16030 3292
rect 16030 3236 16086 3292
rect 16086 3236 16090 3292
rect 16026 3232 16090 3236
rect 20731 3292 20795 3296
rect 20731 3236 20735 3292
rect 20735 3236 20791 3292
rect 20791 3236 20795 3292
rect 20731 3232 20795 3236
rect 20811 3292 20875 3296
rect 20811 3236 20815 3292
rect 20815 3236 20871 3292
rect 20871 3236 20875 3292
rect 20811 3232 20875 3236
rect 20891 3292 20955 3296
rect 20891 3236 20895 3292
rect 20895 3236 20951 3292
rect 20951 3236 20955 3292
rect 20891 3232 20955 3236
rect 20971 3292 21035 3296
rect 20971 3236 20975 3292
rect 20975 3236 21031 3292
rect 21031 3236 21035 3292
rect 20971 3232 21035 3236
rect 9996 2756 10060 2820
rect 12020 2756 12084 2820
rect 12204 2816 12268 2820
rect 12204 2760 12254 2816
rect 12254 2760 12268 2816
rect 12204 2756 12268 2760
rect 13124 2756 13188 2820
rect 14228 2756 14292 2820
rect 8369 2748 8433 2752
rect 8369 2692 8373 2748
rect 8373 2692 8429 2748
rect 8429 2692 8433 2748
rect 8369 2688 8433 2692
rect 8449 2748 8513 2752
rect 8449 2692 8453 2748
rect 8453 2692 8509 2748
rect 8509 2692 8513 2748
rect 8449 2688 8513 2692
rect 8529 2748 8593 2752
rect 8529 2692 8533 2748
rect 8533 2692 8589 2748
rect 8589 2692 8593 2748
rect 8529 2688 8593 2692
rect 8609 2748 8673 2752
rect 8609 2692 8613 2748
rect 8613 2692 8669 2748
rect 8669 2692 8673 2748
rect 8609 2688 8673 2692
rect 4292 2624 4342 2680
rect 4342 2624 4356 2680
rect 4292 2620 4356 2624
rect 1716 2484 1780 2548
rect 13314 2748 13378 2752
rect 13314 2692 13318 2748
rect 13318 2692 13374 2748
rect 13374 2692 13378 2748
rect 13314 2688 13378 2692
rect 13394 2748 13458 2752
rect 13394 2692 13398 2748
rect 13398 2692 13454 2748
rect 13454 2692 13458 2748
rect 13394 2688 13458 2692
rect 13474 2748 13538 2752
rect 13474 2692 13478 2748
rect 13478 2692 13534 2748
rect 13534 2692 13538 2748
rect 13474 2688 13538 2692
rect 13554 2748 13618 2752
rect 13554 2692 13558 2748
rect 13558 2692 13614 2748
rect 13614 2692 13618 2748
rect 13554 2688 13618 2692
rect 12756 2620 12820 2684
rect 13860 2680 13924 2684
rect 13860 2624 13874 2680
rect 13874 2624 13924 2680
rect 13860 2620 13924 2624
rect 18644 2756 18708 2820
rect 19564 2816 19628 2820
rect 19564 2760 19614 2816
rect 19614 2760 19628 2816
rect 19564 2756 19628 2760
rect 18259 2748 18323 2752
rect 18259 2692 18263 2748
rect 18263 2692 18319 2748
rect 18319 2692 18323 2748
rect 18259 2688 18323 2692
rect 18339 2748 18403 2752
rect 18339 2692 18343 2748
rect 18343 2692 18399 2748
rect 18399 2692 18403 2748
rect 18339 2688 18403 2692
rect 18419 2748 18483 2752
rect 18419 2692 18423 2748
rect 18423 2692 18479 2748
rect 18479 2692 18483 2748
rect 18419 2688 18483 2692
rect 18499 2748 18563 2752
rect 18499 2692 18503 2748
rect 18503 2692 18559 2748
rect 18559 2692 18563 2748
rect 18499 2688 18563 2692
rect 796 2348 860 2412
rect 4476 2348 4540 2412
rect 4660 2348 4724 2412
rect 5580 2348 5644 2412
rect 5896 2204 5960 2208
rect 5896 2148 5900 2204
rect 5900 2148 5956 2204
rect 5956 2148 5960 2204
rect 5896 2144 5960 2148
rect 5976 2204 6040 2208
rect 5976 2148 5980 2204
rect 5980 2148 6036 2204
rect 6036 2148 6040 2204
rect 5976 2144 6040 2148
rect 6056 2204 6120 2208
rect 6056 2148 6060 2204
rect 6060 2148 6116 2204
rect 6116 2148 6120 2204
rect 6056 2144 6120 2148
rect 6136 2204 6200 2208
rect 6136 2148 6140 2204
rect 6140 2148 6196 2204
rect 6196 2148 6200 2204
rect 6136 2144 6200 2148
rect 7788 2348 7852 2412
rect 7420 2272 7484 2276
rect 7420 2216 7470 2272
rect 7470 2216 7484 2272
rect 7420 2212 7484 2216
rect 7236 1940 7300 2004
rect 10364 2212 10428 2276
rect 10841 2204 10905 2208
rect 10841 2148 10845 2204
rect 10845 2148 10901 2204
rect 10901 2148 10905 2204
rect 10841 2144 10905 2148
rect 10921 2204 10985 2208
rect 10921 2148 10925 2204
rect 10925 2148 10981 2204
rect 10981 2148 10985 2204
rect 10921 2144 10985 2148
rect 11001 2204 11065 2208
rect 11001 2148 11005 2204
rect 11005 2148 11061 2204
rect 11061 2148 11065 2204
rect 11001 2144 11065 2148
rect 11081 2204 11145 2208
rect 11081 2148 11085 2204
rect 11085 2148 11141 2204
rect 11141 2148 11145 2204
rect 11081 2144 11145 2148
rect 12572 2484 12636 2548
rect 12756 2348 12820 2412
rect 16988 2348 17052 2412
rect 19012 2348 19076 2412
rect 12940 2212 13004 2276
rect 15332 2212 15396 2276
rect 15786 2204 15850 2208
rect 15786 2148 15790 2204
rect 15790 2148 15846 2204
rect 15846 2148 15850 2204
rect 15786 2144 15850 2148
rect 15866 2204 15930 2208
rect 15866 2148 15870 2204
rect 15870 2148 15926 2204
rect 15926 2148 15930 2204
rect 15866 2144 15930 2148
rect 15946 2204 16010 2208
rect 15946 2148 15950 2204
rect 15950 2148 16006 2204
rect 16006 2148 16010 2204
rect 15946 2144 16010 2148
rect 16026 2204 16090 2208
rect 16026 2148 16030 2204
rect 16030 2148 16086 2204
rect 16086 2148 16090 2204
rect 16026 2144 16090 2148
rect 20731 2204 20795 2208
rect 20731 2148 20735 2204
rect 20735 2148 20791 2204
rect 20791 2148 20795 2204
rect 20731 2144 20795 2148
rect 20811 2204 20875 2208
rect 20811 2148 20815 2204
rect 20815 2148 20871 2204
rect 20871 2148 20875 2204
rect 20811 2144 20875 2148
rect 20891 2204 20955 2208
rect 20891 2148 20895 2204
rect 20895 2148 20951 2204
rect 20951 2148 20955 2204
rect 20891 2144 20955 2148
rect 20971 2204 21035 2208
rect 20971 2148 20975 2204
rect 20975 2148 21031 2204
rect 21031 2148 21035 2204
rect 20971 2144 21035 2148
rect 11836 1940 11900 2004
rect 14780 1940 14844 2004
rect 16252 2076 16316 2140
rect 19748 1940 19812 2004
rect 980 1804 1044 1868
rect 7972 1804 8036 1868
rect 6868 1668 6932 1732
rect 3424 1660 3488 1664
rect 3424 1604 3428 1660
rect 3428 1604 3484 1660
rect 3484 1604 3488 1660
rect 3424 1600 3488 1604
rect 3504 1660 3568 1664
rect 3504 1604 3508 1660
rect 3508 1604 3564 1660
rect 3564 1604 3568 1660
rect 3504 1600 3568 1604
rect 3584 1660 3648 1664
rect 3584 1604 3588 1660
rect 3588 1604 3644 1660
rect 3644 1604 3648 1660
rect 3584 1600 3648 1604
rect 3664 1660 3728 1664
rect 3664 1604 3668 1660
rect 3668 1604 3724 1660
rect 3724 1604 3728 1660
rect 3664 1600 3728 1604
rect 8369 1660 8433 1664
rect 8369 1604 8373 1660
rect 8373 1604 8429 1660
rect 8429 1604 8433 1660
rect 8369 1600 8433 1604
rect 8449 1660 8513 1664
rect 8449 1604 8453 1660
rect 8453 1604 8509 1660
rect 8509 1604 8513 1660
rect 8449 1600 8513 1604
rect 8529 1660 8593 1664
rect 8529 1604 8533 1660
rect 8533 1604 8589 1660
rect 8589 1604 8593 1660
rect 8529 1600 8593 1604
rect 8609 1660 8673 1664
rect 8609 1604 8613 1660
rect 8613 1604 8669 1660
rect 8669 1604 8673 1660
rect 8609 1600 8673 1604
rect 12940 1804 13004 1868
rect 9628 1668 9692 1732
rect 13314 1660 13378 1664
rect 13314 1604 13318 1660
rect 13318 1604 13374 1660
rect 13374 1604 13378 1660
rect 13314 1600 13378 1604
rect 13394 1660 13458 1664
rect 13394 1604 13398 1660
rect 13398 1604 13454 1660
rect 13454 1604 13458 1660
rect 13394 1600 13458 1604
rect 13474 1660 13538 1664
rect 13474 1604 13478 1660
rect 13478 1604 13534 1660
rect 13534 1604 13538 1660
rect 13474 1600 13538 1604
rect 13554 1660 13618 1664
rect 13554 1604 13558 1660
rect 13558 1604 13614 1660
rect 13614 1604 13618 1660
rect 13554 1600 13618 1604
rect 1348 1396 1412 1460
rect 6500 1396 6564 1460
rect 9260 1456 9324 1460
rect 9260 1400 9310 1456
rect 9310 1400 9324 1456
rect 9260 1396 9324 1400
rect 12204 1396 12268 1460
rect 14044 1668 14108 1732
rect 14964 1668 15028 1732
rect 18259 1660 18323 1664
rect 18259 1604 18263 1660
rect 18263 1604 18319 1660
rect 18319 1604 18323 1660
rect 18259 1600 18323 1604
rect 18339 1660 18403 1664
rect 18339 1604 18343 1660
rect 18343 1604 18399 1660
rect 18399 1604 18403 1660
rect 18339 1600 18403 1604
rect 18419 1660 18483 1664
rect 18419 1604 18423 1660
rect 18423 1604 18479 1660
rect 18479 1604 18483 1660
rect 18419 1600 18483 1604
rect 18499 1660 18563 1664
rect 18499 1604 18503 1660
rect 18503 1604 18559 1660
rect 18559 1604 18563 1660
rect 18499 1600 18563 1604
rect 2268 1124 2332 1188
rect 7604 1124 7668 1188
rect 14412 1532 14476 1596
rect 12756 1124 12820 1188
rect 14228 1260 14292 1324
rect 16436 1260 16500 1324
rect 20116 1260 20180 1324
rect 15332 1124 15396 1188
rect 17908 1124 17972 1188
rect 5896 1116 5960 1120
rect 5896 1060 5900 1116
rect 5900 1060 5956 1116
rect 5956 1060 5960 1116
rect 5896 1056 5960 1060
rect 5976 1116 6040 1120
rect 5976 1060 5980 1116
rect 5980 1060 6036 1116
rect 6036 1060 6040 1116
rect 5976 1056 6040 1060
rect 6056 1116 6120 1120
rect 6056 1060 6060 1116
rect 6060 1060 6116 1116
rect 6116 1060 6120 1116
rect 6056 1056 6120 1060
rect 6136 1116 6200 1120
rect 6136 1060 6140 1116
rect 6140 1060 6196 1116
rect 6196 1060 6200 1116
rect 6136 1056 6200 1060
rect 10841 1116 10905 1120
rect 10841 1060 10845 1116
rect 10845 1060 10901 1116
rect 10901 1060 10905 1116
rect 10841 1056 10905 1060
rect 10921 1116 10985 1120
rect 10921 1060 10925 1116
rect 10925 1060 10981 1116
rect 10981 1060 10985 1116
rect 10921 1056 10985 1060
rect 11001 1116 11065 1120
rect 11001 1060 11005 1116
rect 11005 1060 11061 1116
rect 11061 1060 11065 1116
rect 11001 1056 11065 1060
rect 11081 1116 11145 1120
rect 11081 1060 11085 1116
rect 11085 1060 11141 1116
rect 11141 1060 11145 1116
rect 11081 1056 11145 1060
rect 15786 1116 15850 1120
rect 15786 1060 15790 1116
rect 15790 1060 15846 1116
rect 15846 1060 15850 1116
rect 15786 1056 15850 1060
rect 15866 1116 15930 1120
rect 15866 1060 15870 1116
rect 15870 1060 15926 1116
rect 15926 1060 15930 1116
rect 15866 1056 15930 1060
rect 15946 1116 16010 1120
rect 15946 1060 15950 1116
rect 15950 1060 16006 1116
rect 16006 1060 16010 1116
rect 15946 1056 16010 1060
rect 16026 1116 16090 1120
rect 16026 1060 16030 1116
rect 16030 1060 16086 1116
rect 16086 1060 16090 1116
rect 16026 1056 16090 1060
rect 20731 1116 20795 1120
rect 20731 1060 20735 1116
rect 20735 1060 20791 1116
rect 20791 1060 20795 1116
rect 20731 1056 20795 1060
rect 20811 1116 20875 1120
rect 20811 1060 20815 1116
rect 20815 1060 20871 1116
rect 20871 1060 20875 1116
rect 20811 1056 20875 1060
rect 20891 1116 20955 1120
rect 20891 1060 20895 1116
rect 20895 1060 20951 1116
rect 20951 1060 20955 1116
rect 20891 1056 20955 1060
rect 20971 1116 21035 1120
rect 20971 1060 20975 1116
rect 20975 1060 21031 1116
rect 21031 1060 21035 1116
rect 20971 1056 21035 1060
rect 15516 988 15580 1052
rect 9812 852 9876 916
rect 10180 852 10244 916
rect 11284 852 11348 916
rect 9996 716 10060 780
rect 10548 716 10612 780
rect 12020 716 12084 780
rect 15700 580 15764 644
rect 12572 444 12636 508
rect 11652 308 11716 372
rect 14090 308 14154 372
rect 14412 444 14476 508
rect 16068 444 16132 508
rect 14780 308 14844 372
rect 12388 172 12452 236
rect 6684 36 6748 100
rect 8156 36 8220 100
rect 12940 36 13004 100
<< metal4 >>
rect 14595 44572 14661 44573
rect 14595 44508 14596 44572
rect 14660 44508 14661 44572
rect 14595 44507 14661 44508
rect 3416 43008 3736 43568
rect 5888 43552 6208 43568
rect 5888 43488 5896 43552
rect 5960 43488 5976 43552
rect 6040 43488 6056 43552
rect 6120 43488 6136 43552
rect 6200 43488 6208 43552
rect 5027 43212 5093 43213
rect 5027 43148 5028 43212
rect 5092 43148 5093 43212
rect 5027 43147 5093 43148
rect 3416 42944 3424 43008
rect 3488 42944 3504 43008
rect 3568 42944 3584 43008
rect 3648 42944 3664 43008
rect 3728 42944 3736 43008
rect 3416 41920 3736 42944
rect 3416 41856 3424 41920
rect 3488 41856 3504 41920
rect 3568 41856 3584 41920
rect 3648 41856 3664 41920
rect 3728 41856 3736 41920
rect 1163 41716 1229 41717
rect 1163 41652 1164 41716
rect 1228 41652 1229 41716
rect 1163 41651 1229 41652
rect 979 38860 1045 38861
rect 979 38796 980 38860
rect 1044 38796 1045 38860
rect 979 38795 1045 38796
rect 795 35324 861 35325
rect 795 35260 796 35324
rect 860 35260 861 35324
rect 795 35259 861 35260
rect 427 33420 493 33421
rect 427 33356 428 33420
rect 492 33356 493 33420
rect 427 33355 493 33356
rect 243 15468 309 15469
rect 243 15404 244 15468
rect 308 15404 309 15468
rect 243 15403 309 15404
rect 246 6221 306 15403
rect 243 6220 309 6221
rect 243 6156 244 6220
rect 308 6156 309 6220
rect 243 6155 309 6156
rect 430 2685 490 33355
rect 798 25533 858 35259
rect 982 30290 1042 38795
rect 1166 31770 1226 41651
rect 2083 41444 2149 41445
rect 2083 41380 2084 41444
rect 2148 41380 2149 41444
rect 2083 41379 2149 41380
rect 1715 40492 1781 40493
rect 1715 40428 1716 40492
rect 1780 40428 1781 40492
rect 1715 40427 1781 40428
rect 1166 31710 1410 31770
rect 982 30230 1226 30290
rect 979 30156 1045 30157
rect 979 30092 980 30156
rect 1044 30092 1045 30156
rect 979 30091 1045 30092
rect 795 25532 861 25533
rect 795 25468 796 25532
rect 860 25468 861 25532
rect 795 25467 861 25468
rect 795 21452 861 21453
rect 795 21388 796 21452
rect 860 21388 861 21452
rect 795 21387 861 21388
rect 798 18189 858 21387
rect 795 18188 861 18189
rect 795 18124 796 18188
rect 860 18124 861 18188
rect 795 18123 861 18124
rect 795 15196 861 15197
rect 795 15132 796 15196
rect 860 15132 861 15196
rect 795 15131 861 15132
rect 611 14516 677 14517
rect 611 14452 612 14516
rect 676 14452 677 14516
rect 611 14451 677 14452
rect 614 2685 674 14451
rect 427 2684 493 2685
rect 427 2620 428 2684
rect 492 2620 493 2684
rect 427 2619 493 2620
rect 611 2684 677 2685
rect 611 2620 612 2684
rect 676 2620 677 2684
rect 611 2619 677 2620
rect 798 2413 858 15131
rect 795 2412 861 2413
rect 795 2348 796 2412
rect 860 2348 861 2412
rect 795 2347 861 2348
rect 982 1869 1042 30091
rect 1166 29069 1226 30230
rect 1163 29068 1229 29069
rect 1163 29004 1164 29068
rect 1228 29004 1229 29068
rect 1163 29003 1229 29004
rect 1350 27570 1410 31710
rect 1531 29068 1597 29069
rect 1531 29004 1532 29068
rect 1596 29004 1597 29068
rect 1531 29003 1597 29004
rect 1166 27510 1410 27570
rect 1166 23901 1226 27510
rect 1347 27436 1413 27437
rect 1347 27372 1348 27436
rect 1412 27372 1413 27436
rect 1347 27371 1413 27372
rect 1163 23900 1229 23901
rect 1163 23836 1164 23900
rect 1228 23836 1229 23900
rect 1163 23835 1229 23836
rect 1163 14516 1229 14517
rect 1163 14452 1164 14516
rect 1228 14452 1229 14516
rect 1163 14451 1229 14452
rect 1166 7581 1226 14451
rect 1350 14245 1410 27371
rect 1534 22110 1594 29003
rect 1718 27165 1778 40427
rect 2086 30157 2146 41379
rect 3187 41036 3253 41037
rect 3187 40972 3188 41036
rect 3252 40972 3253 41036
rect 3187 40971 3253 40972
rect 3003 33964 3069 33965
rect 3003 33900 3004 33964
rect 3068 33900 3069 33964
rect 3003 33899 3069 33900
rect 2451 32876 2517 32877
rect 2451 32812 2452 32876
rect 2516 32812 2517 32876
rect 2451 32811 2517 32812
rect 2267 31380 2333 31381
rect 2267 31316 2268 31380
rect 2332 31316 2333 31380
rect 2267 31315 2333 31316
rect 2083 30156 2149 30157
rect 2083 30092 2084 30156
rect 2148 30092 2149 30156
rect 2083 30091 2149 30092
rect 1899 28932 1965 28933
rect 1899 28868 1900 28932
rect 1964 28868 1965 28932
rect 1899 28867 1965 28868
rect 1715 27164 1781 27165
rect 1715 27100 1716 27164
rect 1780 27100 1781 27164
rect 1715 27099 1781 27100
rect 1715 24172 1781 24173
rect 1715 24108 1716 24172
rect 1780 24108 1781 24172
rect 1715 24107 1781 24108
rect 1718 22810 1778 24107
rect 1902 23493 1962 28867
rect 2270 28661 2330 31315
rect 2267 28660 2333 28661
rect 2267 28596 2268 28660
rect 2332 28596 2333 28660
rect 2267 28595 2333 28596
rect 2083 28252 2149 28253
rect 2083 28188 2084 28252
rect 2148 28188 2149 28252
rect 2083 28187 2149 28188
rect 1899 23492 1965 23493
rect 1899 23428 1900 23492
rect 1964 23428 1965 23492
rect 1899 23427 1965 23428
rect 1718 22750 1962 22810
rect 1534 22050 1778 22110
rect 1718 16013 1778 22050
rect 1902 21997 1962 22750
rect 1899 21996 1965 21997
rect 1899 21932 1900 21996
rect 1964 21932 1965 21996
rect 1899 21931 1965 21932
rect 2086 21181 2146 28187
rect 2454 27845 2514 32811
rect 3006 29341 3066 33899
rect 3003 29340 3069 29341
rect 3003 29276 3004 29340
rect 3068 29276 3069 29340
rect 3003 29275 3069 29276
rect 2819 28252 2885 28253
rect 2819 28188 2820 28252
rect 2884 28188 2885 28252
rect 2819 28187 2885 28188
rect 2635 27980 2701 27981
rect 2635 27916 2636 27980
rect 2700 27916 2701 27980
rect 2635 27915 2701 27916
rect 2267 27844 2333 27845
rect 2267 27780 2268 27844
rect 2332 27780 2333 27844
rect 2267 27779 2333 27780
rect 2451 27844 2517 27845
rect 2451 27780 2452 27844
rect 2516 27780 2517 27844
rect 2451 27779 2517 27780
rect 2083 21180 2149 21181
rect 2083 21116 2084 21180
rect 2148 21116 2149 21180
rect 2083 21115 2149 21116
rect 2270 18325 2330 27779
rect 2451 25668 2517 25669
rect 2451 25604 2452 25668
rect 2516 25604 2517 25668
rect 2451 25603 2517 25604
rect 2454 19410 2514 25603
rect 2638 24173 2698 27915
rect 2822 25397 2882 28187
rect 3003 27708 3069 27709
rect 3003 27644 3004 27708
rect 3068 27644 3069 27708
rect 3003 27643 3069 27644
rect 3006 25805 3066 27643
rect 3003 25804 3069 25805
rect 3003 25740 3004 25804
rect 3068 25740 3069 25804
rect 3003 25739 3069 25740
rect 2819 25396 2885 25397
rect 2819 25332 2820 25396
rect 2884 25332 2885 25396
rect 2819 25331 2885 25332
rect 2635 24172 2701 24173
rect 2635 24108 2636 24172
rect 2700 24108 2701 24172
rect 2635 24107 2701 24108
rect 2819 22812 2885 22813
rect 2819 22748 2820 22812
rect 2884 22748 2885 22812
rect 2819 22747 2885 22748
rect 2822 20093 2882 22747
rect 3006 22110 3066 25739
rect 3190 23085 3250 40971
rect 3416 40832 3736 41856
rect 3923 41580 3989 41581
rect 3923 41516 3924 41580
rect 3988 41516 3989 41580
rect 3923 41515 3989 41516
rect 3416 40768 3424 40832
rect 3488 40768 3504 40832
rect 3568 40768 3584 40832
rect 3648 40768 3664 40832
rect 3728 40768 3736 40832
rect 3416 39744 3736 40768
rect 3416 39680 3424 39744
rect 3488 39680 3504 39744
rect 3568 39680 3584 39744
rect 3648 39680 3664 39744
rect 3728 39680 3736 39744
rect 3416 38656 3736 39680
rect 3416 38592 3424 38656
rect 3488 38592 3504 38656
rect 3568 38592 3584 38656
rect 3648 38592 3664 38656
rect 3728 38592 3736 38656
rect 3416 37568 3736 38592
rect 3416 37504 3424 37568
rect 3488 37504 3504 37568
rect 3568 37504 3584 37568
rect 3648 37504 3664 37568
rect 3728 37504 3736 37568
rect 3416 36480 3736 37504
rect 3416 36416 3424 36480
rect 3488 36416 3504 36480
rect 3568 36416 3584 36480
rect 3648 36416 3664 36480
rect 3728 36416 3736 36480
rect 3416 35392 3736 36416
rect 3416 35328 3424 35392
rect 3488 35328 3504 35392
rect 3568 35328 3584 35392
rect 3648 35328 3664 35392
rect 3728 35328 3736 35392
rect 3416 34304 3736 35328
rect 3416 34240 3424 34304
rect 3488 34240 3504 34304
rect 3568 34240 3584 34304
rect 3648 34240 3664 34304
rect 3728 34240 3736 34304
rect 3416 33216 3736 34240
rect 3416 33152 3424 33216
rect 3488 33152 3504 33216
rect 3568 33152 3584 33216
rect 3648 33152 3664 33216
rect 3728 33152 3736 33216
rect 3416 32128 3736 33152
rect 3416 32064 3424 32128
rect 3488 32064 3504 32128
rect 3568 32064 3584 32128
rect 3648 32064 3664 32128
rect 3728 32064 3736 32128
rect 3416 31040 3736 32064
rect 3416 30976 3424 31040
rect 3488 30976 3504 31040
rect 3568 30976 3584 31040
rect 3648 30976 3664 31040
rect 3728 30976 3736 31040
rect 3416 29952 3736 30976
rect 3926 30021 3986 41515
rect 5030 39133 5090 43147
rect 5579 43076 5645 43077
rect 5579 43012 5580 43076
rect 5644 43012 5645 43076
rect 5579 43011 5645 43012
rect 5395 42124 5461 42125
rect 5395 42060 5396 42124
rect 5460 42060 5461 42124
rect 5395 42059 5461 42060
rect 5027 39132 5093 39133
rect 5027 39068 5028 39132
rect 5092 39068 5093 39132
rect 5027 39067 5093 39068
rect 5398 36685 5458 42059
rect 5395 36684 5461 36685
rect 5395 36620 5396 36684
rect 5460 36620 5461 36684
rect 5395 36619 5461 36620
rect 4475 36004 4541 36005
rect 4475 35940 4476 36004
rect 4540 35940 4541 36004
rect 4475 35939 4541 35940
rect 4107 34236 4173 34237
rect 4107 34172 4108 34236
rect 4172 34172 4173 34236
rect 4107 34171 4173 34172
rect 3923 30020 3989 30021
rect 3923 29956 3924 30020
rect 3988 29956 3989 30020
rect 3923 29955 3989 29956
rect 3416 29888 3424 29952
rect 3488 29888 3504 29952
rect 3568 29888 3584 29952
rect 3648 29888 3664 29952
rect 3728 29888 3736 29952
rect 3416 28864 3736 29888
rect 3416 28800 3424 28864
rect 3488 28800 3504 28864
rect 3568 28800 3584 28864
rect 3648 28800 3664 28864
rect 3728 28800 3736 28864
rect 3416 27776 3736 28800
rect 3416 27712 3424 27776
rect 3488 27712 3504 27776
rect 3568 27712 3584 27776
rect 3648 27712 3664 27776
rect 3728 27712 3736 27776
rect 3416 26688 3736 27712
rect 3923 27708 3989 27709
rect 3923 27644 3924 27708
rect 3988 27644 3989 27708
rect 3923 27643 3989 27644
rect 3416 26624 3424 26688
rect 3488 26624 3504 26688
rect 3568 26624 3584 26688
rect 3648 26624 3664 26688
rect 3728 26624 3736 26688
rect 3416 25600 3736 26624
rect 3416 25536 3424 25600
rect 3488 25536 3504 25600
rect 3568 25536 3584 25600
rect 3648 25536 3664 25600
rect 3728 25536 3736 25600
rect 3416 24512 3736 25536
rect 3416 24448 3424 24512
rect 3488 24448 3504 24512
rect 3568 24448 3584 24512
rect 3648 24448 3664 24512
rect 3728 24448 3736 24512
rect 3416 23424 3736 24448
rect 3926 23626 3986 27643
rect 4110 27573 4170 34171
rect 4478 33557 4538 35939
rect 4843 34372 4909 34373
rect 4843 34308 4844 34372
rect 4908 34308 4909 34372
rect 4843 34307 4909 34308
rect 4475 33556 4541 33557
rect 4475 33492 4476 33556
rect 4540 33492 4541 33556
rect 4475 33491 4541 33492
rect 4291 33420 4357 33421
rect 4291 33356 4292 33420
rect 4356 33356 4357 33420
rect 4291 33355 4357 33356
rect 4294 29885 4354 33355
rect 4291 29884 4357 29885
rect 4291 29820 4292 29884
rect 4356 29820 4357 29884
rect 4291 29819 4357 29820
rect 4107 27572 4173 27573
rect 4107 27508 4108 27572
rect 4172 27508 4173 27572
rect 4107 27507 4173 27508
rect 4291 27300 4357 27301
rect 4291 27236 4292 27300
rect 4356 27236 4357 27300
rect 4291 27235 4357 27236
rect 4107 26348 4173 26349
rect 4107 26284 4108 26348
rect 4172 26284 4173 26348
rect 4107 26283 4173 26284
rect 4110 24309 4170 26283
rect 4107 24308 4173 24309
rect 4107 24244 4108 24308
rect 4172 24244 4173 24308
rect 4107 24243 4173 24244
rect 3926 23566 4170 23626
rect 3416 23360 3424 23424
rect 3488 23360 3504 23424
rect 3568 23360 3584 23424
rect 3648 23360 3664 23424
rect 3728 23360 3736 23424
rect 3187 23084 3253 23085
rect 3187 23020 3188 23084
rect 3252 23020 3253 23084
rect 3187 23019 3253 23020
rect 3416 22336 3736 23360
rect 3416 22272 3424 22336
rect 3488 22272 3504 22336
rect 3568 22272 3584 22336
rect 3648 22272 3664 22336
rect 3728 22272 3736 22336
rect 3006 22050 3250 22110
rect 3003 21724 3069 21725
rect 3003 21660 3004 21724
rect 3068 21660 3069 21724
rect 3003 21659 3069 21660
rect 2819 20092 2885 20093
rect 2819 20028 2820 20092
rect 2884 20028 2885 20092
rect 2819 20027 2885 20028
rect 2454 19350 2882 19410
rect 2451 18460 2517 18461
rect 2451 18396 2452 18460
rect 2516 18396 2517 18460
rect 2451 18395 2517 18396
rect 2635 18460 2701 18461
rect 2635 18396 2636 18460
rect 2700 18396 2701 18460
rect 2635 18395 2701 18396
rect 2267 18324 2333 18325
rect 2267 18260 2268 18324
rect 2332 18260 2333 18324
rect 2267 18259 2333 18260
rect 1899 17644 1965 17645
rect 1899 17580 1900 17644
rect 1964 17580 1965 17644
rect 1899 17579 1965 17580
rect 1715 16012 1781 16013
rect 1715 15948 1716 16012
rect 1780 15948 1781 16012
rect 1715 15947 1781 15948
rect 1902 15058 1962 17579
rect 2083 16556 2149 16557
rect 2083 16492 2084 16556
rect 2148 16492 2149 16556
rect 2083 16491 2149 16492
rect 1718 14998 1962 15058
rect 1347 14244 1413 14245
rect 1347 14180 1348 14244
rect 1412 14180 1413 14244
rect 1347 14179 1413 14180
rect 1531 10980 1597 10981
rect 1531 10916 1532 10980
rect 1596 10916 1597 10980
rect 1531 10915 1597 10916
rect 1347 9484 1413 9485
rect 1347 9420 1348 9484
rect 1412 9420 1413 9484
rect 1347 9419 1413 9420
rect 1350 7853 1410 9419
rect 1347 7852 1413 7853
rect 1347 7788 1348 7852
rect 1412 7788 1413 7852
rect 1347 7787 1413 7788
rect 1163 7580 1229 7581
rect 1163 7516 1164 7580
rect 1228 7516 1229 7580
rect 1163 7515 1229 7516
rect 1347 7308 1413 7309
rect 1347 7244 1348 7308
rect 1412 7244 1413 7308
rect 1347 7243 1413 7244
rect 979 1868 1045 1869
rect 979 1804 980 1868
rect 1044 1804 1045 1868
rect 979 1803 1045 1804
rect 1350 1461 1410 7243
rect 1534 4181 1594 10915
rect 1718 8941 1778 14998
rect 1899 14924 1965 14925
rect 1899 14860 1900 14924
rect 1964 14860 1965 14924
rect 1899 14859 1965 14860
rect 1902 10029 1962 14859
rect 1899 10028 1965 10029
rect 1899 9964 1900 10028
rect 1964 9964 1965 10028
rect 1899 9963 1965 9964
rect 1899 9076 1965 9077
rect 1899 9012 1900 9076
rect 1964 9012 1965 9076
rect 1899 9011 1965 9012
rect 1715 8940 1781 8941
rect 1715 8876 1716 8940
rect 1780 8876 1781 8940
rect 1715 8875 1781 8876
rect 1715 8124 1781 8125
rect 1715 8060 1716 8124
rect 1780 8060 1781 8124
rect 1715 8059 1781 8060
rect 1531 4180 1597 4181
rect 1531 4116 1532 4180
rect 1596 4116 1597 4180
rect 1531 4115 1597 4116
rect 1718 2549 1778 8059
rect 1902 7853 1962 9011
rect 1899 7852 1965 7853
rect 1899 7788 1900 7852
rect 1964 7788 1965 7852
rect 1899 7787 1965 7788
rect 2086 7717 2146 16491
rect 2267 12748 2333 12749
rect 2267 12684 2268 12748
rect 2332 12684 2333 12748
rect 2267 12683 2333 12684
rect 2270 11117 2330 12683
rect 2454 11797 2514 18395
rect 2638 14653 2698 18395
rect 2635 14652 2701 14653
rect 2635 14588 2636 14652
rect 2700 14588 2701 14652
rect 2635 14587 2701 14588
rect 2635 13292 2701 13293
rect 2635 13228 2636 13292
rect 2700 13228 2701 13292
rect 2635 13227 2701 13228
rect 2451 11796 2517 11797
rect 2451 11732 2452 11796
rect 2516 11732 2517 11796
rect 2451 11731 2517 11732
rect 2267 11116 2333 11117
rect 2267 11052 2268 11116
rect 2332 11052 2333 11116
rect 2267 11051 2333 11052
rect 2451 11116 2517 11117
rect 2451 11052 2452 11116
rect 2516 11052 2517 11116
rect 2451 11051 2517 11052
rect 2267 10708 2333 10709
rect 2267 10644 2268 10708
rect 2332 10644 2333 10708
rect 2267 10643 2333 10644
rect 2270 9077 2330 10643
rect 2267 9076 2333 9077
rect 2267 9012 2268 9076
rect 2332 9012 2333 9076
rect 2267 9011 2333 9012
rect 2267 8940 2333 8941
rect 2267 8876 2268 8940
rect 2332 8876 2333 8940
rect 2267 8875 2333 8876
rect 2083 7716 2149 7717
rect 2083 7652 2084 7716
rect 2148 7652 2149 7716
rect 2083 7651 2149 7652
rect 1715 2548 1781 2549
rect 1715 2484 1716 2548
rect 1780 2484 1781 2548
rect 1715 2483 1781 2484
rect 1347 1460 1413 1461
rect 1347 1396 1348 1460
rect 1412 1396 1413 1460
rect 1347 1395 1413 1396
rect 2270 1189 2330 8875
rect 2454 8397 2514 11051
rect 2638 10301 2698 13227
rect 2635 10300 2701 10301
rect 2635 10236 2636 10300
rect 2700 10236 2701 10300
rect 2635 10235 2701 10236
rect 2635 9620 2701 9621
rect 2635 9556 2636 9620
rect 2700 9556 2701 9620
rect 2635 9555 2701 9556
rect 2638 9210 2698 9555
rect 2822 9349 2882 19350
rect 3006 18461 3066 21659
rect 3190 20229 3250 22050
rect 3416 21248 3736 22272
rect 4110 22133 4170 23566
rect 4294 22269 4354 27235
rect 4291 22268 4357 22269
rect 4291 22204 4292 22268
rect 4356 22204 4357 22268
rect 4291 22203 4357 22204
rect 4107 22132 4173 22133
rect 4107 22068 4108 22132
rect 4172 22068 4173 22132
rect 4107 22067 4173 22068
rect 3416 21184 3424 21248
rect 3488 21184 3504 21248
rect 3568 21184 3584 21248
rect 3648 21184 3664 21248
rect 3728 21184 3736 21248
rect 3187 20228 3253 20229
rect 3187 20164 3188 20228
rect 3252 20164 3253 20228
rect 3187 20163 3253 20164
rect 3190 19413 3250 20163
rect 3416 20160 3736 21184
rect 3416 20096 3424 20160
rect 3488 20096 3504 20160
rect 3568 20096 3584 20160
rect 3648 20096 3664 20160
rect 3728 20096 3736 20160
rect 3187 19412 3253 19413
rect 3187 19348 3188 19412
rect 3252 19348 3253 19412
rect 3187 19347 3253 19348
rect 3416 19072 3736 20096
rect 3923 19548 3989 19549
rect 3923 19484 3924 19548
rect 3988 19484 3989 19548
rect 3923 19483 3989 19484
rect 3416 19008 3424 19072
rect 3488 19008 3504 19072
rect 3568 19008 3584 19072
rect 3648 19008 3664 19072
rect 3728 19008 3736 19072
rect 3003 18460 3069 18461
rect 3003 18396 3004 18460
rect 3068 18396 3069 18460
rect 3003 18395 3069 18396
rect 3416 17984 3736 19008
rect 3416 17920 3424 17984
rect 3488 17920 3504 17984
rect 3568 17920 3584 17984
rect 3648 17920 3664 17984
rect 3728 17920 3736 17984
rect 3416 16896 3736 17920
rect 3416 16832 3424 16896
rect 3488 16832 3504 16896
rect 3568 16832 3584 16896
rect 3648 16832 3664 16896
rect 3728 16832 3736 16896
rect 3187 16148 3253 16149
rect 3187 16084 3188 16148
rect 3252 16084 3253 16148
rect 3187 16083 3253 16084
rect 3003 14652 3069 14653
rect 3003 14588 3004 14652
rect 3068 14588 3069 14652
rect 3003 14587 3069 14588
rect 3006 10709 3066 14587
rect 3003 10708 3069 10709
rect 3003 10644 3004 10708
rect 3068 10644 3069 10708
rect 3003 10643 3069 10644
rect 3003 10572 3069 10573
rect 3003 10508 3004 10572
rect 3068 10508 3069 10572
rect 3003 10507 3069 10508
rect 2819 9348 2885 9349
rect 2819 9284 2820 9348
rect 2884 9284 2885 9348
rect 2819 9283 2885 9284
rect 2638 9150 2882 9210
rect 2635 8940 2701 8941
rect 2635 8876 2636 8940
rect 2700 8876 2701 8940
rect 2635 8875 2701 8876
rect 2451 8396 2517 8397
rect 2451 8332 2452 8396
rect 2516 8332 2517 8396
rect 2451 8331 2517 8332
rect 2638 2685 2698 8875
rect 2822 7853 2882 9150
rect 3006 8533 3066 10507
rect 3190 9485 3250 16083
rect 3416 15808 3736 16832
rect 3926 16285 3986 19483
rect 4110 17917 4170 22067
rect 4107 17916 4173 17917
rect 4107 17852 4108 17916
rect 4172 17852 4173 17916
rect 4107 17851 4173 17852
rect 4107 16420 4173 16421
rect 4107 16356 4108 16420
rect 4172 16356 4173 16420
rect 4107 16355 4173 16356
rect 3923 16284 3989 16285
rect 3923 16220 3924 16284
rect 3988 16220 3989 16284
rect 3923 16219 3989 16220
rect 4110 16010 4170 16355
rect 3416 15744 3424 15808
rect 3488 15744 3504 15808
rect 3568 15744 3584 15808
rect 3648 15744 3664 15808
rect 3728 15744 3736 15808
rect 3416 14720 3736 15744
rect 3416 14656 3424 14720
rect 3488 14656 3504 14720
rect 3568 14656 3584 14720
rect 3648 14656 3664 14720
rect 3728 14656 3736 14720
rect 3416 13632 3736 14656
rect 3416 13568 3424 13632
rect 3488 13568 3504 13632
rect 3568 13568 3584 13632
rect 3648 13568 3664 13632
rect 3728 13568 3736 13632
rect 3416 12544 3736 13568
rect 3416 12480 3424 12544
rect 3488 12480 3504 12544
rect 3568 12480 3584 12544
rect 3648 12480 3664 12544
rect 3728 12480 3736 12544
rect 3416 11456 3736 12480
rect 3416 11392 3424 11456
rect 3488 11392 3504 11456
rect 3568 11392 3584 11456
rect 3648 11392 3664 11456
rect 3728 11392 3736 11456
rect 3416 10368 3736 11392
rect 3926 15950 4170 16010
rect 3926 10709 3986 15950
rect 4291 14516 4357 14517
rect 4291 14452 4292 14516
rect 4356 14452 4357 14516
rect 4291 14451 4357 14452
rect 4107 14244 4173 14245
rect 4107 14180 4108 14244
rect 4172 14180 4173 14244
rect 4107 14179 4173 14180
rect 4110 13701 4170 14179
rect 4107 13700 4173 13701
rect 4107 13636 4108 13700
rect 4172 13636 4173 13700
rect 4107 13635 4173 13636
rect 4107 13292 4173 13293
rect 4107 13228 4108 13292
rect 4172 13228 4173 13292
rect 4107 13227 4173 13228
rect 4110 11070 4170 13227
rect 4294 11525 4354 14451
rect 4291 11524 4357 11525
rect 4291 11460 4292 11524
rect 4356 11460 4357 11524
rect 4291 11459 4357 11460
rect 4064 11010 4170 11070
rect 3923 10708 3989 10709
rect 3923 10644 3924 10708
rect 3988 10644 3989 10708
rect 3923 10643 3989 10644
rect 4064 10570 4124 11010
rect 4291 10980 4357 10981
rect 4291 10916 4292 10980
rect 4356 10916 4357 10980
rect 4291 10915 4357 10916
rect 3416 10304 3424 10368
rect 3488 10304 3504 10368
rect 3568 10304 3584 10368
rect 3648 10304 3664 10368
rect 3728 10304 3736 10368
rect 3187 9484 3253 9485
rect 3187 9420 3188 9484
rect 3252 9420 3253 9484
rect 3187 9419 3253 9420
rect 3416 9280 3736 10304
rect 3416 9216 3424 9280
rect 3488 9216 3504 9280
rect 3568 9216 3584 9280
rect 3648 9216 3664 9280
rect 3728 9216 3736 9280
rect 3003 8532 3069 8533
rect 3003 8468 3004 8532
rect 3068 8468 3069 8532
rect 3003 8467 3069 8468
rect 3187 8532 3253 8533
rect 3187 8468 3188 8532
rect 3252 8468 3253 8532
rect 3187 8467 3253 8468
rect 2819 7852 2885 7853
rect 2819 7788 2820 7852
rect 2884 7788 2885 7852
rect 3190 7850 3250 8467
rect 2819 7787 2885 7788
rect 3006 7790 3250 7850
rect 3416 8192 3736 9216
rect 3416 8128 3424 8192
rect 3488 8128 3504 8192
rect 3568 8128 3584 8192
rect 3648 8128 3664 8192
rect 3728 8128 3736 8192
rect 3006 5949 3066 7790
rect 3187 7444 3253 7445
rect 3187 7380 3188 7444
rect 3252 7380 3253 7444
rect 3187 7379 3253 7380
rect 3003 5948 3069 5949
rect 3003 5884 3004 5948
rect 3068 5884 3069 5948
rect 3003 5883 3069 5884
rect 3190 4045 3250 7379
rect 3416 7104 3736 8128
rect 3926 10510 4124 10570
rect 3926 7853 3986 10510
rect 4107 10300 4173 10301
rect 4107 10236 4108 10300
rect 4172 10236 4173 10300
rect 4107 10235 4173 10236
rect 4110 9077 4170 10235
rect 4107 9076 4173 9077
rect 4107 9012 4108 9076
rect 4172 9012 4173 9076
rect 4107 9011 4173 9012
rect 4107 8124 4173 8125
rect 4107 8060 4108 8124
rect 4172 8060 4173 8124
rect 4107 8059 4173 8060
rect 3923 7852 3989 7853
rect 3923 7788 3924 7852
rect 3988 7788 3989 7852
rect 3923 7787 3989 7788
rect 3416 7040 3424 7104
rect 3488 7040 3504 7104
rect 3568 7040 3584 7104
rect 3648 7040 3664 7104
rect 3728 7040 3736 7104
rect 3416 6016 3736 7040
rect 4110 6493 4170 8059
rect 4107 6492 4173 6493
rect 4107 6428 4108 6492
rect 4172 6428 4173 6492
rect 4107 6427 4173 6428
rect 3416 5952 3424 6016
rect 3488 5952 3504 6016
rect 3568 5952 3584 6016
rect 3648 5952 3664 6016
rect 3728 5952 3736 6016
rect 3416 4928 3736 5952
rect 4294 5674 4354 10915
rect 4478 9621 4538 33491
rect 4659 32196 4725 32197
rect 4659 32132 4660 32196
rect 4724 32132 4725 32196
rect 4659 32131 4725 32132
rect 4662 31109 4722 32131
rect 4659 31108 4725 31109
rect 4659 31044 4660 31108
rect 4724 31044 4725 31108
rect 4659 31043 4725 31044
rect 4659 29340 4725 29341
rect 4659 29276 4660 29340
rect 4724 29276 4725 29340
rect 4659 29275 4725 29276
rect 4662 24309 4722 29275
rect 4659 24308 4725 24309
rect 4659 24244 4660 24308
rect 4724 24244 4725 24308
rect 4659 24243 4725 24244
rect 4662 23490 4722 24243
rect 4846 23629 4906 34307
rect 5027 31924 5093 31925
rect 5027 31860 5028 31924
rect 5092 31860 5093 31924
rect 5027 31859 5093 31860
rect 5030 29341 5090 31859
rect 5211 31108 5277 31109
rect 5211 31044 5212 31108
rect 5276 31044 5277 31108
rect 5211 31043 5277 31044
rect 5395 31108 5461 31109
rect 5395 31044 5396 31108
rect 5460 31044 5461 31108
rect 5395 31043 5461 31044
rect 5214 30837 5274 31043
rect 5211 30836 5277 30837
rect 5211 30772 5212 30836
rect 5276 30772 5277 30836
rect 5211 30771 5277 30772
rect 5214 29749 5274 30771
rect 5211 29748 5277 29749
rect 5211 29684 5212 29748
rect 5276 29684 5277 29748
rect 5211 29683 5277 29684
rect 5027 29340 5093 29341
rect 5027 29276 5028 29340
rect 5092 29276 5093 29340
rect 5027 29275 5093 29276
rect 5030 29010 5090 29275
rect 5030 28950 5274 29010
rect 5027 28116 5093 28117
rect 5027 28052 5028 28116
rect 5092 28052 5093 28116
rect 5027 28051 5093 28052
rect 5030 25533 5090 28051
rect 5027 25532 5093 25533
rect 5027 25468 5028 25532
rect 5092 25468 5093 25532
rect 5027 25467 5093 25468
rect 5214 23901 5274 28950
rect 5398 25941 5458 31043
rect 5395 25940 5461 25941
rect 5395 25876 5396 25940
rect 5460 25876 5461 25940
rect 5395 25875 5461 25876
rect 5027 23900 5093 23901
rect 5027 23836 5028 23900
rect 5092 23836 5093 23900
rect 5027 23835 5093 23836
rect 5211 23900 5277 23901
rect 5211 23836 5212 23900
rect 5276 23836 5277 23900
rect 5211 23835 5277 23836
rect 4843 23628 4909 23629
rect 4843 23564 4844 23628
rect 4908 23564 4909 23628
rect 4843 23563 4909 23564
rect 4662 23430 4906 23490
rect 4659 23356 4725 23357
rect 4659 23292 4660 23356
rect 4724 23292 4725 23356
rect 4659 23291 4725 23292
rect 4662 17509 4722 23291
rect 4846 23085 4906 23430
rect 4843 23084 4909 23085
rect 4843 23020 4844 23084
rect 4908 23020 4909 23084
rect 4843 23019 4909 23020
rect 4846 20773 4906 23019
rect 4843 20772 4909 20773
rect 4843 20708 4844 20772
rect 4908 20708 4909 20772
rect 4843 20707 4909 20708
rect 4659 17508 4725 17509
rect 4659 17444 4660 17508
rect 4724 17444 4725 17508
rect 4659 17443 4725 17444
rect 5030 17098 5090 23835
rect 5211 23628 5277 23629
rect 5211 23564 5212 23628
rect 5276 23564 5277 23628
rect 5211 23563 5277 23564
rect 5214 20501 5274 23563
rect 5398 21181 5458 25875
rect 5582 22813 5642 43011
rect 5888 42464 6208 43488
rect 5888 42400 5896 42464
rect 5960 42400 5976 42464
rect 6040 42400 6056 42464
rect 6120 42400 6136 42464
rect 6200 42400 6208 42464
rect 5888 41376 6208 42400
rect 8361 43008 8681 43568
rect 8361 42944 8369 43008
rect 8433 42944 8449 43008
rect 8513 42944 8529 43008
rect 8593 42944 8609 43008
rect 8673 42944 8681 43008
rect 7419 42260 7485 42261
rect 7419 42196 7420 42260
rect 7484 42196 7485 42260
rect 7419 42195 7485 42196
rect 6499 41716 6565 41717
rect 6499 41652 6500 41716
rect 6564 41652 6565 41716
rect 6499 41651 6565 41652
rect 5888 41312 5896 41376
rect 5960 41312 5976 41376
rect 6040 41312 6056 41376
rect 6120 41312 6136 41376
rect 6200 41312 6208 41376
rect 5888 40288 6208 41312
rect 5888 40224 5896 40288
rect 5960 40224 5976 40288
rect 6040 40224 6056 40288
rect 6120 40224 6136 40288
rect 6200 40224 6208 40288
rect 5888 39200 6208 40224
rect 5888 39136 5896 39200
rect 5960 39136 5976 39200
rect 6040 39136 6056 39200
rect 6120 39136 6136 39200
rect 6200 39136 6208 39200
rect 5888 38112 6208 39136
rect 5888 38048 5896 38112
rect 5960 38048 5976 38112
rect 6040 38048 6056 38112
rect 6120 38048 6136 38112
rect 6200 38048 6208 38112
rect 5888 37024 6208 38048
rect 5888 36960 5896 37024
rect 5960 36960 5976 37024
rect 6040 36960 6056 37024
rect 6120 36960 6136 37024
rect 6200 36960 6208 37024
rect 5888 35936 6208 36960
rect 5888 35872 5896 35936
rect 5960 35872 5976 35936
rect 6040 35872 6056 35936
rect 6120 35872 6136 35936
rect 6200 35872 6208 35936
rect 5888 34848 6208 35872
rect 5888 34784 5896 34848
rect 5960 34784 5976 34848
rect 6040 34784 6056 34848
rect 6120 34784 6136 34848
rect 6200 34784 6208 34848
rect 5888 33760 6208 34784
rect 6502 34509 6562 41651
rect 6867 37364 6933 37365
rect 6867 37300 6868 37364
rect 6932 37300 6933 37364
rect 6867 37299 6933 37300
rect 6499 34508 6565 34509
rect 6499 34444 6500 34508
rect 6564 34444 6565 34508
rect 6499 34443 6565 34444
rect 6499 33964 6565 33965
rect 6499 33900 6500 33964
rect 6564 33900 6565 33964
rect 6499 33899 6565 33900
rect 6315 33828 6381 33829
rect 6315 33764 6316 33828
rect 6380 33764 6381 33828
rect 6315 33763 6381 33764
rect 5888 33696 5896 33760
rect 5960 33696 5976 33760
rect 6040 33696 6056 33760
rect 6120 33696 6136 33760
rect 6200 33696 6208 33760
rect 5888 32672 6208 33696
rect 6318 32877 6378 33763
rect 6315 32876 6381 32877
rect 6315 32812 6316 32876
rect 6380 32812 6381 32876
rect 6315 32811 6381 32812
rect 5888 32608 5896 32672
rect 5960 32608 5976 32672
rect 6040 32608 6056 32672
rect 6120 32608 6136 32672
rect 6200 32608 6208 32672
rect 5888 31584 6208 32608
rect 5888 31520 5896 31584
rect 5960 31520 5976 31584
rect 6040 31520 6056 31584
rect 6120 31520 6136 31584
rect 6200 31520 6208 31584
rect 5888 30496 6208 31520
rect 5888 30432 5896 30496
rect 5960 30432 5976 30496
rect 6040 30432 6056 30496
rect 6120 30432 6136 30496
rect 6200 30432 6208 30496
rect 5888 29408 6208 30432
rect 5888 29344 5896 29408
rect 5960 29344 5976 29408
rect 6040 29344 6056 29408
rect 6120 29344 6136 29408
rect 6200 29344 6208 29408
rect 5888 28320 6208 29344
rect 5888 28256 5896 28320
rect 5960 28256 5976 28320
rect 6040 28256 6056 28320
rect 6120 28256 6136 28320
rect 6200 28256 6208 28320
rect 5888 27232 6208 28256
rect 5888 27168 5896 27232
rect 5960 27168 5976 27232
rect 6040 27168 6056 27232
rect 6120 27168 6136 27232
rect 6200 27168 6208 27232
rect 5888 26144 6208 27168
rect 5888 26080 5896 26144
rect 5960 26080 5976 26144
rect 6040 26080 6056 26144
rect 6120 26080 6136 26144
rect 6200 26080 6208 26144
rect 5888 25056 6208 26080
rect 5888 24992 5896 25056
rect 5960 24992 5976 25056
rect 6040 24992 6056 25056
rect 6120 24992 6136 25056
rect 6200 24992 6208 25056
rect 5888 23968 6208 24992
rect 6318 24581 6378 32811
rect 6502 31770 6562 33899
rect 6502 31710 6746 31770
rect 6499 25804 6565 25805
rect 6499 25740 6500 25804
rect 6564 25740 6565 25804
rect 6499 25739 6565 25740
rect 6315 24580 6381 24581
rect 6315 24516 6316 24580
rect 6380 24516 6381 24580
rect 6315 24515 6381 24516
rect 6315 24308 6381 24309
rect 6315 24244 6316 24308
rect 6380 24244 6381 24308
rect 6315 24243 6381 24244
rect 5888 23904 5896 23968
rect 5960 23904 5976 23968
rect 6040 23904 6056 23968
rect 6120 23904 6136 23968
rect 6200 23904 6208 23968
rect 5888 22880 6208 23904
rect 5888 22816 5896 22880
rect 5960 22816 5976 22880
rect 6040 22816 6056 22880
rect 6120 22816 6136 22880
rect 6200 22816 6208 22880
rect 5579 22812 5645 22813
rect 5579 22748 5580 22812
rect 5644 22748 5645 22812
rect 5579 22747 5645 22748
rect 5888 21792 6208 22816
rect 5888 21728 5896 21792
rect 5960 21728 5976 21792
rect 6040 21728 6056 21792
rect 6120 21728 6136 21792
rect 6200 21728 6208 21792
rect 5579 21724 5645 21725
rect 5579 21660 5580 21724
rect 5644 21722 5645 21724
rect 5644 21662 5826 21722
rect 5644 21660 5645 21662
rect 5579 21659 5645 21660
rect 5395 21180 5461 21181
rect 5395 21116 5396 21180
rect 5460 21116 5461 21180
rect 5395 21115 5461 21116
rect 5211 20500 5277 20501
rect 5211 20436 5212 20500
rect 5276 20436 5277 20500
rect 5211 20435 5277 20436
rect 5579 20500 5645 20501
rect 5579 20436 5580 20500
rect 5644 20436 5645 20500
rect 5579 20435 5645 20436
rect 5395 20092 5461 20093
rect 5395 20028 5396 20092
rect 5460 20028 5461 20092
rect 5395 20027 5461 20028
rect 4662 17038 5090 17098
rect 4475 9620 4541 9621
rect 4475 9556 4476 9620
rect 4540 9556 4541 9620
rect 4475 9555 4541 9556
rect 4475 8940 4541 8941
rect 4475 8876 4476 8940
rect 4540 8876 4541 8940
rect 4475 8875 4541 8876
rect 4478 6357 4538 8875
rect 4475 6356 4541 6357
rect 4475 6292 4476 6356
rect 4540 6292 4541 6356
rect 4475 6291 4541 6292
rect 3416 4864 3424 4928
rect 3488 4864 3504 4928
rect 3568 4864 3584 4928
rect 3648 4864 3664 4928
rect 3728 4864 3736 4928
rect 3187 4044 3253 4045
rect 3187 3980 3188 4044
rect 3252 3980 3253 4044
rect 3187 3979 3253 3980
rect 3416 3840 3736 4864
rect 3926 5614 4354 5674
rect 3926 4170 3986 5614
rect 3926 4110 4354 4170
rect 3416 3776 3424 3840
rect 3488 3776 3504 3840
rect 3568 3776 3584 3840
rect 3648 3776 3664 3840
rect 3728 3776 3736 3840
rect 3416 2752 3736 3776
rect 3416 2688 3424 2752
rect 3488 2688 3504 2752
rect 3568 2688 3584 2752
rect 3648 2688 3664 2752
rect 3728 2688 3736 2752
rect 2635 2684 2701 2685
rect 2635 2620 2636 2684
rect 2700 2620 2701 2684
rect 2635 2619 2701 2620
rect 3416 1664 3736 2688
rect 4294 2685 4354 4110
rect 4475 3772 4541 3773
rect 4475 3708 4476 3772
rect 4540 3708 4541 3772
rect 4475 3707 4541 3708
rect 4291 2684 4357 2685
rect 4291 2620 4292 2684
rect 4356 2620 4357 2684
rect 4291 2619 4357 2620
rect 4478 2413 4538 3707
rect 4662 2413 4722 17038
rect 5027 16964 5093 16965
rect 5027 16900 5028 16964
rect 5092 16900 5093 16964
rect 5027 16899 5093 16900
rect 4843 15604 4909 15605
rect 4843 15540 4844 15604
rect 4908 15540 4909 15604
rect 4843 15539 4909 15540
rect 4846 13021 4906 15539
rect 5030 13293 5090 16899
rect 5398 14789 5458 20027
rect 5582 18461 5642 20435
rect 5579 18460 5645 18461
rect 5579 18396 5580 18460
rect 5644 18396 5645 18460
rect 5579 18395 5645 18396
rect 5582 15605 5642 18395
rect 5579 15604 5645 15605
rect 5579 15540 5580 15604
rect 5644 15540 5645 15604
rect 5579 15539 5645 15540
rect 5579 15332 5645 15333
rect 5579 15268 5580 15332
rect 5644 15268 5645 15332
rect 5579 15267 5645 15268
rect 5395 14788 5461 14789
rect 5395 14724 5396 14788
rect 5460 14724 5461 14788
rect 5395 14723 5461 14724
rect 5211 14652 5277 14653
rect 5211 14588 5212 14652
rect 5276 14588 5277 14652
rect 5211 14587 5277 14588
rect 5027 13292 5093 13293
rect 5027 13228 5028 13292
rect 5092 13228 5093 13292
rect 5027 13227 5093 13228
rect 4843 13020 4909 13021
rect 4843 12956 4844 13020
rect 4908 12956 4909 13020
rect 4843 12955 4909 12956
rect 4843 12068 4909 12069
rect 4843 12004 4844 12068
rect 4908 12004 4909 12068
rect 4843 12003 4909 12004
rect 4846 11117 4906 12003
rect 4843 11116 4909 11117
rect 4843 11052 4844 11116
rect 4908 11052 4909 11116
rect 4843 11051 4909 11052
rect 4843 10980 4909 10981
rect 4843 10916 4844 10980
rect 4908 10916 4909 10980
rect 4843 10915 4909 10916
rect 4846 4453 4906 10915
rect 5030 10709 5090 13227
rect 5027 10708 5093 10709
rect 5027 10644 5028 10708
rect 5092 10644 5093 10708
rect 5027 10643 5093 10644
rect 5030 9485 5090 10643
rect 5027 9484 5093 9485
rect 5027 9420 5028 9484
rect 5092 9420 5093 9484
rect 5027 9419 5093 9420
rect 5027 9348 5093 9349
rect 5027 9284 5028 9348
rect 5092 9284 5093 9348
rect 5027 9283 5093 9284
rect 5030 6085 5090 9283
rect 5214 6901 5274 14587
rect 5582 13429 5642 15267
rect 5579 13428 5645 13429
rect 5579 13364 5580 13428
rect 5644 13364 5645 13428
rect 5579 13363 5645 13364
rect 5395 12612 5461 12613
rect 5395 12548 5396 12612
rect 5460 12548 5461 12612
rect 5766 12610 5826 21662
rect 5395 12547 5461 12548
rect 5582 12550 5826 12610
rect 5888 20704 6208 21728
rect 5888 20640 5896 20704
rect 5960 20640 5976 20704
rect 6040 20640 6056 20704
rect 6120 20640 6136 20704
rect 6200 20640 6208 20704
rect 5888 19616 6208 20640
rect 5888 19552 5896 19616
rect 5960 19552 5976 19616
rect 6040 19552 6056 19616
rect 6120 19552 6136 19616
rect 6200 19552 6208 19616
rect 5888 18528 6208 19552
rect 5888 18464 5896 18528
rect 5960 18464 5976 18528
rect 6040 18464 6056 18528
rect 6120 18464 6136 18528
rect 6200 18464 6208 18528
rect 5888 17440 6208 18464
rect 6318 18325 6378 24243
rect 6502 20773 6562 25739
rect 6686 24853 6746 31710
rect 6870 31653 6930 37299
rect 7422 34373 7482 42195
rect 8361 41920 8681 42944
rect 10833 43552 11153 43568
rect 10833 43488 10841 43552
rect 10905 43488 10921 43552
rect 10985 43488 11001 43552
rect 11065 43488 11081 43552
rect 11145 43488 11153 43552
rect 10547 42940 10613 42941
rect 10547 42876 10548 42940
rect 10612 42876 10613 42940
rect 10547 42875 10613 42876
rect 9443 42124 9509 42125
rect 9443 42060 9444 42124
rect 9508 42060 9509 42124
rect 9443 42059 9509 42060
rect 8361 41856 8369 41920
rect 8433 41856 8449 41920
rect 8513 41856 8529 41920
rect 8593 41856 8609 41920
rect 8673 41856 8681 41920
rect 8361 40832 8681 41856
rect 9259 41580 9325 41581
rect 9259 41516 9260 41580
rect 9324 41516 9325 41580
rect 9259 41515 9325 41516
rect 8361 40768 8369 40832
rect 8433 40768 8449 40832
rect 8513 40768 8529 40832
rect 8593 40768 8609 40832
rect 8673 40768 8681 40832
rect 7971 40084 8037 40085
rect 7971 40020 7972 40084
rect 8036 40020 8037 40084
rect 7971 40019 8037 40020
rect 7787 35188 7853 35189
rect 7787 35124 7788 35188
rect 7852 35124 7853 35188
rect 7787 35123 7853 35124
rect 7419 34372 7485 34373
rect 7419 34308 7420 34372
rect 7484 34308 7485 34372
rect 7419 34307 7485 34308
rect 7419 34236 7485 34237
rect 7419 34172 7420 34236
rect 7484 34172 7485 34236
rect 7419 34171 7485 34172
rect 7603 34236 7669 34237
rect 7603 34172 7604 34236
rect 7668 34172 7669 34236
rect 7603 34171 7669 34172
rect 6867 31652 6933 31653
rect 6867 31588 6868 31652
rect 6932 31588 6933 31652
rect 7235 31652 7301 31653
rect 7235 31650 7236 31652
rect 6867 31587 6933 31588
rect 7054 31590 7236 31650
rect 6867 26212 6933 26213
rect 6867 26148 6868 26212
rect 6932 26148 6933 26212
rect 6867 26147 6933 26148
rect 6683 24852 6749 24853
rect 6683 24788 6684 24852
rect 6748 24788 6749 24852
rect 6683 24787 6749 24788
rect 6683 21724 6749 21725
rect 6683 21660 6684 21724
rect 6748 21660 6749 21724
rect 6683 21659 6749 21660
rect 6499 20772 6565 20773
rect 6499 20708 6500 20772
rect 6564 20708 6565 20772
rect 6499 20707 6565 20708
rect 6315 18324 6381 18325
rect 6315 18260 6316 18324
rect 6380 18260 6381 18324
rect 6315 18259 6381 18260
rect 5888 17376 5896 17440
rect 5960 17376 5976 17440
rect 6040 17376 6056 17440
rect 6120 17376 6136 17440
rect 6200 17376 6208 17440
rect 5888 16352 6208 17376
rect 6502 16421 6562 20707
rect 6686 18869 6746 21659
rect 6870 20909 6930 26147
rect 7054 23493 7114 31590
rect 7235 31588 7236 31590
rect 7300 31588 7301 31652
rect 7235 31587 7301 31588
rect 7422 31245 7482 34171
rect 7419 31244 7485 31245
rect 7419 31180 7420 31244
rect 7484 31180 7485 31244
rect 7419 31179 7485 31180
rect 7419 29884 7485 29885
rect 7419 29820 7420 29884
rect 7484 29820 7485 29884
rect 7419 29819 7485 29820
rect 7422 29010 7482 29819
rect 7238 28950 7482 29010
rect 7051 23492 7117 23493
rect 7051 23428 7052 23492
rect 7116 23428 7117 23492
rect 7051 23427 7117 23428
rect 7238 23354 7298 28950
rect 7419 28796 7485 28797
rect 7419 28732 7420 28796
rect 7484 28732 7485 28796
rect 7419 28731 7485 28732
rect 7422 23901 7482 28731
rect 7419 23900 7485 23901
rect 7419 23836 7420 23900
rect 7484 23836 7485 23900
rect 7419 23835 7485 23836
rect 7054 23294 7298 23354
rect 6867 20908 6933 20909
rect 6867 20844 6868 20908
rect 6932 20844 6933 20908
rect 6867 20843 6933 20844
rect 6867 20772 6933 20773
rect 6867 20708 6868 20772
rect 6932 20708 6933 20772
rect 6867 20707 6933 20708
rect 6683 18868 6749 18869
rect 6683 18804 6684 18868
rect 6748 18804 6749 18868
rect 6683 18803 6749 18804
rect 6683 18188 6749 18189
rect 6683 18124 6684 18188
rect 6748 18124 6749 18188
rect 6683 18123 6749 18124
rect 6499 16420 6565 16421
rect 6499 16356 6500 16420
rect 6564 16356 6565 16420
rect 6499 16355 6565 16356
rect 5888 16288 5896 16352
rect 5960 16288 5976 16352
rect 6040 16288 6056 16352
rect 6120 16288 6136 16352
rect 6200 16288 6208 16352
rect 5888 15264 6208 16288
rect 6315 16148 6381 16149
rect 6315 16084 6316 16148
rect 6380 16084 6381 16148
rect 6315 16083 6381 16084
rect 5888 15200 5896 15264
rect 5960 15200 5976 15264
rect 6040 15200 6056 15264
rect 6120 15200 6136 15264
rect 6200 15200 6208 15264
rect 5888 14176 6208 15200
rect 6318 15210 6378 16083
rect 6318 15150 6562 15210
rect 5888 14112 5896 14176
rect 5960 14112 5976 14176
rect 6040 14112 6056 14176
rect 6120 14112 6136 14176
rect 6200 14112 6208 14176
rect 5888 13088 6208 14112
rect 6315 14108 6381 14109
rect 6315 14044 6316 14108
rect 6380 14044 6381 14108
rect 6315 14043 6381 14044
rect 5888 13024 5896 13088
rect 5960 13024 5976 13088
rect 6040 13024 6056 13088
rect 6120 13024 6136 13088
rect 6200 13024 6208 13088
rect 5398 12066 5458 12547
rect 5582 12341 5642 12550
rect 5717 12476 5783 12477
rect 5717 12412 5718 12476
rect 5782 12474 5783 12476
rect 5782 12412 5826 12474
rect 5717 12411 5826 12412
rect 5579 12340 5645 12341
rect 5579 12276 5580 12340
rect 5644 12276 5645 12340
rect 5579 12275 5645 12276
rect 5398 12006 5642 12066
rect 5395 11796 5461 11797
rect 5395 11732 5396 11796
rect 5460 11732 5461 11796
rect 5395 11731 5461 11732
rect 5398 10301 5458 11731
rect 5582 10437 5642 12006
rect 5579 10436 5645 10437
rect 5579 10372 5580 10436
rect 5644 10372 5645 10436
rect 5579 10371 5645 10372
rect 5395 10300 5461 10301
rect 5395 10236 5396 10300
rect 5460 10236 5461 10300
rect 5395 10235 5461 10236
rect 5398 9690 5458 10235
rect 5398 9630 5642 9690
rect 5395 9076 5461 9077
rect 5395 9012 5396 9076
rect 5460 9012 5461 9076
rect 5395 9011 5461 9012
rect 5398 8261 5458 9011
rect 5395 8260 5461 8261
rect 5395 8196 5396 8260
rect 5460 8196 5461 8260
rect 5395 8195 5461 8196
rect 5395 7580 5461 7581
rect 5395 7516 5396 7580
rect 5460 7516 5461 7580
rect 5395 7515 5461 7516
rect 5211 6900 5277 6901
rect 5211 6836 5212 6900
rect 5276 6836 5277 6900
rect 5211 6835 5277 6836
rect 5027 6084 5093 6085
rect 5027 6020 5028 6084
rect 5092 6020 5093 6084
rect 5027 6019 5093 6020
rect 5211 5132 5277 5133
rect 5211 5068 5212 5132
rect 5276 5068 5277 5132
rect 5211 5067 5277 5068
rect 4843 4452 4909 4453
rect 4843 4388 4844 4452
rect 4908 4388 4909 4452
rect 4843 4387 4909 4388
rect 5214 3093 5274 5067
rect 5398 4722 5458 7515
rect 5582 5677 5642 9630
rect 5579 5676 5645 5677
rect 5579 5612 5580 5676
rect 5644 5612 5645 5676
rect 5579 5611 5645 5612
rect 5579 4724 5645 4725
rect 5579 4722 5580 4724
rect 5398 4662 5580 4722
rect 5579 4660 5580 4662
rect 5644 4660 5645 4724
rect 5579 4659 5645 4660
rect 5579 4180 5645 4181
rect 5579 4116 5580 4180
rect 5644 4116 5645 4180
rect 5579 4115 5645 4116
rect 5582 3093 5642 4115
rect 5211 3092 5277 3093
rect 5211 3028 5212 3092
rect 5276 3028 5277 3092
rect 5211 3027 5277 3028
rect 5579 3092 5645 3093
rect 5579 3028 5580 3092
rect 5644 3028 5645 3092
rect 5579 3027 5645 3028
rect 4475 2412 4541 2413
rect 4475 2348 4476 2412
rect 4540 2348 4541 2412
rect 4475 2347 4541 2348
rect 4659 2412 4725 2413
rect 4659 2348 4660 2412
rect 4724 2348 4725 2412
rect 4659 2347 4725 2348
rect 5579 2412 5645 2413
rect 5579 2348 5580 2412
rect 5644 2410 5645 2412
rect 5766 2410 5826 12411
rect 5644 2350 5826 2410
rect 5888 12000 6208 13024
rect 5888 11936 5896 12000
rect 5960 11936 5976 12000
rect 6040 11936 6056 12000
rect 6120 11936 6136 12000
rect 6200 11936 6208 12000
rect 5888 10912 6208 11936
rect 5888 10848 5896 10912
rect 5960 10848 5976 10912
rect 6040 10848 6056 10912
rect 6120 10848 6136 10912
rect 6200 10848 6208 10912
rect 5888 9824 6208 10848
rect 5888 9760 5896 9824
rect 5960 9760 5976 9824
rect 6040 9760 6056 9824
rect 6120 9760 6136 9824
rect 6200 9760 6208 9824
rect 5888 8736 6208 9760
rect 5888 8672 5896 8736
rect 5960 8672 5976 8736
rect 6040 8672 6056 8736
rect 6120 8672 6136 8736
rect 6200 8672 6208 8736
rect 5888 7648 6208 8672
rect 5888 7584 5896 7648
rect 5960 7584 5976 7648
rect 6040 7584 6056 7648
rect 6120 7584 6136 7648
rect 6200 7584 6208 7648
rect 5888 6560 6208 7584
rect 5888 6496 5896 6560
rect 5960 6496 5976 6560
rect 6040 6496 6056 6560
rect 6120 6496 6136 6560
rect 6200 6496 6208 6560
rect 5888 5472 6208 6496
rect 5888 5408 5896 5472
rect 5960 5408 5976 5472
rect 6040 5408 6056 5472
rect 6120 5408 6136 5472
rect 6200 5408 6208 5472
rect 5888 4384 6208 5408
rect 5888 4320 5896 4384
rect 5960 4320 5976 4384
rect 6040 4320 6056 4384
rect 6120 4320 6136 4384
rect 6200 4320 6208 4384
rect 5888 3296 6208 4320
rect 5888 3232 5896 3296
rect 5960 3232 5976 3296
rect 6040 3232 6056 3296
rect 6120 3232 6136 3296
rect 6200 3232 6208 3296
rect 5644 2348 5645 2350
rect 5579 2347 5645 2348
rect 3416 1600 3424 1664
rect 3488 1600 3504 1664
rect 3568 1600 3584 1664
rect 3648 1600 3664 1664
rect 3728 1600 3736 1664
rect 2267 1188 2333 1189
rect 2267 1124 2268 1188
rect 2332 1124 2333 1188
rect 2267 1123 2333 1124
rect 3416 1040 3736 1600
rect 5888 2208 6208 3232
rect 6318 3229 6378 14043
rect 6502 8261 6562 15150
rect 6499 8260 6565 8261
rect 6499 8196 6500 8260
rect 6564 8196 6565 8260
rect 6499 8195 6565 8196
rect 6686 5949 6746 18123
rect 6870 15605 6930 20707
rect 6867 15604 6933 15605
rect 6867 15540 6868 15604
rect 6932 15540 6933 15604
rect 6867 15539 6933 15540
rect 6867 15196 6933 15197
rect 6867 15132 6868 15196
rect 6932 15132 6933 15196
rect 6867 15131 6933 15132
rect 6870 11797 6930 15131
rect 6867 11796 6933 11797
rect 6867 11732 6868 11796
rect 6932 11732 6933 11796
rect 6867 11731 6933 11732
rect 6867 11116 6933 11117
rect 6867 11052 6868 11116
rect 6932 11052 6933 11116
rect 6867 11051 6933 11052
rect 6870 6357 6930 11051
rect 6867 6356 6933 6357
rect 6867 6292 6868 6356
rect 6932 6292 6933 6356
rect 6867 6291 6933 6292
rect 6683 5948 6749 5949
rect 6683 5884 6684 5948
rect 6748 5884 6749 5948
rect 6683 5883 6749 5884
rect 6499 5812 6565 5813
rect 6499 5748 6500 5812
rect 6564 5748 6565 5812
rect 6499 5747 6565 5748
rect 6315 3228 6381 3229
rect 6315 3164 6316 3228
rect 6380 3164 6381 3228
rect 6315 3163 6381 3164
rect 5888 2144 5896 2208
rect 5960 2144 5976 2208
rect 6040 2144 6056 2208
rect 6120 2144 6136 2208
rect 6200 2144 6208 2208
rect 5888 1120 6208 2144
rect 6502 1461 6562 5747
rect 6683 5540 6749 5541
rect 6683 5476 6684 5540
rect 6748 5476 6749 5540
rect 6683 5475 6749 5476
rect 6867 5540 6933 5541
rect 6867 5476 6868 5540
rect 6932 5476 6933 5540
rect 6867 5475 6933 5476
rect 6686 4453 6746 5475
rect 6870 4861 6930 5475
rect 7054 4861 7114 23294
rect 7235 22812 7301 22813
rect 7235 22748 7236 22812
rect 7300 22748 7301 22812
rect 7235 22747 7301 22748
rect 6867 4860 6933 4861
rect 6867 4796 6868 4860
rect 6932 4796 6933 4860
rect 6867 4795 6933 4796
rect 7051 4860 7117 4861
rect 7051 4796 7052 4860
rect 7116 4796 7117 4860
rect 7051 4795 7117 4796
rect 6867 4724 6933 4725
rect 6867 4660 6868 4724
rect 6932 4660 6933 4724
rect 6867 4659 6933 4660
rect 6870 4589 6930 4659
rect 6867 4588 6933 4589
rect 6867 4524 6868 4588
rect 6932 4524 6933 4588
rect 6867 4523 6933 4524
rect 6683 4452 6749 4453
rect 6683 4388 6684 4452
rect 6748 4388 6749 4452
rect 6683 4387 6749 4388
rect 7051 4452 7117 4453
rect 7051 4388 7052 4452
rect 7116 4388 7117 4452
rect 7051 4387 7117 4388
rect 6683 3364 6749 3365
rect 6683 3300 6684 3364
rect 6748 3300 6749 3364
rect 6683 3299 6749 3300
rect 6499 1460 6565 1461
rect 6499 1396 6500 1460
rect 6564 1396 6565 1460
rect 6499 1395 6565 1396
rect 5888 1056 5896 1120
rect 5960 1056 5976 1120
rect 6040 1056 6056 1120
rect 6120 1056 6136 1120
rect 6200 1056 6208 1120
rect 5888 1040 6208 1056
rect 6686 101 6746 3299
rect 7054 2790 7114 4387
rect 6870 2730 7114 2790
rect 6870 1733 6930 2730
rect 7238 2005 7298 22747
rect 7419 22268 7485 22269
rect 7419 22204 7420 22268
rect 7484 22204 7485 22268
rect 7419 22203 7485 22204
rect 7422 18869 7482 22203
rect 7419 18868 7485 18869
rect 7419 18804 7420 18868
rect 7484 18804 7485 18868
rect 7419 18803 7485 18804
rect 7606 16149 7666 34171
rect 7790 29477 7850 35123
rect 7787 29476 7853 29477
rect 7787 29412 7788 29476
rect 7852 29412 7853 29476
rect 7787 29411 7853 29412
rect 7787 20908 7853 20909
rect 7787 20844 7788 20908
rect 7852 20844 7853 20908
rect 7787 20843 7853 20844
rect 7603 16148 7669 16149
rect 7603 16084 7604 16148
rect 7668 16084 7669 16148
rect 7603 16083 7669 16084
rect 7419 14108 7485 14109
rect 7419 14044 7420 14108
rect 7484 14044 7485 14108
rect 7419 14043 7485 14044
rect 7422 13701 7482 14043
rect 7419 13700 7485 13701
rect 7419 13636 7420 13700
rect 7484 13636 7485 13700
rect 7419 13635 7485 13636
rect 7603 12068 7669 12069
rect 7603 12004 7604 12068
rect 7668 12004 7669 12068
rect 7603 12003 7669 12004
rect 7419 11660 7485 11661
rect 7419 11596 7420 11660
rect 7484 11596 7485 11660
rect 7419 11595 7485 11596
rect 7422 5538 7482 11595
rect 7606 6221 7666 12003
rect 7790 9485 7850 20843
rect 7974 20773 8034 40019
rect 8361 39744 8681 40768
rect 8361 39680 8369 39744
rect 8433 39680 8449 39744
rect 8513 39680 8529 39744
rect 8593 39680 8609 39744
rect 8673 39680 8681 39744
rect 8361 38656 8681 39680
rect 8361 38592 8369 38656
rect 8433 38592 8449 38656
rect 8513 38592 8529 38656
rect 8593 38592 8609 38656
rect 8673 38592 8681 38656
rect 8361 37568 8681 38592
rect 8361 37504 8369 37568
rect 8433 37504 8449 37568
rect 8513 37504 8529 37568
rect 8593 37504 8609 37568
rect 8673 37504 8681 37568
rect 8361 36480 8681 37504
rect 8361 36416 8369 36480
rect 8433 36416 8449 36480
rect 8513 36416 8529 36480
rect 8593 36416 8609 36480
rect 8673 36416 8681 36480
rect 8155 36276 8221 36277
rect 8155 36212 8156 36276
rect 8220 36212 8221 36276
rect 8155 36211 8221 36212
rect 8158 30701 8218 36211
rect 8361 35392 8681 36416
rect 9075 35868 9141 35869
rect 9075 35804 9076 35868
rect 9140 35804 9141 35868
rect 9075 35803 9141 35804
rect 8891 35732 8957 35733
rect 8891 35668 8892 35732
rect 8956 35668 8957 35732
rect 8891 35667 8957 35668
rect 8361 35328 8369 35392
rect 8433 35328 8449 35392
rect 8513 35328 8529 35392
rect 8593 35328 8609 35392
rect 8673 35328 8681 35392
rect 8361 34304 8681 35328
rect 8361 34240 8369 34304
rect 8433 34240 8449 34304
rect 8513 34240 8529 34304
rect 8593 34240 8609 34304
rect 8673 34240 8681 34304
rect 8361 33216 8681 34240
rect 8361 33152 8369 33216
rect 8433 33152 8449 33216
rect 8513 33152 8529 33216
rect 8593 33152 8609 33216
rect 8673 33152 8681 33216
rect 8361 32128 8681 33152
rect 8894 32877 8954 35667
rect 8891 32876 8957 32877
rect 8891 32812 8892 32876
rect 8956 32812 8957 32876
rect 8891 32811 8957 32812
rect 8361 32064 8369 32128
rect 8433 32064 8449 32128
rect 8513 32064 8529 32128
rect 8593 32064 8609 32128
rect 8673 32064 8681 32128
rect 8361 31040 8681 32064
rect 8361 30976 8369 31040
rect 8433 30976 8449 31040
rect 8513 30976 8529 31040
rect 8593 30976 8609 31040
rect 8673 30976 8681 31040
rect 8155 30700 8221 30701
rect 8155 30636 8156 30700
rect 8220 30636 8221 30700
rect 8155 30635 8221 30636
rect 8361 29952 8681 30976
rect 8361 29888 8369 29952
rect 8433 29888 8449 29952
rect 8513 29888 8529 29952
rect 8593 29888 8609 29952
rect 8673 29888 8681 29952
rect 8361 28864 8681 29888
rect 8361 28800 8369 28864
rect 8433 28800 8449 28864
rect 8513 28800 8529 28864
rect 8593 28800 8609 28864
rect 8673 28800 8681 28864
rect 8361 27776 8681 28800
rect 8361 27712 8369 27776
rect 8433 27712 8449 27776
rect 8513 27712 8529 27776
rect 8593 27712 8609 27776
rect 8673 27712 8681 27776
rect 8155 27028 8221 27029
rect 8155 26964 8156 27028
rect 8220 26964 8221 27028
rect 8155 26963 8221 26964
rect 7971 20772 8037 20773
rect 7971 20708 7972 20772
rect 8036 20708 8037 20772
rect 7971 20707 8037 20708
rect 8158 20365 8218 26963
rect 8361 26688 8681 27712
rect 8361 26624 8369 26688
rect 8433 26624 8449 26688
rect 8513 26624 8529 26688
rect 8593 26624 8609 26688
rect 8673 26624 8681 26688
rect 8361 25600 8681 26624
rect 8361 25536 8369 25600
rect 8433 25536 8449 25600
rect 8513 25536 8529 25600
rect 8593 25536 8609 25600
rect 8673 25536 8681 25600
rect 8361 24512 8681 25536
rect 8891 24988 8957 24989
rect 8891 24924 8892 24988
rect 8956 24924 8957 24988
rect 8891 24923 8957 24924
rect 8361 24448 8369 24512
rect 8433 24448 8449 24512
rect 8513 24448 8529 24512
rect 8593 24448 8609 24512
rect 8673 24448 8681 24512
rect 8361 23424 8681 24448
rect 8361 23360 8369 23424
rect 8433 23360 8449 23424
rect 8513 23360 8529 23424
rect 8593 23360 8609 23424
rect 8673 23360 8681 23424
rect 8361 22336 8681 23360
rect 8361 22272 8369 22336
rect 8433 22272 8449 22336
rect 8513 22272 8529 22336
rect 8593 22272 8609 22336
rect 8673 22272 8681 22336
rect 8361 21248 8681 22272
rect 8361 21184 8369 21248
rect 8433 21184 8449 21248
rect 8513 21184 8529 21248
rect 8593 21184 8609 21248
rect 8673 21184 8681 21248
rect 8155 20364 8221 20365
rect 8155 20300 8156 20364
rect 8220 20300 8221 20364
rect 8155 20299 8221 20300
rect 8361 20160 8681 21184
rect 8361 20096 8369 20160
rect 8433 20096 8449 20160
rect 8513 20096 8529 20160
rect 8593 20096 8609 20160
rect 8673 20096 8681 20160
rect 8155 19684 8221 19685
rect 8155 19620 8156 19684
rect 8220 19620 8221 19684
rect 8155 19619 8221 19620
rect 7971 18868 8037 18869
rect 7971 18804 7972 18868
rect 8036 18804 8037 18868
rect 7971 18803 8037 18804
rect 7974 10437 8034 18803
rect 7971 10436 8037 10437
rect 7971 10372 7972 10436
rect 8036 10372 8037 10436
rect 7971 10371 8037 10372
rect 7971 10028 8037 10029
rect 7971 9964 7972 10028
rect 8036 9964 8037 10028
rect 7971 9963 8037 9964
rect 7787 9484 7853 9485
rect 7787 9420 7788 9484
rect 7852 9420 7853 9484
rect 7787 9419 7853 9420
rect 7787 8804 7853 8805
rect 7787 8740 7788 8804
rect 7852 8740 7853 8804
rect 7787 8739 7853 8740
rect 7603 6220 7669 6221
rect 7603 6156 7604 6220
rect 7668 6156 7669 6220
rect 7603 6155 7669 6156
rect 7790 5813 7850 8739
rect 7787 5812 7853 5813
rect 7787 5748 7788 5812
rect 7852 5748 7853 5812
rect 7787 5747 7853 5748
rect 7422 5478 7666 5538
rect 7419 5404 7485 5405
rect 7419 5340 7420 5404
rect 7484 5340 7485 5404
rect 7419 5339 7485 5340
rect 7422 2277 7482 5339
rect 7606 3637 7666 5478
rect 7974 5269 8034 9963
rect 8158 9757 8218 19619
rect 8361 19072 8681 20096
rect 8361 19008 8369 19072
rect 8433 19008 8449 19072
rect 8513 19008 8529 19072
rect 8593 19008 8609 19072
rect 8673 19008 8681 19072
rect 8361 17984 8681 19008
rect 8361 17920 8369 17984
rect 8433 17920 8449 17984
rect 8513 17920 8529 17984
rect 8593 17920 8609 17984
rect 8673 17920 8681 17984
rect 8361 16896 8681 17920
rect 8361 16832 8369 16896
rect 8433 16832 8449 16896
rect 8513 16832 8529 16896
rect 8593 16832 8609 16896
rect 8673 16832 8681 16896
rect 8361 15808 8681 16832
rect 8361 15744 8369 15808
rect 8433 15744 8449 15808
rect 8513 15744 8529 15808
rect 8593 15744 8609 15808
rect 8673 15744 8681 15808
rect 8361 14720 8681 15744
rect 8361 14656 8369 14720
rect 8433 14656 8449 14720
rect 8513 14656 8529 14720
rect 8593 14656 8609 14720
rect 8673 14656 8681 14720
rect 8361 13632 8681 14656
rect 8361 13568 8369 13632
rect 8433 13568 8449 13632
rect 8513 13568 8529 13632
rect 8593 13568 8609 13632
rect 8673 13568 8681 13632
rect 8361 12544 8681 13568
rect 8361 12480 8369 12544
rect 8433 12480 8449 12544
rect 8513 12480 8529 12544
rect 8593 12480 8609 12544
rect 8673 12480 8681 12544
rect 8361 11456 8681 12480
rect 8361 11392 8369 11456
rect 8433 11392 8449 11456
rect 8513 11392 8529 11456
rect 8593 11392 8609 11456
rect 8673 11392 8681 11456
rect 8361 10368 8681 11392
rect 8753 11388 8819 11389
rect 8753 11324 8754 11388
rect 8818 11324 8819 11388
rect 8753 11323 8819 11324
rect 8361 10304 8369 10368
rect 8433 10304 8449 10368
rect 8513 10304 8529 10368
rect 8593 10304 8609 10368
rect 8673 10304 8681 10368
rect 8155 9756 8221 9757
rect 8155 9692 8156 9756
rect 8220 9692 8221 9756
rect 8155 9691 8221 9692
rect 8361 9280 8681 10304
rect 8756 10298 8816 11323
rect 8894 10437 8954 24923
rect 9078 22813 9138 35803
rect 9262 29069 9322 41515
rect 9446 29205 9506 42059
rect 9995 39676 10061 39677
rect 9995 39612 9996 39676
rect 10060 39612 10061 39676
rect 9995 39611 10061 39612
rect 9811 31652 9877 31653
rect 9811 31588 9812 31652
rect 9876 31588 9877 31652
rect 9811 31587 9877 31588
rect 9443 29204 9509 29205
rect 9443 29140 9444 29204
rect 9508 29140 9509 29204
rect 9443 29139 9509 29140
rect 9259 29068 9325 29069
rect 9259 29004 9260 29068
rect 9324 29004 9325 29068
rect 9259 29003 9325 29004
rect 9443 29068 9509 29069
rect 9443 29004 9444 29068
rect 9508 29004 9509 29068
rect 9443 29003 9509 29004
rect 9259 25532 9325 25533
rect 9259 25468 9260 25532
rect 9324 25468 9325 25532
rect 9259 25467 9325 25468
rect 9262 23629 9322 25467
rect 9259 23628 9325 23629
rect 9259 23564 9260 23628
rect 9324 23564 9325 23628
rect 9259 23563 9325 23564
rect 9259 23084 9325 23085
rect 9259 23020 9260 23084
rect 9324 23020 9325 23084
rect 9259 23019 9325 23020
rect 9075 22812 9141 22813
rect 9075 22748 9076 22812
rect 9140 22748 9141 22812
rect 9075 22747 9141 22748
rect 9262 19413 9322 23019
rect 9259 19412 9325 19413
rect 9259 19348 9260 19412
rect 9324 19348 9325 19412
rect 9259 19347 9325 19348
rect 9259 18868 9325 18869
rect 9259 18804 9260 18868
rect 9324 18804 9325 18868
rect 9259 18803 9325 18804
rect 8891 10436 8957 10437
rect 8891 10372 8892 10436
rect 8956 10372 8957 10436
rect 8891 10371 8957 10372
rect 8891 10300 8957 10301
rect 8891 10298 8892 10300
rect 8756 10238 8892 10298
rect 8891 10236 8892 10238
rect 8956 10236 8957 10300
rect 8891 10235 8957 10236
rect 9075 10300 9141 10301
rect 9075 10236 9076 10300
rect 9140 10236 9141 10300
rect 9075 10235 9141 10236
rect 8361 9216 8369 9280
rect 8433 9216 8449 9280
rect 8513 9216 8529 9280
rect 8593 9216 8609 9280
rect 8673 9216 8681 9280
rect 8155 9212 8221 9213
rect 8155 9148 8156 9212
rect 8220 9148 8221 9212
rect 8155 9147 8221 9148
rect 7971 5268 8037 5269
rect 7971 5204 7972 5268
rect 8036 5204 8037 5268
rect 7971 5203 8037 5204
rect 8158 5130 8218 9147
rect 7790 5070 8218 5130
rect 8361 8192 8681 9216
rect 8891 9212 8957 9213
rect 8891 9148 8892 9212
rect 8956 9148 8957 9212
rect 8891 9147 8957 9148
rect 8361 8128 8369 8192
rect 8433 8128 8449 8192
rect 8513 8128 8529 8192
rect 8593 8128 8609 8192
rect 8673 8128 8681 8192
rect 8361 7104 8681 8128
rect 8361 7040 8369 7104
rect 8433 7040 8449 7104
rect 8513 7040 8529 7104
rect 8593 7040 8609 7104
rect 8673 7040 8681 7104
rect 8361 6016 8681 7040
rect 8361 5952 8369 6016
rect 8433 5952 8449 6016
rect 8513 5952 8529 6016
rect 8593 5952 8609 6016
rect 8673 5952 8681 6016
rect 7603 3636 7669 3637
rect 7603 3572 7604 3636
rect 7668 3572 7669 3636
rect 7603 3571 7669 3572
rect 7603 2956 7669 2957
rect 7603 2892 7604 2956
rect 7668 2892 7669 2956
rect 7603 2891 7669 2892
rect 7419 2276 7485 2277
rect 7419 2212 7420 2276
rect 7484 2212 7485 2276
rect 7419 2211 7485 2212
rect 7235 2004 7301 2005
rect 7235 1940 7236 2004
rect 7300 1940 7301 2004
rect 7235 1939 7301 1940
rect 6867 1732 6933 1733
rect 6867 1668 6868 1732
rect 6932 1668 6933 1732
rect 6867 1667 6933 1668
rect 7606 1189 7666 2891
rect 7790 2413 7850 5070
rect 8361 4928 8681 5952
rect 8894 5813 8954 9147
rect 8891 5812 8957 5813
rect 8891 5748 8892 5812
rect 8956 5748 8957 5812
rect 8891 5747 8957 5748
rect 9078 5133 9138 10235
rect 9262 5813 9322 18803
rect 9446 10437 9506 29003
rect 9627 27164 9693 27165
rect 9627 27100 9628 27164
rect 9692 27100 9693 27164
rect 9627 27099 9693 27100
rect 9630 25533 9690 27099
rect 9814 27029 9874 31587
rect 9811 27028 9877 27029
rect 9811 26964 9812 27028
rect 9876 26964 9877 27028
rect 9811 26963 9877 26964
rect 9814 26621 9874 26963
rect 9811 26620 9877 26621
rect 9811 26556 9812 26620
rect 9876 26556 9877 26620
rect 9811 26555 9877 26556
rect 9627 25532 9693 25533
rect 9627 25468 9628 25532
rect 9692 25468 9693 25532
rect 9627 25467 9693 25468
rect 9627 24580 9693 24581
rect 9627 24516 9628 24580
rect 9692 24516 9693 24580
rect 9627 24515 9693 24516
rect 9630 23901 9690 24515
rect 9627 23900 9693 23901
rect 9627 23836 9628 23900
rect 9692 23836 9693 23900
rect 9627 23835 9693 23836
rect 9814 23765 9874 26555
rect 9811 23764 9877 23765
rect 9811 23700 9812 23764
rect 9876 23700 9877 23764
rect 9811 23699 9877 23700
rect 9811 23628 9877 23629
rect 9811 23564 9812 23628
rect 9876 23564 9877 23628
rect 9811 23563 9877 23564
rect 9627 23492 9693 23493
rect 9627 23428 9628 23492
rect 9692 23428 9693 23492
rect 9627 23427 9693 23428
rect 9630 18189 9690 23427
rect 9627 18188 9693 18189
rect 9627 18124 9628 18188
rect 9692 18124 9693 18188
rect 9627 18123 9693 18124
rect 9814 17645 9874 23563
rect 9998 22677 10058 39611
rect 10550 36821 10610 42875
rect 10833 42464 11153 43488
rect 10833 42400 10841 42464
rect 10905 42400 10921 42464
rect 10985 42400 11001 42464
rect 11065 42400 11081 42464
rect 11145 42400 11153 42464
rect 10833 41376 11153 42400
rect 13306 43008 13626 43568
rect 13306 42944 13314 43008
rect 13378 42944 13394 43008
rect 13458 42944 13474 43008
rect 13538 42944 13554 43008
rect 13618 42944 13626 43008
rect 12939 42124 13005 42125
rect 12939 42060 12940 42124
rect 13004 42060 13005 42124
rect 12939 42059 13005 42060
rect 11651 41580 11717 41581
rect 11651 41516 11652 41580
rect 11716 41516 11717 41580
rect 11651 41515 11717 41516
rect 10833 41312 10841 41376
rect 10905 41312 10921 41376
rect 10985 41312 11001 41376
rect 11065 41312 11081 41376
rect 11145 41312 11153 41376
rect 10833 40288 11153 41312
rect 10833 40224 10841 40288
rect 10905 40224 10921 40288
rect 10985 40224 11001 40288
rect 11065 40224 11081 40288
rect 11145 40224 11153 40288
rect 10833 39200 11153 40224
rect 10833 39136 10841 39200
rect 10905 39136 10921 39200
rect 10985 39136 11001 39200
rect 11065 39136 11081 39200
rect 11145 39136 11153 39200
rect 10833 38112 11153 39136
rect 10833 38048 10841 38112
rect 10905 38048 10921 38112
rect 10985 38048 11001 38112
rect 11065 38048 11081 38112
rect 11145 38048 11153 38112
rect 10833 37024 11153 38048
rect 10833 36960 10841 37024
rect 10905 36960 10921 37024
rect 10985 36960 11001 37024
rect 11065 36960 11081 37024
rect 11145 36960 11153 37024
rect 10547 36820 10613 36821
rect 10547 36756 10548 36820
rect 10612 36756 10613 36820
rect 10547 36755 10613 36756
rect 10833 35936 11153 36960
rect 10833 35872 10841 35936
rect 10905 35872 10921 35936
rect 10985 35872 11001 35936
rect 11065 35872 11081 35936
rect 11145 35872 11153 35936
rect 10833 34848 11153 35872
rect 11467 35596 11533 35597
rect 11467 35532 11468 35596
rect 11532 35532 11533 35596
rect 11467 35531 11533 35532
rect 11283 35324 11349 35325
rect 11283 35260 11284 35324
rect 11348 35260 11349 35324
rect 11283 35259 11349 35260
rect 10833 34784 10841 34848
rect 10905 34784 10921 34848
rect 10985 34784 11001 34848
rect 11065 34784 11081 34848
rect 11145 34784 11153 34848
rect 10179 34644 10245 34645
rect 10179 34580 10180 34644
rect 10244 34580 10245 34644
rect 10179 34579 10245 34580
rect 10182 22949 10242 34579
rect 10363 34508 10429 34509
rect 10363 34444 10364 34508
rect 10428 34444 10429 34508
rect 10363 34443 10429 34444
rect 10179 22948 10245 22949
rect 10179 22884 10180 22948
rect 10244 22884 10245 22948
rect 10179 22883 10245 22884
rect 9995 22676 10061 22677
rect 9995 22612 9996 22676
rect 10060 22612 10061 22676
rect 9995 22611 10061 22612
rect 10366 22110 10426 34443
rect 10833 33760 11153 34784
rect 10833 33696 10841 33760
rect 10905 33696 10921 33760
rect 10985 33696 11001 33760
rect 11065 33696 11081 33760
rect 11145 33696 11153 33760
rect 10833 32672 11153 33696
rect 10833 32608 10841 32672
rect 10905 32608 10921 32672
rect 10985 32608 11001 32672
rect 11065 32608 11081 32672
rect 11145 32608 11153 32672
rect 10833 31584 11153 32608
rect 10833 31520 10841 31584
rect 10905 31520 10921 31584
rect 10985 31520 11001 31584
rect 11065 31520 11081 31584
rect 11145 31520 11153 31584
rect 10833 30496 11153 31520
rect 11286 31245 11346 35259
rect 11283 31244 11349 31245
rect 11283 31180 11284 31244
rect 11348 31180 11349 31244
rect 11283 31179 11349 31180
rect 10833 30432 10841 30496
rect 10905 30432 10921 30496
rect 10985 30432 11001 30496
rect 11065 30432 11081 30496
rect 11145 30432 11153 30496
rect 10833 29408 11153 30432
rect 10833 29344 10841 29408
rect 10905 29344 10921 29408
rect 10985 29344 11001 29408
rect 11065 29344 11081 29408
rect 11145 29344 11153 29408
rect 10547 29068 10613 29069
rect 10547 29004 10548 29068
rect 10612 29004 10613 29068
rect 10547 29003 10613 29004
rect 10550 22813 10610 29003
rect 10833 28320 11153 29344
rect 10833 28256 10841 28320
rect 10905 28256 10921 28320
rect 10985 28256 11001 28320
rect 11065 28256 11081 28320
rect 11145 28256 11153 28320
rect 10833 27232 11153 28256
rect 10833 27168 10841 27232
rect 10905 27168 10921 27232
rect 10985 27168 11001 27232
rect 11065 27168 11081 27232
rect 11145 27168 11153 27232
rect 10833 26144 11153 27168
rect 10833 26080 10841 26144
rect 10905 26080 10921 26144
rect 10985 26080 11001 26144
rect 11065 26080 11081 26144
rect 11145 26080 11153 26144
rect 10833 25056 11153 26080
rect 10833 24992 10841 25056
rect 10905 24992 10921 25056
rect 10985 24992 11001 25056
rect 11065 24992 11081 25056
rect 11145 24992 11153 25056
rect 10833 23968 11153 24992
rect 11283 24988 11349 24989
rect 11283 24924 11284 24988
rect 11348 24924 11349 24988
rect 11283 24923 11349 24924
rect 10833 23904 10841 23968
rect 10905 23904 10921 23968
rect 10985 23904 11001 23968
rect 11065 23904 11081 23968
rect 11145 23904 11153 23968
rect 10833 22880 11153 23904
rect 10833 22816 10841 22880
rect 10905 22816 10921 22880
rect 10985 22816 11001 22880
rect 11065 22816 11081 22880
rect 11145 22816 11153 22880
rect 10547 22812 10613 22813
rect 10547 22748 10548 22812
rect 10612 22748 10613 22812
rect 10547 22747 10613 22748
rect 10547 22268 10613 22269
rect 10547 22204 10548 22268
rect 10612 22204 10613 22268
rect 10547 22203 10613 22204
rect 10182 22050 10426 22110
rect 9811 17644 9877 17645
rect 9811 17580 9812 17644
rect 9876 17580 9877 17644
rect 9811 17579 9877 17580
rect 10182 17370 10242 22050
rect 10550 20229 10610 22203
rect 10833 21792 11153 22816
rect 10833 21728 10841 21792
rect 10905 21728 10921 21792
rect 10985 21728 11001 21792
rect 11065 21728 11081 21792
rect 11145 21728 11153 21792
rect 10833 20704 11153 21728
rect 10833 20640 10841 20704
rect 10905 20640 10921 20704
rect 10985 20640 11001 20704
rect 11065 20640 11081 20704
rect 11145 20640 11153 20704
rect 10547 20228 10613 20229
rect 10547 20164 10548 20228
rect 10612 20164 10613 20228
rect 10547 20163 10613 20164
rect 10833 19616 11153 20640
rect 10833 19552 10841 19616
rect 10905 19552 10921 19616
rect 10985 19552 11001 19616
rect 11065 19552 11081 19616
rect 11145 19552 11153 19616
rect 10363 19548 10429 19549
rect 10363 19484 10364 19548
rect 10428 19484 10429 19548
rect 10363 19483 10429 19484
rect 9630 17310 10242 17370
rect 9630 16829 9690 17310
rect 10179 17236 10245 17237
rect 10179 17172 10180 17236
rect 10244 17172 10245 17236
rect 10179 17171 10245 17172
rect 9811 17100 9877 17101
rect 9811 17036 9812 17100
rect 9876 17036 9877 17100
rect 9811 17035 9877 17036
rect 9627 16828 9693 16829
rect 9627 16764 9628 16828
rect 9692 16764 9693 16828
rect 9627 16763 9693 16764
rect 9627 14380 9693 14381
rect 9627 14316 9628 14380
rect 9692 14316 9693 14380
rect 9627 14315 9693 14316
rect 9443 10436 9509 10437
rect 9443 10372 9444 10436
rect 9508 10372 9509 10436
rect 9443 10371 9509 10372
rect 9443 10300 9509 10301
rect 9443 10236 9444 10300
rect 9508 10236 9509 10300
rect 9443 10235 9509 10236
rect 9259 5812 9325 5813
rect 9259 5748 9260 5812
rect 9324 5748 9325 5812
rect 9259 5747 9325 5748
rect 9075 5132 9141 5133
rect 9075 5068 9076 5132
rect 9140 5068 9141 5132
rect 9075 5067 9141 5068
rect 8361 4864 8369 4928
rect 8433 4864 8449 4928
rect 8513 4864 8529 4928
rect 8593 4864 8609 4928
rect 8673 4864 8681 4928
rect 7971 4860 8037 4861
rect 7971 4796 7972 4860
rect 8036 4796 8037 4860
rect 7971 4795 8037 4796
rect 7787 2412 7853 2413
rect 7787 2348 7788 2412
rect 7852 2348 7853 2412
rect 7787 2347 7853 2348
rect 7974 1869 8034 4795
rect 8361 3840 8681 4864
rect 8361 3776 8369 3840
rect 8433 3776 8449 3840
rect 8513 3776 8529 3840
rect 8593 3776 8609 3840
rect 8673 3776 8681 3840
rect 8155 3228 8221 3229
rect 8155 3164 8156 3228
rect 8220 3164 8221 3228
rect 8155 3163 8221 3164
rect 7971 1868 8037 1869
rect 7971 1804 7972 1868
rect 8036 1804 8037 1868
rect 7971 1803 8037 1804
rect 7603 1188 7669 1189
rect 7603 1124 7604 1188
rect 7668 1124 7669 1188
rect 7603 1123 7669 1124
rect 8158 101 8218 3163
rect 8361 2752 8681 3776
rect 8361 2688 8369 2752
rect 8433 2688 8449 2752
rect 8513 2688 8529 2752
rect 8593 2688 8609 2752
rect 8673 2688 8681 2752
rect 8361 1664 8681 2688
rect 8361 1600 8369 1664
rect 8433 1600 8449 1664
rect 8513 1600 8529 1664
rect 8593 1600 8609 1664
rect 8673 1600 8681 1664
rect 8361 1040 8681 1600
rect 9262 1461 9322 5747
rect 9446 3093 9506 10235
rect 9630 7986 9690 14315
rect 9814 9077 9874 17035
rect 9995 13564 10061 13565
rect 9995 13500 9996 13564
rect 10060 13500 10061 13564
rect 9995 13499 10061 13500
rect 9811 9076 9877 9077
rect 9811 9012 9812 9076
rect 9876 9012 9877 9076
rect 9811 9011 9877 9012
rect 9630 7926 9874 7986
rect 9627 7852 9693 7853
rect 9627 7788 9628 7852
rect 9692 7788 9693 7852
rect 9627 7787 9693 7788
rect 9630 6357 9690 7787
rect 9627 6356 9693 6357
rect 9627 6292 9628 6356
rect 9692 6292 9693 6356
rect 9627 6291 9693 6292
rect 9443 3092 9509 3093
rect 9443 3028 9444 3092
rect 9508 3028 9509 3092
rect 9443 3027 9509 3028
rect 9630 1733 9690 6291
rect 9814 3770 9874 7926
rect 9998 6629 10058 13499
rect 9995 6628 10061 6629
rect 9995 6564 9996 6628
rect 10060 6564 10061 6628
rect 9995 6563 10061 6564
rect 9995 6492 10061 6493
rect 9995 6428 9996 6492
rect 10060 6428 10061 6492
rect 9995 6427 10061 6428
rect 9998 3909 10058 6427
rect 10182 4586 10242 17171
rect 10366 15333 10426 19483
rect 10547 19276 10613 19277
rect 10547 19212 10548 19276
rect 10612 19212 10613 19276
rect 10547 19211 10613 19212
rect 10363 15332 10429 15333
rect 10363 15268 10364 15332
rect 10428 15268 10429 15332
rect 10363 15267 10429 15268
rect 10363 13156 10429 13157
rect 10363 13092 10364 13156
rect 10428 13092 10429 13156
rect 10363 13091 10429 13092
rect 10366 9349 10426 13091
rect 10363 9348 10429 9349
rect 10363 9284 10364 9348
rect 10428 9284 10429 9348
rect 10363 9283 10429 9284
rect 10363 9076 10429 9077
rect 10363 9012 10364 9076
rect 10428 9012 10429 9076
rect 10363 9011 10429 9012
rect 10366 8805 10426 9011
rect 10550 8805 10610 19211
rect 10833 18528 11153 19552
rect 11286 19413 11346 24923
rect 11283 19412 11349 19413
rect 11283 19348 11284 19412
rect 11348 19348 11349 19412
rect 11283 19347 11349 19348
rect 10833 18464 10841 18528
rect 10905 18464 10921 18528
rect 10985 18464 11001 18528
rect 11065 18464 11081 18528
rect 11145 18464 11153 18528
rect 10833 17440 11153 18464
rect 10833 17376 10841 17440
rect 10905 17376 10921 17440
rect 10985 17376 11001 17440
rect 11065 17376 11081 17440
rect 11145 17376 11153 17440
rect 10833 16352 11153 17376
rect 11283 17372 11349 17373
rect 11283 17308 11284 17372
rect 11348 17308 11349 17372
rect 11283 17307 11349 17308
rect 10833 16288 10841 16352
rect 10905 16288 10921 16352
rect 10985 16288 11001 16352
rect 11065 16288 11081 16352
rect 11145 16288 11153 16352
rect 10833 15264 11153 16288
rect 10833 15200 10841 15264
rect 10905 15200 10921 15264
rect 10985 15200 11001 15264
rect 11065 15200 11081 15264
rect 11145 15200 11153 15264
rect 10833 14176 11153 15200
rect 10833 14112 10841 14176
rect 10905 14112 10921 14176
rect 10985 14112 11001 14176
rect 11065 14112 11081 14176
rect 11145 14112 11153 14176
rect 10833 13088 11153 14112
rect 10833 13024 10841 13088
rect 10905 13024 10921 13088
rect 10985 13024 11001 13088
rect 11065 13024 11081 13088
rect 11145 13024 11153 13088
rect 10833 12000 11153 13024
rect 10833 11936 10841 12000
rect 10905 11936 10921 12000
rect 10985 11936 11001 12000
rect 11065 11936 11081 12000
rect 11145 11936 11153 12000
rect 10833 10912 11153 11936
rect 10833 10848 10841 10912
rect 10905 10848 10921 10912
rect 10985 10848 11001 10912
rect 11065 10848 11081 10912
rect 11145 10848 11153 10912
rect 10685 10436 10751 10437
rect 10685 10372 10686 10436
rect 10750 10372 10751 10436
rect 10685 10371 10751 10372
rect 10363 8804 10429 8805
rect 10363 8740 10364 8804
rect 10428 8740 10429 8804
rect 10363 8739 10429 8740
rect 10547 8804 10613 8805
rect 10547 8740 10548 8804
rect 10612 8740 10613 8804
rect 10547 8739 10613 8740
rect 10366 8198 10610 8258
rect 10366 4725 10426 8198
rect 10550 8125 10610 8198
rect 10547 8124 10613 8125
rect 10547 8060 10548 8124
rect 10612 8060 10613 8124
rect 10547 8059 10613 8060
rect 10547 7988 10613 7989
rect 10547 7924 10548 7988
rect 10612 7924 10613 7988
rect 10547 7923 10613 7924
rect 10550 5269 10610 7923
rect 10547 5268 10613 5269
rect 10547 5204 10548 5268
rect 10612 5204 10613 5268
rect 10547 5203 10613 5204
rect 10688 5130 10748 10371
rect 10550 5070 10748 5130
rect 10833 9824 11153 10848
rect 10833 9760 10841 9824
rect 10905 9760 10921 9824
rect 10985 9760 11001 9824
rect 11065 9760 11081 9824
rect 11145 9760 11153 9824
rect 10833 8736 11153 9760
rect 10833 8672 10841 8736
rect 10905 8672 10921 8736
rect 10985 8672 11001 8736
rect 11065 8672 11081 8736
rect 11145 8672 11153 8736
rect 10833 7648 11153 8672
rect 10833 7584 10841 7648
rect 10905 7584 10921 7648
rect 10985 7584 11001 7648
rect 11065 7584 11081 7648
rect 11145 7584 11153 7648
rect 10833 6560 11153 7584
rect 10833 6496 10841 6560
rect 10905 6496 10921 6560
rect 10985 6496 11001 6560
rect 11065 6496 11081 6560
rect 11145 6496 11153 6560
rect 10833 5472 11153 6496
rect 10833 5408 10841 5472
rect 10905 5408 10921 5472
rect 10985 5408 11001 5472
rect 11065 5408 11081 5472
rect 11145 5408 11153 5472
rect 10550 4997 10610 5070
rect 10547 4996 10613 4997
rect 10547 4932 10548 4996
rect 10612 4932 10613 4996
rect 10547 4931 10613 4932
rect 10363 4724 10429 4725
rect 10363 4660 10364 4724
rect 10428 4660 10429 4724
rect 10363 4659 10429 4660
rect 10182 4526 10426 4586
rect 9995 3908 10061 3909
rect 9995 3844 9996 3908
rect 10060 3844 10061 3908
rect 9995 3843 10061 3844
rect 9814 3710 10058 3770
rect 9811 3364 9877 3365
rect 9811 3300 9812 3364
rect 9876 3300 9877 3364
rect 9811 3299 9877 3300
rect 9627 1732 9693 1733
rect 9627 1668 9628 1732
rect 9692 1668 9693 1732
rect 9627 1667 9693 1668
rect 9259 1460 9325 1461
rect 9259 1396 9260 1460
rect 9324 1396 9325 1460
rect 9259 1395 9325 1396
rect 9814 917 9874 3299
rect 9998 3093 10058 3710
rect 10179 3228 10245 3229
rect 10179 3164 10180 3228
rect 10244 3164 10245 3228
rect 10179 3163 10245 3164
rect 9995 3092 10061 3093
rect 9995 3028 9996 3092
rect 10060 3028 10061 3092
rect 9995 3027 10061 3028
rect 9995 2820 10061 2821
rect 9995 2756 9996 2820
rect 10060 2756 10061 2820
rect 9995 2755 10061 2756
rect 9811 916 9877 917
rect 9811 852 9812 916
rect 9876 852 9877 916
rect 9811 851 9877 852
rect 9998 781 10058 2755
rect 10182 917 10242 3163
rect 10366 2277 10426 4526
rect 10833 4384 11153 5408
rect 11286 5133 11346 17307
rect 11470 13429 11530 35531
rect 11654 34781 11714 41515
rect 12203 40628 12269 40629
rect 12203 40564 12204 40628
rect 12268 40564 12269 40628
rect 12203 40563 12269 40564
rect 12206 37093 12266 40563
rect 12755 40084 12821 40085
rect 12755 40020 12756 40084
rect 12820 40020 12821 40084
rect 12755 40019 12821 40020
rect 12571 38180 12637 38181
rect 12571 38116 12572 38180
rect 12636 38116 12637 38180
rect 12571 38115 12637 38116
rect 12203 37092 12269 37093
rect 12203 37028 12204 37092
rect 12268 37028 12269 37092
rect 12203 37027 12269 37028
rect 11651 34780 11717 34781
rect 11651 34716 11652 34780
rect 11716 34716 11717 34780
rect 11651 34715 11717 34716
rect 11651 34644 11717 34645
rect 11651 34580 11652 34644
rect 11716 34580 11717 34644
rect 11651 34579 11717 34580
rect 12019 34644 12085 34645
rect 12019 34580 12020 34644
rect 12084 34580 12085 34644
rect 12019 34579 12085 34580
rect 11654 31770 11714 34579
rect 11654 31710 11898 31770
rect 11651 26212 11717 26213
rect 11651 26148 11652 26212
rect 11716 26148 11717 26212
rect 11651 26147 11717 26148
rect 11654 19549 11714 26147
rect 11838 21997 11898 31710
rect 12022 23085 12082 34579
rect 12203 34508 12269 34509
rect 12203 34444 12204 34508
rect 12268 34444 12269 34508
rect 12203 34443 12269 34444
rect 12019 23084 12085 23085
rect 12019 23020 12020 23084
rect 12084 23020 12085 23084
rect 12019 23019 12085 23020
rect 11835 21996 11901 21997
rect 11835 21932 11836 21996
rect 11900 21932 11901 21996
rect 11835 21931 11901 21932
rect 12022 21858 12082 23019
rect 12206 22677 12266 34443
rect 12387 27028 12453 27029
rect 12387 26964 12388 27028
rect 12452 26964 12453 27028
rect 12387 26963 12453 26964
rect 12203 22676 12269 22677
rect 12203 22612 12204 22676
rect 12268 22612 12269 22676
rect 12203 22611 12269 22612
rect 11838 21798 12082 21858
rect 11651 19548 11717 19549
rect 11651 19484 11652 19548
rect 11716 19484 11717 19548
rect 11651 19483 11717 19484
rect 11838 18733 11898 21798
rect 12390 21045 12450 26963
rect 12574 24037 12634 38115
rect 12758 28933 12818 40019
rect 12942 28933 13002 42059
rect 13306 41920 13626 42944
rect 13306 41856 13314 41920
rect 13378 41856 13394 41920
rect 13458 41856 13474 41920
rect 13538 41856 13554 41920
rect 13618 41856 13626 41920
rect 13123 41716 13189 41717
rect 13123 41652 13124 41716
rect 13188 41652 13189 41716
rect 13123 41651 13189 41652
rect 13126 37365 13186 41651
rect 13306 40832 13626 41856
rect 14598 41173 14658 44507
rect 16619 43756 16685 43757
rect 16619 43692 16620 43756
rect 16684 43692 16685 43756
rect 16619 43691 16685 43692
rect 15778 43552 16098 43568
rect 15778 43488 15786 43552
rect 15850 43488 15866 43552
rect 15930 43488 15946 43552
rect 16010 43488 16026 43552
rect 16090 43488 16098 43552
rect 15515 42668 15581 42669
rect 15515 42604 15516 42668
rect 15580 42604 15581 42668
rect 15515 42603 15581 42604
rect 15331 41852 15397 41853
rect 15331 41788 15332 41852
rect 15396 41788 15397 41852
rect 15331 41787 15397 41788
rect 14595 41172 14661 41173
rect 14595 41108 14596 41172
rect 14660 41108 14661 41172
rect 14595 41107 14661 41108
rect 14963 41172 15029 41173
rect 14963 41108 14964 41172
rect 15028 41108 15029 41172
rect 14963 41107 15029 41108
rect 13306 40768 13314 40832
rect 13378 40768 13394 40832
rect 13458 40768 13474 40832
rect 13538 40768 13554 40832
rect 13618 40768 13626 40832
rect 13306 39744 13626 40768
rect 13306 39680 13314 39744
rect 13378 39680 13394 39744
rect 13458 39680 13474 39744
rect 13538 39680 13554 39744
rect 13618 39680 13626 39744
rect 13306 38656 13626 39680
rect 13859 39132 13925 39133
rect 13859 39068 13860 39132
rect 13924 39068 13925 39132
rect 13859 39067 13925 39068
rect 13306 38592 13314 38656
rect 13378 38592 13394 38656
rect 13458 38592 13474 38656
rect 13538 38592 13554 38656
rect 13618 38592 13626 38656
rect 13306 37568 13626 38592
rect 13306 37504 13314 37568
rect 13378 37504 13394 37568
rect 13458 37504 13474 37568
rect 13538 37504 13554 37568
rect 13618 37504 13626 37568
rect 13123 37364 13189 37365
rect 13123 37300 13124 37364
rect 13188 37300 13189 37364
rect 13123 37299 13189 37300
rect 13306 36480 13626 37504
rect 13306 36416 13314 36480
rect 13378 36416 13394 36480
rect 13458 36416 13474 36480
rect 13538 36416 13554 36480
rect 13618 36416 13626 36480
rect 13306 35392 13626 36416
rect 13306 35328 13314 35392
rect 13378 35328 13394 35392
rect 13458 35328 13474 35392
rect 13538 35328 13554 35392
rect 13618 35328 13626 35392
rect 13306 34304 13626 35328
rect 13306 34240 13314 34304
rect 13378 34240 13394 34304
rect 13458 34240 13474 34304
rect 13538 34240 13554 34304
rect 13618 34240 13626 34304
rect 13306 33216 13626 34240
rect 13306 33152 13314 33216
rect 13378 33152 13394 33216
rect 13458 33152 13474 33216
rect 13538 33152 13554 33216
rect 13618 33152 13626 33216
rect 13123 32604 13189 32605
rect 13123 32540 13124 32604
rect 13188 32540 13189 32604
rect 13123 32539 13189 32540
rect 13126 29341 13186 32539
rect 13306 32128 13626 33152
rect 13306 32064 13314 32128
rect 13378 32064 13394 32128
rect 13458 32064 13474 32128
rect 13538 32064 13554 32128
rect 13618 32064 13626 32128
rect 13306 31040 13626 32064
rect 13306 30976 13314 31040
rect 13378 30976 13394 31040
rect 13458 30976 13474 31040
rect 13538 30976 13554 31040
rect 13618 30976 13626 31040
rect 13306 29952 13626 30976
rect 13306 29888 13314 29952
rect 13378 29888 13394 29952
rect 13458 29888 13474 29952
rect 13538 29888 13554 29952
rect 13618 29888 13626 29952
rect 13123 29340 13189 29341
rect 13123 29276 13124 29340
rect 13188 29276 13189 29340
rect 13123 29275 13189 29276
rect 12755 28932 12821 28933
rect 12755 28868 12756 28932
rect 12820 28868 12821 28932
rect 12755 28867 12821 28868
rect 12939 28932 13005 28933
rect 12939 28868 12940 28932
rect 13004 28868 13005 28932
rect 12939 28867 13005 28868
rect 12755 28524 12821 28525
rect 12755 28460 12756 28524
rect 12820 28460 12821 28524
rect 12755 28459 12821 28460
rect 12571 24036 12637 24037
rect 12571 23972 12572 24036
rect 12636 23972 12637 24036
rect 12571 23971 12637 23972
rect 12758 23901 12818 28459
rect 13126 26621 13186 29275
rect 13306 28864 13626 29888
rect 13306 28800 13314 28864
rect 13378 28800 13394 28864
rect 13458 28800 13474 28864
rect 13538 28800 13554 28864
rect 13618 28800 13626 28864
rect 13306 27776 13626 28800
rect 13306 27712 13314 27776
rect 13378 27712 13394 27776
rect 13458 27712 13474 27776
rect 13538 27712 13554 27776
rect 13618 27712 13626 27776
rect 13306 26688 13626 27712
rect 13306 26624 13314 26688
rect 13378 26624 13394 26688
rect 13458 26624 13474 26688
rect 13538 26624 13554 26688
rect 13618 26624 13626 26688
rect 13123 26620 13189 26621
rect 13123 26556 13124 26620
rect 13188 26556 13189 26620
rect 13123 26555 13189 26556
rect 12939 25124 13005 25125
rect 12939 25060 12940 25124
rect 13004 25060 13005 25124
rect 12939 25059 13005 25060
rect 12755 23900 12821 23901
rect 12755 23836 12756 23900
rect 12820 23836 12821 23900
rect 12755 23835 12821 23836
rect 12571 23764 12637 23765
rect 12571 23700 12572 23764
rect 12636 23700 12637 23764
rect 12571 23699 12637 23700
rect 12387 21044 12453 21045
rect 12387 20980 12388 21044
rect 12452 20980 12453 21044
rect 12387 20979 12453 20980
rect 12574 20906 12634 23699
rect 12206 20846 12634 20906
rect 12019 19956 12085 19957
rect 12019 19892 12020 19956
rect 12084 19892 12085 19956
rect 12019 19891 12085 19892
rect 11835 18732 11901 18733
rect 11835 18668 11836 18732
rect 11900 18668 11901 18732
rect 11835 18667 11901 18668
rect 11835 17100 11901 17101
rect 11835 17036 11836 17100
rect 11900 17036 11901 17100
rect 11835 17035 11901 17036
rect 11651 16284 11717 16285
rect 11651 16220 11652 16284
rect 11716 16220 11717 16284
rect 11651 16219 11717 16220
rect 11467 13428 11533 13429
rect 11467 13364 11468 13428
rect 11532 13364 11533 13428
rect 11467 13363 11533 13364
rect 11467 12068 11533 12069
rect 11467 12004 11468 12068
rect 11532 12004 11533 12068
rect 11467 12003 11533 12004
rect 11470 10709 11530 12003
rect 11654 10845 11714 16219
rect 11838 15877 11898 17035
rect 11835 15876 11901 15877
rect 11835 15812 11836 15876
rect 11900 15812 11901 15876
rect 11835 15811 11901 15812
rect 12022 11794 12082 19891
rect 12206 15061 12266 20846
rect 12755 20500 12821 20501
rect 12755 20436 12756 20500
rect 12820 20436 12821 20500
rect 12755 20435 12821 20436
rect 12387 19004 12453 19005
rect 12387 18940 12388 19004
rect 12452 18940 12453 19004
rect 12387 18939 12453 18940
rect 12390 18730 12450 18939
rect 12390 18670 12634 18730
rect 12574 15210 12634 18670
rect 12390 15150 12634 15210
rect 12203 15060 12269 15061
rect 12203 14996 12204 15060
rect 12268 14996 12269 15060
rect 12203 14995 12269 14996
rect 12022 11734 12266 11794
rect 12019 11252 12085 11253
rect 12019 11188 12020 11252
rect 12084 11188 12085 11252
rect 12019 11187 12085 11188
rect 11651 10844 11717 10845
rect 11651 10780 11652 10844
rect 11716 10780 11717 10844
rect 11651 10779 11717 10780
rect 11467 10708 11533 10709
rect 11467 10644 11468 10708
rect 11532 10644 11533 10708
rect 11467 10643 11533 10644
rect 11835 10572 11901 10573
rect 11835 10508 11836 10572
rect 11900 10508 11901 10572
rect 11835 10507 11901 10508
rect 11467 10436 11533 10437
rect 11467 10372 11468 10436
rect 11532 10372 11533 10436
rect 11467 10371 11533 10372
rect 11283 5132 11349 5133
rect 11283 5068 11284 5132
rect 11348 5068 11349 5132
rect 11283 5067 11349 5068
rect 11283 4588 11349 4589
rect 11283 4524 11284 4588
rect 11348 4524 11349 4588
rect 11283 4523 11349 4524
rect 10833 4320 10841 4384
rect 10905 4320 10921 4384
rect 10985 4320 11001 4384
rect 11065 4320 11081 4384
rect 11145 4320 11153 4384
rect 10547 3364 10613 3365
rect 10547 3300 10548 3364
rect 10612 3300 10613 3364
rect 10547 3299 10613 3300
rect 10363 2276 10429 2277
rect 10363 2212 10364 2276
rect 10428 2212 10429 2276
rect 10363 2211 10429 2212
rect 10179 916 10245 917
rect 10179 852 10180 916
rect 10244 852 10245 916
rect 10179 851 10245 852
rect 10550 781 10610 3299
rect 10833 3296 11153 4320
rect 11286 3365 11346 4523
rect 11283 3364 11349 3365
rect 11283 3300 11284 3364
rect 11348 3300 11349 3364
rect 11283 3299 11349 3300
rect 10833 3232 10841 3296
rect 10905 3232 10921 3296
rect 10985 3232 11001 3296
rect 11065 3232 11081 3296
rect 11145 3232 11153 3296
rect 10833 2208 11153 3232
rect 11283 3228 11349 3229
rect 11283 3164 11284 3228
rect 11348 3164 11349 3228
rect 11283 3163 11349 3164
rect 10833 2144 10841 2208
rect 10905 2144 10921 2208
rect 10985 2144 11001 2208
rect 11065 2144 11081 2208
rect 11145 2144 11153 2208
rect 10833 1120 11153 2144
rect 10833 1056 10841 1120
rect 10905 1056 10921 1120
rect 10985 1056 11001 1120
rect 11065 1056 11081 1120
rect 11145 1056 11153 1120
rect 10833 1040 11153 1056
rect 11286 917 11346 3163
rect 11470 3093 11530 10371
rect 11651 9756 11717 9757
rect 11651 9692 11652 9756
rect 11716 9692 11717 9756
rect 11651 9691 11717 9692
rect 11654 5541 11714 9691
rect 11651 5540 11717 5541
rect 11651 5476 11652 5540
rect 11716 5476 11717 5540
rect 11651 5475 11717 5476
rect 11651 5132 11717 5133
rect 11651 5068 11652 5132
rect 11716 5068 11717 5132
rect 11651 5067 11717 5068
rect 11654 4861 11714 5067
rect 11838 4861 11898 10507
rect 12022 5813 12082 11187
rect 12206 9213 12266 11734
rect 12203 9212 12269 9213
rect 12203 9148 12204 9212
rect 12268 9148 12269 9212
rect 12203 9147 12269 9148
rect 12390 9074 12450 15150
rect 12571 13428 12637 13429
rect 12571 13364 12572 13428
rect 12636 13364 12637 13428
rect 12571 13363 12637 13364
rect 12206 9014 12450 9074
rect 12206 5949 12266 9014
rect 12387 8804 12453 8805
rect 12387 8740 12388 8804
rect 12452 8740 12453 8804
rect 12387 8739 12453 8740
rect 12203 5948 12269 5949
rect 12203 5884 12204 5948
rect 12268 5884 12269 5948
rect 12203 5883 12269 5884
rect 12019 5812 12085 5813
rect 12019 5748 12020 5812
rect 12084 5748 12085 5812
rect 12019 5747 12085 5748
rect 12390 5674 12450 8739
rect 12022 5614 12450 5674
rect 11651 4860 11717 4861
rect 11651 4796 11652 4860
rect 11716 4796 11717 4860
rect 11651 4795 11717 4796
rect 11835 4860 11901 4861
rect 11835 4796 11836 4860
rect 11900 4796 11901 4860
rect 11835 4795 11901 4796
rect 12022 4725 12082 5614
rect 12574 5538 12634 13363
rect 12758 10301 12818 20435
rect 12942 15877 13002 25059
rect 13126 20909 13186 26555
rect 13306 25600 13626 26624
rect 13306 25536 13314 25600
rect 13378 25536 13394 25600
rect 13458 25536 13474 25600
rect 13538 25536 13554 25600
rect 13618 25536 13626 25600
rect 13306 24512 13626 25536
rect 13306 24448 13314 24512
rect 13378 24448 13394 24512
rect 13458 24448 13474 24512
rect 13538 24448 13554 24512
rect 13618 24448 13626 24512
rect 13306 23424 13626 24448
rect 13306 23360 13314 23424
rect 13378 23360 13394 23424
rect 13458 23360 13474 23424
rect 13538 23360 13554 23424
rect 13618 23360 13626 23424
rect 13306 22336 13626 23360
rect 13306 22272 13314 22336
rect 13378 22272 13394 22336
rect 13458 22272 13474 22336
rect 13538 22272 13554 22336
rect 13618 22272 13626 22336
rect 13306 21248 13626 22272
rect 13306 21184 13314 21248
rect 13378 21184 13394 21248
rect 13458 21184 13474 21248
rect 13538 21184 13554 21248
rect 13618 21184 13626 21248
rect 13123 20908 13189 20909
rect 13123 20844 13124 20908
rect 13188 20844 13189 20908
rect 13123 20843 13189 20844
rect 13306 20160 13626 21184
rect 13306 20096 13314 20160
rect 13378 20096 13394 20160
rect 13458 20096 13474 20160
rect 13538 20096 13554 20160
rect 13618 20096 13626 20160
rect 13306 19072 13626 20096
rect 13862 19957 13922 39067
rect 14411 35868 14477 35869
rect 14411 35804 14412 35868
rect 14476 35804 14477 35868
rect 14411 35803 14477 35804
rect 14043 35324 14109 35325
rect 14043 35260 14044 35324
rect 14108 35260 14109 35324
rect 14043 35259 14109 35260
rect 14046 30565 14106 35259
rect 14043 30564 14109 30565
rect 14043 30500 14044 30564
rect 14108 30500 14109 30564
rect 14043 30499 14109 30500
rect 14227 29748 14293 29749
rect 14227 29684 14228 29748
rect 14292 29684 14293 29748
rect 14227 29683 14293 29684
rect 14230 29205 14290 29683
rect 14227 29204 14293 29205
rect 14227 29140 14228 29204
rect 14292 29140 14293 29204
rect 14227 29139 14293 29140
rect 14043 28660 14109 28661
rect 14043 28596 14044 28660
rect 14108 28596 14109 28660
rect 14043 28595 14109 28596
rect 14046 20229 14106 28595
rect 14230 22110 14290 29139
rect 14414 29069 14474 35803
rect 14595 35188 14661 35189
rect 14595 35124 14596 35188
rect 14660 35124 14661 35188
rect 14595 35123 14661 35124
rect 14411 29068 14477 29069
rect 14411 29004 14412 29068
rect 14476 29004 14477 29068
rect 14411 29003 14477 29004
rect 14598 23629 14658 35123
rect 14966 31770 15026 41107
rect 15334 40357 15394 41787
rect 15518 41445 15578 42603
rect 15778 42464 16098 43488
rect 16251 43212 16317 43213
rect 16251 43148 16252 43212
rect 16316 43210 16317 43212
rect 16316 43150 16498 43210
rect 16316 43148 16317 43150
rect 16251 43147 16317 43148
rect 15778 42400 15786 42464
rect 15850 42400 15866 42464
rect 15930 42400 15946 42464
rect 16010 42400 16026 42464
rect 16090 42400 16098 42464
rect 15515 41444 15581 41445
rect 15515 41380 15516 41444
rect 15580 41380 15581 41444
rect 15515 41379 15581 41380
rect 15778 41376 16098 42400
rect 15778 41312 15786 41376
rect 15850 41312 15866 41376
rect 15930 41312 15946 41376
rect 16010 41312 16026 41376
rect 16090 41312 16098 41376
rect 15331 40356 15397 40357
rect 15331 40292 15332 40356
rect 15396 40292 15397 40356
rect 15331 40291 15397 40292
rect 15778 40288 16098 41312
rect 16438 41309 16498 43150
rect 16435 41308 16501 41309
rect 16435 41244 16436 41308
rect 16500 41244 16501 41308
rect 16435 41243 16501 41244
rect 16622 40765 16682 43691
rect 18251 43008 18571 43568
rect 18251 42944 18259 43008
rect 18323 42944 18339 43008
rect 18403 42944 18419 43008
rect 18483 42944 18499 43008
rect 18563 42944 18571 43008
rect 18091 42124 18157 42125
rect 18091 42060 18092 42124
rect 18156 42060 18157 42124
rect 18091 42059 18157 42060
rect 18094 40901 18154 42059
rect 18251 41920 18571 42944
rect 18251 41856 18259 41920
rect 18323 41856 18339 41920
rect 18403 41856 18419 41920
rect 18483 41856 18499 41920
rect 18563 41856 18571 41920
rect 18091 40900 18157 40901
rect 18091 40836 18092 40900
rect 18156 40836 18157 40900
rect 18091 40835 18157 40836
rect 18251 40832 18571 41856
rect 18251 40768 18259 40832
rect 18323 40768 18339 40832
rect 18403 40768 18419 40832
rect 18483 40768 18499 40832
rect 18563 40768 18571 40832
rect 16619 40764 16685 40765
rect 16619 40700 16620 40764
rect 16684 40700 16685 40764
rect 16619 40699 16685 40700
rect 15778 40224 15786 40288
rect 15850 40224 15866 40288
rect 15930 40224 15946 40288
rect 16010 40224 16026 40288
rect 16090 40224 16098 40288
rect 15778 39200 16098 40224
rect 16987 40084 17053 40085
rect 16987 40020 16988 40084
rect 17052 40020 17053 40084
rect 16987 40019 17053 40020
rect 17907 40084 17973 40085
rect 17907 40020 17908 40084
rect 17972 40020 17973 40084
rect 17907 40019 17973 40020
rect 16251 39268 16317 39269
rect 16251 39204 16252 39268
rect 16316 39204 16317 39268
rect 16251 39203 16317 39204
rect 15778 39136 15786 39200
rect 15850 39136 15866 39200
rect 15930 39136 15946 39200
rect 16010 39136 16026 39200
rect 16090 39136 16098 39200
rect 15778 38112 16098 39136
rect 15778 38048 15786 38112
rect 15850 38048 15866 38112
rect 15930 38048 15946 38112
rect 16010 38048 16026 38112
rect 16090 38048 16098 38112
rect 15778 37024 16098 38048
rect 15778 36960 15786 37024
rect 15850 36960 15866 37024
rect 15930 36960 15946 37024
rect 16010 36960 16026 37024
rect 16090 36960 16098 37024
rect 15778 35936 16098 36960
rect 15778 35872 15786 35936
rect 15850 35872 15866 35936
rect 15930 35872 15946 35936
rect 16010 35872 16026 35936
rect 16090 35872 16098 35936
rect 15778 34848 16098 35872
rect 15778 34784 15786 34848
rect 15850 34784 15866 34848
rect 15930 34784 15946 34848
rect 16010 34784 16026 34848
rect 16090 34784 16098 34848
rect 15147 34780 15213 34781
rect 15147 34716 15148 34780
rect 15212 34716 15213 34780
rect 15147 34715 15213 34716
rect 15515 34780 15581 34781
rect 15515 34716 15516 34780
rect 15580 34716 15581 34780
rect 15515 34715 15581 34716
rect 14782 31710 15026 31770
rect 14595 23628 14661 23629
rect 14595 23564 14596 23628
rect 14660 23564 14661 23628
rect 14595 23563 14661 23564
rect 14782 22677 14842 31710
rect 15150 29069 15210 34715
rect 15147 29068 15213 29069
rect 15147 29004 15148 29068
rect 15212 29004 15213 29068
rect 15147 29003 15213 29004
rect 15147 28252 15213 28253
rect 15147 28188 15148 28252
rect 15212 28188 15213 28252
rect 15147 28187 15213 28188
rect 14963 27708 15029 27709
rect 14963 27644 14964 27708
rect 15028 27644 15029 27708
rect 14963 27643 15029 27644
rect 14595 22676 14661 22677
rect 14595 22612 14596 22676
rect 14660 22612 14661 22676
rect 14595 22611 14661 22612
rect 14779 22676 14845 22677
rect 14779 22612 14780 22676
rect 14844 22612 14845 22676
rect 14779 22611 14845 22612
rect 14230 22050 14474 22110
rect 14227 21588 14293 21589
rect 14227 21524 14228 21588
rect 14292 21524 14293 21588
rect 14227 21523 14293 21524
rect 14043 20228 14109 20229
rect 14043 20164 14044 20228
rect 14108 20164 14109 20228
rect 14043 20163 14109 20164
rect 13859 19956 13925 19957
rect 13859 19892 13860 19956
rect 13924 19892 13925 19956
rect 13859 19891 13925 19892
rect 13306 19008 13314 19072
rect 13378 19008 13394 19072
rect 13458 19008 13474 19072
rect 13538 19008 13554 19072
rect 13618 19008 13626 19072
rect 13123 18188 13189 18189
rect 13123 18124 13124 18188
rect 13188 18124 13189 18188
rect 13123 18123 13189 18124
rect 12939 15876 13005 15877
rect 12939 15812 12940 15876
rect 13004 15812 13005 15876
rect 12939 15811 13005 15812
rect 13126 15210 13186 18123
rect 12942 15150 13186 15210
rect 13306 17984 13626 19008
rect 13306 17920 13314 17984
rect 13378 17920 13394 17984
rect 13458 17920 13474 17984
rect 13538 17920 13554 17984
rect 13618 17920 13626 17984
rect 13306 16896 13626 17920
rect 14230 17781 14290 21523
rect 14414 18461 14474 22050
rect 14598 18869 14658 22611
rect 14966 22110 15026 27643
rect 14782 22050 15026 22110
rect 14782 20501 14842 22050
rect 14963 20772 15029 20773
rect 14963 20708 14964 20772
rect 15028 20708 15029 20772
rect 14963 20707 15029 20708
rect 14779 20500 14845 20501
rect 14779 20436 14780 20500
rect 14844 20436 14845 20500
rect 14779 20435 14845 20436
rect 14595 18868 14661 18869
rect 14595 18804 14596 18868
rect 14660 18804 14661 18868
rect 14595 18803 14661 18804
rect 14411 18460 14477 18461
rect 14411 18396 14412 18460
rect 14476 18396 14477 18460
rect 14411 18395 14477 18396
rect 14227 17780 14293 17781
rect 14227 17716 14228 17780
rect 14292 17716 14293 17780
rect 14227 17715 14293 17716
rect 13306 16832 13314 16896
rect 13378 16832 13394 16896
rect 13458 16832 13474 16896
rect 13538 16832 13554 16896
rect 13618 16832 13626 16896
rect 13306 15808 13626 16832
rect 14043 16828 14109 16829
rect 14043 16764 14044 16828
rect 14108 16764 14109 16828
rect 14043 16763 14109 16764
rect 13306 15744 13314 15808
rect 13378 15744 13394 15808
rect 13458 15744 13474 15808
rect 13538 15744 13554 15808
rect 13618 15744 13626 15808
rect 12755 10300 12821 10301
rect 12755 10236 12756 10300
rect 12820 10236 12821 10300
rect 12755 10235 12821 10236
rect 12755 9892 12821 9893
rect 12755 9828 12756 9892
rect 12820 9828 12821 9892
rect 12755 9827 12821 9828
rect 12758 7581 12818 9827
rect 12942 9349 13002 15150
rect 13306 14720 13626 15744
rect 13859 15060 13925 15061
rect 13859 14996 13860 15060
rect 13924 14996 13925 15060
rect 13859 14995 13925 14996
rect 13306 14656 13314 14720
rect 13378 14656 13394 14720
rect 13458 14656 13474 14720
rect 13538 14656 13554 14720
rect 13618 14656 13626 14720
rect 13123 14244 13189 14245
rect 13123 14180 13124 14244
rect 13188 14180 13189 14244
rect 13123 14179 13189 14180
rect 12939 9348 13005 9349
rect 12939 9284 12940 9348
rect 13004 9284 13005 9348
rect 12939 9283 13005 9284
rect 12755 7580 12821 7581
rect 12755 7516 12756 7580
rect 12820 7516 12821 7580
rect 12755 7515 12821 7516
rect 12939 7580 13005 7581
rect 12939 7516 12940 7580
rect 13004 7516 13005 7580
rect 12939 7515 13005 7516
rect 12755 7308 12821 7309
rect 12755 7244 12756 7308
rect 12820 7244 12821 7308
rect 12755 7243 12821 7244
rect 12206 5478 12634 5538
rect 12206 4861 12266 5478
rect 12758 5405 12818 7243
rect 12942 7037 13002 7515
rect 12939 7036 13005 7037
rect 12939 6972 12940 7036
rect 13004 6972 13005 7036
rect 12939 6971 13005 6972
rect 12939 6900 13005 6901
rect 12939 6836 12940 6900
rect 13004 6836 13005 6900
rect 12939 6835 13005 6836
rect 12755 5404 12821 5405
rect 12755 5340 12756 5404
rect 12820 5340 12821 5404
rect 12755 5339 12821 5340
rect 12942 5266 13002 6835
rect 13126 5949 13186 14179
rect 13306 13632 13626 14656
rect 13306 13568 13314 13632
rect 13378 13568 13394 13632
rect 13458 13568 13474 13632
rect 13538 13568 13554 13632
rect 13618 13568 13626 13632
rect 13306 12544 13626 13568
rect 13306 12480 13314 12544
rect 13378 12480 13394 12544
rect 13458 12480 13474 12544
rect 13538 12480 13554 12544
rect 13618 12480 13626 12544
rect 13306 11456 13626 12480
rect 13862 12069 13922 14995
rect 13859 12068 13925 12069
rect 13859 12004 13860 12068
rect 13924 12004 13925 12068
rect 13859 12003 13925 12004
rect 13306 11392 13314 11456
rect 13378 11392 13394 11456
rect 13458 11392 13474 11456
rect 13538 11392 13554 11456
rect 13618 11392 13626 11456
rect 13306 10368 13626 11392
rect 13859 10844 13925 10845
rect 13859 10780 13860 10844
rect 13924 10780 13925 10844
rect 13859 10779 13925 10780
rect 13306 10304 13314 10368
rect 13378 10304 13394 10368
rect 13458 10304 13474 10368
rect 13538 10304 13554 10368
rect 13618 10304 13626 10368
rect 13306 9280 13626 10304
rect 13862 9890 13922 10779
rect 14046 10573 14106 16763
rect 14230 15210 14290 17715
rect 14966 15605 15026 20707
rect 14963 15604 15029 15605
rect 14963 15540 14964 15604
rect 15028 15540 15029 15604
rect 14963 15539 15029 15540
rect 14230 15150 14474 15210
rect 14227 14652 14293 14653
rect 14227 14588 14228 14652
rect 14292 14588 14293 14652
rect 14227 14587 14293 14588
rect 14230 11933 14290 14587
rect 14414 14381 14474 15150
rect 15150 14517 15210 28187
rect 15518 25125 15578 34715
rect 15778 33760 16098 34784
rect 15778 33696 15786 33760
rect 15850 33696 15866 33760
rect 15930 33696 15946 33760
rect 16010 33696 16026 33760
rect 16090 33696 16098 33760
rect 15778 32672 16098 33696
rect 15778 32608 15786 32672
rect 15850 32608 15866 32672
rect 15930 32608 15946 32672
rect 16010 32608 16026 32672
rect 16090 32608 16098 32672
rect 15778 31584 16098 32608
rect 15778 31520 15786 31584
rect 15850 31520 15866 31584
rect 15930 31520 15946 31584
rect 16010 31520 16026 31584
rect 16090 31520 16098 31584
rect 15778 30496 16098 31520
rect 15778 30432 15786 30496
rect 15850 30432 15866 30496
rect 15930 30432 15946 30496
rect 16010 30432 16026 30496
rect 16090 30432 16098 30496
rect 15778 29408 16098 30432
rect 15778 29344 15786 29408
rect 15850 29344 15866 29408
rect 15930 29344 15946 29408
rect 16010 29344 16026 29408
rect 16090 29344 16098 29408
rect 15778 28320 16098 29344
rect 15778 28256 15786 28320
rect 15850 28256 15866 28320
rect 15930 28256 15946 28320
rect 16010 28256 16026 28320
rect 16090 28256 16098 28320
rect 15778 27232 16098 28256
rect 15778 27168 15786 27232
rect 15850 27168 15866 27232
rect 15930 27168 15946 27232
rect 16010 27168 16026 27232
rect 16090 27168 16098 27232
rect 15778 26144 16098 27168
rect 15778 26080 15786 26144
rect 15850 26080 15866 26144
rect 15930 26080 15946 26144
rect 16010 26080 16026 26144
rect 16090 26080 16098 26144
rect 15515 25124 15581 25125
rect 15515 25060 15516 25124
rect 15580 25060 15581 25124
rect 15515 25059 15581 25060
rect 15518 22405 15578 25059
rect 15778 25056 16098 26080
rect 15778 24992 15786 25056
rect 15850 24992 15866 25056
rect 15930 24992 15946 25056
rect 16010 24992 16026 25056
rect 16090 24992 16098 25056
rect 15778 23968 16098 24992
rect 15778 23904 15786 23968
rect 15850 23904 15866 23968
rect 15930 23904 15946 23968
rect 16010 23904 16026 23968
rect 16090 23904 16098 23968
rect 15778 22880 16098 23904
rect 16254 23493 16314 39203
rect 16435 37908 16501 37909
rect 16435 37844 16436 37908
rect 16500 37844 16501 37908
rect 16435 37843 16501 37844
rect 16438 31517 16498 37843
rect 16803 37500 16869 37501
rect 16803 37436 16804 37500
rect 16868 37436 16869 37500
rect 16803 37435 16869 37436
rect 16619 33964 16685 33965
rect 16619 33900 16620 33964
rect 16684 33900 16685 33964
rect 16619 33899 16685 33900
rect 16435 31516 16501 31517
rect 16435 31452 16436 31516
rect 16500 31452 16501 31516
rect 16435 31451 16501 31452
rect 16435 31380 16501 31381
rect 16435 31316 16436 31380
rect 16500 31316 16501 31380
rect 16435 31315 16501 31316
rect 16438 30426 16498 31315
rect 16622 30701 16682 33899
rect 16806 31109 16866 37435
rect 16803 31108 16869 31109
rect 16803 31044 16804 31108
rect 16868 31044 16869 31108
rect 16803 31043 16869 31044
rect 16619 30700 16685 30701
rect 16619 30636 16620 30700
rect 16684 30636 16685 30700
rect 16619 30635 16685 30636
rect 16438 30366 16682 30426
rect 16435 29204 16501 29205
rect 16435 29140 16436 29204
rect 16500 29140 16501 29204
rect 16435 29139 16501 29140
rect 16251 23492 16317 23493
rect 16251 23428 16252 23492
rect 16316 23428 16317 23492
rect 16251 23427 16317 23428
rect 15778 22816 15786 22880
rect 15850 22816 15866 22880
rect 15930 22816 15946 22880
rect 16010 22816 16026 22880
rect 16090 22816 16098 22880
rect 15515 22404 15581 22405
rect 15515 22340 15516 22404
rect 15580 22340 15581 22404
rect 15515 22339 15581 22340
rect 15331 22132 15397 22133
rect 15331 22068 15332 22132
rect 15396 22068 15397 22132
rect 15331 22067 15397 22068
rect 15147 14516 15213 14517
rect 15147 14452 15148 14516
rect 15212 14452 15213 14516
rect 15147 14451 15213 14452
rect 14411 14380 14477 14381
rect 14411 14316 14412 14380
rect 14476 14316 14477 14380
rect 14411 14315 14477 14316
rect 15147 14380 15213 14381
rect 15147 14316 15148 14380
rect 15212 14316 15213 14380
rect 15147 14315 15213 14316
rect 14779 14108 14845 14109
rect 14779 14044 14780 14108
rect 14844 14044 14845 14108
rect 14779 14043 14845 14044
rect 14782 13837 14842 14043
rect 14779 13836 14845 13837
rect 14779 13772 14780 13836
rect 14844 13772 14845 13836
rect 14779 13771 14845 13772
rect 14595 13428 14661 13429
rect 14595 13364 14596 13428
rect 14660 13364 14661 13428
rect 14595 13363 14661 13364
rect 14411 13156 14477 13157
rect 14411 13092 14412 13156
rect 14476 13092 14477 13156
rect 14411 13091 14477 13092
rect 14414 12069 14474 13091
rect 14411 12068 14477 12069
rect 14411 12004 14412 12068
rect 14476 12004 14477 12068
rect 14411 12003 14477 12004
rect 14227 11932 14293 11933
rect 14227 11868 14228 11932
rect 14292 11868 14293 11932
rect 14227 11867 14293 11868
rect 14043 10572 14109 10573
rect 14043 10508 14044 10572
rect 14108 10508 14109 10572
rect 14043 10507 14109 10508
rect 14411 10572 14477 10573
rect 14411 10508 14412 10572
rect 14476 10508 14477 10572
rect 14411 10507 14477 10508
rect 14414 10165 14474 10507
rect 14411 10164 14477 10165
rect 14411 10100 14412 10164
rect 14476 10100 14477 10164
rect 14411 10099 14477 10100
rect 13862 9830 14106 9890
rect 13306 9216 13314 9280
rect 13378 9216 13394 9280
rect 13458 9216 13474 9280
rect 13538 9216 13554 9280
rect 13618 9216 13626 9280
rect 13306 8192 13626 9216
rect 13859 8804 13925 8805
rect 13859 8740 13860 8804
rect 13924 8740 13925 8804
rect 13859 8739 13925 8740
rect 13306 8128 13314 8192
rect 13378 8128 13394 8192
rect 13458 8128 13474 8192
rect 13538 8128 13554 8192
rect 13618 8128 13626 8192
rect 13306 7104 13626 8128
rect 13862 7989 13922 8739
rect 13859 7988 13925 7989
rect 13859 7924 13860 7988
rect 13924 7924 13925 7988
rect 13859 7923 13925 7924
rect 13306 7040 13314 7104
rect 13378 7040 13394 7104
rect 13458 7040 13474 7104
rect 13538 7040 13554 7104
rect 13618 7040 13626 7104
rect 13306 6016 13626 7040
rect 13306 5952 13314 6016
rect 13378 5952 13394 6016
rect 13458 5952 13474 6016
rect 13538 5952 13554 6016
rect 13618 5952 13626 6016
rect 13123 5948 13189 5949
rect 13123 5884 13124 5948
rect 13188 5884 13189 5948
rect 13123 5883 13189 5884
rect 12390 5206 13002 5266
rect 12203 4860 12269 4861
rect 12203 4796 12204 4860
rect 12268 4796 12269 4860
rect 12203 4795 12269 4796
rect 12019 4724 12085 4725
rect 12019 4660 12020 4724
rect 12084 4660 12085 4724
rect 12019 4659 12085 4660
rect 12203 4588 12269 4589
rect 12203 4524 12204 4588
rect 12268 4524 12269 4588
rect 12203 4523 12269 4524
rect 12019 4044 12085 4045
rect 12019 3980 12020 4044
rect 12084 3980 12085 4044
rect 12019 3979 12085 3980
rect 11651 3908 11717 3909
rect 11651 3844 11652 3908
rect 11716 3844 11717 3908
rect 11651 3843 11717 3844
rect 11467 3092 11533 3093
rect 11467 3028 11468 3092
rect 11532 3028 11533 3092
rect 11467 3027 11533 3028
rect 11283 916 11349 917
rect 11283 852 11284 916
rect 11348 852 11349 916
rect 11283 851 11349 852
rect 9995 780 10061 781
rect 9995 716 9996 780
rect 10060 716 10061 780
rect 9995 715 10061 716
rect 10547 780 10613 781
rect 10547 716 10548 780
rect 10612 716 10613 780
rect 10547 715 10613 716
rect 11654 373 11714 3843
rect 12022 3226 12082 3979
rect 12206 3634 12266 4523
rect 12390 4317 12450 5206
rect 13123 5132 13189 5133
rect 13123 5130 13124 5132
rect 12758 5070 13124 5130
rect 12571 4724 12637 4725
rect 12571 4660 12572 4724
rect 12636 4660 12637 4724
rect 12571 4659 12637 4660
rect 12387 4316 12453 4317
rect 12387 4252 12388 4316
rect 12452 4252 12453 4316
rect 12387 4251 12453 4252
rect 12574 3773 12634 4659
rect 12758 4453 12818 5070
rect 13123 5068 13124 5070
rect 13188 5068 13189 5132
rect 13123 5067 13189 5068
rect 13306 4928 13626 5952
rect 13859 5948 13925 5949
rect 13859 5884 13860 5948
rect 13924 5884 13925 5948
rect 13859 5883 13925 5884
rect 13306 4864 13314 4928
rect 13378 4864 13394 4928
rect 13458 4864 13474 4928
rect 13538 4864 13554 4928
rect 13618 4864 13626 4928
rect 12755 4452 12821 4453
rect 12755 4388 12756 4452
rect 12820 4388 12821 4452
rect 13123 4452 13189 4453
rect 13123 4450 13124 4452
rect 12755 4387 12821 4388
rect 12942 4390 13124 4450
rect 12755 4316 12821 4317
rect 12755 4252 12756 4316
rect 12820 4252 12821 4316
rect 12755 4251 12821 4252
rect 12571 3772 12637 3773
rect 12571 3708 12572 3772
rect 12636 3708 12637 3772
rect 12571 3707 12637 3708
rect 12571 3636 12637 3637
rect 12571 3634 12572 3636
rect 12206 3574 12572 3634
rect 12571 3572 12572 3574
rect 12636 3572 12637 3636
rect 12571 3571 12637 3572
rect 12387 3364 12453 3365
rect 12387 3300 12388 3364
rect 12452 3300 12453 3364
rect 12387 3299 12453 3300
rect 11838 3166 12082 3226
rect 11838 2005 11898 3166
rect 12019 2820 12085 2821
rect 12019 2756 12020 2820
rect 12084 2756 12085 2820
rect 12019 2755 12085 2756
rect 12203 2820 12269 2821
rect 12203 2756 12204 2820
rect 12268 2756 12269 2820
rect 12203 2755 12269 2756
rect 11835 2004 11901 2005
rect 11835 1940 11836 2004
rect 11900 1940 11901 2004
rect 11835 1939 11901 1940
rect 12022 781 12082 2755
rect 12206 1461 12266 2755
rect 12203 1460 12269 1461
rect 12203 1396 12204 1460
rect 12268 1396 12269 1460
rect 12203 1395 12269 1396
rect 12019 780 12085 781
rect 12019 716 12020 780
rect 12084 716 12085 780
rect 12019 715 12085 716
rect 11651 372 11717 373
rect 11651 308 11652 372
rect 11716 308 11717 372
rect 11651 307 11717 308
rect 12390 237 12450 3299
rect 12758 2685 12818 4251
rect 12755 2684 12821 2685
rect 12755 2620 12756 2684
rect 12820 2620 12821 2684
rect 12755 2619 12821 2620
rect 12571 2548 12637 2549
rect 12571 2484 12572 2548
rect 12636 2484 12637 2548
rect 12571 2483 12637 2484
rect 12574 509 12634 2483
rect 12755 2412 12821 2413
rect 12755 2348 12756 2412
rect 12820 2348 12821 2412
rect 12755 2347 12821 2348
rect 12758 1189 12818 2347
rect 12942 2277 13002 4390
rect 13123 4388 13124 4390
rect 13188 4388 13189 4452
rect 13123 4387 13189 4388
rect 13306 3840 13626 4864
rect 13306 3776 13314 3840
rect 13378 3776 13394 3840
rect 13458 3776 13474 3840
rect 13538 3776 13554 3840
rect 13618 3776 13626 3840
rect 13123 3772 13189 3773
rect 13123 3708 13124 3772
rect 13188 3708 13189 3772
rect 13123 3707 13189 3708
rect 13126 3229 13186 3707
rect 13123 3228 13189 3229
rect 13123 3164 13124 3228
rect 13188 3164 13189 3228
rect 13123 3163 13189 3164
rect 13123 2820 13189 2821
rect 13123 2756 13124 2820
rect 13188 2756 13189 2820
rect 13123 2755 13189 2756
rect 12939 2276 13005 2277
rect 12939 2212 12940 2276
rect 13004 2212 13005 2276
rect 12939 2211 13005 2212
rect 12939 1868 13005 1869
rect 12939 1804 12940 1868
rect 13004 1804 13005 1868
rect 12939 1803 13005 1804
rect 12755 1188 12821 1189
rect 12755 1124 12756 1188
rect 12820 1124 12821 1188
rect 12755 1123 12821 1124
rect 12571 508 12637 509
rect 12571 444 12572 508
rect 12636 444 12637 508
rect 12571 443 12637 444
rect 12387 236 12453 237
rect 12387 172 12388 236
rect 12452 172 12453 236
rect 12387 171 12453 172
rect 12942 101 13002 1803
rect 13126 506 13186 2755
rect 13306 2752 13626 3776
rect 13862 3773 13922 5883
rect 14046 3906 14106 9830
rect 14227 6628 14293 6629
rect 14227 6564 14228 6628
rect 14292 6564 14293 6628
rect 14227 6563 14293 6564
rect 14230 4589 14290 6563
rect 14411 5948 14477 5949
rect 14411 5884 14412 5948
rect 14476 5884 14477 5948
rect 14411 5883 14477 5884
rect 14227 4588 14293 4589
rect 14227 4524 14228 4588
rect 14292 4524 14293 4588
rect 14227 4523 14293 4524
rect 14414 4450 14474 5883
rect 14230 4390 14474 4450
rect 14046 3846 14152 3906
rect 13862 3772 13971 3773
rect 13862 3710 13906 3772
rect 13905 3708 13906 3710
rect 13970 3708 13971 3772
rect 13905 3707 13971 3708
rect 14092 3090 14152 3846
rect 14230 3773 14290 4390
rect 14598 4314 14658 13363
rect 15150 13157 15210 14315
rect 15334 13973 15394 22067
rect 15778 21792 16098 22816
rect 16251 22404 16317 22405
rect 16251 22340 16252 22404
rect 16316 22340 16317 22404
rect 16251 22339 16317 22340
rect 15778 21728 15786 21792
rect 15850 21728 15866 21792
rect 15930 21728 15946 21792
rect 16010 21728 16026 21792
rect 16090 21728 16098 21792
rect 15515 21180 15581 21181
rect 15515 21116 15516 21180
rect 15580 21116 15581 21180
rect 15515 21115 15581 21116
rect 15518 16285 15578 21115
rect 15778 20704 16098 21728
rect 15778 20640 15786 20704
rect 15850 20640 15866 20704
rect 15930 20640 15946 20704
rect 16010 20640 16026 20704
rect 16090 20640 16098 20704
rect 15778 19616 16098 20640
rect 15778 19552 15786 19616
rect 15850 19552 15866 19616
rect 15930 19552 15946 19616
rect 16010 19552 16026 19616
rect 16090 19552 16098 19616
rect 15778 18528 16098 19552
rect 15778 18464 15786 18528
rect 15850 18464 15866 18528
rect 15930 18464 15946 18528
rect 16010 18464 16026 18528
rect 16090 18464 16098 18528
rect 15778 17440 16098 18464
rect 15778 17376 15786 17440
rect 15850 17376 15866 17440
rect 15930 17376 15946 17440
rect 16010 17376 16026 17440
rect 16090 17376 16098 17440
rect 15778 16352 16098 17376
rect 15778 16288 15786 16352
rect 15850 16288 15866 16352
rect 15930 16288 15946 16352
rect 16010 16288 16026 16352
rect 16090 16288 16098 16352
rect 15515 16284 15581 16285
rect 15515 16220 15516 16284
rect 15580 16220 15581 16284
rect 15515 16219 15581 16220
rect 15515 16148 15581 16149
rect 15515 16084 15516 16148
rect 15580 16084 15581 16148
rect 15515 16083 15581 16084
rect 15331 13972 15397 13973
rect 15331 13908 15332 13972
rect 15396 13908 15397 13972
rect 15331 13907 15397 13908
rect 15518 13157 15578 16083
rect 15778 15264 16098 16288
rect 15778 15200 15786 15264
rect 15850 15200 15866 15264
rect 15930 15200 15946 15264
rect 16010 15200 16026 15264
rect 16090 15200 16098 15264
rect 15778 14176 16098 15200
rect 15778 14112 15786 14176
rect 15850 14112 15866 14176
rect 15930 14112 15946 14176
rect 16010 14112 16026 14176
rect 16090 14112 16098 14176
rect 15147 13156 15213 13157
rect 15147 13092 15148 13156
rect 15212 13092 15213 13156
rect 15147 13091 15213 13092
rect 15515 13156 15581 13157
rect 15515 13092 15516 13156
rect 15580 13092 15581 13156
rect 15515 13091 15581 13092
rect 15518 11797 15578 13091
rect 15778 13088 16098 14112
rect 16254 13293 16314 22339
rect 16438 21181 16498 29139
rect 16622 26621 16682 30366
rect 16803 30156 16869 30157
rect 16803 30092 16804 30156
rect 16868 30092 16869 30156
rect 16803 30091 16869 30092
rect 16619 26620 16685 26621
rect 16619 26556 16620 26620
rect 16684 26556 16685 26620
rect 16619 26555 16685 26556
rect 16619 24172 16685 24173
rect 16619 24108 16620 24172
rect 16684 24108 16685 24172
rect 16619 24107 16685 24108
rect 16435 21180 16501 21181
rect 16435 21116 16436 21180
rect 16500 21116 16501 21180
rect 16435 21115 16501 21116
rect 16435 20772 16501 20773
rect 16435 20708 16436 20772
rect 16500 20708 16501 20772
rect 16435 20707 16501 20708
rect 16438 13565 16498 20707
rect 16435 13564 16501 13565
rect 16435 13500 16436 13564
rect 16500 13500 16501 13564
rect 16435 13499 16501 13500
rect 16622 13429 16682 24107
rect 16806 22110 16866 30091
rect 16990 29069 17050 40019
rect 17539 39812 17605 39813
rect 17539 39748 17540 39812
rect 17604 39748 17605 39812
rect 17539 39747 17605 39748
rect 17171 38724 17237 38725
rect 17171 38660 17172 38724
rect 17236 38660 17237 38724
rect 17171 38659 17237 38660
rect 16987 29068 17053 29069
rect 16987 29004 16988 29068
rect 17052 29004 17053 29068
rect 16987 29003 17053 29004
rect 16806 22050 17050 22110
rect 16803 15468 16869 15469
rect 16803 15404 16804 15468
rect 16868 15404 16869 15468
rect 16803 15403 16869 15404
rect 16619 13428 16685 13429
rect 16619 13364 16620 13428
rect 16684 13364 16685 13428
rect 16619 13363 16685 13364
rect 16251 13292 16317 13293
rect 16251 13228 16252 13292
rect 16316 13228 16317 13292
rect 16251 13227 16317 13228
rect 15778 13024 15786 13088
rect 15850 13024 15866 13088
rect 15930 13024 15946 13088
rect 16010 13024 16026 13088
rect 16090 13024 16098 13088
rect 15778 12000 16098 13024
rect 16254 12477 16314 13227
rect 16806 12749 16866 15403
rect 16990 15061 17050 22050
rect 16987 15060 17053 15061
rect 16987 14996 16988 15060
rect 17052 14996 17053 15060
rect 16987 14995 17053 14996
rect 16803 12748 16869 12749
rect 16803 12684 16804 12748
rect 16868 12684 16869 12748
rect 16803 12683 16869 12684
rect 16251 12476 16317 12477
rect 16251 12412 16252 12476
rect 16316 12412 16317 12476
rect 16251 12411 16317 12412
rect 17174 12338 17234 38659
rect 17355 34236 17421 34237
rect 17355 34172 17356 34236
rect 17420 34172 17421 34236
rect 17355 34171 17421 34172
rect 17358 30429 17418 34171
rect 17355 30428 17421 30429
rect 17355 30364 17356 30428
rect 17420 30364 17421 30428
rect 17355 30363 17421 30364
rect 17542 23629 17602 39747
rect 17723 32604 17789 32605
rect 17723 32540 17724 32604
rect 17788 32540 17789 32604
rect 17723 32539 17789 32540
rect 17726 29069 17786 32539
rect 17723 29068 17789 29069
rect 17723 29004 17724 29068
rect 17788 29004 17789 29068
rect 17723 29003 17789 29004
rect 17723 27028 17789 27029
rect 17723 26964 17724 27028
rect 17788 26964 17789 27028
rect 17723 26963 17789 26964
rect 17539 23628 17605 23629
rect 17539 23564 17540 23628
rect 17604 23564 17605 23628
rect 17539 23563 17605 23564
rect 17355 23492 17421 23493
rect 17355 23428 17356 23492
rect 17420 23428 17421 23492
rect 17355 23427 17421 23428
rect 17358 16557 17418 23427
rect 17726 19821 17786 26963
rect 17723 19820 17789 19821
rect 17723 19756 17724 19820
rect 17788 19756 17789 19820
rect 17723 19755 17789 19756
rect 17910 17970 17970 40019
rect 18251 39744 18571 40768
rect 20723 43552 21043 43568
rect 20723 43488 20731 43552
rect 20795 43488 20811 43552
rect 20875 43488 20891 43552
rect 20955 43488 20971 43552
rect 21035 43488 21043 43552
rect 20723 42464 21043 43488
rect 20723 42400 20731 42464
rect 20795 42400 20811 42464
rect 20875 42400 20891 42464
rect 20955 42400 20971 42464
rect 21035 42400 21043 42464
rect 20723 41376 21043 42400
rect 20723 41312 20731 41376
rect 20795 41312 20811 41376
rect 20875 41312 20891 41376
rect 20955 41312 20971 41376
rect 21035 41312 21043 41376
rect 20723 40288 21043 41312
rect 20723 40224 20731 40288
rect 20795 40224 20811 40288
rect 20875 40224 20891 40288
rect 20955 40224 20971 40288
rect 21035 40224 21043 40288
rect 18643 40084 18709 40085
rect 18643 40020 18644 40084
rect 18708 40020 18709 40084
rect 18643 40019 18709 40020
rect 18251 39680 18259 39744
rect 18323 39680 18339 39744
rect 18403 39680 18419 39744
rect 18483 39680 18499 39744
rect 18563 39680 18571 39744
rect 18251 38656 18571 39680
rect 18646 39269 18706 40019
rect 18643 39268 18709 39269
rect 18643 39204 18644 39268
rect 18708 39204 18709 39268
rect 18643 39203 18709 39204
rect 18251 38592 18259 38656
rect 18323 38592 18339 38656
rect 18403 38592 18419 38656
rect 18483 38592 18499 38656
rect 18563 38592 18571 38656
rect 18251 37568 18571 38592
rect 20723 39200 21043 40224
rect 20723 39136 20731 39200
rect 20795 39136 20811 39200
rect 20875 39136 20891 39200
rect 20955 39136 20971 39200
rect 21035 39136 21043 39200
rect 20723 38112 21043 39136
rect 20723 38048 20731 38112
rect 20795 38048 20811 38112
rect 20875 38048 20891 38112
rect 20955 38048 20971 38112
rect 21035 38048 21043 38112
rect 19011 37908 19077 37909
rect 19011 37844 19012 37908
rect 19076 37844 19077 37908
rect 19011 37843 19077 37844
rect 18251 37504 18259 37568
rect 18323 37504 18339 37568
rect 18403 37504 18419 37568
rect 18483 37504 18499 37568
rect 18563 37504 18571 37568
rect 18091 36956 18157 36957
rect 18091 36892 18092 36956
rect 18156 36892 18157 36956
rect 18091 36891 18157 36892
rect 18094 31381 18154 36891
rect 18251 36480 18571 37504
rect 18251 36416 18259 36480
rect 18323 36416 18339 36480
rect 18403 36416 18419 36480
rect 18483 36416 18499 36480
rect 18563 36416 18571 36480
rect 18251 35392 18571 36416
rect 18643 36412 18709 36413
rect 18643 36348 18644 36412
rect 18708 36348 18709 36412
rect 18643 36347 18709 36348
rect 18251 35328 18259 35392
rect 18323 35328 18339 35392
rect 18403 35328 18419 35392
rect 18483 35328 18499 35392
rect 18563 35328 18571 35392
rect 18251 34304 18571 35328
rect 18251 34240 18259 34304
rect 18323 34240 18339 34304
rect 18403 34240 18419 34304
rect 18483 34240 18499 34304
rect 18563 34240 18571 34304
rect 18251 33216 18571 34240
rect 18251 33152 18259 33216
rect 18323 33152 18339 33216
rect 18403 33152 18419 33216
rect 18483 33152 18499 33216
rect 18563 33152 18571 33216
rect 18251 32128 18571 33152
rect 18251 32064 18259 32128
rect 18323 32064 18339 32128
rect 18403 32064 18419 32128
rect 18483 32064 18499 32128
rect 18563 32064 18571 32128
rect 18091 31380 18157 31381
rect 18091 31316 18092 31380
rect 18156 31316 18157 31380
rect 18091 31315 18157 31316
rect 18251 31040 18571 32064
rect 18251 30976 18259 31040
rect 18323 30976 18339 31040
rect 18403 30976 18419 31040
rect 18483 30976 18499 31040
rect 18563 30976 18571 31040
rect 18251 29952 18571 30976
rect 18251 29888 18259 29952
rect 18323 29888 18339 29952
rect 18403 29888 18419 29952
rect 18483 29888 18499 29952
rect 18563 29888 18571 29952
rect 18251 28864 18571 29888
rect 18646 29205 18706 36347
rect 19014 36277 19074 37843
rect 19931 37364 19997 37365
rect 19931 37300 19932 37364
rect 19996 37300 19997 37364
rect 19931 37299 19997 37300
rect 19011 36276 19077 36277
rect 19011 36212 19012 36276
rect 19076 36212 19077 36276
rect 19011 36211 19077 36212
rect 18827 36140 18893 36141
rect 18827 36076 18828 36140
rect 18892 36076 18893 36140
rect 18827 36075 18893 36076
rect 18830 33285 18890 36075
rect 18827 33284 18893 33285
rect 18827 33220 18828 33284
rect 18892 33220 18893 33284
rect 18827 33219 18893 33220
rect 18827 33012 18893 33013
rect 18827 32948 18828 33012
rect 18892 32948 18893 33012
rect 18827 32947 18893 32948
rect 18643 29204 18709 29205
rect 18643 29140 18644 29204
rect 18708 29140 18709 29204
rect 18643 29139 18709 29140
rect 18251 28800 18259 28864
rect 18323 28800 18339 28864
rect 18403 28800 18419 28864
rect 18483 28800 18499 28864
rect 18563 28800 18571 28864
rect 18251 27776 18571 28800
rect 18251 27712 18259 27776
rect 18323 27712 18339 27776
rect 18403 27712 18419 27776
rect 18483 27712 18499 27776
rect 18563 27712 18571 27776
rect 18251 26688 18571 27712
rect 18251 26624 18259 26688
rect 18323 26624 18339 26688
rect 18403 26624 18419 26688
rect 18483 26624 18499 26688
rect 18563 26624 18571 26688
rect 18251 25600 18571 26624
rect 18251 25536 18259 25600
rect 18323 25536 18339 25600
rect 18403 25536 18419 25600
rect 18483 25536 18499 25600
rect 18563 25536 18571 25600
rect 18251 24512 18571 25536
rect 18251 24448 18259 24512
rect 18323 24448 18339 24512
rect 18403 24448 18419 24512
rect 18483 24448 18499 24512
rect 18563 24448 18571 24512
rect 18251 23424 18571 24448
rect 18251 23360 18259 23424
rect 18323 23360 18339 23424
rect 18403 23360 18419 23424
rect 18483 23360 18499 23424
rect 18563 23360 18571 23424
rect 18091 22540 18157 22541
rect 18091 22476 18092 22540
rect 18156 22476 18157 22540
rect 18091 22475 18157 22476
rect 18094 20637 18154 22475
rect 18251 22336 18571 23360
rect 18251 22272 18259 22336
rect 18323 22272 18339 22336
rect 18403 22272 18419 22336
rect 18483 22272 18499 22336
rect 18563 22272 18571 22336
rect 18251 21248 18571 22272
rect 18830 22110 18890 32947
rect 19014 30565 19074 36211
rect 19195 35868 19261 35869
rect 19195 35804 19196 35868
rect 19260 35804 19261 35868
rect 19195 35803 19261 35804
rect 19011 30564 19077 30565
rect 19011 30500 19012 30564
rect 19076 30500 19077 30564
rect 19011 30499 19077 30500
rect 19011 30428 19077 30429
rect 19011 30364 19012 30428
rect 19076 30364 19077 30428
rect 19011 30363 19077 30364
rect 18251 21184 18259 21248
rect 18323 21184 18339 21248
rect 18403 21184 18419 21248
rect 18483 21184 18499 21248
rect 18563 21184 18571 21248
rect 18091 20636 18157 20637
rect 18091 20572 18092 20636
rect 18156 20572 18157 20636
rect 18091 20571 18157 20572
rect 17726 17910 17970 17970
rect 18251 20160 18571 21184
rect 18251 20096 18259 20160
rect 18323 20096 18339 20160
rect 18403 20096 18419 20160
rect 18483 20096 18499 20160
rect 18563 20096 18571 20160
rect 18251 19072 18571 20096
rect 18251 19008 18259 19072
rect 18323 19008 18339 19072
rect 18403 19008 18419 19072
rect 18483 19008 18499 19072
rect 18563 19008 18571 19072
rect 18251 17984 18571 19008
rect 18251 17920 18259 17984
rect 18323 17920 18339 17984
rect 18403 17920 18419 17984
rect 18483 17920 18499 17984
rect 18563 17920 18571 17984
rect 17355 16556 17421 16557
rect 17355 16492 17356 16556
rect 17420 16492 17421 16556
rect 17355 16491 17421 16492
rect 17355 15060 17421 15061
rect 17355 14996 17356 15060
rect 17420 14996 17421 15060
rect 17355 14995 17421 14996
rect 15778 11936 15786 12000
rect 15850 11936 15866 12000
rect 15930 11936 15946 12000
rect 16010 11936 16026 12000
rect 16090 11936 16098 12000
rect 14963 11796 15029 11797
rect 14963 11732 14964 11796
rect 15028 11732 15029 11796
rect 14963 11731 15029 11732
rect 15331 11796 15397 11797
rect 15331 11732 15332 11796
rect 15396 11732 15397 11796
rect 15331 11731 15397 11732
rect 15515 11796 15581 11797
rect 15515 11732 15516 11796
rect 15580 11732 15581 11796
rect 15515 11731 15581 11732
rect 14966 9213 15026 11731
rect 15147 9484 15213 9485
rect 15147 9420 15148 9484
rect 15212 9420 15213 9484
rect 15147 9419 15213 9420
rect 14963 9212 15029 9213
rect 14963 9148 14964 9212
rect 15028 9148 15029 9212
rect 14963 9147 15029 9148
rect 14963 6764 15029 6765
rect 14963 6762 14964 6764
rect 14414 4254 14658 4314
rect 14782 6702 14964 6762
rect 14227 3772 14293 3773
rect 14227 3708 14228 3772
rect 14292 3708 14293 3772
rect 14227 3707 14293 3708
rect 13306 2688 13314 2752
rect 13378 2688 13394 2752
rect 13458 2688 13474 2752
rect 13538 2688 13554 2752
rect 13618 2688 13626 2752
rect 13306 1664 13626 2688
rect 14046 3030 14152 3090
rect 13859 2684 13925 2685
rect 13859 2620 13860 2684
rect 13924 2620 13925 2684
rect 13859 2619 13925 2620
rect 13306 1600 13314 1664
rect 13378 1600 13394 1664
rect 13458 1600 13474 1664
rect 13538 1600 13554 1664
rect 13618 1600 13626 1664
rect 13306 1040 13626 1600
rect 13862 1322 13922 2619
rect 14046 2410 14106 3030
rect 14227 2820 14293 2821
rect 14227 2756 14228 2820
rect 14292 2818 14293 2820
rect 14414 2818 14474 4254
rect 14782 4181 14842 6702
rect 14963 6700 14964 6702
rect 15028 6700 15029 6764
rect 14963 6699 15029 6700
rect 15150 6626 15210 9419
rect 14966 6566 15210 6626
rect 14779 4180 14845 4181
rect 14779 4116 14780 4180
rect 14844 4116 14845 4180
rect 14779 4115 14845 4116
rect 14966 3773 15026 6566
rect 15147 5268 15213 5269
rect 15147 5204 15148 5268
rect 15212 5204 15213 5268
rect 15147 5203 15213 5204
rect 15150 4725 15210 5203
rect 15147 4724 15213 4725
rect 15147 4660 15148 4724
rect 15212 4660 15213 4724
rect 15147 4659 15213 4660
rect 14595 3772 14661 3773
rect 14595 3708 14596 3772
rect 14660 3708 14661 3772
rect 14595 3707 14661 3708
rect 14963 3772 15029 3773
rect 14963 3708 14964 3772
rect 15028 3708 15029 3772
rect 14963 3707 15029 3708
rect 15147 3772 15213 3773
rect 15147 3708 15148 3772
rect 15212 3708 15213 3772
rect 15147 3707 15213 3708
rect 14292 2758 14474 2818
rect 14292 2756 14293 2758
rect 14227 2755 14293 2756
rect 14046 2350 14474 2410
rect 14043 1732 14109 1733
rect 14043 1668 14044 1732
rect 14108 1730 14109 1732
rect 14108 1670 14290 1730
rect 14108 1668 14109 1670
rect 14043 1667 14109 1668
rect 14230 1458 14290 1670
rect 14414 1597 14474 2350
rect 14598 2002 14658 3707
rect 14963 3636 15029 3637
rect 14963 3572 14964 3636
rect 15028 3572 15029 3636
rect 14963 3571 15029 3572
rect 14779 2004 14845 2005
rect 14779 2002 14780 2004
rect 14598 1942 14780 2002
rect 14779 1940 14780 1942
rect 14844 1940 14845 2004
rect 14779 1939 14845 1940
rect 14966 1733 15026 3571
rect 14963 1732 15029 1733
rect 14963 1668 14964 1732
rect 15028 1668 15029 1732
rect 14963 1667 15029 1668
rect 14411 1596 14477 1597
rect 14411 1532 14412 1596
rect 14476 1532 14477 1596
rect 14411 1531 14477 1532
rect 14230 1398 14474 1458
rect 14227 1324 14293 1325
rect 14227 1322 14228 1324
rect 13862 1262 14228 1322
rect 14227 1260 14228 1262
rect 14292 1260 14293 1324
rect 14227 1259 14293 1260
rect 14414 509 14474 1398
rect 14411 508 14477 509
rect 13126 446 14290 506
rect 14089 372 14155 373
rect 14089 308 14090 372
rect 14154 308 14155 372
rect 14230 370 14290 446
rect 14411 444 14412 508
rect 14476 444 14477 508
rect 14411 443 14477 444
rect 14779 372 14845 373
rect 14779 370 14780 372
rect 14230 310 14780 370
rect 14089 307 14155 308
rect 14779 308 14780 310
rect 14844 308 14845 372
rect 14779 307 14845 308
rect 14092 234 14152 307
rect 15150 234 15210 3707
rect 15334 2277 15394 11731
rect 15778 10912 16098 11936
rect 16438 12278 17234 12338
rect 16251 11524 16317 11525
rect 16251 11460 16252 11524
rect 16316 11460 16317 11524
rect 16251 11459 16317 11460
rect 15778 10848 15786 10912
rect 15850 10848 15866 10912
rect 15930 10848 15946 10912
rect 16010 10848 16026 10912
rect 16090 10848 16098 10912
rect 15515 10572 15581 10573
rect 15515 10508 15516 10572
rect 15580 10508 15581 10572
rect 15515 10507 15581 10508
rect 15518 6493 15578 10507
rect 15778 9824 16098 10848
rect 15778 9760 15786 9824
rect 15850 9760 15866 9824
rect 15930 9760 15946 9824
rect 16010 9760 16026 9824
rect 16090 9760 16098 9824
rect 15778 8736 16098 9760
rect 15778 8672 15786 8736
rect 15850 8672 15866 8736
rect 15930 8672 15946 8736
rect 16010 8672 16026 8736
rect 16090 8672 16098 8736
rect 15778 7648 16098 8672
rect 15778 7584 15786 7648
rect 15850 7584 15866 7648
rect 15930 7584 15946 7648
rect 16010 7584 16026 7648
rect 16090 7584 16098 7648
rect 15778 6560 16098 7584
rect 15778 6496 15786 6560
rect 15850 6496 15866 6560
rect 15930 6496 15946 6560
rect 16010 6496 16026 6560
rect 16090 6496 16098 6560
rect 15515 6492 15581 6493
rect 15515 6428 15516 6492
rect 15580 6428 15581 6492
rect 15515 6427 15581 6428
rect 15778 5472 16098 6496
rect 15778 5408 15786 5472
rect 15850 5408 15866 5472
rect 15930 5408 15946 5472
rect 16010 5408 16026 5472
rect 16090 5408 16098 5472
rect 15778 4384 16098 5408
rect 15778 4320 15786 4384
rect 15850 4320 15866 4384
rect 15930 4320 15946 4384
rect 16010 4320 16026 4384
rect 16090 4320 16098 4384
rect 15515 3908 15581 3909
rect 15515 3844 15516 3908
rect 15580 3844 15581 3908
rect 15515 3843 15581 3844
rect 15331 2276 15397 2277
rect 15331 2212 15332 2276
rect 15396 2212 15397 2276
rect 15331 2211 15397 2212
rect 15331 1188 15397 1189
rect 15331 1124 15332 1188
rect 15396 1124 15397 1188
rect 15331 1123 15397 1124
rect 15334 778 15394 1123
rect 15518 1053 15578 3843
rect 15778 3296 16098 4320
rect 15778 3232 15786 3296
rect 15850 3232 15866 3296
rect 15930 3232 15946 3296
rect 16010 3232 16026 3296
rect 16090 3232 16098 3296
rect 15778 2208 16098 3232
rect 16254 2790 16314 11459
rect 16438 3090 16498 12278
rect 17171 11932 17237 11933
rect 17171 11868 17172 11932
rect 17236 11868 17237 11932
rect 17171 11867 17237 11868
rect 16619 11524 16685 11525
rect 16619 11460 16620 11524
rect 16684 11460 16685 11524
rect 16619 11459 16685 11460
rect 16622 3365 16682 11459
rect 17174 10165 17234 11867
rect 17171 10164 17237 10165
rect 17171 10100 17172 10164
rect 17236 10100 17237 10164
rect 17171 10099 17237 10100
rect 16803 9348 16869 9349
rect 16803 9284 16804 9348
rect 16868 9284 16869 9348
rect 16803 9283 16869 9284
rect 16806 8125 16866 9283
rect 16987 8940 17053 8941
rect 16987 8876 16988 8940
rect 17052 8876 17053 8940
rect 16987 8875 17053 8876
rect 16803 8124 16869 8125
rect 16803 8060 16804 8124
rect 16868 8060 16869 8124
rect 16803 8059 16869 8060
rect 16990 4725 17050 8875
rect 17174 7309 17234 10099
rect 17171 7308 17237 7309
rect 17171 7244 17172 7308
rect 17236 7244 17237 7308
rect 17171 7243 17237 7244
rect 16987 4724 17053 4725
rect 16987 4660 16988 4724
rect 17052 4660 17053 4724
rect 16987 4659 17053 4660
rect 17358 4045 17418 14995
rect 17539 14652 17605 14653
rect 17539 14588 17540 14652
rect 17604 14588 17605 14652
rect 17539 14587 17605 14588
rect 17542 12341 17602 14587
rect 17726 13565 17786 17910
rect 18251 16896 18571 17920
rect 18251 16832 18259 16896
rect 18323 16832 18339 16896
rect 18403 16832 18419 16896
rect 18483 16832 18499 16896
rect 18563 16832 18571 16896
rect 18091 16556 18157 16557
rect 18091 16492 18092 16556
rect 18156 16492 18157 16556
rect 18091 16491 18157 16492
rect 17907 16012 17973 16013
rect 17907 15948 17908 16012
rect 17972 15948 17973 16012
rect 17907 15947 17973 15948
rect 17723 13564 17789 13565
rect 17723 13500 17724 13564
rect 17788 13500 17789 13564
rect 17723 13499 17789 13500
rect 17910 13426 17970 15947
rect 17726 13366 17970 13426
rect 17539 12340 17605 12341
rect 17539 12276 17540 12340
rect 17604 12276 17605 12340
rect 17539 12275 17605 12276
rect 17539 10708 17605 10709
rect 17539 10644 17540 10708
rect 17604 10644 17605 10708
rect 17539 10643 17605 10644
rect 17355 4044 17421 4045
rect 17355 3980 17356 4044
rect 17420 3980 17421 4044
rect 17355 3979 17421 3980
rect 17542 3773 17602 10643
rect 17726 7309 17786 13366
rect 18094 10029 18154 16491
rect 18251 15808 18571 16832
rect 18251 15744 18259 15808
rect 18323 15744 18339 15808
rect 18403 15744 18419 15808
rect 18483 15744 18499 15808
rect 18563 15744 18571 15808
rect 18251 14720 18571 15744
rect 18646 22050 18890 22110
rect 18646 15061 18706 22050
rect 19014 20909 19074 30363
rect 19198 27709 19258 35803
rect 19379 34100 19445 34101
rect 19379 34036 19380 34100
rect 19444 34036 19445 34100
rect 19379 34035 19445 34036
rect 19382 33285 19442 34035
rect 19747 33828 19813 33829
rect 19747 33764 19748 33828
rect 19812 33764 19813 33828
rect 19747 33763 19813 33764
rect 19750 33285 19810 33763
rect 19379 33284 19445 33285
rect 19379 33220 19380 33284
rect 19444 33220 19445 33284
rect 19379 33219 19445 33220
rect 19747 33284 19813 33285
rect 19747 33220 19748 33284
rect 19812 33220 19813 33284
rect 19747 33219 19813 33220
rect 19379 33012 19445 33013
rect 19379 32948 19380 33012
rect 19444 32948 19445 33012
rect 19379 32947 19445 32948
rect 19382 29613 19442 32947
rect 19747 31516 19813 31517
rect 19747 31452 19748 31516
rect 19812 31452 19813 31516
rect 19747 31451 19813 31452
rect 19379 29612 19445 29613
rect 19379 29548 19380 29612
rect 19444 29548 19445 29612
rect 19379 29547 19445 29548
rect 19379 28252 19445 28253
rect 19379 28188 19380 28252
rect 19444 28188 19445 28252
rect 19379 28187 19445 28188
rect 19195 27708 19261 27709
rect 19195 27644 19196 27708
rect 19260 27644 19261 27708
rect 19195 27643 19261 27644
rect 19195 24852 19261 24853
rect 19195 24788 19196 24852
rect 19260 24788 19261 24852
rect 19195 24787 19261 24788
rect 19011 20908 19077 20909
rect 19011 20844 19012 20908
rect 19076 20844 19077 20908
rect 19011 20843 19077 20844
rect 19198 18325 19258 24787
rect 19382 22405 19442 28187
rect 19563 25124 19629 25125
rect 19563 25060 19564 25124
rect 19628 25060 19629 25124
rect 19563 25059 19629 25060
rect 19379 22404 19445 22405
rect 19379 22340 19380 22404
rect 19444 22340 19445 22404
rect 19379 22339 19445 22340
rect 19566 22110 19626 25059
rect 19750 22541 19810 31451
rect 19934 31245 19994 37299
rect 20723 37024 21043 38048
rect 20723 36960 20731 37024
rect 20795 36960 20811 37024
rect 20875 36960 20891 37024
rect 20955 36960 20971 37024
rect 21035 36960 21043 37024
rect 20723 35936 21043 36960
rect 20723 35872 20731 35936
rect 20795 35872 20811 35936
rect 20875 35872 20891 35936
rect 20955 35872 20971 35936
rect 21035 35872 21043 35936
rect 20723 34848 21043 35872
rect 20723 34784 20731 34848
rect 20795 34784 20811 34848
rect 20875 34784 20891 34848
rect 20955 34784 20971 34848
rect 21035 34784 21043 34848
rect 20723 33760 21043 34784
rect 20723 33696 20731 33760
rect 20795 33696 20811 33760
rect 20875 33696 20891 33760
rect 20955 33696 20971 33760
rect 21035 33696 21043 33760
rect 20723 32672 21043 33696
rect 20723 32608 20731 32672
rect 20795 32608 20811 32672
rect 20875 32608 20891 32672
rect 20955 32608 20971 32672
rect 21035 32608 21043 32672
rect 20723 31584 21043 32608
rect 20723 31520 20731 31584
rect 20795 31520 20811 31584
rect 20875 31520 20891 31584
rect 20955 31520 20971 31584
rect 21035 31520 21043 31584
rect 19931 31244 19997 31245
rect 19931 31180 19932 31244
rect 19996 31180 19997 31244
rect 19931 31179 19997 31180
rect 20723 30496 21043 31520
rect 20723 30432 20731 30496
rect 20795 30432 20811 30496
rect 20875 30432 20891 30496
rect 20955 30432 20971 30496
rect 21035 30432 21043 30496
rect 20723 29408 21043 30432
rect 20723 29344 20731 29408
rect 20795 29344 20811 29408
rect 20875 29344 20891 29408
rect 20955 29344 20971 29408
rect 21035 29344 21043 29408
rect 20723 28320 21043 29344
rect 20723 28256 20731 28320
rect 20795 28256 20811 28320
rect 20875 28256 20891 28320
rect 20955 28256 20971 28320
rect 21035 28256 21043 28320
rect 20723 27232 21043 28256
rect 20723 27168 20731 27232
rect 20795 27168 20811 27232
rect 20875 27168 20891 27232
rect 20955 27168 20971 27232
rect 21035 27168 21043 27232
rect 20723 26144 21043 27168
rect 20723 26080 20731 26144
rect 20795 26080 20811 26144
rect 20875 26080 20891 26144
rect 20955 26080 20971 26144
rect 21035 26080 21043 26144
rect 20723 25056 21043 26080
rect 20723 24992 20731 25056
rect 20795 24992 20811 25056
rect 20875 24992 20891 25056
rect 20955 24992 20971 25056
rect 21035 24992 21043 25056
rect 20723 23968 21043 24992
rect 20723 23904 20731 23968
rect 20795 23904 20811 23968
rect 20875 23904 20891 23968
rect 20955 23904 20971 23968
rect 21035 23904 21043 23968
rect 20723 22880 21043 23904
rect 20723 22816 20731 22880
rect 20795 22816 20811 22880
rect 20875 22816 20891 22880
rect 20955 22816 20971 22880
rect 21035 22816 21043 22880
rect 19931 22676 19997 22677
rect 19931 22612 19932 22676
rect 19996 22612 19997 22676
rect 19931 22611 19997 22612
rect 19747 22540 19813 22541
rect 19747 22476 19748 22540
rect 19812 22476 19813 22540
rect 19747 22475 19813 22476
rect 19382 22050 19626 22110
rect 19195 18324 19261 18325
rect 19195 18260 19196 18324
rect 19260 18260 19261 18324
rect 19195 18259 19261 18260
rect 19382 16421 19442 22050
rect 19934 16826 19994 22611
rect 20723 21792 21043 22816
rect 20723 21728 20731 21792
rect 20795 21728 20811 21792
rect 20875 21728 20891 21792
rect 20955 21728 20971 21792
rect 21035 21728 21043 21792
rect 20723 20704 21043 21728
rect 20723 20640 20731 20704
rect 20795 20640 20811 20704
rect 20875 20640 20891 20704
rect 20955 20640 20971 20704
rect 21035 20640 21043 20704
rect 20723 19616 21043 20640
rect 20723 19552 20731 19616
rect 20795 19552 20811 19616
rect 20875 19552 20891 19616
rect 20955 19552 20971 19616
rect 21035 19552 21043 19616
rect 20723 18528 21043 19552
rect 20723 18464 20731 18528
rect 20795 18464 20811 18528
rect 20875 18464 20891 18528
rect 20955 18464 20971 18528
rect 21035 18464 21043 18528
rect 20115 18188 20181 18189
rect 20115 18124 20116 18188
rect 20180 18124 20181 18188
rect 20115 18123 20181 18124
rect 19566 16766 19994 16826
rect 19379 16420 19445 16421
rect 19379 16356 19380 16420
rect 19444 16356 19445 16420
rect 19379 16355 19445 16356
rect 18827 15196 18893 15197
rect 18827 15132 18828 15196
rect 18892 15132 18893 15196
rect 18827 15131 18893 15132
rect 18643 15060 18709 15061
rect 18643 14996 18644 15060
rect 18708 14996 18709 15060
rect 18643 14995 18709 14996
rect 18643 14924 18709 14925
rect 18643 14860 18644 14924
rect 18708 14860 18709 14924
rect 18643 14859 18709 14860
rect 18251 14656 18259 14720
rect 18323 14656 18339 14720
rect 18403 14656 18419 14720
rect 18483 14656 18499 14720
rect 18563 14656 18571 14720
rect 18251 13632 18571 14656
rect 18251 13568 18259 13632
rect 18323 13568 18339 13632
rect 18403 13568 18419 13632
rect 18483 13568 18499 13632
rect 18563 13568 18571 13632
rect 18251 12544 18571 13568
rect 18251 12480 18259 12544
rect 18323 12480 18339 12544
rect 18403 12480 18419 12544
rect 18483 12480 18499 12544
rect 18563 12480 18571 12544
rect 18251 11456 18571 12480
rect 18251 11392 18259 11456
rect 18323 11392 18339 11456
rect 18403 11392 18419 11456
rect 18483 11392 18499 11456
rect 18563 11392 18571 11456
rect 18251 10368 18571 11392
rect 18251 10304 18259 10368
rect 18323 10304 18339 10368
rect 18403 10304 18419 10368
rect 18483 10304 18499 10368
rect 18563 10304 18571 10368
rect 17907 10028 17973 10029
rect 17907 9964 17908 10028
rect 17972 9964 17973 10028
rect 17907 9963 17973 9964
rect 18091 10028 18157 10029
rect 18091 9964 18092 10028
rect 18156 9964 18157 10028
rect 18091 9963 18157 9964
rect 17723 7308 17789 7309
rect 17723 7244 17724 7308
rect 17788 7244 17789 7308
rect 17723 7243 17789 7244
rect 17539 3772 17605 3773
rect 17539 3708 17540 3772
rect 17604 3708 17605 3772
rect 17539 3707 17605 3708
rect 16619 3364 16685 3365
rect 16619 3300 16620 3364
rect 16684 3300 16685 3364
rect 16619 3299 16685 3300
rect 16438 3030 17050 3090
rect 16254 2730 16498 2790
rect 15778 2144 15786 2208
rect 15850 2144 15866 2208
rect 15930 2144 15946 2208
rect 16010 2144 16026 2208
rect 16090 2144 16098 2208
rect 15778 1120 16098 2144
rect 16251 2140 16317 2141
rect 16251 2076 16252 2140
rect 16316 2076 16317 2140
rect 16251 2075 16317 2076
rect 15778 1056 15786 1120
rect 15850 1056 15866 1120
rect 15930 1056 15946 1120
rect 16010 1056 16026 1120
rect 16090 1056 16098 1120
rect 15515 1052 15581 1053
rect 15515 988 15516 1052
rect 15580 988 15581 1052
rect 15778 1040 16098 1056
rect 15515 987 15581 988
rect 16254 778 16314 2075
rect 16438 1325 16498 2730
rect 16990 2413 17050 3030
rect 16987 2412 17053 2413
rect 16987 2348 16988 2412
rect 17052 2348 17053 2412
rect 16987 2347 17053 2348
rect 16435 1324 16501 1325
rect 16435 1260 16436 1324
rect 16500 1260 16501 1324
rect 16435 1259 16501 1260
rect 17910 1189 17970 9963
rect 18091 9348 18157 9349
rect 18091 9284 18092 9348
rect 18156 9284 18157 9348
rect 18091 9283 18157 9284
rect 18094 7037 18154 9283
rect 18251 9280 18571 10304
rect 18251 9216 18259 9280
rect 18323 9216 18339 9280
rect 18403 9216 18419 9280
rect 18483 9216 18499 9280
rect 18563 9216 18571 9280
rect 18251 8192 18571 9216
rect 18251 8128 18259 8192
rect 18323 8128 18339 8192
rect 18403 8128 18419 8192
rect 18483 8128 18499 8192
rect 18563 8128 18571 8192
rect 18251 7104 18571 8128
rect 18251 7040 18259 7104
rect 18323 7040 18339 7104
rect 18403 7040 18419 7104
rect 18483 7040 18499 7104
rect 18563 7040 18571 7104
rect 18091 7036 18157 7037
rect 18091 6972 18092 7036
rect 18156 6972 18157 7036
rect 18091 6971 18157 6972
rect 18251 6016 18571 7040
rect 18251 5952 18259 6016
rect 18323 5952 18339 6016
rect 18403 5952 18419 6016
rect 18483 5952 18499 6016
rect 18563 5952 18571 6016
rect 18251 4928 18571 5952
rect 18251 4864 18259 4928
rect 18323 4864 18339 4928
rect 18403 4864 18419 4928
rect 18483 4864 18499 4928
rect 18563 4864 18571 4928
rect 18251 3840 18571 4864
rect 18251 3776 18259 3840
rect 18323 3776 18339 3840
rect 18403 3776 18419 3840
rect 18483 3776 18499 3840
rect 18563 3776 18571 3840
rect 18251 2752 18571 3776
rect 18646 2821 18706 14859
rect 18830 10981 18890 15131
rect 19382 14650 19442 16355
rect 19014 14590 19442 14650
rect 18827 10980 18893 10981
rect 18827 10916 18828 10980
rect 18892 10916 18893 10980
rect 18827 10915 18893 10916
rect 18827 10164 18893 10165
rect 18827 10100 18828 10164
rect 18892 10100 18893 10164
rect 18827 10099 18893 10100
rect 18830 9213 18890 10099
rect 18827 9212 18893 9213
rect 18827 9148 18828 9212
rect 18892 9148 18893 9212
rect 18827 9147 18893 9148
rect 18643 2820 18709 2821
rect 18643 2756 18644 2820
rect 18708 2756 18709 2820
rect 18643 2755 18709 2756
rect 18251 2688 18259 2752
rect 18323 2688 18339 2752
rect 18403 2688 18419 2752
rect 18483 2688 18499 2752
rect 18563 2688 18571 2752
rect 18251 1664 18571 2688
rect 19014 2413 19074 14590
rect 19195 14516 19261 14517
rect 19195 14452 19196 14516
rect 19260 14452 19261 14516
rect 19195 14451 19261 14452
rect 19198 4317 19258 14451
rect 19566 12069 19626 16766
rect 19747 16692 19813 16693
rect 19747 16628 19748 16692
rect 19812 16628 19813 16692
rect 19747 16627 19813 16628
rect 19563 12068 19629 12069
rect 19563 12004 19564 12068
rect 19628 12004 19629 12068
rect 19563 12003 19629 12004
rect 19379 9348 19445 9349
rect 19379 9284 19380 9348
rect 19444 9284 19445 9348
rect 19379 9283 19445 9284
rect 19382 5541 19442 9283
rect 19563 8124 19629 8125
rect 19563 8060 19564 8124
rect 19628 8060 19629 8124
rect 19563 8059 19629 8060
rect 19379 5540 19445 5541
rect 19379 5476 19380 5540
rect 19444 5476 19445 5540
rect 19379 5475 19445 5476
rect 19195 4316 19261 4317
rect 19195 4252 19196 4316
rect 19260 4252 19261 4316
rect 19195 4251 19261 4252
rect 19566 2821 19626 8059
rect 19563 2820 19629 2821
rect 19563 2756 19564 2820
rect 19628 2756 19629 2820
rect 19563 2755 19629 2756
rect 19011 2412 19077 2413
rect 19011 2348 19012 2412
rect 19076 2348 19077 2412
rect 19011 2347 19077 2348
rect 19750 2005 19810 16627
rect 20118 14106 20178 18123
rect 19934 14046 20178 14106
rect 20723 17440 21043 18464
rect 20723 17376 20731 17440
rect 20795 17376 20811 17440
rect 20875 17376 20891 17440
rect 20955 17376 20971 17440
rect 21035 17376 21043 17440
rect 20723 16352 21043 17376
rect 20723 16288 20731 16352
rect 20795 16288 20811 16352
rect 20875 16288 20891 16352
rect 20955 16288 20971 16352
rect 21035 16288 21043 16352
rect 20723 15264 21043 16288
rect 20723 15200 20731 15264
rect 20795 15200 20811 15264
rect 20875 15200 20891 15264
rect 20955 15200 20971 15264
rect 21035 15200 21043 15264
rect 20723 14176 21043 15200
rect 20723 14112 20731 14176
rect 20795 14112 20811 14176
rect 20875 14112 20891 14176
rect 20955 14112 20971 14176
rect 21035 14112 21043 14176
rect 19934 9077 19994 14046
rect 20115 13972 20181 13973
rect 20115 13908 20116 13972
rect 20180 13908 20181 13972
rect 20115 13907 20181 13908
rect 19931 9076 19997 9077
rect 19931 9012 19932 9076
rect 19996 9012 19997 9076
rect 19931 9011 19997 9012
rect 19934 4453 19994 9011
rect 19931 4452 19997 4453
rect 19931 4388 19932 4452
rect 19996 4388 19997 4452
rect 19931 4387 19997 4388
rect 19747 2004 19813 2005
rect 19747 1940 19748 2004
rect 19812 1940 19813 2004
rect 19747 1939 19813 1940
rect 18251 1600 18259 1664
rect 18323 1600 18339 1664
rect 18403 1600 18419 1664
rect 18483 1600 18499 1664
rect 18563 1600 18571 1664
rect 17907 1188 17973 1189
rect 17907 1124 17908 1188
rect 17972 1124 17973 1188
rect 17907 1123 17973 1124
rect 18251 1040 18571 1600
rect 20118 1325 20178 13907
rect 20723 13088 21043 14112
rect 20723 13024 20731 13088
rect 20795 13024 20811 13088
rect 20875 13024 20891 13088
rect 20955 13024 20971 13088
rect 21035 13024 21043 13088
rect 20299 12748 20365 12749
rect 20299 12684 20300 12748
rect 20364 12684 20365 12748
rect 20299 12683 20365 12684
rect 20302 9213 20362 12683
rect 20723 12000 21043 13024
rect 20723 11936 20731 12000
rect 20795 11936 20811 12000
rect 20875 11936 20891 12000
rect 20955 11936 20971 12000
rect 21035 11936 21043 12000
rect 20723 10912 21043 11936
rect 20723 10848 20731 10912
rect 20795 10848 20811 10912
rect 20875 10848 20891 10912
rect 20955 10848 20971 10912
rect 21035 10848 21043 10912
rect 20723 9824 21043 10848
rect 20723 9760 20731 9824
rect 20795 9760 20811 9824
rect 20875 9760 20891 9824
rect 20955 9760 20971 9824
rect 21035 9760 21043 9824
rect 20299 9212 20365 9213
rect 20299 9148 20300 9212
rect 20364 9148 20365 9212
rect 20299 9147 20365 9148
rect 20723 8736 21043 9760
rect 20723 8672 20731 8736
rect 20795 8672 20811 8736
rect 20875 8672 20891 8736
rect 20955 8672 20971 8736
rect 21035 8672 21043 8736
rect 20723 7648 21043 8672
rect 20723 7584 20731 7648
rect 20795 7584 20811 7648
rect 20875 7584 20891 7648
rect 20955 7584 20971 7648
rect 21035 7584 21043 7648
rect 20723 6560 21043 7584
rect 20723 6496 20731 6560
rect 20795 6496 20811 6560
rect 20875 6496 20891 6560
rect 20955 6496 20971 6560
rect 21035 6496 21043 6560
rect 20723 5472 21043 6496
rect 20723 5408 20731 5472
rect 20795 5408 20811 5472
rect 20875 5408 20891 5472
rect 20955 5408 20971 5472
rect 21035 5408 21043 5472
rect 20723 4384 21043 5408
rect 20723 4320 20731 4384
rect 20795 4320 20811 4384
rect 20875 4320 20891 4384
rect 20955 4320 20971 4384
rect 21035 4320 21043 4384
rect 20723 3296 21043 4320
rect 20723 3232 20731 3296
rect 20795 3232 20811 3296
rect 20875 3232 20891 3296
rect 20955 3232 20971 3296
rect 21035 3232 21043 3296
rect 20723 2208 21043 3232
rect 20723 2144 20731 2208
rect 20795 2144 20811 2208
rect 20875 2144 20891 2208
rect 20955 2144 20971 2208
rect 21035 2144 21043 2208
rect 20115 1324 20181 1325
rect 20115 1260 20116 1324
rect 20180 1260 20181 1324
rect 20115 1259 20181 1260
rect 20723 1120 21043 2144
rect 20723 1056 20731 1120
rect 20795 1056 20811 1120
rect 20875 1056 20891 1120
rect 20955 1056 20971 1120
rect 21035 1056 21043 1120
rect 20723 1040 21043 1056
rect 15334 718 16314 778
rect 15699 644 15765 645
rect 15699 580 15700 644
rect 15764 580 15765 644
rect 15699 579 15765 580
rect 15702 506 15762 579
rect 16067 508 16133 509
rect 16067 506 16068 508
rect 15702 446 16068 506
rect 16067 444 16068 446
rect 16132 444 16133 508
rect 16067 443 16133 444
rect 14092 174 15210 234
rect 6683 100 6749 101
rect 6683 36 6684 100
rect 6748 36 6749 100
rect 6683 35 6749 36
rect 8155 100 8221 101
rect 8155 36 8156 100
rect 8220 36 8221 100
rect 8155 35 8221 36
rect 12939 100 13005 101
rect 12939 36 12940 100
rect 13004 36 13005 100
rect 12939 35 13005 36
use sky130_fd_sc_hd__clkbuf_1  _000_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19596 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _001_
timestamp 1688980957
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _002_
timestamp 1688980957
transform 1 0 19780 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _003_
timestamp 1688980957
transform 1 0 19780 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _004_
timestamp 1688980957
transform 1 0 19412 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp 1688980957
transform 1 0 17848 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _006_
timestamp 1688980957
transform 1 0 18768 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _007_
timestamp 1688980957
transform 1 0 18860 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _008_
timestamp 1688980957
transform 1 0 18124 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _009_
timestamp 1688980957
transform 1 0 19780 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _010_
timestamp 1688980957
transform 1 0 18032 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _011_
timestamp 1688980957
transform 1 0 20332 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _012_
timestamp 1688980957
transform 1 0 18584 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _013_
timestamp 1688980957
transform 1 0 18308 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _014_
timestamp 1688980957
transform 1 0 18032 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _015_
timestamp 1688980957
transform 1 0 17664 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _016_
timestamp 1688980957
transform 1 0 18676 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _017_
timestamp 1688980957
transform 1 0 18584 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _018_
timestamp 1688980957
transform 1 0 19780 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _019_
timestamp 1688980957
transform 1 0 18216 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _020_
timestamp 1688980957
transform 1 0 17940 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _021_
timestamp 1688980957
transform 1 0 19780 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _022_
timestamp 1688980957
transform 1 0 19596 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _023_
timestamp 1688980957
transform 1 0 18768 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _024_
timestamp 1688980957
transform 1 0 19780 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp 1688980957
transform 1 0 17940 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp 1688980957
transform 1 0 16376 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _027_
timestamp 1688980957
transform 1 0 18584 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _028_
timestamp 1688980957
transform 1 0 17296 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_
timestamp 1688980957
transform 1 0 18032 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform 1 0 17756 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform 1 0 18216 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform 1 0 15824 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp 1688980957
transform 1 0 19504 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform 1 0 12144 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform 1 0 13708 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp 1688980957
transform 1 0 17572 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp 1688980957
transform 1 0 16560 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform 1 0 17388 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform 1 0 13432 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform 1 0 12696 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform 1 0 14076 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform 1 0 13156 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform 1 0 17572 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp 1688980957
transform 1 0 17664 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform 1 0 18308 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform 1 0 17112 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp 1688980957
transform 1 0 18492 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp 1688980957
transform 1 0 17480 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _052_
timestamp 1688980957
transform 1 0 10396 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp 1688980957
transform 1 0 1472 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp 1688980957
transform 1 0 2852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1688980957
transform 1 0 12328 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1688980957
transform 1 0 2576 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1688980957
transform 1 0 2300 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform 1 0 3680 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform 1 0 3404 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 3128 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1688980957
transform 1 0 12604 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1688980957
transform 1 0 1748 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1688980957
transform 1 0 3956 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 3864 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform 1 0 4232 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform 1 0 5060 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1688980957
transform 1 0 4784 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1688980957
transform 1 0 4692 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform 1 0 3680 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 5796 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform 1 0 4140 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 6532 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform 1 0 4416 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform 1 0 5520 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform 1 0 4876 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 6808 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 7912 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform 1 0 9200 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform 1 0 8280 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 11868 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform 1 0 8556 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1688980957
transform 1 0 9844 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform 1 0 8924 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform 1 0 6440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform 1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform 1 0 6992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1688980957
transform 1 0 9476 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _098_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1688980957
transform 1 0 20332 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1688980957
transform 1 0 8648 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1688980957
transform 1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1688980957
transform 1 0 9568 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1688980957
transform 1 0 9752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1688980957
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1688980957
transform 1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1688980957
transform 1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1688980957
transform 1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1688980957
transform 1 0 12144 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1688980957
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1688980957
transform 1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1688980957
transform 1 0 10856 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1688980957
transform 1 0 9292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _124_
timestamp 1688980957
transform 1 0 10212 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1688980957
transform 1 0 4600 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _127_
timestamp 1688980957
transform 1 0 13064 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp 1688980957
transform 1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1688980957
transform 1 0 5888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1688980957
transform 1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1688980957
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1688980957
transform 1 0 4324 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1688980957
transform 1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _136_
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1688980957
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1688980957
transform 1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _145_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3864 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1688980957
transform 1 0 3312 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1688980957
transform 1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1688980957
transform 1 0 4324 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform 1 0 1564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1688980957
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1688980957
transform 1 0 4232 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1688980957
transform 1 0 3036 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1688980957
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _155_
timestamp 1688980957
transform 1 0 1472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1688980957
transform 1 0 4324 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1688980957
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1688980957
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1688980957
transform 1 0 6532 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1688980957
transform 1 0 1472 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1688980957
transform 1 0 2024 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1688980957
transform 1 0 6808 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1688980957
transform 1 0 4324 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1688980957
transform 1 0 4508 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1688980957
transform 1 0 1564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1688980957
transform 1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _171_
timestamp 1688980957
transform 1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9844 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 10120 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 6348 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 7728 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 9752 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 16192 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 4508 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1688980957
transform 1 0 4232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1688980957
transform 1 0 8280 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1688980957
transform 1 0 19688 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1688980957
transform 1 0 6348 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1688980957
transform 1 0 14536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1688980957
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1688980957
transform 1 0 11868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1688980957
transform 1 0 9108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1688980957
transform 1 0 9384 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1688980957
transform 1 0 19412 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1688980957
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1688980957
transform 1 0 2300 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0._0_
timestamp 1688980957
transform 1 0 18308 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1._0_
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2._0_
timestamp 1688980957
transform 1 0 18124 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3._0_
timestamp 1688980957
transform 1 0 18400 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4._0_
timestamp 1688980957
transform 1 0 18952 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5._0_
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6._0_
timestamp 1688980957
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7._0_
timestamp 1688980957
transform 1 0 19044 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8._0_
timestamp 1688980957
transform 1 0 17940 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9._0_
timestamp 1688980957
transform 1 0 17572 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10._0_
timestamp 1688980957
transform 1 0 17112 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11._0_
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12._0_
timestamp 1688980957
transform 1 0 18860 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13._0_
timestamp 1688980957
transform 1 0 18584 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14._0_
timestamp 1688980957
transform 1 0 19136 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15._0_
timestamp 1688980957
transform 1 0 17756 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16._0_
timestamp 1688980957
transform 1 0 17940 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17._0_
timestamp 1688980957
transform 1 0 15548 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18._0_
timestamp 1688980957
transform 1 0 18308 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19._0_
timestamp 1688980957
transform 1 0 18216 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20._0_
timestamp 1688980957
transform 1 0 17940 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21._0_
timestamp 1688980957
transform 1 0 18768 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22._0_
timestamp 1688980957
transform 1 0 18676 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23._0_
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24._0_
timestamp 1688980957
transform 1 0 18216 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25._0_
timestamp 1688980957
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26._0_
timestamp 1688980957
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27._0_
timestamp 1688980957
transform 1 0 17940 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28._0_
timestamp 1688980957
transform 1 0 19596 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29._0_
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30._0_
timestamp 1688980957
transform 1 0 18400 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31._0_
timestamp 1688980957
transform 1 0 18124 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0._0_
timestamp 1688980957
transform 1 0 19136 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1._0_
timestamp 1688980957
transform 1 0 18584 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2._0_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3._0_
timestamp 1688980957
transform 1 0 19228 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4._0_
timestamp 1688980957
transform 1 0 19412 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5._0_
timestamp 1688980957
transform 1 0 19504 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6._0_
timestamp 1688980957
transform 1 0 18584 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7._0_
timestamp 1688980957
transform 1 0 18584 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8._0_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9._0_
timestamp 1688980957
transform 1 0 18308 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10._0_
timestamp 1688980957
transform 1 0 19596 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11._0_
timestamp 1688980957
transform 1 0 19412 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12._0_
timestamp 1688980957
transform 1 0 19412 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13._0_
timestamp 1688980957
transform 1 0 19136 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14._0_
timestamp 1688980957
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15._0_
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16._0_
timestamp 1688980957
transform 1 0 18400 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17._0_
timestamp 1688980957
transform 1 0 17112 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18._0_
timestamp 1688980957
transform 1 0 19504 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19._0_
timestamp 1688980957
transform 1 0 19780 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20._0_
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21._0_
timestamp 1688980957
transform 1 0 18952 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22._0_
timestamp 1688980957
transform 1 0 19412 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23._0_
timestamp 1688980957
transform 1 0 19044 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24._0_
timestamp 1688980957
transform 1 0 19320 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25._0_
timestamp 1688980957
transform 1 0 19504 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26._0_
timestamp 1688980957
transform 1 0 19228 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27._0_
timestamp 1688980957
transform 1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28._0_
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29._0_
timestamp 1688980957
transform 1 0 17664 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30._0_
timestamp 1688980957
transform 1 0 10856 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31._0_
timestamp 1688980957
transform 1 0 14904 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_11
timestamp 1688980957
transform 1 0 2116 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_21
timestamp 1688980957
transform 1 0 3036 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_35
timestamp 1688980957
transform 1 0 4324 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_155
timestamp 1688980957
transform 1 0 15364 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_23
timestamp 1688980957
transform 1 0 3220 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_32
timestamp 1688980957
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_51
timestamp 1688980957
transform 1 0 5796 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_66
timestamp 1688980957
transform 1 0 7176 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_71
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_75
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_108
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_128
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_132
timestamp 1688980957
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_144
timestamp 1688980957
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_168
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_187
timestamp 1688980957
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_191
timestamp 1688980957
transform 1 0 18676 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_203
timestamp 1688980957
transform 1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_207
timestamp 1688980957
transform 1 0 20148 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_32
timestamp 1688980957
transform 1 0 4048 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_36 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_48
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_54
timestamp 1688980957
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_129
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_211
timestamp 1688980957
transform 1 0 20516 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_26
timestamp 1688980957
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_68
timestamp 1688980957
transform 1 0 7360 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_75
timestamp 1688980957
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_80
timestamp 1688980957
transform 1 0 8464 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_88
timestamp 1688980957
transform 1 0 9200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_92
timestamp 1688980957
transform 1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_101
timestamp 1688980957
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_106
timestamp 1688980957
transform 1 0 10856 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_131
timestamp 1688980957
transform 1 0 13156 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_138
timestamp 1688980957
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_159
timestamp 1688980957
transform 1 0 15732 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_210
timestamp 1688980957
transform 1 0 20424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_12
timestamp 1688980957
transform 1 0 2208 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_37
timestamp 1688980957
transform 1 0 4508 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_85
timestamp 1688980957
transform 1 0 8924 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_89
timestamp 1688980957
transform 1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_129
timestamp 1688980957
transform 1 0 12972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_140
timestamp 1688980957
transform 1 0 13984 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_157
timestamp 1688980957
transform 1 0 15548 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_12
timestamp 1688980957
transform 1 0 2208 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_76 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8096 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_85 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_89
timestamp 1688980957
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_92
timestamp 1688980957
transform 1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_96
timestamp 1688980957
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_112
timestamp 1688980957
transform 1 0 11408 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_154
timestamp 1688980957
transform 1 0 15272 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_210
timestamp 1688980957
transform 1 0 20424 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_33
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_75
timestamp 1688980957
transform 1 0 8004 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_118
timestamp 1688980957
transform 1 0 11960 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_128
timestamp 1688980957
transform 1 0 12880 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_136
timestamp 1688980957
transform 1 0 13616 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_166
timestamp 1688980957
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_195
timestamp 1688980957
transform 1 0 19044 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_9
timestamp 1688980957
transform 1 0 1932 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_68
timestamp 1688980957
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_80
timestamp 1688980957
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_115
timestamp 1688980957
transform 1 0 11684 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_119
timestamp 1688980957
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_172
timestamp 1688980957
transform 1 0 16928 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_190
timestamp 1688980957
transform 1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_60
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_102
timestamp 1688980957
transform 1 0 10488 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_128
timestamp 1688980957
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_164
timestamp 1688980957
transform 1 0 16192 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_89
timestamp 1688980957
transform 1 0 9292 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_210
timestamp 1688980957
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_21
timestamp 1688980957
transform 1 0 3036 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_60
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_68
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_73
timestamp 1688980957
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_140
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_184
timestamp 1688980957
transform 1 0 18032 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_204
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_12
timestamp 1688980957
transform 1 0 2208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_100
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_117
timestamp 1688980957
transform 1 0 11868 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_159
timestamp 1688980957
transform 1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_210
timestamp 1688980957
transform 1 0 20424 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_54
timestamp 1688980957
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_90
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_151
timestamp 1688980957
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_175
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_179
timestamp 1688980957
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_11
timestamp 1688980957
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_174
timestamp 1688980957
transform 1 0 17112 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_60
timestamp 1688980957
transform 1 0 6624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_130
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_185
timestamp 1688980957
transform 1 0 18124 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_210
timestamp 1688980957
transform 1 0 20424 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_23
timestamp 1688980957
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_38
timestamp 1688980957
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_91
timestamp 1688980957
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_128
timestamp 1688980957
transform 1 0 12880 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_9
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_106
timestamp 1688980957
transform 1 0 10856 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_128
timestamp 1688980957
transform 1 0 12880 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_135
timestamp 1688980957
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_171
timestamp 1688980957
transform 1 0 16836 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_9
timestamp 1688980957
transform 1 0 1932 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_11
timestamp 1688980957
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_89
timestamp 1688980957
transform 1 0 9292 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_111
timestamp 1688980957
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_181
timestamp 1688980957
transform 1 0 17756 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_185
timestamp 1688980957
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_35
timestamp 1688980957
transform 1 0 4324 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_63
timestamp 1688980957
transform 1 0 6900 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_135
timestamp 1688980957
transform 1 0 13524 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_164
timestamp 1688980957
transform 1 0 16192 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_188
timestamp 1688980957
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_9
timestamp 1688980957
transform 1 0 1932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_26
timestamp 1688980957
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_74
timestamp 1688980957
transform 1 0 7912 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_93
timestamp 1688980957
transform 1 0 9660 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_115
timestamp 1688980957
transform 1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_135
timestamp 1688980957
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_192
timestamp 1688980957
transform 1 0 18768 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_11
timestamp 1688980957
transform 1 0 2116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_40
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_78
timestamp 1688980957
transform 1 0 8280 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_90
timestamp 1688980957
transform 1 0 9384 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_121
timestamp 1688980957
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_155
timestamp 1688980957
transform 1 0 15364 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_191
timestamp 1688980957
transform 1 0 18676 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_195
timestamp 1688980957
transform 1 0 19044 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_50
timestamp 1688980957
transform 1 0 5704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_110
timestamp 1688980957
transform 1 0 11224 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_132
timestamp 1688980957
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_78
timestamp 1688980957
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_155
timestamp 1688980957
transform 1 0 15364 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_204
timestamp 1688980957
transform 1 0 19872 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_38
timestamp 1688980957
transform 1 0 4600 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_131
timestamp 1688980957
transform 1 0 13156 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_192
timestamp 1688980957
transform 1 0 18768 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_18
timestamp 1688980957
transform 1 0 2760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_79
timestamp 1688980957
transform 1 0 8372 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_104
timestamp 1688980957
transform 1 0 10672 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_121
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_139
timestamp 1688980957
transform 1 0 13892 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_162
timestamp 1688980957
transform 1 0 16008 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_190
timestamp 1688980957
transform 1 0 18584 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_11
timestamp 1688980957
transform 1 0 2116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_65
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_93
timestamp 1688980957
transform 1 0 9660 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_112
timestamp 1688980957
transform 1 0 11408 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 1688980957
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_191
timestamp 1688980957
transform 1 0 18676 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_201
timestamp 1688980957
transform 1 0 19596 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_9
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_40
timestamp 1688980957
transform 1 0 4784 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_106
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_159
timestamp 1688980957
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_184
timestamp 1688980957
transform 1 0 18032 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_7
timestamp 1688980957
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_47
timestamp 1688980957
transform 1 0 5428 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_76
timestamp 1688980957
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_114
timestamp 1688980957
transform 1 0 11592 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_120
timestamp 1688980957
transform 1 0 12144 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_136
timestamp 1688980957
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_147
timestamp 1688980957
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_178
timestamp 1688980957
transform 1 0 17480 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_190
timestamp 1688980957
transform 1 0 18584 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_7
timestamp 1688980957
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_23
timestamp 1688980957
transform 1 0 3220 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_42
timestamp 1688980957
transform 1 0 4968 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1688980957
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_65
timestamp 1688980957
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_130
timestamp 1688980957
transform 1 0 13064 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_157
timestamp 1688980957
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1688980957
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_187
timestamp 1688980957
transform 1 0 18308 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_204
timestamp 1688980957
transform 1 0 19872 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_11
timestamp 1688980957
transform 1 0 2116 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_26
timestamp 1688980957
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_68
timestamp 1688980957
transform 1 0 7360 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_93
timestamp 1688980957
transform 1 0 9660 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_113
timestamp 1688980957
transform 1 0 11500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1688980957
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_149
timestamp 1688980957
transform 1 0 14812 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_186
timestamp 1688980957
transform 1 0 18216 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_192
timestamp 1688980957
transform 1 0 18768 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_7
timestamp 1688980957
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_42
timestamp 1688980957
transform 1 0 4968 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_54
timestamp 1688980957
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_110
timestamp 1688980957
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 1688980957
transform 1 0 11868 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_136
timestamp 1688980957
transform 1 0 13616 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_163
timestamp 1688980957
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 1688980957
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_194
timestamp 1688980957
transform 1 0 18952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_198
timestamp 1688980957
transform 1 0 19320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_63
timestamp 1688980957
transform 1 0 6900 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_136
timestamp 1688980957
transform 1 0 13616 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_171
timestamp 1688980957
transform 1 0 16836 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_175
timestamp 1688980957
transform 1 0 17204 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_181
timestamp 1688980957
transform 1 0 17756 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_185
timestamp 1688980957
transform 1 0 18124 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_20
timestamp 1688980957
transform 1 0 2944 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_40
timestamp 1688980957
transform 1 0 4784 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_80
timestamp 1688980957
transform 1 0 8464 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_100
timestamp 1688980957
transform 1 0 10304 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_130
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_185
timestamp 1688980957
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_189
timestamp 1688980957
transform 1 0 18492 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_210
timestamp 1688980957
transform 1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_66
timestamp 1688980957
transform 1 0 7176 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_100
timestamp 1688980957
transform 1 0 10304 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_127
timestamp 1688980957
transform 1 0 12788 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_132
timestamp 1688980957
transform 1 0 13248 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_172
timestamp 1688980957
transform 1 0 16928 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_184
timestamp 1688980957
transform 1 0 18032 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_210
timestamp 1688980957
transform 1 0 20424 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_19
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_36
timestamp 1688980957
transform 1 0 4416 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_72
timestamp 1688980957
transform 1 0 7728 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_91
timestamp 1688980957
transform 1 0 9476 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_164
timestamp 1688980957
transform 1 0 16192 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_175
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_201
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_9
timestamp 1688980957
transform 1 0 1932 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_33
timestamp 1688980957
transform 1 0 4140 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_55
timestamp 1688980957
transform 1 0 6164 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_59
timestamp 1688980957
transform 1 0 6532 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_76
timestamp 1688980957
transform 1 0 8096 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_91
timestamp 1688980957
transform 1 0 9476 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_97
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_116
timestamp 1688980957
transform 1 0 11776 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1688980957
transform 1 0 13708 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_159
timestamp 1688980957
transform 1 0 15732 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_192
timestamp 1688980957
transform 1 0 18768 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_6
timestamp 1688980957
transform 1 0 1656 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_54
timestamp 1688980957
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_60
timestamp 1688980957
transform 1 0 6624 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_72
timestamp 1688980957
transform 1 0 7728 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_128
timestamp 1688980957
transform 1 0 12880 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_140
timestamp 1688980957
transform 1 0 13984 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_144
timestamp 1688980957
transform 1 0 14352 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_166
timestamp 1688980957
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_184
timestamp 1688980957
transform 1 0 18032 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_204
timestamp 1688980957
transform 1 0 19872 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_24
timestamp 1688980957
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_44
timestamp 1688980957
transform 1 0 5152 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_56
timestamp 1688980957
transform 1 0 6256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_82
timestamp 1688980957
transform 1 0 8648 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_88
timestamp 1688980957
transform 1 0 9200 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_107
timestamp 1688980957
transform 1 0 10948 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_125
timestamp 1688980957
transform 1 0 12604 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_137
timestamp 1688980957
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_166
timestamp 1688980957
transform 1 0 16376 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_178
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_186
timestamp 1688980957
transform 1 0 18216 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_201
timestamp 1688980957
transform 1 0 19596 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_78
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_86
timestamp 1688980957
transform 1 0 9016 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_107
timestamp 1688980957
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_134
timestamp 1688980957
transform 1 0 13432 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_157
timestamp 1688980957
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_165
timestamp 1688980957
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_184
timestamp 1688980957
transform 1 0 18032 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_192
timestamp 1688980957
transform 1 0 18768 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_201
timestamp 1688980957
transform 1 0 19596 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_22
timestamp 1688980957
transform 1 0 3128 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_44
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_81
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_107
timestamp 1688980957
transform 1 0 10948 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_111
timestamp 1688980957
transform 1 0 11316 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 1688980957
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_159
timestamp 1688980957
transform 1 0 15732 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_19
timestamp 1688980957
transform 1 0 2852 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_53
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_72
timestamp 1688980957
transform 1 0 7728 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_107
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_158
timestamp 1688980957
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_202
timestamp 1688980957
transform 1 0 19688 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_210
timestamp 1688980957
transform 1 0 20424 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_6
timestamp 1688980957
transform 1 0 1656 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_25
timestamp 1688980957
transform 1 0 3404 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_47
timestamp 1688980957
transform 1 0 5428 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_70
timestamp 1688980957
transform 1 0 7544 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_100
timestamp 1688980957
transform 1 0 10304 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_112
timestamp 1688980957
transform 1 0 11408 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_118
timestamp 1688980957
transform 1 0 11960 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_174
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_186
timestamp 1688980957
transform 1 0 18216 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_24
timestamp 1688980957
transform 1 0 3312 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_84
timestamp 1688980957
transform 1 0 8832 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_106
timestamp 1688980957
transform 1 0 10856 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_152
timestamp 1688980957
transform 1 0 15088 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_184
timestamp 1688980957
transform 1 0 18032 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_204
timestamp 1688980957
transform 1 0 19872 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_52
timestamp 1688980957
transform 1 0 5888 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_64
timestamp 1688980957
transform 1 0 6992 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_120
timestamp 1688980957
transform 1 0 12144 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_124
timestamp 1688980957
transform 1 0 12512 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_149
timestamp 1688980957
transform 1 0 14812 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_168
timestamp 1688980957
transform 1 0 16560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_173
timestamp 1688980957
transform 1 0 17020 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_179
timestamp 1688980957
transform 1 0 17572 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_183
timestamp 1688980957
transform 1 0 17940 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_29
timestamp 1688980957
transform 1 0 3772 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_48
timestamp 1688980957
transform 1 0 5520 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_63
timestamp 1688980957
transform 1 0 6900 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_82
timestamp 1688980957
transform 1 0 8648 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_94
timestamp 1688980957
transform 1 0 9752 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_128
timestamp 1688980957
transform 1 0 12880 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_150
timestamp 1688980957
transform 1 0 14904 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_191
timestamp 1688980957
transform 1 0 18676 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_199
timestamp 1688980957
transform 1 0 19412 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_24
timestamp 1688980957
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_61
timestamp 1688980957
transform 1 0 6716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_80
timestamp 1688980957
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_100
timestamp 1688980957
transform 1 0 10304 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_112
timestamp 1688980957
transform 1 0 11408 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_124
timestamp 1688980957
transform 1 0 12512 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_136
timestamp 1688980957
transform 1 0 13616 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_171
timestamp 1688980957
transform 1 0 16836 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_188
timestamp 1688980957
transform 1 0 18400 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_52
timestamp 1688980957
transform 1 0 5888 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_81
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_100
timestamp 1688980957
transform 1 0 10304 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_134
timestamp 1688980957
transform 1 0 13432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_142
timestamp 1688980957
transform 1 0 14168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_164
timestamp 1688980957
transform 1 0 16192 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_187
timestamp 1688980957
transform 1 0 18308 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_204
timestamp 1688980957
transform 1 0 19872 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_7
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_26
timestamp 1688980957
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_46
timestamp 1688980957
transform 1 0 5336 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_69
timestamp 1688980957
transform 1 0 7452 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_78
timestamp 1688980957
transform 1 0 8280 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_106
timestamp 1688980957
transform 1 0 10856 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_112
timestamp 1688980957
transform 1 0 11408 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_128
timestamp 1688980957
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_178
timestamp 1688980957
transform 1 0 17480 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_200
timestamp 1688980957
transform 1 0 19504 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_18
timestamp 1688980957
transform 1 0 2760 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_40
timestamp 1688980957
transform 1 0 4784 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_61
timestamp 1688980957
transform 1 0 6716 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_102
timestamp 1688980957
transform 1 0 10488 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_110
timestamp 1688980957
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_128
timestamp 1688980957
transform 1 0 12880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_187
timestamp 1688980957
transform 1 0 18308 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_7
timestamp 1688980957
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_44
timestamp 1688980957
transform 1 0 5152 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_82
timestamp 1688980957
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_119
timestamp 1688980957
transform 1 0 12052 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_158
timestamp 1688980957
transform 1 0 15640 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_185
timestamp 1688980957
transform 1 0 18124 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_200
timestamp 1688980957
transform 1 0 19504 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_204
timestamp 1688980957
transform 1 0 19872 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_9
timestamp 1688980957
transform 1 0 1932 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_52
timestamp 1688980957
transform 1 0 5888 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_97
timestamp 1688980957
transform 1 0 10028 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_109
timestamp 1688980957
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_125
timestamp 1688980957
transform 1 0 12604 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_198
timestamp 1688980957
transform 1 0 19320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_26
timestamp 1688980957
transform 1 0 3496 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_47
timestamp 1688980957
transform 1 0 5428 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_59
timestamp 1688980957
transform 1 0 6532 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 1688980957
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_89
timestamp 1688980957
transform 1 0 9292 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_120
timestamp 1688980957
transform 1 0 12144 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_132
timestamp 1688980957
transform 1 0 13248 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_178
timestamp 1688980957
transform 1 0 17480 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_182
timestamp 1688980957
transform 1 0 17848 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_186
timestamp 1688980957
transform 1 0 18216 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_13
timestamp 1688980957
transform 1 0 2300 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_40
timestamp 1688980957
transform 1 0 4784 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_65
timestamp 1688980957
transform 1 0 7084 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_82
timestamp 1688980957
transform 1 0 8648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_86
timestamp 1688980957
transform 1 0 9016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_108
timestamp 1688980957
transform 1 0 11040 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_172
timestamp 1688980957
transform 1 0 16928 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_180
timestamp 1688980957
transform 1 0 17664 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_194
timestamp 1688980957
transform 1 0 18952 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_19
timestamp 1688980957
transform 1 0 2852 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_40
timestamp 1688980957
transform 1 0 4784 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_60
timestamp 1688980957
transform 1 0 6624 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_78
timestamp 1688980957
transform 1 0 8280 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_93
timestamp 1688980957
transform 1 0 9660 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_127
timestamp 1688980957
transform 1 0 12788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_182
timestamp 1688980957
transform 1 0 17848 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_9
timestamp 1688980957
transform 1 0 1932 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_34
timestamp 1688980957
transform 1 0 4232 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 1688980957
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_80
timestamp 1688980957
transform 1 0 8464 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_86
timestamp 1688980957
transform 1 0 9016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_106
timestamp 1688980957
transform 1 0 10856 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_121
timestamp 1688980957
transform 1 0 12236 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_173
timestamp 1688980957
transform 1 0 17020 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_24
timestamp 1688980957
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_60
timestamp 1688980957
transform 1 0 6624 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_66
timestamp 1688980957
transform 1 0 7176 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_82
timestamp 1688980957
transform 1 0 8648 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_100
timestamp 1688980957
transform 1 0 10304 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_108
timestamp 1688980957
transform 1 0 11040 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_130
timestamp 1688980957
transform 1 0 13064 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_138
timestamp 1688980957
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_162
timestamp 1688980957
transform 1 0 16008 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_174
timestamp 1688980957
transform 1 0 17112 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_180
timestamp 1688980957
transform 1 0 17664 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_201
timestamp 1688980957
transform 1 0 19596 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_24
timestamp 1688980957
transform 1 0 3312 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_44
timestamp 1688980957
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_99
timestamp 1688980957
transform 1 0 10212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_128
timestamp 1688980957
transform 1 0 12880 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_164
timestamp 1688980957
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_189
timestamp 1688980957
transform 1 0 18492 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_199
timestamp 1688980957
transform 1 0 19412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_204
timestamp 1688980957
transform 1 0 19872 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_9
timestamp 1688980957
transform 1 0 1932 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_35
timestamp 1688980957
transform 1 0 4324 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_57
timestamp 1688980957
transform 1 0 6348 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_80
timestamp 1688980957
transform 1 0 8464 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_104
timestamp 1688980957
transform 1 0 10672 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_120
timestamp 1688980957
transform 1 0 12144 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_132
timestamp 1688980957
transform 1 0 13248 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_174
timestamp 1688980957
transform 1 0 17112 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_202
timestamp 1688980957
transform 1 0 19688 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_206
timestamp 1688980957
transform 1 0 20056 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_85
timestamp 1688980957
transform 1 0 8924 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_109
timestamp 1688980957
transform 1 0 11132 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_131
timestamp 1688980957
transform 1 0 13156 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_154
timestamp 1688980957
transform 1 0 15272 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_166
timestamp 1688980957
transform 1 0 16376 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_195
timestamp 1688980957
transform 1 0 19044 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_24
timestamp 1688980957
transform 1 0 3312 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_35
timestamp 1688980957
transform 1 0 4324 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_39
timestamp 1688980957
transform 1 0 4692 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_73
timestamp 1688980957
transform 1 0 7820 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_82
timestamp 1688980957
transform 1 0 8648 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_106
timestamp 1688980957
transform 1 0 10856 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_112
timestamp 1688980957
transform 1 0 11408 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_137
timestamp 1688980957
transform 1 0 13708 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_159
timestamp 1688980957
transform 1 0 15732 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_210
timestamp 1688980957
transform 1 0 20424 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_34
timestamp 1688980957
transform 1 0 4232 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_50
timestamp 1688980957
transform 1 0 5704 0 -1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 1688980957
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_81
timestamp 1688980957
transform 1 0 8556 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_87
timestamp 1688980957
transform 1 0 9108 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_110
timestamp 1688980957
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_134
timestamp 1688980957
transform 1 0 13432 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_142
timestamp 1688980957
transform 1 0 14168 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_158
timestamp 1688980957
transform 1 0 15640 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_162
timestamp 1688980957
transform 1 0 16008 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_166
timestamp 1688980957
transform 1 0 16376 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_186
timestamp 1688980957
transform 1 0 18216 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_194
timestamp 1688980957
transform 1 0 18952 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_26
timestamp 1688980957
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_50
timestamp 1688980957
transform 1 0 5704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_58
timestamp 1688980957
transform 1 0 6440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_80
timestamp 1688980957
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_106
timestamp 1688980957
transform 1 0 10856 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1688980957
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_157
timestamp 1688980957
transform 1 0 15548 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_183
timestamp 1688980957
transform 1 0 17940 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_20
timestamp 1688980957
transform 1 0 2944 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_109
timestamp 1688980957
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_128
timestamp 1688980957
transform 1 0 12880 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_136
timestamp 1688980957
transform 1 0 13616 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_155
timestamp 1688980957
transform 1 0 15364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_160
timestamp 1688980957
transform 1 0 15824 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_35
timestamp 1688980957
transform 1 0 4324 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_47
timestamp 1688980957
transform 1 0 5428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_51
timestamp 1688980957
transform 1 0 5796 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_67
timestamp 1688980957
transform 1 0 7268 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_100
timestamp 1688980957
transform 1 0 10304 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_123
timestamp 1688980957
transform 1 0 12420 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_135
timestamp 1688980957
transform 1 0 13524 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_139
timestamp 1688980957
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_156
timestamp 1688980957
transform 1 0 15456 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_168
timestamp 1688980957
transform 1 0 16560 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_180
timestamp 1688980957
transform 1 0 17664 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_210
timestamp 1688980957
transform 1 0 20424 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_35
timestamp 1688980957
transform 1 0 4324 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_43
timestamp 1688980957
transform 1 0 5060 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_49
timestamp 1688980957
transform 1 0 5612 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_63
timestamp 1688980957
transform 1 0 6900 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_79
timestamp 1688980957
transform 1 0 8372 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_86
timestamp 1688980957
transform 1 0 9016 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_128
timestamp 1688980957
transform 1 0 12880 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_140
timestamp 1688980957
transform 1 0 13984 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_144
timestamp 1688980957
transform 1 0 14352 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_148
timestamp 1688980957
transform 1 0 14720 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_159
timestamp 1688980957
transform 1 0 15732 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_184
timestamp 1688980957
transform 1 0 18032 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_190
timestamp 1688980957
transform 1 0 18584 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_9
timestamp 1688980957
transform 1 0 1932 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_47
timestamp 1688980957
transform 1 0 5428 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_59
timestamp 1688980957
transform 1 0 6532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_71
timestamp 1688980957
transform 1 0 7636 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_101
timestamp 1688980957
transform 1 0 10396 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_160
timestamp 1688980957
transform 1 0 15824 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_169
timestamp 1688980957
transform 1 0 16652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_173
timestamp 1688980957
transform 1 0 17020 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_192
timestamp 1688980957
transform 1 0 18768 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_15
timestamp 1688980957
transform 1 0 2484 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_53
timestamp 1688980957
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_82
timestamp 1688980957
transform 1 0 8648 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_94
timestamp 1688980957
transform 1 0 9752 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_106
timestamp 1688980957
transform 1 0 10856 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_179
timestamp 1688980957
transform 1 0 17572 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_198
timestamp 1688980957
transform 1 0 19320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_202
timestamp 1688980957
transform 1 0 19688 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_70_24
timestamp 1688980957
transform 1 0 3312 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_44
timestamp 1688980957
transform 1 0 5152 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_56
timestamp 1688980957
transform 1 0 6256 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_72
timestamp 1688980957
transform 1 0 7728 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1688980957
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1688980957
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1688980957
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_157
timestamp 1688980957
transform 1 0 15548 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_163
timestamp 1688980957
transform 1 0 16100 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_204
timestamp 1688980957
transform 1 0 19872 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_14
timestamp 1688980957
transform 1 0 2392 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_35
timestamp 1688980957
transform 1 0 4324 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_52
timestamp 1688980957
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_86
timestamp 1688980957
transform 1 0 9016 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_98
timestamp 1688980957
transform 1 0 10120 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_110
timestamp 1688980957
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_145
timestamp 1688980957
transform 1 0 14444 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_186
timestamp 1688980957
transform 1 0 18216 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_191
timestamp 1688980957
transform 1 0 18676 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_196
timestamp 1688980957
transform 1 0 19136 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_20
timestamp 1688980957
transform 1 0 2944 0 1 40256
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_149
timestamp 1688980957
transform 1 0 14812 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_169
timestamp 1688980957
transform 1 0 16652 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_174
timestamp 1688980957
transform 1 0 17112 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_188
timestamp 1688980957
transform 1 0 18400 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_14
timestamp 1688980957
transform 1 0 2392 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_22
timestamp 1688980957
transform 1 0 3128 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_37
timestamp 1688980957
transform 1 0 4508 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_46
timestamp 1688980957
transform 1 0 5336 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_54
timestamp 1688980957
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_65
timestamp 1688980957
transform 1 0 7084 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_75
timestamp 1688980957
transform 1 0 8004 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_87
timestamp 1688980957
transform 1 0 9108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_99
timestamp 1688980957
transform 1 0 10212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_156
timestamp 1688980957
transform 1 0 15456 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_166
timestamp 1688980957
transform 1 0 16376 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_172
timestamp 1688980957
transform 1 0 16928 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_182
timestamp 1688980957
transform 1 0 17848 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_196
timestamp 1688980957
transform 1 0 19136 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_201
timestamp 1688980957
transform 1 0 19596 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_11
timestamp 1688980957
transform 1 0 2116 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_55
timestamp 1688980957
transform 1 0 6164 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_59
timestamp 1688980957
transform 1 0 6532 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_70
timestamp 1688980957
transform 1 0 7544 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_88
timestamp 1688980957
transform 1 0 9200 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_100
timestamp 1688980957
transform 1 0 10304 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_112
timestamp 1688980957
transform 1 0 11408 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_124
timestamp 1688980957
transform 1 0 12512 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_130
timestamp 1688980957
transform 1 0 13064 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_145
timestamp 1688980957
transform 1 0 14444 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_167
timestamp 1688980957
transform 1 0 16468 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_183
timestamp 1688980957
transform 1 0 17940 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_204
timestamp 1688980957
transform 1 0 19872 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_18
timestamp 1688980957
transform 1 0 2760 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_45
timestamp 1688980957
transform 1 0 5244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_75_94
timestamp 1688980957
transform 1 0 9752 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_100
timestamp 1688980957
transform 1 0 10304 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_107
timestamp 1688980957
transform 1 0 10948 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_119
timestamp 1688980957
transform 1 0 12052 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_172
timestamp 1688980957
transform 1 0 16928 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_200
timestamp 1688980957
transform 1 0 19504 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_210
timestamp 1688980957
transform 1 0 20424 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1688980957
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_120
timestamp 1688980957
transform 1 0 12144 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_138
timestamp 1688980957
transform 1 0 13800 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 1688980957
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_26
timestamp 1688980957
transform 1 0 3496 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_29
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_66
timestamp 1688980957
transform 1 0 7176 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_85
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_119
timestamp 1688980957
transform 1 0 12052 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_157
timestamp 1688980957
transform 1 0 15548 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_195
timestamp 1688980957
transform 1 0 19044 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2300 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 3312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 1656 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 3220 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 2944 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 2668 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1688980957
transform 1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 1688980957
transform 1 0 4508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1688980957
transform 1 0 5152 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1688980957
transform 1 0 2760 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1688980957
transform 1 0 3220 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 4508 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input25
timestamp 1688980957
transform 1 0 4048 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 3036 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1688980957
transform 1 0 2300 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1688980957
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 3404 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 2944 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 3220 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 3496 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 3220 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 2852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input42
timestamp 1688980957
transform 1 0 2300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 2576 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 3128 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 3128 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input51
timestamp 1688980957
transform 1 0 3864 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input52
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input53
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input54 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1688980957
transform 1 0 4140 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input56
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input57
timestamp 1688980957
transform 1 0 1932 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input58
timestamp 1688980957
transform 1 0 3036 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input59
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input60
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input61
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input62
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input63
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input64
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input65
timestamp 1688980957
transform 1 0 1932 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input66
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input67
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input68
timestamp 1688980957
transform 1 0 3036 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input69
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input70
timestamp 1688980957
transform 1 0 1932 0 1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input71
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input72
timestamp 1688980957
transform 1 0 2484 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input73
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input74
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input75
timestamp 1688980957
transform 1 0 3680 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input76
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1688980957
transform 1 0 2760 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1688980957
transform 1 0 1932 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input80
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1688980957
transform 1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input85
timestamp 1688980957
transform 1 0 12144 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input86
timestamp 1688980957
transform 1 0 11868 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1688980957
transform 1 0 12328 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1688980957
transform 1 0 11592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1688980957
transform 1 0 12052 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input90
timestamp 1688980957
transform 1 0 11132 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1688980957
transform 1 0 12420 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input92
timestamp 1688980957
transform 1 0 15456 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input93 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input94
timestamp 1688980957
transform 1 0 18032 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input95
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input96
timestamp 1688980957
transform 1 0 18032 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input97
timestamp 1688980957
transform 1 0 18492 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input98
timestamp 1688980957
transform 1 0 14352 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input99
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input100
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input102
timestamp 1688980957
transform 1 0 2024 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input103
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input104
timestamp 1688980957
transform 1 0 1472 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input105
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input106
timestamp 1688980957
transform 1 0 4784 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input107
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1688980957
transform 1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input111
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input112
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input113
timestamp 1688980957
transform 1 0 3220 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input115
timestamp 1688980957
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1688980957
transform 1 0 2944 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input117
timestamp 1688980957
transform 1 0 3956 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1688980957
transform 1 0 4600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1688980957
transform 1 0 4416 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1688980957
transform 1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1688980957
transform 1 0 5612 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1688980957
transform 1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1688980957
transform 1 0 8096 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1688980957
transform 1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1688980957
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input128
timestamp 1688980957
transform 1 0 6808 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 1688980957
transform 1 0 5520 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1688980957
transform 1 0 4416 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1688980957
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1688980957
transform 1 0 6716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1688980957
transform 1 0 6808 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1688980957
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input137
timestamp 1688980957
transform 1 0 11776 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1688980957
transform 1 0 10120 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input139
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1688980957
transform 1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1688980957
transform 1 0 12328 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input143
timestamp 1688980957
transform 1 0 14720 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input144
timestamp 1688980957
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input145
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1688980957
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input147
timestamp 1688980957
transform 1 0 13248 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1688980957
transform 1 0 13156 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1688980957
transform 1 0 13432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1688980957
transform 1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1688980957
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input152
timestamp 1688980957
transform 1 0 11776 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1688980957
transform 1 0 8464 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input154
timestamp 1688980957
transform 1 0 9476 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input155
timestamp 1688980957
transform 1 0 9108 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1688980957
transform 1 0 9476 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input157
timestamp 1688980957
transform 1 0 10672 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input158
timestamp 1688980957
transform 1 0 10028 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1688980957
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1688980957
transform 1 0 10396 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1688980957
transform 1 0 10120 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1688980957
transform 1 0 9844 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input163
timestamp 1688980957
transform 1 0 10948 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1688980957
transform 1 0 11132 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input165
timestamp 1688980957
transform 1 0 10672 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1688980957
transform 1 0 11316 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input167
timestamp 1688980957
transform 1 0 11684 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1688980957
transform 1 0 11592 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input169
timestamp 1688980957
transform 1 0 11132 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input170
timestamp 1688980957
transform 1 0 12236 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input171
timestamp 1688980957
transform 1 0 12604 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input172
timestamp 1688980957
transform 1 0 12880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input173
timestamp 1688980957
transform 1 0 12972 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1688980957
transform 1 0 14628 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1688980957
transform 1 0 14904 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1688980957
transform 1 0 15180 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1688980957
transform 1 0 18676 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1688980957
transform 1 0 12420 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input179
timestamp 1688980957
transform 1 0 14352 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1688980957
transform 1 0 13340 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input181
timestamp 1688980957
transform 1 0 13156 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input182
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1688980957
transform 1 0 14720 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1688980957
transform 1 0 14996 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1688980957
transform 1 0 15272 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1688980957
transform 1 0 19780 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1688980957
transform 1 0 16192 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf
timestamp 1688980957
transform 1 0 14628 0 -1 40256
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._0_
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._1_
timestamp 1688980957
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._2_
timestamp 1688980957
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._3_
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16376 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 18216 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 18400 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._2_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17848 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18216 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16100 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18124 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 19320 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 19504 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18768 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19780 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20240 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 14444 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 15088 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15364 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18400 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 18584 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 16744 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 15088 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18768 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20148 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 18584 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18216 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19044 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 16928 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 17664 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 18308 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17296 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 16744 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 18492 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 17848 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18216 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17480 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18768 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 19504 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 19780 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 19688 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 18400 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 18032 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 18584 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 16376 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 15640 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 15088 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17664 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18216 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18768 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 17848 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16100 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18492 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 17388 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 17020 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16100 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17664 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 16744 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15640 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 19504 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 19688 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19872 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18676 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 18400 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 17388 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 18216 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19320 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19688 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18768 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 18676 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 19412 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18032 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19136 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 19688 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18768 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 18032 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 17572 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 17204 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17848 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 15088 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 18400 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 16744 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 17940 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 17296 0 1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16008 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17296 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 14444 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 15456 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 13708 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15548 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 19412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20240 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18124 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 17204 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18492 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 18124 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17572 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 18584 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 17480 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18676 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16928 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17848 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 19136 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 18400 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 19688 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20332 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19688 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18584 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19320 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 17480 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18768 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 18124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16836 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18492 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 15640 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 16468 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 20332 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16652 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 17940 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 16836 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19412 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17296 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19136 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 17112 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 12328 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 13340 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 12880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 12512 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 11684 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 11500 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 10856 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 19412 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 10580 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 14444 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 15364 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 18492 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 15456 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 15456 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15180 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 14996 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 15456 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 10028 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 12052 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 18216 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 13432 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 14720 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 16836 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 18676 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 11592 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 14444 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 10948 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 17756 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 12420 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 13524 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 13064 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 13156 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit1
timestamp 1688980957
transform 1 0 7268 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit2
timestamp 1688980957
transform 1 0 1932 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit3
timestamp 1688980957
transform 1 0 2668 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit4
timestamp 1688980957
transform 1 0 1840 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit5
timestamp 1688980957
transform 1 0 3404 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit6
timestamp 1688980957
transform 1 0 8648 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit7
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit8
timestamp 1688980957
transform 1 0 7084 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit9
timestamp 1688980957
transform 1 0 8648 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit10
timestamp 1688980957
transform 1 0 4416 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit11
timestamp 1688980957
transform 1 0 4968 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit12
timestamp 1688980957
transform 1 0 6716 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit13
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit14
timestamp 1688980957
transform 1 0 9016 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit15
timestamp 1688980957
transform 1 0 9476 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit16
timestamp 1688980957
transform 1 0 9752 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit17
timestamp 1688980957
transform 1 0 9476 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit18
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit19
timestamp 1688980957
transform 1 0 7452 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit20
timestamp 1688980957
transform 1 0 5336 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit21
timestamp 1688980957
transform 1 0 6716 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit22
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit23
timestamp 1688980957
transform 1 0 10488 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit24
timestamp 1688980957
transform 1 0 8924 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit25
timestamp 1688980957
transform 1 0 9200 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit26
timestamp 1688980957
transform 1 0 1656 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit27
timestamp 1688980957
transform 1 0 2300 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit28
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit30
timestamp 1688980957
transform 1 0 11960 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit31
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit0
timestamp 1688980957
transform 1 0 14720 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit1
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit2
timestamp 1688980957
transform 1 0 7452 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit3
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit4
timestamp 1688980957
transform 1 0 4600 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit5
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit6
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit7
timestamp 1688980957
transform 1 0 14168 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit8
timestamp 1688980957
transform 1 0 8648 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit9
timestamp 1688980957
transform 1 0 10028 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit10
timestamp 1688980957
transform 1 0 2852 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit11
timestamp 1688980957
transform 1 0 4324 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit12
timestamp 1688980957
transform 1 0 3128 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit13
timestamp 1688980957
transform 1 0 5520 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit14
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit15
timestamp 1688980957
transform 1 0 12144 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit16
timestamp 1688980957
transform 1 0 9016 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit17
timestamp 1688980957
transform 1 0 7452 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit18
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit19
timestamp 1688980957
transform 1 0 2300 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit20
timestamp 1688980957
transform 1 0 1932 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit21
timestamp 1688980957
transform 1 0 2300 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit22
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit23
timestamp 1688980957
transform 1 0 12328 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit24
timestamp 1688980957
transform 1 0 7820 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit25
timestamp 1688980957
transform 1 0 10396 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit26
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit27
timestamp 1688980957
transform 1 0 4508 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit28
timestamp 1688980957
transform 1 0 2300 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit29
timestamp 1688980957
transform 1 0 2024 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit30
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit31
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit0
timestamp 1688980957
transform 1 0 12604 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit1
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit2
timestamp 1688980957
transform 1 0 6348 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit3
timestamp 1688980957
transform 1 0 7636 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit4
timestamp 1688980957
transform 1 0 2852 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit5
timestamp 1688980957
transform 1 0 3128 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit6
timestamp 1688980957
transform 1 0 12420 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit7
timestamp 1688980957
transform 1 0 14904 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit8
timestamp 1688980957
transform 1 0 14352 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit9
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit10
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit11
timestamp 1688980957
transform 1 0 1932 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit12
timestamp 1688980957
transform 1 0 2944 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit13
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit14
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit15
timestamp 1688980957
transform 1 0 15456 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit16
timestamp 1688980957
transform 1 0 11684 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit17
timestamp 1688980957
transform 1 0 12328 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit18
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit19
timestamp 1688980957
transform 1 0 1564 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit20
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit21
timestamp 1688980957
transform 1 0 7452 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit22
timestamp 1688980957
transform 1 0 11224 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit23
timestamp 1688980957
transform 1 0 11776 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit24
timestamp 1688980957
transform 1 0 10580 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit25
timestamp 1688980957
transform 1 0 10028 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit26
timestamp 1688980957
transform 1 0 8372 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit27
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit28
timestamp 1688980957
transform 1 0 6808 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit29
timestamp 1688980957
transform 1 0 7176 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit30
timestamp 1688980957
transform 1 0 12604 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit31
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit0
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit1
timestamp 1688980957
transform 1 0 13984 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit2
timestamp 1688980957
transform 1 0 2300 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit3
timestamp 1688980957
transform 1 0 2944 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit4
timestamp 1688980957
transform 1 0 4692 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit5
timestamp 1688980957
transform 1 0 4876 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit6
timestamp 1688980957
transform 1 0 11960 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit7
timestamp 1688980957
transform 1 0 12512 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit8
timestamp 1688980957
transform 1 0 13984 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit9
timestamp 1688980957
transform 1 0 16100 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit10
timestamp 1688980957
transform 1 0 3496 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit11
timestamp 1688980957
transform 1 0 2852 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit12
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit13
timestamp 1688980957
transform 1 0 6440 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit14
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit15
timestamp 1688980957
transform 1 0 16008 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit16
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit17
timestamp 1688980957
transform 1 0 15456 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit18
timestamp 1688980957
transform 1 0 5888 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit19
timestamp 1688980957
transform 1 0 6992 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit20
timestamp 1688980957
transform 1 0 3956 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit21
timestamp 1688980957
transform 1 0 4508 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit22
timestamp 1688980957
transform 1 0 13156 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit23
timestamp 1688980957
transform 1 0 14536 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit24
timestamp 1688980957
transform 1 0 14168 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit25
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit26
timestamp 1688980957
transform 1 0 4416 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit27
timestamp 1688980957
transform 1 0 4876 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit28
timestamp 1688980957
transform 1 0 3496 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit29
timestamp 1688980957
transform 1 0 4508 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit30
timestamp 1688980957
transform 1 0 14260 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit31
timestamp 1688980957
transform 1 0 15456 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit0
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit1
timestamp 1688980957
transform 1 0 14904 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit2
timestamp 1688980957
transform 1 0 2300 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit3
timestamp 1688980957
transform 1 0 2024 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit4
timestamp 1688980957
transform 1 0 4876 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit5
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit6
timestamp 1688980957
transform 1 0 7452 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit7
timestamp 1688980957
transform 1 0 9752 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit8
timestamp 1688980957
transform 1 0 15088 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit9
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit10
timestamp 1688980957
transform 1 0 2116 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit11
timestamp 1688980957
transform 1 0 3496 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit12
timestamp 1688980957
transform 1 0 5704 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit13
timestamp 1688980957
transform 1 0 4600 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit14
timestamp 1688980957
transform 1 0 7268 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit15
timestamp 1688980957
transform 1 0 9936 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit16
timestamp 1688980957
transform 1 0 15456 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit17
timestamp 1688980957
transform 1 0 16008 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit18
timestamp 1688980957
transform 1 0 2116 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit19
timestamp 1688980957
transform 1 0 2300 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit20
timestamp 1688980957
transform 1 0 4324 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit21
timestamp 1688980957
transform 1 0 6072 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit22
timestamp 1688980957
transform 1 0 6072 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit23
timestamp 1688980957
transform 1 0 8648 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit24
timestamp 1688980957
transform 1 0 11684 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit25
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit26
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit27
timestamp 1688980957
transform 1 0 4048 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit28
timestamp 1688980957
transform 1 0 4048 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit29
timestamp 1688980957
transform 1 0 5704 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit30
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit31
timestamp 1688980957
transform 1 0 12328 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit0
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit1
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit2
timestamp 1688980957
transform 1 0 2024 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit3
timestamp 1688980957
transform 1 0 2300 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit4
timestamp 1688980957
transform 1 0 1840 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit5
timestamp 1688980957
transform 1 0 2668 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit6
timestamp 1688980957
transform 1 0 9752 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit7
timestamp 1688980957
transform 1 0 10304 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit8
timestamp 1688980957
transform 1 0 13616 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit9
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit10
timestamp 1688980957
transform 1 0 1840 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit11
timestamp 1688980957
transform 1 0 2300 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit12
timestamp 1688980957
transform 1 0 4692 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit13
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit14
timestamp 1688980957
transform 1 0 7452 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit15
timestamp 1688980957
transform 1 0 9844 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit16
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit17
timestamp 1688980957
transform 1 0 16008 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit18
timestamp 1688980957
transform 1 0 1656 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit19
timestamp 1688980957
transform 1 0 2300 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit20
timestamp 1688980957
transform 1 0 1564 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit21
timestamp 1688980957
transform 1 0 2300 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit22
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit23
timestamp 1688980957
transform 1 0 10488 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit24
timestamp 1688980957
transform 1 0 16100 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit25
timestamp 1688980957
transform 1 0 15456 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit26
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit27
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit28
timestamp 1688980957
transform 1 0 4876 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit29
timestamp 1688980957
transform 1 0 6072 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit30
timestamp 1688980957
transform 1 0 8096 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit31
timestamp 1688980957
transform 1 0 9476 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit0
timestamp 1688980957
transform 1 0 1472 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit1
timestamp 1688980957
transform 1 0 1748 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit2
timestamp 1688980957
transform 1 0 10028 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit3
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit4
timestamp 1688980957
transform 1 0 13248 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit5
timestamp 1688980957
transform 1 0 14628 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit6
timestamp 1688980957
transform 1 0 15456 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit7
timestamp 1688980957
transform 1 0 4876 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit8
timestamp 1688980957
transform 1 0 7176 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit9
timestamp 1688980957
transform 1 0 8004 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit10
timestamp 1688980957
transform 1 0 4876 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit11
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit12
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit13
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit14
timestamp 1688980957
transform 1 0 14352 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit15
timestamp 1688980957
transform 1 0 16008 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit16
timestamp 1688980957
transform 1 0 7452 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit17
timestamp 1688980957
transform 1 0 7452 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit18
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit19
timestamp 1688980957
transform 1 0 4692 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit20
timestamp 1688980957
transform 1 0 4508 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit21
timestamp 1688980957
transform 1 0 4600 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit22
timestamp 1688980957
transform 1 0 11684 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit23
timestamp 1688980957
transform 1 0 12236 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit24
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit25
timestamp 1688980957
transform 1 0 12052 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit26
timestamp 1688980957
transform 1 0 4600 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit27
timestamp 1688980957
transform 1 0 4600 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit28
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit29
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit30
timestamp 1688980957
transform 1 0 7452 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit31
timestamp 1688980957
transform 1 0 8096 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit0
timestamp 1688980957
transform 1 0 11224 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit1
timestamp 1688980957
transform 1 0 11776 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit2
timestamp 1688980957
transform 1 0 11684 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit3
timestamp 1688980957
transform 1 0 5060 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit4
timestamp 1688980957
transform 1 0 7084 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit5
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit6
timestamp 1688980957
transform 1 0 7268 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit7
timestamp 1688980957
transform 1 0 4876 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit8
timestamp 1688980957
transform 1 0 6900 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit9
timestamp 1688980957
transform 1 0 12328 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit10
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit11
timestamp 1688980957
transform 1 0 13892 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit12
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit13
timestamp 1688980957
transform 1 0 9568 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit14
timestamp 1688980957
transform 1 0 6440 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit15
timestamp 1688980957
transform 1 0 7268 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit16
timestamp 1688980957
transform 1 0 4876 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit17
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit18
timestamp 1688980957
transform 1 0 9752 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit19
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit20
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit21
timestamp 1688980957
transform 1 0 9108 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit22
timestamp 1688980957
transform 1 0 6900 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit23
timestamp 1688980957
transform 1 0 7268 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit24
timestamp 1688980957
transform 1 0 7176 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit25
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit26
timestamp 1688980957
transform 1 0 9384 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit27
timestamp 1688980957
transform 1 0 10764 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit28
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit29
timestamp 1688980957
transform 1 0 10028 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit30
timestamp 1688980957
transform 1 0 7452 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit31
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit0
timestamp 1688980957
transform 1 0 17296 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit1
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit2
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit3
timestamp 1688980957
transform 1 0 16836 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit4
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit5
timestamp 1688980957
transform 1 0 18768 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit6
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit7
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit8
timestamp 1688980957
transform 1 0 8188 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit9
timestamp 1688980957
transform 1 0 9568 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit10
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit11
timestamp 1688980957
transform 1 0 1472 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit12
timestamp 1688980957
transform 1 0 1840 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit13
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit14
timestamp 1688980957
transform 1 0 10764 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit15
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit16
timestamp 1688980957
transform 1 0 8924 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit17
timestamp 1688980957
transform 1 0 9016 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit18
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit19
timestamp 1688980957
transform 1 0 1472 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit20
timestamp 1688980957
transform 1 0 1472 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit21
timestamp 1688980957
transform 1 0 1932 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit22
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit23
timestamp 1688980957
transform 1 0 9476 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit24
timestamp 1688980957
transform 1 0 11040 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit25
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit26
timestamp 1688980957
transform 1 0 1472 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit27
timestamp 1688980957
transform 1 0 2024 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit28
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit29
timestamp 1688980957
transform 1 0 1564 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit30
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit31
timestamp 1688980957
transform 1 0 11500 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit0
timestamp 1688980957
transform 1 0 14076 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit1
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit2
timestamp 1688980957
transform 1 0 14260 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit3
timestamp 1688980957
transform 1 0 17664 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit4
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit5
timestamp 1688980957
transform 1 0 16376 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit6
timestamp 1688980957
transform 1 0 17112 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit7
timestamp 1688980957
transform 1 0 13064 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit8
timestamp 1688980957
transform 1 0 16836 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit9
timestamp 1688980957
transform 1 0 16100 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit10
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit11
timestamp 1688980957
transform 1 0 18492 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit12
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit13
timestamp 1688980957
transform 1 0 17756 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit14
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit15
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit16
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit17
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit18
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit19
timestamp 1688980957
transform 1 0 16744 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit20
timestamp 1688980957
transform 1 0 16928 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit21
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit22
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit23
timestamp 1688980957
transform 1 0 17480 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit24
timestamp 1688980957
transform 1 0 16836 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit25
timestamp 1688980957
transform 1 0 18676 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit26
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit27
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit28
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit29
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit30
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit31
timestamp 1688980957
transform 1 0 16928 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit24
timestamp 1688980957
transform 1 0 17112 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit25
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit26
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit27
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit28
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit29
timestamp 1688980957
transform 1 0 16836 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit30
timestamp 1688980957
transform 1 0 18032 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit31
timestamp 1688980957
transform 1 0 17204 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform 1 0 4232 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform 1 0 4692 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform 1 0 4600 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._36_
timestamp 1688980957
transform 1 0 4784 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._37_
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._38_
timestamp 1688980957
transform 1 0 4968 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._39_
timestamp 1688980957
transform 1 0 5336 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._40_
timestamp 1688980957
transform 1 0 10120 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._41_
timestamp 1688980957
transform 1 0 9108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._42_
timestamp 1688980957
transform 1 0 9476 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._43_
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._44_
timestamp 1688980957
transform 1 0 10856 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._45_
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._46_
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._47_
timestamp 1688980957
transform 1 0 11868 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0_395 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12972 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1_396
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2_397
timestamp 1688980957
transform 1 0 8648 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2
timestamp 1688980957
transform 1 0 7636 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3_398
timestamp 1688980957
transform 1 0 13432 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3
timestamp 1688980957
transform 1 0 11500 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0_399
timestamp 1688980957
transform 1 0 11776 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0
timestamp 1688980957
transform 1 0 10856 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1_400
timestamp 1688980957
transform 1 0 9016 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2_401
timestamp 1688980957
transform 1 0 8188 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2
timestamp 1688980957
transform 1 0 6992 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3_402
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3
timestamp 1688980957
transform 1 0 12972 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0_403
timestamp 1688980957
transform 1 0 15824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0
timestamp 1688980957
transform 1 0 14904 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1_404
timestamp 1688980957
transform 1 0 8740 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1
timestamp 1688980957
transform 1 0 7820 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2_405
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3_409
timestamp 1688980957
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3
timestamp 1688980957
transform 1 0 13892 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I0
timestamp 1688980957
transform 1 0 13708 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I1
timestamp 1688980957
transform 1 0 6532 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I2
timestamp 1688980957
transform 1 0 4324 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I3
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I0
timestamp 1688980957
transform 1 0 14444 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I1
timestamp 1688980957
transform 1 0 4968 0 1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I2
timestamp 1688980957
transform 1 0 4324 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I3
timestamp 1688980957
transform 1 0 14260 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I0
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I1
timestamp 1688980957
transform 1 0 6716 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I2
timestamp 1688980957
transform 1 0 3864 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I3
timestamp 1688980957
transform 1 0 12972 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I0
timestamp 1688980957
transform 1 0 14444 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I1
timestamp 1688980957
transform 1 0 2024 0 -1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I2
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I3
timestamp 1688980957
transform 1 0 13984 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0
timestamp 1688980957
transform 1 0 9568 0 -1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0_406
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1_407
timestamp 1688980957
transform 1 0 4048 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1
timestamp 1688980957
transform 1 0 2668 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2
timestamp 1688980957
transform 1 0 3496 0 -1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2_408
timestamp 1688980957
transform 1 0 4232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3_394
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3
timestamp 1688980957
transform 1 0 11960 0 -1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG0
timestamp 1688980957
transform 1 0 8464 0 -1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG1
timestamp 1688980957
transform 1 0 4968 0 1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG2
timestamp 1688980957
transform 1 0 8280 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG3
timestamp 1688980957
transform 1 0 9108 0 -1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG4
timestamp 1688980957
transform 1 0 9200 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG5
timestamp 1688980957
transform 1 0 7728 0 -1 8704
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG6
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG7
timestamp 1688980957
transform 1 0 9752 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG0
timestamp 1688980957
transform 1 0 9844 0 1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG1
timestamp 1688980957
transform 1 0 4048 0 1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG2
timestamp 1688980957
transform 1 0 3864 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG3
timestamp 1688980957
transform 1 0 11868 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG4
timestamp 1688980957
transform 1 0 9752 0 1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG5
timestamp 1688980957
transform 1 0 3496 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG6
timestamp 1688980957
transform 1 0 3312 0 -1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG7
timestamp 1688980957
transform 1 0 11868 0 1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG8
timestamp 1688980957
transform 1 0 9936 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG9
timestamp 1688980957
transform 1 0 4324 0 -1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG10
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG11
timestamp 1688980957
transform 1 0 11684 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG12
timestamp 1688980957
transform 1 0 9200 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG13
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG14
timestamp 1688980957
transform 1 0 3312 0 -1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG15
timestamp 1688980957
transform 1 0 11592 0 1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG0
timestamp 1688980957
transform 1 0 9292 0 1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG1
timestamp 1688980957
transform 1 0 1564 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG2
timestamp 1688980957
transform 1 0 2024 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG3
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG0
timestamp 1688980957
transform 1 0 9200 0 1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG1
timestamp 1688980957
transform 1 0 1564 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG2
timestamp 1688980957
transform 1 0 1932 0 -1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG3
timestamp 1688980957
transform 1 0 9108 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG4
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG5
timestamp 1688980957
transform 1 0 1840 0 -1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG6
timestamp 1688980957
transform 1 0 1656 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG7
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG0
timestamp 1688980957
transform 1 0 9292 0 -1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG1
timestamp 1688980957
transform 1 0 6900 0 -1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG2
timestamp 1688980957
transform 1 0 5520 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG3
timestamp 1688980957
transform 1 0 11132 0 1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG0
timestamp 1688980957
transform 1 0 9200 0 -1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG1
timestamp 1688980957
transform 1 0 6808 0 1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG2
timestamp 1688980957
transform 1 0 8004 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG3
timestamp 1688980957
transform 1 0 10396 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG4
timestamp 1688980957
transform 1 0 10120 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG5
timestamp 1688980957
transform 1 0 7820 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG6
timestamp 1688980957
transform 1 0 1656 0 -1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG7
timestamp 1688980957
transform 1 0 10488 0 1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG0
timestamp 1688980957
transform 1 0 8740 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG1
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG2
timestamp 1688980957
transform 1 0 4324 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG3
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG0
timestamp 1688980957
transform 1 0 11776 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG1
timestamp 1688980957
transform 1 0 4324 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG2
timestamp 1688980957
transform 1 0 6256 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG3
timestamp 1688980957
transform 1 0 9476 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG4
timestamp 1688980957
transform 1 0 13800 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG5
timestamp 1688980957
transform 1 0 2576 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG6
timestamp 1688980957
transform 1 0 2300 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG7
timestamp 1688980957
transform 1 0 10120 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb0
timestamp 1688980957
transform 1 0 12052 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb1
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb2
timestamp 1688980957
transform 1 0 6256 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb3
timestamp 1688980957
transform 1 0 9568 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb4
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb5
timestamp 1688980957
transform 1 0 2392 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb6
timestamp 1688980957
transform 1 0 2208 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb7
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG0
timestamp 1688980957
transform 1 0 11868 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG1
timestamp 1688980957
transform 1 0 3956 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG2
timestamp 1688980957
transform 1 0 5428 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG3
timestamp 1688980957
transform 1 0 12052 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG4
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG5
timestamp 1688980957
transform 1 0 4600 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG6
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG7
timestamp 1688980957
transform 1 0 13800 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG8
timestamp 1688980957
transform 1 0 14076 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG9
timestamp 1688980957
transform 1 0 4232 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG10
timestamp 1688980957
transform 1 0 6164 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG11
timestamp 1688980957
transform 1 0 14168 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG0
timestamp 1688980957
transform 1 0 14168 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG1
timestamp 1688980957
transform 1 0 2300 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG2
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG3
timestamp 1688980957
transform 1 0 9384 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG4
timestamp 1688980957
transform 1 0 12972 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG5
timestamp 1688980957
transform 1 0 3404 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG6
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG7
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG8
timestamp 1688980957
transform 1 0 14260 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG9
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG10
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG11
timestamp 1688980957
transform 1 0 9476 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG12
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG13
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG14
timestamp 1688980957
transform 1 0 6440 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG15
timestamp 1688980957
transform 1 0 9292 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 12328 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 12052 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 13064 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 13156 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 13432 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 10396 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 8372 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 9936 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6532 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6624 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 8004 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 8464 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 8280 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6808 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7728 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 5336 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5520 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 15732 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 13616 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 13800 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15456 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 12880 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 16008 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16008 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 13984 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 9200 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 9384 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6440 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 6900 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 7176 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 7636 0 1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6624 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7912 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5612 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 16284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 16008 0 1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16008 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16192 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 14076 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 4968 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 5244 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 5520 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 6716 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 6992 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 7268 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 7176 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 7728 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 9476 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 8648 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 6440 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 5888 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  N4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 6808 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 6440 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 6440 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 6808 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 7360 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 7176 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 7544 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 7912 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 8280 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output189
timestamp 1688980957
transform 1 0 18584 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output190
timestamp 1688980957
transform 1 0 18216 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output191
timestamp 1688980957
transform 1 0 20056 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 20056 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output193
timestamp 1688980957
transform 1 0 20056 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output194
timestamp 1688980957
transform 1 0 20056 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1688980957
transform 1 0 19688 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output196
timestamp 1688980957
transform 1 0 20056 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output197
timestamp 1688980957
transform 1 0 19136 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output198
timestamp 1688980957
transform 1 0 20056 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output199
timestamp 1688980957
transform 1 0 20056 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output200
timestamp 1688980957
transform 1 0 20056 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output201
timestamp 1688980957
transform 1 0 18952 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output202
timestamp 1688980957
transform 1 0 19504 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output203
timestamp 1688980957
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output204
timestamp 1688980957
transform 1 0 20056 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 19872 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output206
timestamp 1688980957
transform 1 0 20056 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output207
timestamp 1688980957
transform 1 0 19504 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output208
timestamp 1688980957
transform 1 0 19688 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output209
timestamp 1688980957
transform 1 0 20056 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output210
timestamp 1688980957
transform 1 0 20056 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output211
timestamp 1688980957
transform 1 0 20056 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output212
timestamp 1688980957
transform 1 0 20056 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output213
timestamp 1688980957
transform 1 0 19872 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output214
timestamp 1688980957
transform 1 0 19320 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1688980957
transform 1 0 19688 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output216
timestamp 1688980957
transform 1 0 20056 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output217
timestamp 1688980957
transform 1 0 20056 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output218
timestamp 1688980957
transform 1 0 19504 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output219
timestamp 1688980957
transform 1 0 19688 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output220
timestamp 1688980957
transform 1 0 20056 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output221
timestamp 1688980957
transform 1 0 20056 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output222
timestamp 1688980957
transform 1 0 20056 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1688980957
transform 1 0 19688 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output224
timestamp 1688980957
transform 1 0 20056 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1688980957
transform 1 0 20240 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output226
timestamp 1688980957
transform 1 0 20056 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output227
timestamp 1688980957
transform 1 0 19320 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output228
timestamp 1688980957
transform 1 0 19872 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output229
timestamp 1688980957
transform 1 0 20056 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output230
timestamp 1688980957
transform 1 0 19320 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output231
timestamp 1688980957
transform 1 0 19872 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output232
timestamp 1688980957
transform 1 0 19504 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output233
timestamp 1688980957
transform 1 0 20056 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output234
timestamp 1688980957
transform 1 0 20056 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output235
timestamp 1688980957
transform 1 0 20056 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output236
timestamp 1688980957
transform 1 0 20056 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output237
timestamp 1688980957
transform 1 0 20056 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output238
timestamp 1688980957
transform 1 0 20056 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output239
timestamp 1688980957
transform 1 0 20056 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output240
timestamp 1688980957
transform 1 0 19320 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output241
timestamp 1688980957
transform 1 0 18952 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output242
timestamp 1688980957
transform 1 0 20056 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output243
timestamp 1688980957
transform 1 0 20056 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output244
timestamp 1688980957
transform 1 0 19504 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output245
timestamp 1688980957
transform 1 0 19872 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1688980957
transform 1 0 20240 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output247
timestamp 1688980957
transform 1 0 20056 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output248
timestamp 1688980957
transform 1 0 20056 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output249
timestamp 1688980957
transform 1 0 20056 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output250
timestamp 1688980957
transform 1 0 20056 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output251
timestamp 1688980957
transform 1 0 20056 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output252
timestamp 1688980957
transform 1 0 18584 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1688980957
transform 1 0 15640 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output254
timestamp 1688980957
transform 1 0 19228 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output255
timestamp 1688980957
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output256
timestamp 1688980957
transform 1 0 18124 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output257
timestamp 1688980957
transform 1 0 20056 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output258
timestamp 1688980957
transform 1 0 20056 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output259
timestamp 1688980957
transform 1 0 16008 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output260
timestamp 1688980957
transform 1 0 18032 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output261
timestamp 1688980957
transform 1 0 17572 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output262
timestamp 1688980957
transform 1 0 17020 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output263
timestamp 1688980957
transform 1 0 18584 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output264
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output265
timestamp 1688980957
transform 1 0 17204 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output266
timestamp 1688980957
transform 1 0 16284 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output267
timestamp 1688980957
transform 1 0 17756 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output268
timestamp 1688980957
transform 1 0 16836 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output269
timestamp 1688980957
transform 1 0 18676 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output270
timestamp 1688980957
transform 1 0 17388 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output271
timestamp 1688980957
transform 1 0 18124 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output272
timestamp 1688980957
transform 1 0 17940 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output273
timestamp 1688980957
transform 1 0 1472 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output274
timestamp 1688980957
transform 1 0 2208 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output275
timestamp 1688980957
transform 1 0 2944 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output276
timestamp 1688980957
transform 1 0 2024 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output277
timestamp 1688980957
transform 1 0 1840 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output278
timestamp 1688980957
transform 1 0 2576 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output279
timestamp 1688980957
transform 1 0 2392 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output280
timestamp 1688980957
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output281
timestamp 1688980957
transform 1 0 2944 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output282
timestamp 1688980957
transform 1 0 3312 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output283
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output284
timestamp 1688980957
transform 1 0 4324 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output285
timestamp 1688980957
transform 1 0 4324 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output286
timestamp 1688980957
transform 1 0 3956 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output287
timestamp 1688980957
transform 1 0 4324 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output288
timestamp 1688980957
transform 1 0 4876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output289
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output290
timestamp 1688980957
transform 1 0 5704 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output291
timestamp 1688980957
transform 1 0 5428 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output292
timestamp 1688980957
transform 1 0 5152 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output293
timestamp 1688980957
transform 1 0 5428 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output294
timestamp 1688980957
transform 1 0 7636 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output295
timestamp 1688980957
transform 1 0 8188 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output296
timestamp 1688980957
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output297
timestamp 1688980957
transform 1 0 7360 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output298
timestamp 1688980957
transform 1 0 7912 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output299
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output300
timestamp 1688980957
transform 1 0 3956 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output301
timestamp 1688980957
transform 1 0 5980 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output302
timestamp 1688980957
transform 1 0 5796 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output303
timestamp 1688980957
transform 1 0 6532 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output304
timestamp 1688980957
transform 1 0 6532 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output305
timestamp 1688980957
transform 1 0 7084 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output306
timestamp 1688980957
transform 1 0 6624 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output307
timestamp 1688980957
transform 1 0 7636 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output308
timestamp 1688980957
transform 1 0 7084 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output309
timestamp 1688980957
transform 1 0 7728 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output310
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output311
timestamp 1688980957
transform 1 0 8648 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output312
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output313
timestamp 1688980957
transform 1 0 10488 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output314
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output315
timestamp 1688980957
transform 1 0 11684 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output316
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output317
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output318
timestamp 1688980957
transform 1 0 12420 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output319
timestamp 1688980957
transform 1 0 12972 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output320
timestamp 1688980957
transform 1 0 13524 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output321
timestamp 1688980957
transform 1 0 9844 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output322
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output323
timestamp 1688980957
transform 1 0 9752 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output324
timestamp 1688980957
transform 1 0 9568 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output325
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output326
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output327
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output328
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output329
timestamp 1688980957
transform 1 0 14996 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output330
timestamp 1688980957
transform 1 0 12236 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output331
timestamp 1688980957
transform 1 0 15088 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output332
timestamp 1688980957
transform 1 0 15640 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output333
timestamp 1688980957
transform 1 0 15640 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output334
timestamp 1688980957
transform 1 0 16836 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output335
timestamp 1688980957
transform 1 0 15824 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output336
timestamp 1688980957
transform 1 0 12788 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output337
timestamp 1688980957
transform 1 0 13340 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output338
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output339
timestamp 1688980957
transform 1 0 13892 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output340
timestamp 1688980957
transform 1 0 11868 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output341
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output342
timestamp 1688980957
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output343
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output344
timestamp 1688980957
transform 1 0 17756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output345
timestamp 1688980957
transform 1 0 16008 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output346
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output347
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output348
timestamp 1688980957
transform 1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output349
timestamp 1688980957
transform 1 0 1564 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output350
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output351
timestamp 1688980957
transform 1 0 1656 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output352
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output353
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output354
timestamp 1688980957
transform 1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output355
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output356
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output357
timestamp 1688980957
transform 1 0 4140 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output358
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output359
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output360
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output361
timestamp 1688980957
transform 1 0 3220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output362
timestamp 1688980957
transform 1 0 1748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output363
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output364
timestamp 1688980957
transform 1 0 4324 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output365
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output366
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output367
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output368
timestamp 1688980957
transform 1 0 2484 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output369
timestamp 1688980957
transform 1 0 1564 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output370
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output371
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output372
timestamp 1688980957
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output373
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output374
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output375
timestamp 1688980957
transform 1 0 1564 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output376
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output377
timestamp 1688980957
transform 1 0 1932 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output378
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output379
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output380
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output381
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output382
timestamp 1688980957
transform 1 0 1840 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output383
timestamp 1688980957
transform 1 0 2392 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output384
timestamp 1688980957
transform 1 0 1564 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output385
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output386
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output387
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output388
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output389
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output390
timestamp 1688980957
transform 1 0 1564 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output391
timestamp 1688980957
transform 1 0 1472 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output392
timestamp 1688980957
transform 1 0 5336 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output393
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 20884 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 20884 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 20884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 20884 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 20884 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 20884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 20884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 20884 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 20884 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 20884 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 20884 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 20884 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 20884 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 20884 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 20884 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 20884 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 20884 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 20884 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 20884 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 20884 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 20884 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 20884 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 20884 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 20884 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 20884 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 20884 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 20884 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 20884 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 20884 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 20884 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 20884 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 20884 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 20884 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 20884 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 20884 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 20884 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 20884 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 20884 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 20884 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 20884 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 20884 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 20884 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 20884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 20884 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 20884 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 20884 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 20884 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 20884 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 20884 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 20884 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 20884 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 20884 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 20884 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 20884 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 20884 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 12972 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 13340 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 14076 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 14444 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 14260 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 15180 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 14628 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 15548 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 14996 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 13524 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 13708 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 14628 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 14904 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 14444 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 15180 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 15456 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 15732 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 16008 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 15364 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 17664 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 15272 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 15732 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 15548 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 16100 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 16376 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 15824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 16836 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 17020 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 16928 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 16744 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 17296 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 16928 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 15456 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 15640 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 15916 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 16192 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 16836 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 17112 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 18584 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 17020 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 17204 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 17296 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 10580 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 16836 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 16928 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 18308 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 16652 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 19780 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 18032 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 17848 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 18584 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s 21840 9256 22300 9376 0 FreeSans 480 0 0 0 Config_accessC_bit0
port 0 nsew signal tristate
flabel metal3 s 21840 9800 22300 9920 0 FreeSans 480 0 0 0 Config_accessC_bit1
port 1 nsew signal tristate
flabel metal3 s 21840 10344 22300 10464 0 FreeSans 480 0 0 0 Config_accessC_bit2
port 2 nsew signal tristate
flabel metal3 s 21840 10888 22300 11008 0 FreeSans 480 0 0 0 Config_accessC_bit3
port 3 nsew signal tristate
flabel metal3 s -300 17960 160 18080 0 FreeSans 480 0 0 0 E1END[0]
port 4 nsew signal input
flabel metal3 s -300 18232 160 18352 0 FreeSans 480 0 0 0 E1END[1]
port 5 nsew signal input
flabel metal3 s -300 18504 160 18624 0 FreeSans 480 0 0 0 E1END[2]
port 6 nsew signal input
flabel metal3 s -300 18776 160 18896 0 FreeSans 480 0 0 0 E1END[3]
port 7 nsew signal input
flabel metal3 s -300 21224 160 21344 0 FreeSans 480 0 0 0 E2END[0]
port 8 nsew signal input
flabel metal3 s -300 21496 160 21616 0 FreeSans 480 0 0 0 E2END[1]
port 9 nsew signal input
flabel metal3 s -300 21768 160 21888 0 FreeSans 480 0 0 0 E2END[2]
port 10 nsew signal input
flabel metal3 s -300 22040 160 22160 0 FreeSans 480 0 0 0 E2END[3]
port 11 nsew signal input
flabel metal3 s -300 22312 160 22432 0 FreeSans 480 0 0 0 E2END[4]
port 12 nsew signal input
flabel metal3 s -300 22584 160 22704 0 FreeSans 480 0 0 0 E2END[5]
port 13 nsew signal input
flabel metal3 s -300 22856 160 22976 0 FreeSans 480 0 0 0 E2END[6]
port 14 nsew signal input
flabel metal3 s -300 23128 160 23248 0 FreeSans 480 0 0 0 E2END[7]
port 15 nsew signal input
flabel metal3 s -300 19048 160 19168 0 FreeSans 480 0 0 0 E2MID[0]
port 16 nsew signal input
flabel metal3 s -300 19320 160 19440 0 FreeSans 480 0 0 0 E2MID[1]
port 17 nsew signal input
flabel metal3 s -300 19592 160 19712 0 FreeSans 480 0 0 0 E2MID[2]
port 18 nsew signal input
flabel metal3 s -300 19864 160 19984 0 FreeSans 480 0 0 0 E2MID[3]
port 19 nsew signal input
flabel metal3 s -300 20136 160 20256 0 FreeSans 480 0 0 0 E2MID[4]
port 20 nsew signal input
flabel metal3 s -300 20408 160 20528 0 FreeSans 480 0 0 0 E2MID[5]
port 21 nsew signal input
flabel metal3 s -300 20680 160 20800 0 FreeSans 480 0 0 0 E2MID[6]
port 22 nsew signal input
flabel metal3 s -300 20952 160 21072 0 FreeSans 480 0 0 0 E2MID[7]
port 23 nsew signal input
flabel metal3 s -300 27752 160 27872 0 FreeSans 480 0 0 0 E6END[0]
port 24 nsew signal input
flabel metal3 s -300 30472 160 30592 0 FreeSans 480 0 0 0 E6END[10]
port 25 nsew signal input
flabel metal3 s -300 30744 160 30864 0 FreeSans 480 0 0 0 E6END[11]
port 26 nsew signal input
flabel metal3 s -300 28024 160 28144 0 FreeSans 480 0 0 0 E6END[1]
port 27 nsew signal input
flabel metal3 s -300 28296 160 28416 0 FreeSans 480 0 0 0 E6END[2]
port 28 nsew signal input
flabel metal3 s -300 28568 160 28688 0 FreeSans 480 0 0 0 E6END[3]
port 29 nsew signal input
flabel metal3 s -300 28840 160 28960 0 FreeSans 480 0 0 0 E6END[4]
port 30 nsew signal input
flabel metal3 s -300 29112 160 29232 0 FreeSans 480 0 0 0 E6END[5]
port 31 nsew signal input
flabel metal3 s -300 29384 160 29504 0 FreeSans 480 0 0 0 E6END[6]
port 32 nsew signal input
flabel metal3 s -300 29656 160 29776 0 FreeSans 480 0 0 0 E6END[7]
port 33 nsew signal input
flabel metal3 s -300 29928 160 30048 0 FreeSans 480 0 0 0 E6END[8]
port 34 nsew signal input
flabel metal3 s -300 30200 160 30320 0 FreeSans 480 0 0 0 E6END[9]
port 35 nsew signal input
flabel metal3 s -300 23400 160 23520 0 FreeSans 480 0 0 0 EE4END[0]
port 36 nsew signal input
flabel metal3 s -300 26120 160 26240 0 FreeSans 480 0 0 0 EE4END[10]
port 37 nsew signal input
flabel metal3 s -300 26392 160 26512 0 FreeSans 480 0 0 0 EE4END[11]
port 38 nsew signal input
flabel metal3 s -300 26664 160 26784 0 FreeSans 480 0 0 0 EE4END[12]
port 39 nsew signal input
flabel metal3 s -300 26936 160 27056 0 FreeSans 480 0 0 0 EE4END[13]
port 40 nsew signal input
flabel metal3 s -300 27208 160 27328 0 FreeSans 480 0 0 0 EE4END[14]
port 41 nsew signal input
flabel metal3 s -300 27480 160 27600 0 FreeSans 480 0 0 0 EE4END[15]
port 42 nsew signal input
flabel metal3 s -300 23672 160 23792 0 FreeSans 480 0 0 0 EE4END[1]
port 43 nsew signal input
flabel metal3 s -300 23944 160 24064 0 FreeSans 480 0 0 0 EE4END[2]
port 44 nsew signal input
flabel metal3 s -300 24216 160 24336 0 FreeSans 480 0 0 0 EE4END[3]
port 45 nsew signal input
flabel metal3 s -300 24488 160 24608 0 FreeSans 480 0 0 0 EE4END[4]
port 46 nsew signal input
flabel metal3 s -300 24760 160 24880 0 FreeSans 480 0 0 0 EE4END[5]
port 47 nsew signal input
flabel metal3 s -300 25032 160 25152 0 FreeSans 480 0 0 0 EE4END[6]
port 48 nsew signal input
flabel metal3 s -300 25304 160 25424 0 FreeSans 480 0 0 0 EE4END[7]
port 49 nsew signal input
flabel metal3 s -300 25576 160 25696 0 FreeSans 480 0 0 0 EE4END[8]
port 50 nsew signal input
flabel metal3 s -300 25848 160 25968 0 FreeSans 480 0 0 0 EE4END[9]
port 51 nsew signal input
flabel metal3 s 21840 15784 22300 15904 0 FreeSans 480 0 0 0 FAB2RAM_A0_O0
port 52 nsew signal tristate
flabel metal3 s 21840 16328 22300 16448 0 FreeSans 480 0 0 0 FAB2RAM_A0_O1
port 53 nsew signal tristate
flabel metal3 s 21840 16872 22300 16992 0 FreeSans 480 0 0 0 FAB2RAM_A0_O2
port 54 nsew signal tristate
flabel metal3 s 21840 17416 22300 17536 0 FreeSans 480 0 0 0 FAB2RAM_A0_O3
port 55 nsew signal tristate
flabel metal3 s 21840 13608 22300 13728 0 FreeSans 480 0 0 0 FAB2RAM_A1_O0
port 56 nsew signal tristate
flabel metal3 s 21840 14152 22300 14272 0 FreeSans 480 0 0 0 FAB2RAM_A1_O1
port 57 nsew signal tristate
flabel metal3 s 21840 14696 22300 14816 0 FreeSans 480 0 0 0 FAB2RAM_A1_O2
port 58 nsew signal tristate
flabel metal3 s 21840 15240 22300 15360 0 FreeSans 480 0 0 0 FAB2RAM_A1_O3
port 59 nsew signal tristate
flabel metal3 s 21840 11432 22300 11552 0 FreeSans 480 0 0 0 FAB2RAM_C_O0
port 60 nsew signal tristate
flabel metal3 s 21840 11976 22300 12096 0 FreeSans 480 0 0 0 FAB2RAM_C_O1
port 61 nsew signal tristate
flabel metal3 s 21840 12520 22300 12640 0 FreeSans 480 0 0 0 FAB2RAM_C_O2
port 62 nsew signal tristate
flabel metal3 s 21840 13064 22300 13184 0 FreeSans 480 0 0 0 FAB2RAM_C_O3
port 63 nsew signal tristate
flabel metal3 s 21840 24488 22300 24608 0 FreeSans 480 0 0 0 FAB2RAM_D0_O0
port 64 nsew signal tristate
flabel metal3 s 21840 25032 22300 25152 0 FreeSans 480 0 0 0 FAB2RAM_D0_O1
port 65 nsew signal tristate
flabel metal3 s 21840 25576 22300 25696 0 FreeSans 480 0 0 0 FAB2RAM_D0_O2
port 66 nsew signal tristate
flabel metal3 s 21840 26120 22300 26240 0 FreeSans 480 0 0 0 FAB2RAM_D0_O3
port 67 nsew signal tristate
flabel metal3 s 21840 22312 22300 22432 0 FreeSans 480 0 0 0 FAB2RAM_D1_O0
port 68 nsew signal tristate
flabel metal3 s 21840 22856 22300 22976 0 FreeSans 480 0 0 0 FAB2RAM_D1_O1
port 69 nsew signal tristate
flabel metal3 s 21840 23400 22300 23520 0 FreeSans 480 0 0 0 FAB2RAM_D1_O2
port 70 nsew signal tristate
flabel metal3 s 21840 23944 22300 24064 0 FreeSans 480 0 0 0 FAB2RAM_D1_O3
port 71 nsew signal tristate
flabel metal3 s 21840 20136 22300 20256 0 FreeSans 480 0 0 0 FAB2RAM_D2_O0
port 72 nsew signal tristate
flabel metal3 s 21840 20680 22300 20800 0 FreeSans 480 0 0 0 FAB2RAM_D2_O1
port 73 nsew signal tristate
flabel metal3 s 21840 21224 22300 21344 0 FreeSans 480 0 0 0 FAB2RAM_D2_O2
port 74 nsew signal tristate
flabel metal3 s 21840 21768 22300 21888 0 FreeSans 480 0 0 0 FAB2RAM_D2_O3
port 75 nsew signal tristate
flabel metal3 s 21840 17960 22300 18080 0 FreeSans 480 0 0 0 FAB2RAM_D3_O0
port 76 nsew signal tristate
flabel metal3 s 21840 18504 22300 18624 0 FreeSans 480 0 0 0 FAB2RAM_D3_O1
port 77 nsew signal tristate
flabel metal3 s 21840 19048 22300 19168 0 FreeSans 480 0 0 0 FAB2RAM_D3_O2
port 78 nsew signal tristate
flabel metal3 s 21840 19592 22300 19712 0 FreeSans 480 0 0 0 FAB2RAM_D3_O3
port 79 nsew signal tristate
flabel metal3 s -300 31016 160 31136 0 FreeSans 480 0 0 0 FrameData[0]
port 80 nsew signal input
flabel metal3 s -300 33736 160 33856 0 FreeSans 480 0 0 0 FrameData[10]
port 81 nsew signal input
flabel metal3 s -300 34008 160 34128 0 FreeSans 480 0 0 0 FrameData[11]
port 82 nsew signal input
flabel metal3 s -300 34280 160 34400 0 FreeSans 480 0 0 0 FrameData[12]
port 83 nsew signal input
flabel metal3 s -300 34552 160 34672 0 FreeSans 480 0 0 0 FrameData[13]
port 84 nsew signal input
flabel metal3 s -300 34824 160 34944 0 FreeSans 480 0 0 0 FrameData[14]
port 85 nsew signal input
flabel metal3 s -300 35096 160 35216 0 FreeSans 480 0 0 0 FrameData[15]
port 86 nsew signal input
flabel metal3 s -300 35368 160 35488 0 FreeSans 480 0 0 0 FrameData[16]
port 87 nsew signal input
flabel metal3 s -300 35640 160 35760 0 FreeSans 480 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s -300 35912 160 36032 0 FreeSans 480 0 0 0 FrameData[18]
port 89 nsew signal input
flabel metal3 s -300 36184 160 36304 0 FreeSans 480 0 0 0 FrameData[19]
port 90 nsew signal input
flabel metal3 s -300 31288 160 31408 0 FreeSans 480 0 0 0 FrameData[1]
port 91 nsew signal input
flabel metal3 s -300 36456 160 36576 0 FreeSans 480 0 0 0 FrameData[20]
port 92 nsew signal input
flabel metal3 s -300 36728 160 36848 0 FreeSans 480 0 0 0 FrameData[21]
port 93 nsew signal input
flabel metal3 s -300 37000 160 37120 0 FreeSans 480 0 0 0 FrameData[22]
port 94 nsew signal input
flabel metal3 s -300 37272 160 37392 0 FreeSans 480 0 0 0 FrameData[23]
port 95 nsew signal input
flabel metal3 s -300 37544 160 37664 0 FreeSans 480 0 0 0 FrameData[24]
port 96 nsew signal input
flabel metal3 s -300 37816 160 37936 0 FreeSans 480 0 0 0 FrameData[25]
port 97 nsew signal input
flabel metal3 s -300 38088 160 38208 0 FreeSans 480 0 0 0 FrameData[26]
port 98 nsew signal input
flabel metal3 s -300 38360 160 38480 0 FreeSans 480 0 0 0 FrameData[27]
port 99 nsew signal input
flabel metal3 s -300 38632 160 38752 0 FreeSans 480 0 0 0 FrameData[28]
port 100 nsew signal input
flabel metal3 s -300 38904 160 39024 0 FreeSans 480 0 0 0 FrameData[29]
port 101 nsew signal input
flabel metal3 s -300 31560 160 31680 0 FreeSans 480 0 0 0 FrameData[2]
port 102 nsew signal input
flabel metal3 s -300 39176 160 39296 0 FreeSans 480 0 0 0 FrameData[30]
port 103 nsew signal input
flabel metal3 s -300 39448 160 39568 0 FreeSans 480 0 0 0 FrameData[31]
port 104 nsew signal input
flabel metal3 s -300 31832 160 31952 0 FreeSans 480 0 0 0 FrameData[3]
port 105 nsew signal input
flabel metal3 s -300 32104 160 32224 0 FreeSans 480 0 0 0 FrameData[4]
port 106 nsew signal input
flabel metal3 s -300 32376 160 32496 0 FreeSans 480 0 0 0 FrameData[5]
port 107 nsew signal input
flabel metal3 s -300 32648 160 32768 0 FreeSans 480 0 0 0 FrameData[6]
port 108 nsew signal input
flabel metal3 s -300 32920 160 33040 0 FreeSans 480 0 0 0 FrameData[7]
port 109 nsew signal input
flabel metal3 s -300 33192 160 33312 0 FreeSans 480 0 0 0 FrameData[8]
port 110 nsew signal input
flabel metal3 s -300 33464 160 33584 0 FreeSans 480 0 0 0 FrameData[9]
port 111 nsew signal input
flabel metal3 s 21840 26664 22300 26784 0 FreeSans 480 0 0 0 FrameData_O[0]
port 112 nsew signal tristate
flabel metal3 s 21840 32104 22300 32224 0 FreeSans 480 0 0 0 FrameData_O[10]
port 113 nsew signal tristate
flabel metal3 s 21840 32648 22300 32768 0 FreeSans 480 0 0 0 FrameData_O[11]
port 114 nsew signal tristate
flabel metal3 s 21840 33192 22300 33312 0 FreeSans 480 0 0 0 FrameData_O[12]
port 115 nsew signal tristate
flabel metal3 s 21840 33736 22300 33856 0 FreeSans 480 0 0 0 FrameData_O[13]
port 116 nsew signal tristate
flabel metal3 s 21840 34280 22300 34400 0 FreeSans 480 0 0 0 FrameData_O[14]
port 117 nsew signal tristate
flabel metal3 s 21840 34824 22300 34944 0 FreeSans 480 0 0 0 FrameData_O[15]
port 118 nsew signal tristate
flabel metal3 s 21840 35368 22300 35488 0 FreeSans 480 0 0 0 FrameData_O[16]
port 119 nsew signal tristate
flabel metal3 s 21840 35912 22300 36032 0 FreeSans 480 0 0 0 FrameData_O[17]
port 120 nsew signal tristate
flabel metal3 s 21840 36456 22300 36576 0 FreeSans 480 0 0 0 FrameData_O[18]
port 121 nsew signal tristate
flabel metal3 s 21840 37000 22300 37120 0 FreeSans 480 0 0 0 FrameData_O[19]
port 122 nsew signal tristate
flabel metal3 s 21840 27208 22300 27328 0 FreeSans 480 0 0 0 FrameData_O[1]
port 123 nsew signal tristate
flabel metal3 s 21840 37544 22300 37664 0 FreeSans 480 0 0 0 FrameData_O[20]
port 124 nsew signal tristate
flabel metal3 s 21840 38088 22300 38208 0 FreeSans 480 0 0 0 FrameData_O[21]
port 125 nsew signal tristate
flabel metal3 s 21840 38632 22300 38752 0 FreeSans 480 0 0 0 FrameData_O[22]
port 126 nsew signal tristate
flabel metal3 s 21840 39176 22300 39296 0 FreeSans 480 0 0 0 FrameData_O[23]
port 127 nsew signal tristate
flabel metal3 s 21840 39720 22300 39840 0 FreeSans 480 0 0 0 FrameData_O[24]
port 128 nsew signal tristate
flabel metal3 s 21840 40264 22300 40384 0 FreeSans 480 0 0 0 FrameData_O[25]
port 129 nsew signal tristate
flabel metal3 s 21840 40808 22300 40928 0 FreeSans 480 0 0 0 FrameData_O[26]
port 130 nsew signal tristate
flabel metal3 s 21840 41352 22300 41472 0 FreeSans 480 0 0 0 FrameData_O[27]
port 131 nsew signal tristate
flabel metal3 s 21840 41896 22300 42016 0 FreeSans 480 0 0 0 FrameData_O[28]
port 132 nsew signal tristate
flabel metal3 s 21840 42440 22300 42560 0 FreeSans 480 0 0 0 FrameData_O[29]
port 133 nsew signal tristate
flabel metal3 s 21840 27752 22300 27872 0 FreeSans 480 0 0 0 FrameData_O[2]
port 134 nsew signal tristate
flabel metal3 s 21840 42984 22300 43104 0 FreeSans 480 0 0 0 FrameData_O[30]
port 135 nsew signal tristate
flabel metal3 s 21840 43528 22300 43648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 136 nsew signal tristate
flabel metal3 s 21840 28296 22300 28416 0 FreeSans 480 0 0 0 FrameData_O[3]
port 137 nsew signal tristate
flabel metal3 s 21840 28840 22300 28960 0 FreeSans 480 0 0 0 FrameData_O[4]
port 138 nsew signal tristate
flabel metal3 s 21840 29384 22300 29504 0 FreeSans 480 0 0 0 FrameData_O[5]
port 139 nsew signal tristate
flabel metal3 s 21840 29928 22300 30048 0 FreeSans 480 0 0 0 FrameData_O[6]
port 140 nsew signal tristate
flabel metal3 s 21840 30472 22300 30592 0 FreeSans 480 0 0 0 FrameData_O[7]
port 141 nsew signal tristate
flabel metal3 s 21840 31016 22300 31136 0 FreeSans 480 0 0 0 FrameData_O[8]
port 142 nsew signal tristate
flabel metal3 s 21840 31560 22300 31680 0 FreeSans 480 0 0 0 FrameData_O[9]
port 143 nsew signal tristate
flabel metal2 s 15842 -300 15898 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 144 nsew signal input
flabel metal2 s 17682 -300 17738 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 145 nsew signal input
flabel metal2 s 17866 -300 17922 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 146 nsew signal input
flabel metal2 s 18050 -300 18106 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 147 nsew signal input
flabel metal2 s 18234 -300 18290 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 148 nsew signal input
flabel metal2 s 18418 -300 18474 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 149 nsew signal input
flabel metal2 s 18602 -300 18658 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 150 nsew signal input
flabel metal2 s 18786 -300 18842 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 151 nsew signal input
flabel metal2 s 18970 -300 19026 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 152 nsew signal input
flabel metal2 s 19154 -300 19210 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 153 nsew signal input
flabel metal2 s 19338 -300 19394 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 154 nsew signal input
flabel metal2 s 16026 -300 16082 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 155 nsew signal input
flabel metal2 s 16210 -300 16266 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 156 nsew signal input
flabel metal2 s 16394 -300 16450 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 157 nsew signal input
flabel metal2 s 16578 -300 16634 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 158 nsew signal input
flabel metal2 s 16762 -300 16818 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 159 nsew signal input
flabel metal2 s 16946 -300 17002 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 160 nsew signal input
flabel metal2 s 17130 -300 17186 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 161 nsew signal input
flabel metal2 s 17314 -300 17370 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 162 nsew signal input
flabel metal2 s 17498 -300 17554 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 163 nsew signal input
flabel metal2 s 15842 44540 15898 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 164 nsew signal tristate
flabel metal2 s 17682 44540 17738 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 165 nsew signal tristate
flabel metal2 s 17866 44540 17922 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 166 nsew signal tristate
flabel metal2 s 18050 44540 18106 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 167 nsew signal tristate
flabel metal2 s 18234 44540 18290 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 168 nsew signal tristate
flabel metal2 s 18418 44540 18474 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 169 nsew signal tristate
flabel metal2 s 18602 44540 18658 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 170 nsew signal tristate
flabel metal2 s 18786 44540 18842 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 171 nsew signal tristate
flabel metal2 s 18970 44540 19026 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 172 nsew signal tristate
flabel metal2 s 19154 44540 19210 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 173 nsew signal tristate
flabel metal2 s 19338 44540 19394 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 174 nsew signal tristate
flabel metal2 s 16026 44540 16082 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 175 nsew signal tristate
flabel metal2 s 16210 44540 16266 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 176 nsew signal tristate
flabel metal2 s 16394 44540 16450 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 177 nsew signal tristate
flabel metal2 s 16578 44540 16634 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 178 nsew signal tristate
flabel metal2 s 16762 44540 16818 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 179 nsew signal tristate
flabel metal2 s 16946 44540 17002 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 180 nsew signal tristate
flabel metal2 s 17130 44540 17186 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 181 nsew signal tristate
flabel metal2 s 17314 44540 17370 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 182 nsew signal tristate
flabel metal2 s 17498 44540 17554 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 183 nsew signal tristate
flabel metal2 s 2410 44540 2466 45000 0 FreeSans 224 90 0 0 N1BEG[0]
port 184 nsew signal tristate
flabel metal2 s 2594 44540 2650 45000 0 FreeSans 224 90 0 0 N1BEG[1]
port 185 nsew signal tristate
flabel metal2 s 2778 44540 2834 45000 0 FreeSans 224 90 0 0 N1BEG[2]
port 186 nsew signal tristate
flabel metal2 s 2962 44540 3018 45000 0 FreeSans 224 90 0 0 N1BEG[3]
port 187 nsew signal tristate
flabel metal2 s 2410 -300 2466 160 0 FreeSans 224 90 0 0 N1END[0]
port 188 nsew signal input
flabel metal2 s 2594 -300 2650 160 0 FreeSans 224 90 0 0 N1END[1]
port 189 nsew signal input
flabel metal2 s 2778 -300 2834 160 0 FreeSans 224 90 0 0 N1END[2]
port 190 nsew signal input
flabel metal2 s 2962 -300 3018 160 0 FreeSans 224 90 0 0 N1END[3]
port 191 nsew signal input
flabel metal2 s 3146 44540 3202 45000 0 FreeSans 224 90 0 0 N2BEG[0]
port 192 nsew signal tristate
flabel metal2 s 3330 44540 3386 45000 0 FreeSans 224 90 0 0 N2BEG[1]
port 193 nsew signal tristate
flabel metal2 s 3514 44540 3570 45000 0 FreeSans 224 90 0 0 N2BEG[2]
port 194 nsew signal tristate
flabel metal2 s 3698 44540 3754 45000 0 FreeSans 224 90 0 0 N2BEG[3]
port 195 nsew signal tristate
flabel metal2 s 3882 44540 3938 45000 0 FreeSans 224 90 0 0 N2BEG[4]
port 196 nsew signal tristate
flabel metal2 s 4066 44540 4122 45000 0 FreeSans 224 90 0 0 N2BEG[5]
port 197 nsew signal tristate
flabel metal2 s 4250 44540 4306 45000 0 FreeSans 224 90 0 0 N2BEG[6]
port 198 nsew signal tristate
flabel metal2 s 4434 44540 4490 45000 0 FreeSans 224 90 0 0 N2BEG[7]
port 199 nsew signal tristate
flabel metal2 s 4618 44540 4674 45000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 200 nsew signal tristate
flabel metal2 s 4802 44540 4858 45000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 201 nsew signal tristate
flabel metal2 s 4986 44540 5042 45000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 202 nsew signal tristate
flabel metal2 s 5170 44540 5226 45000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 203 nsew signal tristate
flabel metal2 s 5354 44540 5410 45000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 204 nsew signal tristate
flabel metal2 s 5538 44540 5594 45000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 205 nsew signal tristate
flabel metal2 s 5722 44540 5778 45000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 206 nsew signal tristate
flabel metal2 s 5906 44540 5962 45000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 207 nsew signal tristate
flabel metal2 s 4618 -300 4674 160 0 FreeSans 224 90 0 0 N2END[0]
port 208 nsew signal input
flabel metal2 s 4802 -300 4858 160 0 FreeSans 224 90 0 0 N2END[1]
port 209 nsew signal input
flabel metal2 s 4986 -300 5042 160 0 FreeSans 224 90 0 0 N2END[2]
port 210 nsew signal input
flabel metal2 s 5170 -300 5226 160 0 FreeSans 224 90 0 0 N2END[3]
port 211 nsew signal input
flabel metal2 s 5354 -300 5410 160 0 FreeSans 224 90 0 0 N2END[4]
port 212 nsew signal input
flabel metal2 s 5538 -300 5594 160 0 FreeSans 224 90 0 0 N2END[5]
port 213 nsew signal input
flabel metal2 s 5722 -300 5778 160 0 FreeSans 224 90 0 0 N2END[6]
port 214 nsew signal input
flabel metal2 s 5906 -300 5962 160 0 FreeSans 224 90 0 0 N2END[7]
port 215 nsew signal input
flabel metal2 s 3146 -300 3202 160 0 FreeSans 224 90 0 0 N2MID[0]
port 216 nsew signal input
flabel metal2 s 3330 -300 3386 160 0 FreeSans 224 90 0 0 N2MID[1]
port 217 nsew signal input
flabel metal2 s 3514 -300 3570 160 0 FreeSans 224 90 0 0 N2MID[2]
port 218 nsew signal input
flabel metal2 s 3698 -300 3754 160 0 FreeSans 224 90 0 0 N2MID[3]
port 219 nsew signal input
flabel metal2 s 3882 -300 3938 160 0 FreeSans 224 90 0 0 N2MID[4]
port 220 nsew signal input
flabel metal2 s 4066 -300 4122 160 0 FreeSans 224 90 0 0 N2MID[5]
port 221 nsew signal input
flabel metal2 s 4250 -300 4306 160 0 FreeSans 224 90 0 0 N2MID[6]
port 222 nsew signal input
flabel metal2 s 4434 -300 4490 160 0 FreeSans 224 90 0 0 N2MID[7]
port 223 nsew signal input
flabel metal2 s 6090 44540 6146 45000 0 FreeSans 224 90 0 0 N4BEG[0]
port 224 nsew signal tristate
flabel metal2 s 7930 44540 7986 45000 0 FreeSans 224 90 0 0 N4BEG[10]
port 225 nsew signal tristate
flabel metal2 s 8114 44540 8170 45000 0 FreeSans 224 90 0 0 N4BEG[11]
port 226 nsew signal tristate
flabel metal2 s 8298 44540 8354 45000 0 FreeSans 224 90 0 0 N4BEG[12]
port 227 nsew signal tristate
flabel metal2 s 8482 44540 8538 45000 0 FreeSans 224 90 0 0 N4BEG[13]
port 228 nsew signal tristate
flabel metal2 s 8666 44540 8722 45000 0 FreeSans 224 90 0 0 N4BEG[14]
port 229 nsew signal tristate
flabel metal2 s 8850 44540 8906 45000 0 FreeSans 224 90 0 0 N4BEG[15]
port 230 nsew signal tristate
flabel metal2 s 6274 44540 6330 45000 0 FreeSans 224 90 0 0 N4BEG[1]
port 231 nsew signal tristate
flabel metal2 s 6458 44540 6514 45000 0 FreeSans 224 90 0 0 N4BEG[2]
port 232 nsew signal tristate
flabel metal2 s 6642 44540 6698 45000 0 FreeSans 224 90 0 0 N4BEG[3]
port 233 nsew signal tristate
flabel metal2 s 6826 44540 6882 45000 0 FreeSans 224 90 0 0 N4BEG[4]
port 234 nsew signal tristate
flabel metal2 s 7010 44540 7066 45000 0 FreeSans 224 90 0 0 N4BEG[5]
port 235 nsew signal tristate
flabel metal2 s 7194 44540 7250 45000 0 FreeSans 224 90 0 0 N4BEG[6]
port 236 nsew signal tristate
flabel metal2 s 7378 44540 7434 45000 0 FreeSans 224 90 0 0 N4BEG[7]
port 237 nsew signal tristate
flabel metal2 s 7562 44540 7618 45000 0 FreeSans 224 90 0 0 N4BEG[8]
port 238 nsew signal tristate
flabel metal2 s 7746 44540 7802 45000 0 FreeSans 224 90 0 0 N4BEG[9]
port 239 nsew signal tristate
flabel metal2 s 6090 -300 6146 160 0 FreeSans 224 90 0 0 N4END[0]
port 240 nsew signal input
flabel metal2 s 7930 -300 7986 160 0 FreeSans 224 90 0 0 N4END[10]
port 241 nsew signal input
flabel metal2 s 8114 -300 8170 160 0 FreeSans 224 90 0 0 N4END[11]
port 242 nsew signal input
flabel metal2 s 8298 -300 8354 160 0 FreeSans 224 90 0 0 N4END[12]
port 243 nsew signal input
flabel metal2 s 8482 -300 8538 160 0 FreeSans 224 90 0 0 N4END[13]
port 244 nsew signal input
flabel metal2 s 8666 -300 8722 160 0 FreeSans 224 90 0 0 N4END[14]
port 245 nsew signal input
flabel metal2 s 8850 -300 8906 160 0 FreeSans 224 90 0 0 N4END[15]
port 246 nsew signal input
flabel metal2 s 6274 -300 6330 160 0 FreeSans 224 90 0 0 N4END[1]
port 247 nsew signal input
flabel metal2 s 6458 -300 6514 160 0 FreeSans 224 90 0 0 N4END[2]
port 248 nsew signal input
flabel metal2 s 6642 -300 6698 160 0 FreeSans 224 90 0 0 N4END[3]
port 249 nsew signal input
flabel metal2 s 6826 -300 6882 160 0 FreeSans 224 90 0 0 N4END[4]
port 250 nsew signal input
flabel metal2 s 7010 -300 7066 160 0 FreeSans 224 90 0 0 N4END[5]
port 251 nsew signal input
flabel metal2 s 7194 -300 7250 160 0 FreeSans 224 90 0 0 N4END[6]
port 252 nsew signal input
flabel metal2 s 7378 -300 7434 160 0 FreeSans 224 90 0 0 N4END[7]
port 253 nsew signal input
flabel metal2 s 7562 -300 7618 160 0 FreeSans 224 90 0 0 N4END[8]
port 254 nsew signal input
flabel metal2 s 7746 -300 7802 160 0 FreeSans 224 90 0 0 N4END[9]
port 255 nsew signal input
flabel metal3 s 21840 7080 22300 7200 0 FreeSans 480 0 0 0 RAM2FAB_D0_I0
port 256 nsew signal input
flabel metal3 s 21840 7624 22300 7744 0 FreeSans 480 0 0 0 RAM2FAB_D0_I1
port 257 nsew signal input
flabel metal3 s 21840 8168 22300 8288 0 FreeSans 480 0 0 0 RAM2FAB_D0_I2
port 258 nsew signal input
flabel metal3 s 21840 8712 22300 8832 0 FreeSans 480 0 0 0 RAM2FAB_D0_I3
port 259 nsew signal input
flabel metal3 s 21840 4904 22300 5024 0 FreeSans 480 0 0 0 RAM2FAB_D1_I0
port 260 nsew signal input
flabel metal3 s 21840 5448 22300 5568 0 FreeSans 480 0 0 0 RAM2FAB_D1_I1
port 261 nsew signal input
flabel metal3 s 21840 5992 22300 6112 0 FreeSans 480 0 0 0 RAM2FAB_D1_I2
port 262 nsew signal input
flabel metal3 s 21840 6536 22300 6656 0 FreeSans 480 0 0 0 RAM2FAB_D1_I3
port 263 nsew signal input
flabel metal3 s 21840 2728 22300 2848 0 FreeSans 480 0 0 0 RAM2FAB_D2_I0
port 264 nsew signal input
flabel metal3 s 21840 3272 22300 3392 0 FreeSans 480 0 0 0 RAM2FAB_D2_I1
port 265 nsew signal input
flabel metal3 s 21840 3816 22300 3936 0 FreeSans 480 0 0 0 RAM2FAB_D2_I2
port 266 nsew signal input
flabel metal3 s 21840 4360 22300 4480 0 FreeSans 480 0 0 0 RAM2FAB_D2_I3
port 267 nsew signal input
flabel metal3 s 21840 552 22300 672 0 FreeSans 480 0 0 0 RAM2FAB_D3_I0
port 268 nsew signal input
flabel metal3 s 21840 1096 22300 1216 0 FreeSans 480 0 0 0 RAM2FAB_D3_I1
port 269 nsew signal input
flabel metal3 s 21840 1640 22300 1760 0 FreeSans 480 0 0 0 RAM2FAB_D3_I2
port 270 nsew signal input
flabel metal3 s 21840 2184 22300 2304 0 FreeSans 480 0 0 0 RAM2FAB_D3_I3
port 271 nsew signal input
flabel metal2 s 9034 -300 9090 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 272 nsew signal tristate
flabel metal2 s 9218 -300 9274 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 273 nsew signal tristate
flabel metal2 s 9402 -300 9458 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 274 nsew signal tristate
flabel metal2 s 9586 -300 9642 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 275 nsew signal tristate
flabel metal2 s 9034 44540 9090 45000 0 FreeSans 224 90 0 0 S1END[0]
port 276 nsew signal input
flabel metal2 s 9218 44540 9274 45000 0 FreeSans 224 90 0 0 S1END[1]
port 277 nsew signal input
flabel metal2 s 9402 44540 9458 45000 0 FreeSans 224 90 0 0 S1END[2]
port 278 nsew signal input
flabel metal2 s 9586 44540 9642 45000 0 FreeSans 224 90 0 0 S1END[3]
port 279 nsew signal input
flabel metal2 s 11242 -300 11298 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 280 nsew signal tristate
flabel metal2 s 11426 -300 11482 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 281 nsew signal tristate
flabel metal2 s 11610 -300 11666 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 282 nsew signal tristate
flabel metal2 s 11794 -300 11850 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 283 nsew signal tristate
flabel metal2 s 11978 -300 12034 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 284 nsew signal tristate
flabel metal2 s 12162 -300 12218 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 285 nsew signal tristate
flabel metal2 s 12346 -300 12402 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 286 nsew signal tristate
flabel metal2 s 12530 -300 12586 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 287 nsew signal tristate
flabel metal2 s 9770 -300 9826 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 288 nsew signal tristate
flabel metal2 s 9954 -300 10010 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 289 nsew signal tristate
flabel metal2 s 10138 -300 10194 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 290 nsew signal tristate
flabel metal2 s 10322 -300 10378 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 291 nsew signal tristate
flabel metal2 s 10506 -300 10562 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 292 nsew signal tristate
flabel metal2 s 10690 -300 10746 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 293 nsew signal tristate
flabel metal2 s 10874 -300 10930 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 294 nsew signal tristate
flabel metal2 s 11058 -300 11114 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 295 nsew signal tristate
flabel metal2 s 9770 44540 9826 45000 0 FreeSans 224 90 0 0 S2END[0]
port 296 nsew signal input
flabel metal2 s 9954 44540 10010 45000 0 FreeSans 224 90 0 0 S2END[1]
port 297 nsew signal input
flabel metal2 s 10138 44540 10194 45000 0 FreeSans 224 90 0 0 S2END[2]
port 298 nsew signal input
flabel metal2 s 10322 44540 10378 45000 0 FreeSans 224 90 0 0 S2END[3]
port 299 nsew signal input
flabel metal2 s 10506 44540 10562 45000 0 FreeSans 224 90 0 0 S2END[4]
port 300 nsew signal input
flabel metal2 s 10690 44540 10746 45000 0 FreeSans 224 90 0 0 S2END[5]
port 301 nsew signal input
flabel metal2 s 10874 44540 10930 45000 0 FreeSans 224 90 0 0 S2END[6]
port 302 nsew signal input
flabel metal2 s 11058 44540 11114 45000 0 FreeSans 224 90 0 0 S2END[7]
port 303 nsew signal input
flabel metal2 s 11242 44540 11298 45000 0 FreeSans 224 90 0 0 S2MID[0]
port 304 nsew signal input
flabel metal2 s 11426 44540 11482 45000 0 FreeSans 224 90 0 0 S2MID[1]
port 305 nsew signal input
flabel metal2 s 11610 44540 11666 45000 0 FreeSans 224 90 0 0 S2MID[2]
port 306 nsew signal input
flabel metal2 s 11794 44540 11850 45000 0 FreeSans 224 90 0 0 S2MID[3]
port 307 nsew signal input
flabel metal2 s 11978 44540 12034 45000 0 FreeSans 224 90 0 0 S2MID[4]
port 308 nsew signal input
flabel metal2 s 12162 44540 12218 45000 0 FreeSans 224 90 0 0 S2MID[5]
port 309 nsew signal input
flabel metal2 s 12346 44540 12402 45000 0 FreeSans 224 90 0 0 S2MID[6]
port 310 nsew signal input
flabel metal2 s 12530 44540 12586 45000 0 FreeSans 224 90 0 0 S2MID[7]
port 311 nsew signal input
flabel metal2 s 12714 -300 12770 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 312 nsew signal tristate
flabel metal2 s 14554 -300 14610 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 313 nsew signal tristate
flabel metal2 s 14738 -300 14794 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 314 nsew signal tristate
flabel metal2 s 14922 -300 14978 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 315 nsew signal tristate
flabel metal2 s 15106 -300 15162 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 316 nsew signal tristate
flabel metal2 s 15290 -300 15346 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 317 nsew signal tristate
flabel metal2 s 15474 -300 15530 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 318 nsew signal tristate
flabel metal2 s 12898 -300 12954 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 319 nsew signal tristate
flabel metal2 s 13082 -300 13138 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 320 nsew signal tristate
flabel metal2 s 13266 -300 13322 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 321 nsew signal tristate
flabel metal2 s 13450 -300 13506 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 322 nsew signal tristate
flabel metal2 s 13634 -300 13690 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 323 nsew signal tristate
flabel metal2 s 13818 -300 13874 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 324 nsew signal tristate
flabel metal2 s 14002 -300 14058 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 325 nsew signal tristate
flabel metal2 s 14186 -300 14242 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 326 nsew signal tristate
flabel metal2 s 14370 -300 14426 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 327 nsew signal tristate
flabel metal2 s 12714 44540 12770 45000 0 FreeSans 224 90 0 0 S4END[0]
port 328 nsew signal input
flabel metal2 s 14554 44540 14610 45000 0 FreeSans 224 90 0 0 S4END[10]
port 329 nsew signal input
flabel metal2 s 14738 44540 14794 45000 0 FreeSans 224 90 0 0 S4END[11]
port 330 nsew signal input
flabel metal2 s 14922 44540 14978 45000 0 FreeSans 224 90 0 0 S4END[12]
port 331 nsew signal input
flabel metal2 s 15106 44540 15162 45000 0 FreeSans 224 90 0 0 S4END[13]
port 332 nsew signal input
flabel metal2 s 15290 44540 15346 45000 0 FreeSans 224 90 0 0 S4END[14]
port 333 nsew signal input
flabel metal2 s 15474 44540 15530 45000 0 FreeSans 224 90 0 0 S4END[15]
port 334 nsew signal input
flabel metal2 s 12898 44540 12954 45000 0 FreeSans 224 90 0 0 S4END[1]
port 335 nsew signal input
flabel metal2 s 13082 44540 13138 45000 0 FreeSans 224 90 0 0 S4END[2]
port 336 nsew signal input
flabel metal2 s 13266 44540 13322 45000 0 FreeSans 224 90 0 0 S4END[3]
port 337 nsew signal input
flabel metal2 s 13450 44540 13506 45000 0 FreeSans 224 90 0 0 S4END[4]
port 338 nsew signal input
flabel metal2 s 13634 44540 13690 45000 0 FreeSans 224 90 0 0 S4END[5]
port 339 nsew signal input
flabel metal2 s 13818 44540 13874 45000 0 FreeSans 224 90 0 0 S4END[6]
port 340 nsew signal input
flabel metal2 s 14002 44540 14058 45000 0 FreeSans 224 90 0 0 S4END[7]
port 341 nsew signal input
flabel metal2 s 14186 44540 14242 45000 0 FreeSans 224 90 0 0 S4END[8]
port 342 nsew signal input
flabel metal2 s 14370 44540 14426 45000 0 FreeSans 224 90 0 0 S4END[9]
port 343 nsew signal input
flabel metal2 s 15658 -300 15714 160 0 FreeSans 224 90 0 0 UserCLK
port 344 nsew signal input
flabel metal2 s 15658 44540 15714 45000 0 FreeSans 224 90 0 0 UserCLKo
port 345 nsew signal tristate
flabel metal4 s 5888 1040 6208 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 10833 1040 11153 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 15778 1040 16098 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 20723 1040 21043 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 3416 1040 3736 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 8361 1040 8681 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 13306 1040 13626 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 18251 1040 18571 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal3 s -300 4904 160 5024 0 FreeSans 480 0 0 0 W1BEG[0]
port 348 nsew signal tristate
flabel metal3 s -300 5176 160 5296 0 FreeSans 480 0 0 0 W1BEG[1]
port 349 nsew signal tristate
flabel metal3 s -300 5448 160 5568 0 FreeSans 480 0 0 0 W1BEG[2]
port 350 nsew signal tristate
flabel metal3 s -300 5720 160 5840 0 FreeSans 480 0 0 0 W1BEG[3]
port 351 nsew signal tristate
flabel metal3 s -300 5992 160 6112 0 FreeSans 480 0 0 0 W2BEG[0]
port 352 nsew signal tristate
flabel metal3 s -300 6264 160 6384 0 FreeSans 480 0 0 0 W2BEG[1]
port 353 nsew signal tristate
flabel metal3 s -300 6536 160 6656 0 FreeSans 480 0 0 0 W2BEG[2]
port 354 nsew signal tristate
flabel metal3 s -300 6808 160 6928 0 FreeSans 480 0 0 0 W2BEG[3]
port 355 nsew signal tristate
flabel metal3 s -300 7080 160 7200 0 FreeSans 480 0 0 0 W2BEG[4]
port 356 nsew signal tristate
flabel metal3 s -300 7352 160 7472 0 FreeSans 480 0 0 0 W2BEG[5]
port 357 nsew signal tristate
flabel metal3 s -300 7624 160 7744 0 FreeSans 480 0 0 0 W2BEG[6]
port 358 nsew signal tristate
flabel metal3 s -300 7896 160 8016 0 FreeSans 480 0 0 0 W2BEG[7]
port 359 nsew signal tristate
flabel metal3 s -300 8168 160 8288 0 FreeSans 480 0 0 0 W2BEGb[0]
port 360 nsew signal tristate
flabel metal3 s -300 8440 160 8560 0 FreeSans 480 0 0 0 W2BEGb[1]
port 361 nsew signal tristate
flabel metal3 s -300 8712 160 8832 0 FreeSans 480 0 0 0 W2BEGb[2]
port 362 nsew signal tristate
flabel metal3 s -300 8984 160 9104 0 FreeSans 480 0 0 0 W2BEGb[3]
port 363 nsew signal tristate
flabel metal3 s -300 9256 160 9376 0 FreeSans 480 0 0 0 W2BEGb[4]
port 364 nsew signal tristate
flabel metal3 s -300 9528 160 9648 0 FreeSans 480 0 0 0 W2BEGb[5]
port 365 nsew signal tristate
flabel metal3 s -300 9800 160 9920 0 FreeSans 480 0 0 0 W2BEGb[6]
port 366 nsew signal tristate
flabel metal3 s -300 10072 160 10192 0 FreeSans 480 0 0 0 W2BEGb[7]
port 367 nsew signal tristate
flabel metal3 s -300 14696 160 14816 0 FreeSans 480 0 0 0 W6BEG[0]
port 368 nsew signal tristate
flabel metal3 s -300 17416 160 17536 0 FreeSans 480 0 0 0 W6BEG[10]
port 369 nsew signal tristate
flabel metal3 s -300 17688 160 17808 0 FreeSans 480 0 0 0 W6BEG[11]
port 370 nsew signal tristate
flabel metal3 s -300 14968 160 15088 0 FreeSans 480 0 0 0 W6BEG[1]
port 371 nsew signal tristate
flabel metal3 s -300 15240 160 15360 0 FreeSans 480 0 0 0 W6BEG[2]
port 372 nsew signal tristate
flabel metal3 s -300 15512 160 15632 0 FreeSans 480 0 0 0 W6BEG[3]
port 373 nsew signal tristate
flabel metal3 s -300 15784 160 15904 0 FreeSans 480 0 0 0 W6BEG[4]
port 374 nsew signal tristate
flabel metal3 s -300 16056 160 16176 0 FreeSans 480 0 0 0 W6BEG[5]
port 375 nsew signal tristate
flabel metal3 s -300 16328 160 16448 0 FreeSans 480 0 0 0 W6BEG[6]
port 376 nsew signal tristate
flabel metal3 s -300 16600 160 16720 0 FreeSans 480 0 0 0 W6BEG[7]
port 377 nsew signal tristate
flabel metal3 s -300 16872 160 16992 0 FreeSans 480 0 0 0 W6BEG[8]
port 378 nsew signal tristate
flabel metal3 s -300 17144 160 17264 0 FreeSans 480 0 0 0 W6BEG[9]
port 379 nsew signal tristate
flabel metal3 s -300 10344 160 10464 0 FreeSans 480 0 0 0 WW4BEG[0]
port 380 nsew signal tristate
flabel metal3 s -300 13064 160 13184 0 FreeSans 480 0 0 0 WW4BEG[10]
port 381 nsew signal tristate
flabel metal3 s -300 13336 160 13456 0 FreeSans 480 0 0 0 WW4BEG[11]
port 382 nsew signal tristate
flabel metal3 s -300 13608 160 13728 0 FreeSans 480 0 0 0 WW4BEG[12]
port 383 nsew signal tristate
flabel metal3 s -300 13880 160 14000 0 FreeSans 480 0 0 0 WW4BEG[13]
port 384 nsew signal tristate
flabel metal3 s -300 14152 160 14272 0 FreeSans 480 0 0 0 WW4BEG[14]
port 385 nsew signal tristate
flabel metal3 s -300 14424 160 14544 0 FreeSans 480 0 0 0 WW4BEG[15]
port 386 nsew signal tristate
flabel metal3 s -300 10616 160 10736 0 FreeSans 480 0 0 0 WW4BEG[1]
port 387 nsew signal tristate
flabel metal3 s -300 10888 160 11008 0 FreeSans 480 0 0 0 WW4BEG[2]
port 388 nsew signal tristate
flabel metal3 s -300 11160 160 11280 0 FreeSans 480 0 0 0 WW4BEG[3]
port 389 nsew signal tristate
flabel metal3 s -300 11432 160 11552 0 FreeSans 480 0 0 0 WW4BEG[4]
port 390 nsew signal tristate
flabel metal3 s -300 11704 160 11824 0 FreeSans 480 0 0 0 WW4BEG[5]
port 391 nsew signal tristate
flabel metal3 s -300 11976 160 12096 0 FreeSans 480 0 0 0 WW4BEG[6]
port 392 nsew signal tristate
flabel metal3 s -300 12248 160 12368 0 FreeSans 480 0 0 0 WW4BEG[7]
port 393 nsew signal tristate
flabel metal3 s -300 12520 160 12640 0 FreeSans 480 0 0 0 WW4BEG[8]
port 394 nsew signal tristate
flabel metal3 s -300 12792 160 12912 0 FreeSans 480 0 0 0 WW4BEG[9]
port 395 nsew signal tristate
rlabel via1 11073 43520 11073 43520 0 VGND
rlabel metal1 10994 42976 10994 42976 0 VPWR
rlabel metal1 19688 9146 19688 9146 0 Config_accessC_bit0
rlabel metal1 18676 9486 18676 9486 0 Config_accessC_bit1
rlabel metal1 20516 7514 20516 7514 0 Config_accessC_bit2
rlabel metal3 21594 10948 21594 10948 0 Config_accessC_bit3
rlabel metal3 820 18020 820 18020 0 E1END[0]
rlabel metal3 682 18292 682 18292 0 E1END[1]
rlabel metal3 452 18564 452 18564 0 E1END[2]
rlabel metal3 452 18836 452 18836 0 E1END[3]
rlabel metal3 1050 21284 1050 21284 0 E2END[0]
rlabel metal3 544 21556 544 21556 0 E2END[1]
rlabel metal3 498 21828 498 21828 0 E2END[2]
rlabel metal3 774 22100 774 22100 0 E2END[3]
rlabel metal3 452 22372 452 22372 0 E2END[4]
rlabel metal3 774 22644 774 22644 0 E2END[5]
rlabel metal3 452 22916 452 22916 0 E2END[6]
rlabel metal3 912 23188 912 23188 0 E2END[7]
rlabel metal3 1027 19108 1027 19108 0 E2MID[0]
rlabel metal3 682 19380 682 19380 0 E2MID[1]
rlabel metal3 751 19652 751 19652 0 E2MID[2]
rlabel metal3 1004 19924 1004 19924 0 E2MID[3]
rlabel metal3 1441 20196 1441 20196 0 E2MID[4]
rlabel metal3 452 20468 452 20468 0 E2MID[5]
rlabel metal3 1441 20740 1441 20740 0 E2MID[6]
rlabel metal3 636 21012 636 21012 0 E2MID[7]
rlabel metal3 728 27812 728 27812 0 E6END[0]
rlabel metal3 1464 30532 1464 30532 0 E6END[10]
rlabel metal1 3358 32878 3358 32878 0 E6END[11]
rlabel metal2 3818 28577 3818 28577 0 E6END[1]
rlabel metal2 4646 27897 4646 27897 0 E6END[2]
rlabel metal3 820 28628 820 28628 0 E6END[3]
rlabel metal3 452 28900 452 28900 0 E6END[4]
rlabel metal3 866 29172 866 29172 0 E6END[5]
rlabel metal3 360 29444 360 29444 0 E6END[6]
rlabel metal3 682 29716 682 29716 0 E6END[7]
rlabel metal3 935 29988 935 29988 0 E6END[8]
rlabel metal2 3450 30481 3450 30481 0 E6END[9]
rlabel metal3 452 23460 452 23460 0 EE4END[0]
rlabel via2 3634 26197 3634 26197 0 EE4END[10]
rlabel metal3 682 26452 682 26452 0 EE4END[11]
rlabel metal3 728 26724 728 26724 0 EE4END[12]
rlabel metal3 636 26996 636 26996 0 EE4END[13]
rlabel metal3 728 27268 728 27268 0 EE4END[14]
rlabel metal2 3266 28033 3266 28033 0 EE4END[15]
rlabel metal3 728 23732 728 23732 0 EE4END[1]
rlabel metal3 406 24004 406 24004 0 EE4END[2]
rlabel metal3 682 24276 682 24276 0 EE4END[3]
rlabel metal3 728 24548 728 24548 0 EE4END[4]
rlabel metal3 452 24820 452 24820 0 EE4END[5]
rlabel metal3 728 25092 728 25092 0 EE4END[6]
rlabel metal3 682 25364 682 25364 0 EE4END[7]
rlabel metal3 452 25636 452 25636 0 EE4END[8]
rlabel metal2 3174 26129 3174 26129 0 EE4END[9]
rlabel metal3 21180 15844 21180 15844 0 FAB2RAM_A0_O0
rlabel metal3 21571 16388 21571 16388 0 FAB2RAM_A0_O1
rlabel metal3 21410 16932 21410 16932 0 FAB2RAM_A0_O2
rlabel metal1 20884 17306 20884 17306 0 FAB2RAM_A0_O3
rlabel metal3 20720 13668 20720 13668 0 FAB2RAM_A1_O0
rlabel metal1 20884 14042 20884 14042 0 FAB2RAM_A1_O1
rlabel metal3 21180 14756 21180 14756 0 FAB2RAM_A1_O2
rlabel metal3 21594 15300 21594 15300 0 FAB2RAM_A1_O3
rlabel metal2 19366 12517 19366 12517 0 FAB2RAM_C_O0
rlabel metal3 21571 12036 21571 12036 0 FAB2RAM_C_O1
rlabel metal3 20490 12580 20490 12580 0 FAB2RAM_C_O2
rlabel metal1 20884 12954 20884 12954 0 FAB2RAM_C_O3
rlabel metal3 21088 24548 21088 24548 0 FAB2RAM_D0_O0
rlabel metal3 21571 25092 21571 25092 0 FAB2RAM_D0_O1
rlabel metal3 20904 25636 20904 25636 0 FAB2RAM_D0_O2
rlabel metal3 21594 26180 21594 26180 0 FAB2RAM_D0_O3
rlabel metal3 21180 22372 21180 22372 0 FAB2RAM_D1_O0
rlabel metal3 21594 22916 21594 22916 0 FAB2RAM_D1_O1
rlabel metal3 21180 23460 21180 23460 0 FAB2RAM_D1_O2
rlabel metal3 21571 24004 21571 24004 0 FAB2RAM_D1_O3
rlabel metal3 21732 20196 21732 20196 0 FAB2RAM_D2_O0
rlabel metal3 21594 20740 21594 20740 0 FAB2RAM_D2_O1
rlabel metal3 20904 21284 20904 21284 0 FAB2RAM_D2_O2
rlabel metal1 20884 21658 20884 21658 0 FAB2RAM_D2_O3
rlabel metal3 21456 18020 21456 18020 0 FAB2RAM_D3_O0
rlabel metal3 21594 18564 21594 18564 0 FAB2RAM_D3_O1
rlabel metal3 20996 19108 20996 19108 0 FAB2RAM_D3_O2
rlabel metal1 21022 18870 21022 18870 0 FAB2RAM_D3_O3
rlabel metal1 1472 30294 1472 30294 0 FrameData[0]
rlabel metal2 2806 34425 2806 34425 0 FrameData[10]
rlabel metal2 3358 34323 3358 34323 0 FrameData[11]
rlabel metal3 1441 34340 1441 34340 0 FrameData[12]
rlabel metal3 475 34612 475 34612 0 FrameData[13]
rlabel metal3 1050 34884 1050 34884 0 FrameData[14]
rlabel metal3 2200 35156 2200 35156 0 FrameData[15]
rlabel metal3 774 35428 774 35428 0 FrameData[16]
rlabel metal3 682 35700 682 35700 0 FrameData[17]
rlabel metal3 682 35972 682 35972 0 FrameData[18]
rlabel metal3 728 36244 728 36244 0 FrameData[19]
rlabel metal3 452 31348 452 31348 0 FrameData[1]
rlabel metal3 475 36516 475 36516 0 FrameData[20]
rlabel metal3 682 36788 682 36788 0 FrameData[21]
rlabel metal3 728 37060 728 37060 0 FrameData[22]
rlabel metal3 820 37332 820 37332 0 FrameData[23]
rlabel metal3 1050 37604 1050 37604 0 FrameData[24]
rlabel metal3 774 37876 774 37876 0 FrameData[25]
rlabel metal3 475 38148 475 38148 0 FrameData[26]
rlabel metal2 3082 39219 3082 39219 0 FrameData[27]
rlabel metal2 2806 39899 2806 39899 0 FrameData[28]
rlabel metal3 1050 38964 1050 38964 0 FrameData[29]
rlabel metal3 1104 31756 1104 31756 0 FrameData[2]
rlabel metal3 728 39236 728 39236 0 FrameData[30]
rlabel metal3 199 39508 199 39508 0 FrameData[31]
rlabel metal3 452 31892 452 31892 0 FrameData[3]
rlabel metal3 728 32164 728 32164 0 FrameData[4]
rlabel metal3 774 32436 774 32436 0 FrameData[5]
rlabel metal2 2806 33099 2806 33099 0 FrameData[6]
rlabel metal3 475 32980 475 32980 0 FrameData[7]
rlabel metal3 1050 33252 1050 33252 0 FrameData[8]
rlabel metal3 728 33524 728 33524 0 FrameData[9]
rlabel metal3 21226 26724 21226 26724 0 FrameData_O[0]
rlabel metal3 21226 32164 21226 32164 0 FrameData_O[10]
rlabel metal3 21594 32708 21594 32708 0 FrameData_O[11]
rlabel metal3 21180 33252 21180 33252 0 FrameData_O[12]
rlabel metal3 21548 33796 21548 33796 0 FrameData_O[13]
rlabel metal3 21180 34340 21180 34340 0 FrameData_O[14]
rlabel metal3 21594 34884 21594 34884 0 FrameData_O[15]
rlabel metal1 20332 35258 20332 35258 0 FrameData_O[16]
rlabel metal3 21594 35972 21594 35972 0 FrameData_O[17]
rlabel metal3 20858 36516 20858 36516 0 FrameData_O[18]
rlabel metal3 21571 37060 21571 37060 0 FrameData_O[19]
rlabel metal3 21594 27268 21594 27268 0 FrameData_O[1]
rlabel metal3 21180 37604 21180 37604 0 FrameData_O[20]
rlabel metal3 21594 38148 21594 38148 0 FrameData_O[21]
rlabel metal3 21180 38692 21180 38692 0 FrameData_O[22]
rlabel metal3 21594 39236 21594 39236 0 FrameData_O[23]
rlabel metal3 21456 39780 21456 39780 0 FrameData_O[24]
rlabel metal3 21594 40324 21594 40324 0 FrameData_O[25]
rlabel metal3 21226 40868 21226 40868 0 FrameData_O[26]
rlabel metal3 21594 41412 21594 41412 0 FrameData_O[27]
rlabel metal3 20628 41956 20628 41956 0 FrameData_O[28]
rlabel metal3 21594 42500 21594 42500 0 FrameData_O[29]
rlabel metal3 21180 27812 21180 27812 0 FrameData_O[2]
rlabel metal1 19964 42874 19964 42874 0 FrameData_O[30]
rlabel metal1 20746 42330 20746 42330 0 FrameData_O[31]
rlabel metal3 21571 28356 21571 28356 0 FrameData_O[3]
rlabel metal3 21180 28900 21180 28900 0 FrameData_O[4]
rlabel metal3 21594 29444 21594 29444 0 FrameData_O[5]
rlabel metal3 21180 29988 21180 29988 0 FrameData_O[6]
rlabel metal3 21594 30532 21594 30532 0 FrameData_O[7]
rlabel metal3 21180 31076 21180 31076 0 FrameData_O[8]
rlabel metal3 21548 31620 21548 31620 0 FrameData_O[9]
rlabel metal2 15923 68 15923 68 0 FrameStrobe[0]
rlabel metal2 17710 1421 17710 1421 0 FrameStrobe[10]
rlabel metal2 17894 330 17894 330 0 FrameStrobe[11]
rlabel metal2 18078 126 18078 126 0 FrameStrobe[12]
rlabel metal2 18262 262 18262 262 0 FrameStrobe[13]
rlabel metal2 18446 483 18446 483 0 FrameStrobe[14]
rlabel metal2 18577 68 18577 68 0 FrameStrobe[15]
rlabel metal2 18814 211 18814 211 0 FrameStrobe[16]
rlabel metal2 18998 551 18998 551 0 FrameStrobe[17]
rlabel metal2 19182 160 19182 160 0 FrameStrobe[18]
rlabel metal1 12650 4148 12650 4148 0 FrameStrobe[19]
rlabel metal1 15916 1326 15916 1326 0 FrameStrobe[1]
rlabel metal2 16238 500 16238 500 0 FrameStrobe[2]
rlabel metal2 16422 398 16422 398 0 FrameStrobe[3]
rlabel metal2 16659 68 16659 68 0 FrameStrobe[4]
rlabel metal2 16843 68 16843 68 0 FrameStrobe[5]
rlabel metal2 17027 68 17027 68 0 FrameStrobe[6]
rlabel viali 14583 1326 14583 1326 0 FrameStrobe[7]
rlabel metal2 17342 738 17342 738 0 FrameStrobe[8]
rlabel metal1 15916 1938 15916 1938 0 FrameStrobe[9]
rlabel metal1 16008 43418 16008 43418 0 FrameStrobe_O[0]
rlabel metal2 17710 44261 17710 44261 0 FrameStrobe_O[10]
rlabel metal2 17894 43632 17894 43632 0 FrameStrobe_O[11]
rlabel metal2 18078 43802 18078 43802 0 FrameStrobe_O[12]
rlabel metal2 18262 43853 18262 43853 0 FrameStrobe_O[13]
rlabel metal1 19780 41242 19780 41242 0 FrameStrobe_O[14]
rlabel metal1 17526 43214 17526 43214 0 FrameStrobe_O[15]
rlabel metal1 18630 41786 18630 41786 0 FrameStrobe_O[16]
rlabel metal1 18078 42296 18078 42296 0 FrameStrobe_O[17]
rlabel metal1 18308 41990 18308 41990 0 FrameStrobe_O[18]
rlabel metal1 19228 41786 19228 41786 0 FrameStrobe_O[19]
rlabel metal2 16054 44261 16054 44261 0 FrameStrobe_O[1]
rlabel metal2 16238 44329 16238 44329 0 FrameStrobe_O[2]
rlabel metal2 16422 44057 16422 44057 0 FrameStrobe_O[3]
rlabel metal1 17296 43078 17296 43078 0 FrameStrobe_O[4]
rlabel metal2 16790 43632 16790 43632 0 FrameStrobe_O[5]
rlabel metal1 17940 43146 17940 43146 0 FrameStrobe_O[6]
rlabel metal2 17158 44057 17158 44057 0 FrameStrobe_O[7]
rlabel metal2 17342 44193 17342 44193 0 FrameStrobe_O[8]
rlabel metal2 17526 44057 17526 44057 0 FrameStrobe_O[9]
rlabel metal1 20194 9078 20194 9078 0 Inst_Config_accessConfig_access.ConfigBits\[0\]
rlabel metal1 19458 9690 19458 9690 0 Inst_Config_accessConfig_access.ConfigBits\[1\]
rlabel metal1 19596 10234 19596 10234 0 Inst_Config_accessConfig_access.ConfigBits\[2\]
rlabel metal1 19872 14858 19872 14858 0 Inst_Config_accessConfig_access.ConfigBits\[3\]
rlabel metal1 18262 16048 18262 16048 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 19734 16388 19734 16388 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal2 20286 18598 20286 18598 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 14766 36074 14766 36074 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 16146 16524 16146 16524 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 18298 17170 18298 17170 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 16866 18326 16866 18326 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 13892 36142 13892 36142 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 18216 16558 18216 16558 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 20010 15504 20010 15504 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 19734 18394 19734 18394 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 15548 35666 15548 35666 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 17894 16592 17894 16592 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18630 16524 18630 16524 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 18354 16116 18354 16116 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 18538 16116 18538 16116 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 19366 16592 19366 16592 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 19780 15470 19780 15470 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 19642 16626 19642 16626 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 19642 16184 19642 16184 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 19274 18700 19274 18700 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 19090 17680 19090 17680 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 19872 18938 19872 18938 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19780 17578 19780 17578 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 14122 35666 14122 35666 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal2 15410 36278 15410 36278 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 14766 35666 14766 35666 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 15272 35734 15272 35734 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 19918 13906 19918 13906 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 18446 12818 18446 12818 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18538 21522 18538 21522 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 17848 26758 17848 26758 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal3 14283 20740 14283 20740 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 18487 11798 18487 11798 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 16698 21964 16698 21964 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 16141 26962 16141 26962 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[3\]
rlabel viali 19089 13310 19089 13310 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 18584 15130 18584 15130 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 18584 21998 18584 21998 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 17296 26350 17296 26350 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19090 14586 19090 14586 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18952 13498 18952 13498 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19596 13770 19596 13770 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19826 13838 19826 13838 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20654 14586 20654 14586 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 13938 12240 13938 12240 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 19136 12682 19136 12682 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 18446 12954 18446 12954 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 17388 21862 17388 21862 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 18906 21862 18906 21862 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18814 21556 18814 21556 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19090 21454 19090 21454 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 16836 27098 16836 27098 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 17894 26316 17894 26316 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 18446 26996 18446 26996 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 17940 26214 17940 26214 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 18860 15402 18860 15402 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20194 36278 20194 36278 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18308 13498 18308 13498 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 18216 14382 18216 14382 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal2 16836 13668 16836 13668 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 17107 36822 17107 36822 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 16872 13906 16872 13906 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 16146 15062 16146 15062 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 18584 10030 18584 10030 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 19688 36890 19688 36890 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[1\]
rlabel metal2 19044 12886 19044 12886 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 18216 13906 18216 13906 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 17894 12172 17894 12172 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal3 18791 15164 18791 15164 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 18354 11900 18354 11900 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal2 18860 15334 18860 15334 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 19412 37978 19412 37978 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 20010 38284 20010 38284 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 19918 35700 19918 35700 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 20148 35734 20148 35734 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 17204 12954 17204 12954 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 18676 13804 18676 13804 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18308 12410 18308 12410 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal2 18354 13073 18354 13073 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18538 14382 18538 14382 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 18216 13702 18216 13702 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 18538 14314 18538 14314 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 18584 14450 18584 14450 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 18814 24208 18814 24208 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 17066 35462 17066 35462 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal2 16790 26180 16790 26180 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19918 28560 19918 28560 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 15962 24174 15962 24174 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 15624 36074 15624 36074 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 14980 26282 14980 26282 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 17884 28526 17884 28526 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 18722 24140 18722 24140 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 17894 36108 17894 36108 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 16790 25262 16790 25262 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 18998 28730 18998 28730 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 18124 24174 18124 24174 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18952 24174 18952 24174 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 18170 24310 18170 24310 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel viali 18170 24246 18170 24246 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 16790 35802 16790 35802 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 17664 35666 17664 35666 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 17204 35598 17204 35598 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 17434 35598 17434 35598 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 15962 25908 15962 25908 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 16928 25466 16928 25466 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 16192 25670 16192 25670 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 16468 25806 16468 25806 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal2 19274 28900 19274 28900 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19918 30158 19918 30158 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 19826 28730 19826 28730 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20148 28594 20148 28594 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 18170 22678 18170 22678 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 19458 33524 19458 33524 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19734 23766 19734 23766 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 17618 27642 17618 27642 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18906 23086 18906 23086 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 6716 31994 6716 31994 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 18223 24854 18223 24854 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[2\]
rlabel via1 16330 28050 16330 28050 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 19458 22406 19458 22406 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 18952 32538 18952 32538 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 19274 23732 19274 23732 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 18078 27506 18078 27506 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19366 23018 19366 23018 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18768 22202 18768 22202 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19642 23154 19642 23154 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 18446 22678 18446 22678 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal2 18722 31484 18722 31484 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal2 19642 33796 19642 33796 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 18768 31110 18768 31110 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 19550 32980 19550 32980 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 19366 24412 19366 24412 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 18722 23120 18722 23120 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 19642 23494 19642 23494 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 18676 23290 18676 23290 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18078 28084 18078 28084 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 17848 27438 17848 27438 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 17572 27574 17572 27574 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 17618 27506 17618 27506 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 17848 38318 17848 38318 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 15226 37876 15226 37876 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18630 26316 18630 26316 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 18170 30022 18170 30022 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 15308 38930 15308 38930 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 13892 38318 13892 38318 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 18998 26350 18998 26350 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 16514 30260 16514 30260 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 17526 38964 17526 38964 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 15640 38318 15640 38318 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 18354 25908 18354 25908 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 17940 30362 17940 30362 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 16790 38284 16790 38284 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 18170 38556 18170 38556 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 17526 38352 17526 38352 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 17986 38250 17986 38250 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 14122 37842 14122 37842 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 15640 37842 15640 37842 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 14812 37842 14812 37842 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 15410 37808 15410 37808 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 19458 26384 19458 26384 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 18492 26010 18492 26010 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 19550 26452 19550 26452 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 20562 26486 20562 26486 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal2 16330 30498 16330 30498 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 18722 30260 18722 30260 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 18032 30158 18032 30158 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 18538 30158 18538 30158 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 18170 19346 18170 19346 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20010 31314 20010 31314 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19872 20434 19872 20434 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 18814 34612 18814 34612 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 16918 20434 16918 20434 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 19080 32402 19080 32402 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 19550 21556 19550 21556 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 16836 33966 16836 33966 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 17940 19822 17940 19822 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 20102 32266 20102 32266 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 19090 19924 19090 19924 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 18538 34578 18538 34578 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 17526 19788 17526 19788 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18906 19380 18906 19380 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 18032 19278 18032 19278 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 18722 19278 18722 19278 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel viali 19182 31319 19182 31319 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 18584 31314 18584 31314 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 19596 31178 19596 31178 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 20010 31450 20010 31450 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 18630 20944 18630 20944 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 18952 20026 18952 20026 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 20194 20468 20194 20468 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 20056 20366 20056 20366 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 17526 33932 17526 33932 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 18998 34510 18998 34510 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 17618 34272 17618 34272 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 18676 34510 18676 34510 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 16376 6290 16376 6290 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 17526 7956 17526 7956 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19504 7922 19504 7922 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19090 9894 19090 9894 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 11500 7310 11500 7310 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
rlabel metal2 18906 8517 18906 8517 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
rlabel metal1 20010 7990 20010 7990 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
rlabel metal1 14398 16490 14398 16490 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
rlabel metal2 17802 5678 17802 5678 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 17986 7752 17986 7752 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[1\]
rlabel metal2 17434 8500 17434 8500 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[2\]
rlabel metal2 18170 8806 18170 8806 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 19090 4148 19090 4148 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 18078 3944 18078 3944 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 18170 5083 18170 5083 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 16468 5678 16468 5678 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 16192 8058 16192 8058 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 15916 8058 15916 8058 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 18308 7854 18308 7854 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 18814 7888 18814 7888 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 15778 8500 15778 8500 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 11362 6256 11362 6256 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18897 8976 18897 8976 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 11868 6086 11868 6086 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 16744 8942 16744 8942 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 17296 8602 17296 8602 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 17066 9146 17066 9146 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal2 20194 10659 20194 10659 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 17204 4658 17204 4658 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 17388 6086 17388 6086 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel via2 17802 10421 17802 10421 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 19688 7378 19688 7378 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 17480 4726 17480 4726 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
rlabel metal2 5290 7667 5290 7667 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
rlabel metal2 18078 7973 18078 7973 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
rlabel metal2 19826 11067 19826 11067 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
rlabel metal1 13110 4624 13110 4624 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 12834 5236 12834 5236 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 18745 7514 18745 7514 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[2\]
rlabel metal2 16422 7344 16422 7344 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 13478 5066 13478 5066 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 12650 4590 12650 4590 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 17112 4590 17112 4590 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 17894 4522 17894 4522 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 12190 5338 12190 5338 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 11914 5168 11914 5168 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 12696 5882 12696 5882 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 17802 6902 17802 6902 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 11546 4488 11546 4488 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 10810 4148 10810 4148 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 19274 8296 19274 8296 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal2 10718 3621 10718 3621 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 15870 8874 15870 8874 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal2 17158 7854 17158 7854 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 18722 10438 18722 10438 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20056 7514 20056 7514 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 15502 7582 15502 7582 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 15042 4624 15042 4624 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 15870 6630 15870 6630 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 18676 6290 18676 6290 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 15548 7242 15548 7242 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\]
rlabel metal1 4278 5134 4278 5134 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\]
rlabel metal3 15548 5372 15548 5372 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\]
rlabel metal1 18262 6766 18262 6766 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\]
rlabel metal2 15962 6426 15962 6426 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 15824 3978 15824 3978 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[1\]
rlabel metal2 10258 3995 10258 3995 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 13662 4148 13662 4148 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 15180 5338 15180 5338 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 16146 7684 16146 7684 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 15686 7412 15686 7412 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 15916 7378 15916 7378 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 15870 3638 15870 3638 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 15276 4590 15276 4590 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 14306 4658 14306 4658 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 14766 4522 14766 4522 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 20470 1431 20470 1431 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal3 15502 6664 15502 6664 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 20470 5236 20470 5236 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 16420 5270 16420 5270 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel via1 11190 4250 11190 4250 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 13616 4250 13616 4250 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 12236 4658 12236 4658 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 18676 6358 18676 6358 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 14490 2992 14490 2992 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 17342 3638 17342 3638 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 18078 3910 18078 3910 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 13754 5950 13754 5950 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 14030 9554 14030 9554 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\]
rlabel metal3 12374 1496 12374 1496 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\]
rlabel metal2 14306 544 14306 544 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\]
rlabel metal3 10833 7004 10833 7004 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\]
rlabel metal1 15548 2278 15548 2278 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 12642 3060 12642 3060 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 20102 2856 20102 2856 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 16698 5202 16698 5202 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 11270 3468 11270 3468 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 11362 3706 11362 3706 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 14573 3026 14573 3026 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 15042 3128 15042 3128 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 12556 3026 12556 3026 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal2 10902 2516 10902 2516 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal4 15732 544 15732 544 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 18492 3502 18492 3502 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 13800 3026 13800 3026 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 13386 3094 13386 3094 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal3 16100 2720 16100 2720 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 13156 2890 13156 2890 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 13202 4760 13202 4760 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 14077 4590 14077 4590 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 13570 5644 13570 5644 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal2 13846 5083 13846 5083 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 11829 22066 11829 22066 0 Inst_RAM_IO_ConfigMem.ConfigBits\[100\]
rlabel metal1 10948 21998 10948 21998 0 Inst_RAM_IO_ConfigMem.ConfigBits\[101\]
rlabel metal1 8372 21114 8372 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[102\]
rlabel metal1 9522 21114 9522 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[103\]
rlabel metal1 2530 25847 2530 25847 0 Inst_RAM_IO_ConfigMem.ConfigBits\[104\]
rlabel metal1 2530 25466 2530 25466 0 Inst_RAM_IO_ConfigMem.ConfigBits\[105\]
rlabel metal2 11086 26588 11086 26588 0 Inst_RAM_IO_ConfigMem.ConfigBits\[106\]
rlabel metal1 11086 26316 11086 26316 0 Inst_RAM_IO_ConfigMem.ConfigBits\[107\]
rlabel metal1 14628 20978 14628 20978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[108\]
rlabel metal2 15318 20740 15318 20740 0 Inst_RAM_IO_ConfigMem.ConfigBits\[109\]
rlabel metal1 16376 20434 16376 20434 0 Inst_RAM_IO_ConfigMem.ConfigBits\[110\]
rlabel metal1 6486 23562 6486 23562 0 Inst_RAM_IO_ConfigMem.ConfigBits\[111\]
rlabel metal2 7590 23868 7590 23868 0 Inst_RAM_IO_ConfigMem.ConfigBits\[112\]
rlabel via1 9246 22474 9246 22474 0 Inst_RAM_IO_ConfigMem.ConfigBits\[113\]
rlabel metal1 5888 24310 5888 24310 0 Inst_RAM_IO_ConfigMem.ConfigBits\[114\]
rlabel metal1 7130 24922 7130 24922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[115\]
rlabel metal1 7222 25942 7222 25942 0 Inst_RAM_IO_ConfigMem.ConfigBits\[116\]
rlabel metal1 14812 32266 14812 32266 0 Inst_RAM_IO_ConfigMem.ConfigBits\[117\]
rlabel metal2 15318 33660 15318 33660 0 Inst_RAM_IO_ConfigMem.ConfigBits\[118\]
rlabel metal1 16652 31314 16652 31314 0 Inst_RAM_IO_ConfigMem.ConfigBits\[119\]
rlabel metal1 8970 14518 8970 14518 0 Inst_RAM_IO_ConfigMem.ConfigBits\[120\]
rlabel metal1 9108 15674 9108 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[121\]
rlabel metal1 5244 8602 5244 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[122\]
rlabel metal2 5566 9554 5566 9554 0 Inst_RAM_IO_ConfigMem.ConfigBits\[123\]
rlabel metal2 5014 6834 5014 6834 0 Inst_RAM_IO_ConfigMem.ConfigBits\[124\]
rlabel metal1 5612 6970 5612 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[125\]
rlabel metal1 12696 9078 12696 9078 0 Inst_RAM_IO_ConfigMem.ConfigBits\[126\]
rlabel metal1 13248 8330 13248 8330 0 Inst_RAM_IO_ConfigMem.ConfigBits\[127\]
rlabel metal1 12466 6426 12466 6426 0 Inst_RAM_IO_ConfigMem.ConfigBits\[128\]
rlabel metal1 13064 6970 13064 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[129\]
rlabel metal2 5382 4624 5382 4624 0 Inst_RAM_IO_ConfigMem.ConfigBits\[130\]
rlabel metal1 5612 5542 5612 5542 0 Inst_RAM_IO_ConfigMem.ConfigBits\[131\]
rlabel metal1 6992 5882 6992 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[132\]
rlabel via1 7497 6766 7497 6766 0 Inst_RAM_IO_ConfigMem.ConfigBits\[133\]
rlabel metal1 9798 9418 9798 9418 0 Inst_RAM_IO_ConfigMem.ConfigBits\[134\]
rlabel metal1 10902 9486 10902 9486 0 Inst_RAM_IO_ConfigMem.ConfigBits\[135\]
rlabel metal1 14812 9146 14812 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[136\]
rlabel metal1 16376 9146 16376 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[137\]
rlabel metal1 3174 5882 3174 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[138\]
rlabel metal2 3818 6460 3818 6460 0 Inst_RAM_IO_ConfigMem.ConfigBits\[139\]
rlabel metal1 2944 2618 2944 2618 0 Inst_RAM_IO_ConfigMem.ConfigBits\[140\]
rlabel metal1 3818 3162 3818 3162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[141\]
rlabel metal1 10764 5338 10764 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[142\]
rlabel metal2 11362 6324 11362 6324 0 Inst_RAM_IO_ConfigMem.ConfigBits\[143\]
rlabel metal2 12742 8449 12742 8449 0 Inst_RAM_IO_ConfigMem.ConfigBits\[144\]
rlabel metal1 13524 7922 13524 7922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[145\]
rlabel metal1 3036 8398 3036 8398 0 Inst_RAM_IO_ConfigMem.ConfigBits\[146\]
rlabel metal2 3726 8636 3726 8636 0 Inst_RAM_IO_ConfigMem.ConfigBits\[147\]
rlabel metal4 5428 8636 5428 8636 0 Inst_RAM_IO_ConfigMem.ConfigBits\[148\]
rlabel metal1 7774 9010 7774 9010 0 Inst_RAM_IO_ConfigMem.ConfigBits\[149\]
rlabel metal1 9844 10166 9844 10166 0 Inst_RAM_IO_ConfigMem.ConfigBits\[150\]
rlabel metal1 10810 8602 10810 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[151\]
rlabel metal2 15870 10370 15870 10370 0 Inst_RAM_IO_ConfigMem.ConfigBits\[152\]
rlabel metal1 15686 10098 15686 10098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[153\]
rlabel metal1 2898 7514 2898 7514 0 Inst_RAM_IO_ConfigMem.ConfigBits\[154\]
rlabel metal2 4186 8772 4186 8772 0 Inst_RAM_IO_ConfigMem.ConfigBits\[155\]
rlabel metal1 2760 5066 2760 5066 0 Inst_RAM_IO_ConfigMem.ConfigBits\[156\]
rlabel metal2 3358 4947 3358 4947 0 Inst_RAM_IO_ConfigMem.ConfigBits\[157\]
rlabel metal1 10810 7514 10810 7514 0 Inst_RAM_IO_ConfigMem.ConfigBits\[158\]
rlabel metal1 11408 8058 11408 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[159\]
rlabel metal1 14858 12376 14858 12376 0 Inst_RAM_IO_ConfigMem.ConfigBits\[160\]
rlabel metal1 16514 11016 16514 11016 0 Inst_RAM_IO_ConfigMem.ConfigBits\[161\]
rlabel metal1 2944 13838 2944 13838 0 Inst_RAM_IO_ConfigMem.ConfigBits\[162\]
rlabel metal1 3266 13498 3266 13498 0 Inst_RAM_IO_ConfigMem.ConfigBits\[163\]
rlabel metal1 6440 10778 6440 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[164\]
rlabel metal1 7038 10234 7038 10234 0 Inst_RAM_IO_ConfigMem.ConfigBits\[165\]
rlabel metal1 9614 10778 9614 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[166\]
rlabel metal1 10580 10778 10580 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[167\]
rlabel metal1 13708 10574 13708 10574 0 Inst_RAM_IO_ConfigMem.ConfigBits\[168\]
rlabel metal1 14950 10472 14950 10472 0 Inst_RAM_IO_ConfigMem.ConfigBits\[169\]
rlabel metal1 3726 11322 3726 11322 0 Inst_RAM_IO_ConfigMem.ConfigBits\[170\]
rlabel metal1 4646 11696 4646 11696 0 Inst_RAM_IO_ConfigMem.ConfigBits\[171\]
rlabel metal1 5934 12648 5934 12648 0 Inst_RAM_IO_ConfigMem.ConfigBits\[172\]
rlabel metal1 7774 13838 7774 13838 0 Inst_RAM_IO_ConfigMem.ConfigBits\[173\]
rlabel metal1 8970 12410 8970 12410 0 Inst_RAM_IO_ConfigMem.ConfigBits\[174\]
rlabel metal1 11086 11322 11086 11322 0 Inst_RAM_IO_ConfigMem.ConfigBits\[175\]
rlabel metal1 15870 11866 15870 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[176\]
rlabel metal1 15778 12750 15778 12750 0 Inst_RAM_IO_ConfigMem.ConfigBits\[177\]
rlabel metal2 4462 10982 4462 10982 0 Inst_RAM_IO_ConfigMem.ConfigBits\[178\]
rlabel metal1 4784 10778 4784 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[179\]
rlabel metal1 6716 11322 6716 11322 0 Inst_RAM_IO_ConfigMem.ConfigBits\[180\]
rlabel metal1 7497 13362 7497 13362 0 Inst_RAM_IO_ConfigMem.ConfigBits\[181\]
rlabel metal2 8326 13039 8326 13039 0 Inst_RAM_IO_ConfigMem.ConfigBits\[182\]
rlabel metal1 10856 11866 10856 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[183\]
rlabel metal2 14766 13838 14766 13838 0 Inst_RAM_IO_ConfigMem.ConfigBits\[184\]
rlabel metal1 15686 13362 15686 13362 0 Inst_RAM_IO_ConfigMem.ConfigBits\[185\]
rlabel metal2 3174 14654 3174 14654 0 Inst_RAM_IO_ConfigMem.ConfigBits\[186\]
rlabel metal1 5014 14416 5014 14416 0 Inst_RAM_IO_ConfigMem.ConfigBits\[187\]
rlabel metal1 7084 15946 7084 15946 0 Inst_RAM_IO_ConfigMem.ConfigBits\[188\]
rlabel metal1 7360 15674 7360 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[189\]
rlabel metal1 9292 14450 9292 14450 0 Inst_RAM_IO_ConfigMem.ConfigBits\[190\]
rlabel metal1 10120 12954 10120 12954 0 Inst_RAM_IO_ConfigMem.ConfigBits\[191\]
rlabel metal1 12328 17034 12328 17034 0 Inst_RAM_IO_ConfigMem.ConfigBits\[192\]
rlabel metal2 13110 17340 13110 17340 0 Inst_RAM_IO_ConfigMem.ConfigBits\[193\]
rlabel metal1 4738 29818 4738 29818 0 Inst_RAM_IO_ConfigMem.ConfigBits\[194\]
rlabel metal2 5198 30396 5198 30396 0 Inst_RAM_IO_ConfigMem.ConfigBits\[195\]
rlabel metal1 5612 18870 5612 18870 0 Inst_RAM_IO_ConfigMem.ConfigBits\[196\]
rlabel metal1 6716 16762 6716 16762 0 Inst_RAM_IO_ConfigMem.ConfigBits\[197\]
rlabel metal1 12466 14858 12466 14858 0 Inst_RAM_IO_ConfigMem.ConfigBits\[198\]
rlabel metal1 13294 14042 13294 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[199\]
rlabel metal3 14766 15300 14766 15300 0 Inst_RAM_IO_ConfigMem.ConfigBits\[200\]
rlabel metal1 15180 13770 15180 13770 0 Inst_RAM_IO_ConfigMem.ConfigBits\[201\]
rlabel metal1 4324 12342 4324 12342 0 Inst_RAM_IO_ConfigMem.ConfigBits\[202\]
rlabel metal1 4922 12614 4922 12614 0 Inst_RAM_IO_ConfigMem.ConfigBits\[203\]
rlabel metal1 6210 15334 6210 15334 0 Inst_RAM_IO_ConfigMem.ConfigBits\[204\]
rlabel metal1 7774 14926 7774 14926 0 Inst_RAM_IO_ConfigMem.ConfigBits\[205\]
rlabel metal1 13018 16728 13018 16728 0 Inst_RAM_IO_ConfigMem.ConfigBits\[206\]
rlabel metal1 13800 16218 13800 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[207\]
rlabel metal1 14904 15130 14904 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[208\]
rlabel metal2 15318 16796 15318 16796 0 Inst_RAM_IO_ConfigMem.ConfigBits\[209\]
rlabel metal1 4646 14858 4646 14858 0 Inst_RAM_IO_ConfigMem.ConfigBits\[210\]
rlabel metal1 5474 16048 5474 16048 0 Inst_RAM_IO_ConfigMem.ConfigBits\[211\]
rlabel metal1 6394 17306 6394 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[212\]
rlabel metal1 7452 17306 7452 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[213\]
rlabel metal1 14858 16728 14858 16728 0 Inst_RAM_IO_ConfigMem.ConfigBits\[214\]
rlabel metal1 16238 15674 16238 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[215\]
rlabel metal1 14398 24616 14398 24616 0 Inst_RAM_IO_ConfigMem.ConfigBits\[216\]
rlabel metal1 15778 24718 15778 24718 0 Inst_RAM_IO_ConfigMem.ConfigBits\[217\]
rlabel metal1 7222 36312 7222 36312 0 Inst_RAM_IO_ConfigMem.ConfigBits\[218\]
rlabel metal1 7866 36210 7866 36210 0 Inst_RAM_IO_ConfigMem.ConfigBits\[219\]
rlabel metal2 5014 27948 5014 27948 0 Inst_RAM_IO_ConfigMem.ConfigBits\[220\]
rlabel metal1 5014 27438 5014 27438 0 Inst_RAM_IO_ConfigMem.ConfigBits\[221\]
rlabel metal1 14490 28662 14490 28662 0 Inst_RAM_IO_ConfigMem.ConfigBits\[222\]
rlabel metal1 15410 28594 15410 28594 0 Inst_RAM_IO_ConfigMem.ConfigBits\[223\]
rlabel metal2 15226 23392 15226 23392 0 Inst_RAM_IO_ConfigMem.ConfigBits\[224\]
rlabel metal2 15686 23290 15686 23290 0 Inst_RAM_IO_ConfigMem.ConfigBits\[225\]
rlabel metal2 5474 32028 5474 32028 0 Inst_RAM_IO_ConfigMem.ConfigBits\[226\]
rlabel metal1 5474 31790 5474 31790 0 Inst_RAM_IO_ConfigMem.ConfigBits\[227\]
rlabel metal2 4554 25194 4554 25194 0 Inst_RAM_IO_ConfigMem.ConfigBits\[228\]
rlabel metal2 4922 25670 4922 25670 0 Inst_RAM_IO_ConfigMem.ConfigBits\[229\]
rlabel metal1 15180 29478 15180 29478 0 Inst_RAM_IO_ConfigMem.ConfigBits\[230\]
rlabel metal1 16008 27642 16008 27642 0 Inst_RAM_IO_ConfigMem.ConfigBits\[231\]
rlabel metal1 13892 25126 13892 25126 0 Inst_RAM_IO_ConfigMem.ConfigBits\[232\]
rlabel metal1 14720 24174 14720 24174 0 Inst_RAM_IO_ConfigMem.ConfigBits\[233\]
rlabel metal2 7406 39202 7406 39202 0 Inst_RAM_IO_ConfigMem.ConfigBits\[234\]
rlabel metal2 7958 39372 7958 39372 0 Inst_RAM_IO_ConfigMem.ConfigBits\[235\]
rlabel metal2 3910 27948 3910 27948 0 Inst_RAM_IO_ConfigMem.ConfigBits\[236\]
rlabel metal1 4324 27030 4324 27030 0 Inst_RAM_IO_ConfigMem.ConfigBits\[237\]
rlabel metal1 13570 29818 13570 29818 0 Inst_RAM_IO_ConfigMem.ConfigBits\[238\]
rlabel metal1 14536 30158 14536 30158 0 Inst_RAM_IO_ConfigMem.ConfigBits\[239\]
rlabel metal1 15272 22202 15272 22202 0 Inst_RAM_IO_ConfigMem.ConfigBits\[240\]
rlabel metal1 16192 22542 16192 22542 0 Inst_RAM_IO_ConfigMem.ConfigBits\[241\]
rlabel metal2 2438 32810 2438 32810 0 Inst_RAM_IO_ConfigMem.ConfigBits\[242\]
rlabel metal2 3082 32606 3082 32606 0 Inst_RAM_IO_ConfigMem.ConfigBits\[243\]
rlabel metal2 4002 25126 4002 25126 0 Inst_RAM_IO_ConfigMem.ConfigBits\[244\]
rlabel metal1 4738 24378 4738 24378 0 Inst_RAM_IO_ConfigMem.ConfigBits\[245\]
rlabel metal1 14536 33422 14536 33422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[246\]
rlabel metal2 15226 33660 15226 33660 0 Inst_RAM_IO_ConfigMem.ConfigBits\[247\]
rlabel metal2 12742 20978 12742 20978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[248\]
rlabel metal2 13294 21828 13294 21828 0 Inst_RAM_IO_ConfigMem.ConfigBits\[249\]
rlabel metal1 3365 20978 3365 20978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[250\]
rlabel metal1 2438 20570 2438 20570 0 Inst_RAM_IO_ConfigMem.ConfigBits\[251\]
rlabel metal2 8326 19669 8326 19669 0 Inst_RAM_IO_ConfigMem.ConfigBits\[252\]
rlabel metal2 8878 19516 8878 19516 0 Inst_RAM_IO_ConfigMem.ConfigBits\[253\]
rlabel metal1 12190 35224 12190 35224 0 Inst_RAM_IO_ConfigMem.ConfigBits\[254\]
rlabel metal1 12788 34714 12788 34714 0 Inst_RAM_IO_ConfigMem.ConfigBits\[255\]
rlabel metal1 11592 20026 11592 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[256\]
rlabel metal2 12098 21148 12098 21148 0 Inst_RAM_IO_ConfigMem.ConfigBits\[257\]
rlabel metal2 9430 5780 9430 5780 0 Inst_RAM_IO_ConfigMem.ConfigBits\[258\]
rlabel metal2 9982 6052 9982 6052 0 Inst_RAM_IO_ConfigMem.ConfigBits\[259\]
rlabel metal2 7866 27268 7866 27268 0 Inst_RAM_IO_ConfigMem.ConfigBits\[260\]
rlabel metal1 7912 26554 7912 26554 0 Inst_RAM_IO_ConfigMem.ConfigBits\[261\]
rlabel metal2 13662 26690 13662 26690 0 Inst_RAM_IO_ConfigMem.ConfigBits\[262\]
rlabel metal2 14214 27132 14214 27132 0 Inst_RAM_IO_ConfigMem.ConfigBits\[263\]
rlabel metal1 15686 17850 15686 17850 0 Inst_RAM_IO_ConfigMem.ConfigBits\[264\]
rlabel metal1 16514 18802 16514 18802 0 Inst_RAM_IO_ConfigMem.ConfigBits\[265\]
rlabel metal2 8510 36890 8510 36890 0 Inst_RAM_IO_ConfigMem.ConfigBits\[266\]
rlabel metal2 9062 36924 9062 36924 0 Inst_RAM_IO_ConfigMem.ConfigBits\[267\]
rlabel metal1 5612 21658 5612 21658 0 Inst_RAM_IO_ConfigMem.ConfigBits\[268\]
rlabel metal1 5658 21998 5658 21998 0 Inst_RAM_IO_ConfigMem.ConfigBits\[269\]
rlabel metal1 14628 19278 14628 19278 0 Inst_RAM_IO_ConfigMem.ConfigBits\[270\]
rlabel metal1 15180 18394 15180 18394 0 Inst_RAM_IO_ConfigMem.ConfigBits\[271\]
rlabel metal2 9706 18598 9706 18598 0 Inst_RAM_IO_ConfigMem.ConfigBits\[272\]
rlabel metal1 10764 18394 10764 18394 0 Inst_RAM_IO_ConfigMem.ConfigBits\[273\]
rlabel metal2 3910 36006 3910 36006 0 Inst_RAM_IO_ConfigMem.ConfigBits\[274\]
rlabel metal1 5014 35802 5014 35802 0 Inst_RAM_IO_ConfigMem.ConfigBits\[275\]
rlabel metal1 4140 20230 4140 20230 0 Inst_RAM_IO_ConfigMem.ConfigBits\[276\]
rlabel metal1 4968 19822 4968 19822 0 Inst_RAM_IO_ConfigMem.ConfigBits\[277\]
rlabel metal2 12558 11764 12558 11764 0 Inst_RAM_IO_ConfigMem.ConfigBits\[278\]
rlabel metal1 12834 11322 12834 11322 0 Inst_RAM_IO_ConfigMem.ConfigBits\[279\]
rlabel metal1 10028 15674 10028 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[280\]
rlabel metal1 8510 16660 8510 16660 0 Inst_RAM_IO_ConfigMem.ConfigBits\[281\]
rlabel metal1 3726 34374 3726 34374 0 Inst_RAM_IO_ConfigMem.ConfigBits\[282\]
rlabel metal1 4094 33592 4094 33592 0 Inst_RAM_IO_ConfigMem.ConfigBits\[283\]
rlabel metal1 2990 19244 2990 19244 0 Inst_RAM_IO_ConfigMem.ConfigBits\[284\]
rlabel metal1 3772 19346 3772 19346 0 Inst_RAM_IO_ConfigMem.ConfigBits\[285\]
rlabel metal1 11500 12954 11500 12954 0 Inst_RAM_IO_ConfigMem.ConfigBits\[286\]
rlabel metal1 13064 11526 13064 11526 0 Inst_RAM_IO_ConfigMem.ConfigBits\[287\]
rlabel metal2 8878 17510 8878 17510 0 Inst_RAM_IO_ConfigMem.ConfigBits\[288\]
rlabel metal1 10994 15674 10994 15674 0 Inst_RAM_IO_ConfigMem.ConfigBits\[289\]
rlabel metal1 4784 39270 4784 39270 0 Inst_RAM_IO_ConfigMem.ConfigBits\[290\]
rlabel metal1 5244 38998 5244 38998 0 Inst_RAM_IO_ConfigMem.ConfigBits\[291\]
rlabel metal2 3358 17204 3358 17204 0 Inst_RAM_IO_ConfigMem.ConfigBits\[292\]
rlabel metal1 3358 17306 3358 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[293\]
rlabel metal1 12604 10234 12604 10234 0 Inst_RAM_IO_ConfigMem.ConfigBits\[294\]
rlabel metal1 13524 11866 13524 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[295\]
rlabel metal1 8878 18598 8878 18598 0 Inst_RAM_IO_ConfigMem.ConfigBits\[296\]
rlabel metal1 9890 17170 9890 17170 0 Inst_RAM_IO_ConfigMem.ConfigBits\[297\]
rlabel metal1 3404 39270 3404 39270 0 Inst_RAM_IO_ConfigMem.ConfigBits\[298\]
rlabel metal1 4278 38318 4278 38318 0 Inst_RAM_IO_ConfigMem.ConfigBits\[299\]
rlabel metal1 3128 18122 3128 18122 0 Inst_RAM_IO_ConfigMem.ConfigBits\[300\]
rlabel metal2 3910 17782 3910 17782 0 Inst_RAM_IO_ConfigMem.ConfigBits\[301\]
rlabel metal1 10672 14790 10672 14790 0 Inst_RAM_IO_ConfigMem.ConfigBits\[302\]
rlabel metal1 12052 15334 12052 15334 0 Inst_RAM_IO_ConfigMem.ConfigBits\[303\]
rlabel metal1 8326 29002 8326 29002 0 Inst_RAM_IO_ConfigMem.ConfigBits\[304\]
rlabel metal1 9200 29206 9200 29206 0 Inst_RAM_IO_ConfigMem.ConfigBits\[305\]
rlabel metal2 5474 33830 5474 33830 0 Inst_RAM_IO_ConfigMem.ConfigBits\[306\]
rlabel metal2 5566 33354 5566 33354 0 Inst_RAM_IO_ConfigMem.ConfigBits\[307\]
rlabel metal2 7774 10676 7774 10676 0 Inst_RAM_IO_ConfigMem.ConfigBits\[308\]
rlabel metal1 8326 10778 8326 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[309\]
rlabel metal1 10028 34170 10028 34170 0 Inst_RAM_IO_ConfigMem.ConfigBits\[310\]
rlabel metal1 9706 34680 9706 34680 0 Inst_RAM_IO_ConfigMem.ConfigBits\[311\]
rlabel metal2 9614 36074 9614 36074 0 Inst_RAM_IO_ConfigMem.ConfigBits\[312\]
rlabel metal2 9798 35785 9798 35785 0 Inst_RAM_IO_ConfigMem.ConfigBits\[313\]
rlabel metal1 7590 8330 7590 8330 0 Inst_RAM_IO_ConfigMem.ConfigBits\[314\]
rlabel metal1 8418 8058 8418 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[315\]
rlabel metal2 6394 4964 6394 4964 0 Inst_RAM_IO_ConfigMem.ConfigBits\[316\]
rlabel metal1 7498 4794 7498 4794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[317\]
rlabel metal1 10994 37815 10994 37815 0 Inst_RAM_IO_ConfigMem.ConfigBits\[318\]
rlabel metal1 10488 37842 10488 37842 0 Inst_RAM_IO_ConfigMem.ConfigBits\[319\]
rlabel metal2 9982 19754 9982 19754 0 Inst_RAM_IO_ConfigMem.ConfigBits\[320\]
rlabel metal1 10212 19414 10212 19414 0 Inst_RAM_IO_ConfigMem.ConfigBits\[321\]
rlabel metal2 2806 37604 2806 37604 0 Inst_RAM_IO_ConfigMem.ConfigBits\[322\]
rlabel metal1 3312 37910 3312 37910 0 Inst_RAM_IO_ConfigMem.ConfigBits\[323\]
rlabel metal1 4094 21624 4094 21624 0 Inst_RAM_IO_ConfigMem.ConfigBits\[324\]
rlabel metal2 4094 22780 4094 22780 0 Inst_RAM_IO_ConfigMem.ConfigBits\[325\]
rlabel metal2 13018 19482 13018 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[326\]
rlabel metal1 12926 18938 12926 18938 0 Inst_RAM_IO_ConfigMem.ConfigBits\[327\]
rlabel metal1 9246 24888 9246 24888 0 Inst_RAM_IO_ConfigMem.ConfigBits\[48\]
rlabel metal1 10120 24174 10120 24174 0 Inst_RAM_IO_ConfigMem.ConfigBits\[49\]
rlabel metal1 2346 35258 2346 35258 0 Inst_RAM_IO_ConfigMem.ConfigBits\[50\]
rlabel metal2 2806 35972 2806 35972 0 Inst_RAM_IO_ConfigMem.ConfigBits\[51\]
rlabel metal2 2714 29954 2714 29954 0 Inst_RAM_IO_ConfigMem.ConfigBits\[52\]
rlabel via1 3250 30158 3250 30158 0 Inst_RAM_IO_ConfigMem.ConfigBits\[53\]
rlabel metal2 11822 33422 11822 33422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[54\]
rlabel metal2 12374 33116 12374 33116 0 Inst_RAM_IO_ConfigMem.ConfigBits\[55\]
rlabel metal1 9338 28186 9338 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[56\]
rlabel metal1 9936 28458 9936 28458 0 Inst_RAM_IO_ConfigMem.ConfigBits\[57\]
rlabel metal1 1886 29274 1886 29274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[58\]
rlabel metal2 2760 30702 2760 30702 0 Inst_RAM_IO_ConfigMem.ConfigBits\[59\]
rlabel metal1 2484 24038 2484 24038 0 Inst_RAM_IO_ConfigMem.ConfigBits\[60\]
rlabel metal2 2714 23494 2714 23494 0 Inst_RAM_IO_ConfigMem.ConfigBits\[61\]
rlabel metal2 9798 31246 9798 31246 0 Inst_RAM_IO_ConfigMem.ConfigBits\[62\]
rlabel metal2 10534 31969 10534 31969 0 Inst_RAM_IO_ConfigMem.ConfigBits\[63\]
rlabel metal1 12144 35598 12144 35598 0 Inst_RAM_IO_ConfigMem.ConfigBits\[64\]
rlabel metal2 12742 36108 12742 36108 0 Inst_RAM_IO_ConfigMem.ConfigBits\[65\]
rlabel metal2 2530 22100 2530 22100 0 Inst_RAM_IO_ConfigMem.ConfigBits\[66\]
rlabel metal2 2438 22236 2438 22236 0 Inst_RAM_IO_ConfigMem.ConfigBits\[67\]
rlabel metal2 2438 27676 2438 27676 0 Inst_RAM_IO_ConfigMem.ConfigBits\[68\]
rlabel metal1 2438 27098 2438 27098 0 Inst_RAM_IO_ConfigMem.ConfigBits\[69\]
rlabel metal2 12282 28492 12282 28492 0 Inst_RAM_IO_ConfigMem.ConfigBits\[70\]
rlabel metal2 12742 28220 12742 28220 0 Inst_RAM_IO_ConfigMem.ConfigBits\[71\]
rlabel metal1 12190 23290 12190 23290 0 Inst_RAM_IO_ConfigMem.ConfigBits\[72\]
rlabel metal1 12742 24242 12742 24242 0 Inst_RAM_IO_ConfigMem.ConfigBits\[73\]
rlabel metal1 12926 25738 12926 25738 0 Inst_RAM_IO_ConfigMem.ConfigBits\[74\]
rlabel metal1 7038 34102 7038 34102 0 Inst_RAM_IO_ConfigMem.ConfigBits\[75\]
rlabel metal1 7958 33422 7958 33422 0 Inst_RAM_IO_ConfigMem.ConfigBits\[76\]
rlabel metal1 8602 33898 8602 33898 0 Inst_RAM_IO_ConfigMem.ConfigBits\[77\]
rlabel metal1 6210 28696 6210 28696 0 Inst_RAM_IO_ConfigMem.ConfigBits\[78\]
rlabel metal1 6532 28934 6532 28934 0 Inst_RAM_IO_ConfigMem.ConfigBits\[79\]
rlabel metal1 8326 30192 8326 30192 0 Inst_RAM_IO_ConfigMem.ConfigBits\[80\]
rlabel metal1 13386 31246 13386 31246 0 Inst_RAM_IO_ConfigMem.ConfigBits\[81\]
rlabel metal1 15410 31858 15410 31858 0 Inst_RAM_IO_ConfigMem.ConfigBits\[82\]
rlabel metal1 14996 34374 14996 34374 0 Inst_RAM_IO_ConfigMem.ConfigBits\[83\]
rlabel via1 10073 23630 10073 23630 0 Inst_RAM_IO_ConfigMem.ConfigBits\[84\]
rlabel metal1 10304 23290 10304 23290 0 Inst_RAM_IO_ConfigMem.ConfigBits\[85\]
rlabel metal1 7544 34918 7544 34918 0 Inst_RAM_IO_ConfigMem.ConfigBits\[86\]
rlabel metal1 8280 33082 8280 33082 0 Inst_RAM_IO_ConfigMem.ConfigBits\[87\]
rlabel metal1 5888 20298 5888 20298 0 Inst_RAM_IO_ConfigMem.ConfigBits\[88\]
rlabel metal1 6762 20910 6762 20910 0 Inst_RAM_IO_ConfigMem.ConfigBits\[89\]
rlabel metal1 10810 31892 10810 31892 0 Inst_RAM_IO_ConfigMem.ConfigBits\[90\]
rlabel metal2 12558 31620 12558 31620 0 Inst_RAM_IO_ConfigMem.ConfigBits\[91\]
rlabel metal1 9154 27302 9154 27302 0 Inst_RAM_IO_ConfigMem.ConfigBits\[92\]
rlabel metal1 9798 25976 9798 25976 0 Inst_RAM_IO_ConfigMem.ConfigBits\[93\]
rlabel metal1 7912 31654 7912 31654 0 Inst_RAM_IO_ConfigMem.ConfigBits\[94\]
rlabel metal1 7820 30702 7820 30702 0 Inst_RAM_IO_ConfigMem.ConfigBits\[95\]
rlabel metal1 8464 7174 8464 7174 0 Inst_RAM_IO_ConfigMem.ConfigBits\[96\]
rlabel metal2 9246 7548 9246 7548 0 Inst_RAM_IO_ConfigMem.ConfigBits\[97\]
rlabel metal2 10442 30124 10442 30124 0 Inst_RAM_IO_ConfigMem.ConfigBits\[98\]
rlabel metal1 11408 29614 11408 29614 0 Inst_RAM_IO_ConfigMem.ConfigBits\[99\]
rlabel metal2 11086 18938 11086 18938 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG0
rlabel metal2 7406 35632 7406 35632 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG1
rlabel metal1 4692 22746 4692 22746 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG2
rlabel metal2 11684 31790 11684 31790 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG3
rlabel metal2 12328 24174 12328 24174 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
rlabel metal1 1564 28934 1564 28934 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
rlabel metal2 7314 15980 7314 15980 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
rlabel metal1 16100 26554 16100 26554 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
rlabel metal1 10488 35802 10488 35802 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
rlabel metal1 7313 23154 7313 23154 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
rlabel metal1 4186 13872 4186 13872 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
rlabel metal1 14374 26894 14374 26894 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
rlabel metal1 14490 24718 14490 24718 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG0
rlabel metal1 6210 17782 6210 17782 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG1
rlabel metal1 5221 30158 5221 30158 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG10
rlabel metal2 13984 20332 13984 20332 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG11
rlabel metal1 15318 22542 15318 22542 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG12
rlabel via1 7510 23154 7510 23154 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG13
rlabel metal2 4278 25347 4278 25347 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG14
rlabel metal2 12236 27540 12236 27540 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG15
rlabel metal1 5520 19686 5520 19686 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG2
rlabel metal1 14950 28594 14950 28594 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG3
rlabel metal1 14766 23188 14766 23188 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG4
rlabel metal1 6394 14892 6394 14892 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG5
rlabel metal2 4830 24735 4830 24735 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG6
rlabel metal1 14306 31926 14306 31926 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG7
rlabel metal2 14582 24225 14582 24225 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG8
rlabel metal1 7590 38862 7590 38862 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG9
rlabel metal2 10810 24582 10810 24582 0 Inst_RAM_IO_switch_matrix.N1BEG0
rlabel metal2 1702 42398 1702 42398 0 Inst_RAM_IO_switch_matrix.N1BEG1
rlabel metal1 3956 30090 3956 30090 0 Inst_RAM_IO_switch_matrix.N1BEG2
rlabel metal2 12558 39965 12558 39965 0 Inst_RAM_IO_switch_matrix.N1BEG3
rlabel metal2 2300 41106 2300 41106 0 Inst_RAM_IO_switch_matrix.N2BEG0
rlabel metal2 2530 41491 2530 41491 0 Inst_RAM_IO_switch_matrix.N2BEG1
rlabel metal1 1564 42194 1564 42194 0 Inst_RAM_IO_switch_matrix.N2BEG2
rlabel metal2 7636 39916 7636 39916 0 Inst_RAM_IO_switch_matrix.N2BEG3
rlabel metal2 3956 38964 3956 38964 0 Inst_RAM_IO_switch_matrix.N2BEG4
rlabel metal3 3427 41004 3427 41004 0 Inst_RAM_IO_switch_matrix.N2BEG5
rlabel metal3 1495 32844 1495 32844 0 Inst_RAM_IO_switch_matrix.N2BEG6
rlabel metal1 13294 27914 13294 27914 0 Inst_RAM_IO_switch_matrix.N2BEG7
rlabel metal3 2047 41412 2047 41412 0 Inst_RAM_IO_switch_matrix.N2BEGb0
rlabel metal1 4554 33082 4554 33082 0 Inst_RAM_IO_switch_matrix.N2BEGb1
rlabel metal2 184 27404 184 27404 0 Inst_RAM_IO_switch_matrix.N2BEGb2
rlabel metal1 4554 34170 4554 34170 0 Inst_RAM_IO_switch_matrix.N2BEGb3
rlabel metal1 4968 35258 4968 35258 0 Inst_RAM_IO_switch_matrix.N2BEGb4
rlabel metal4 1104 30260 1104 30260 0 Inst_RAM_IO_switch_matrix.N2BEGb5
rlabel metal2 13110 39899 13110 39899 0 Inst_RAM_IO_switch_matrix.N2BEGb6
rlabel metal1 4968 37978 4968 37978 0 Inst_RAM_IO_switch_matrix.N2BEGb7
rlabel metal1 13662 25942 13662 25942 0 Inst_RAM_IO_switch_matrix.N4BEG0
rlabel metal1 8924 34714 8924 34714 0 Inst_RAM_IO_switch_matrix.N4BEG1
rlabel metal2 9016 34612 9016 34612 0 Inst_RAM_IO_switch_matrix.N4BEG2
rlabel metal1 12052 41514 12052 41514 0 Inst_RAM_IO_switch_matrix.N4BEG3
rlabel metal3 9131 19380 9131 19380 0 Inst_RAM_IO_switch_matrix.S1BEG0
rlabel metal1 7774 15334 7774 15334 0 Inst_RAM_IO_switch_matrix.S1BEG1
rlabel metal1 7544 20774 7544 20774 0 Inst_RAM_IO_switch_matrix.S1BEG2
rlabel metal1 12880 31654 12880 31654 0 Inst_RAM_IO_switch_matrix.S1BEG3
rlabel metal3 10649 19244 10649 19244 0 Inst_RAM_IO_switch_matrix.S2BEG0
rlabel metal1 8602 30838 8602 30838 0 Inst_RAM_IO_switch_matrix.S2BEG1
rlabel metal1 9798 6630 9798 6630 0 Inst_RAM_IO_switch_matrix.S2BEG2
rlabel metal2 12466 28917 12466 28917 0 Inst_RAM_IO_switch_matrix.S2BEG3
rlabel metal3 15065 22100 15065 22100 0 Inst_RAM_IO_switch_matrix.S2BEG4
rlabel via3 805 18156 805 18156 0 Inst_RAM_IO_switch_matrix.S2BEG5
rlabel metal2 2162 19924 2162 19924 0 Inst_RAM_IO_switch_matrix.S2BEG6
rlabel metal3 18446 21420 18446 21420 0 Inst_RAM_IO_switch_matrix.S2BEG7
rlabel metal2 10304 22508 10304 22508 0 Inst_RAM_IO_switch_matrix.S2BEGb0
rlabel metal3 1725 23460 1725 23460 0 Inst_RAM_IO_switch_matrix.S2BEGb1
rlabel metal1 9660 8466 9660 8466 0 Inst_RAM_IO_switch_matrix.S2BEGb2
rlabel metal3 13800 20468 13800 20468 0 Inst_RAM_IO_switch_matrix.S2BEGb3
rlabel metal2 8004 22542 8004 22542 0 Inst_RAM_IO_switch_matrix.S2BEGb4
rlabel metal2 9568 8364 9568 8364 0 Inst_RAM_IO_switch_matrix.S2BEGb5
rlabel metal1 9936 4726 9936 4726 0 Inst_RAM_IO_switch_matrix.S2BEGb6
rlabel metal2 15410 35156 15410 35156 0 Inst_RAM_IO_switch_matrix.S2BEGb7
rlabel via3 16491 20740 16491 20740 0 Inst_RAM_IO_switch_matrix.S4BEG0
rlabel metal3 11661 20196 11661 20196 0 Inst_RAM_IO_switch_matrix.S4BEG1
rlabel metal3 8855 24956 8855 24956 0 Inst_RAM_IO_switch_matrix.S4BEG2
rlabel metal2 19366 17408 19366 17408 0 Inst_RAM_IO_switch_matrix.S4BEG3
rlabel metal1 10212 15878 10212 15878 0 Inst_RAM_IO_switch_matrix.W1BEG0
rlabel metal1 6578 6358 6578 6358 0 Inst_RAM_IO_switch_matrix.W1BEG1
rlabel metal1 5980 7174 5980 7174 0 Inst_RAM_IO_switch_matrix.W1BEG2
rlabel metal2 13110 5445 13110 5445 0 Inst_RAM_IO_switch_matrix.W1BEG3
rlabel metal1 13570 6766 13570 6766 0 Inst_RAM_IO_switch_matrix.W2BEG0
rlabel metal1 6256 5338 6256 5338 0 Inst_RAM_IO_switch_matrix.W2BEG1
rlabel metal1 4554 5780 4554 5780 0 Inst_RAM_IO_switch_matrix.W2BEG2
rlabel metal3 5106 6868 5106 6868 0 Inst_RAM_IO_switch_matrix.W2BEG3
rlabel metal2 4186 6443 4186 6443 0 Inst_RAM_IO_switch_matrix.W2BEG4
rlabel metal1 4508 6426 4508 6426 0 Inst_RAM_IO_switch_matrix.W2BEG5
rlabel metal1 4324 4114 4324 4114 0 Inst_RAM_IO_switch_matrix.W2BEG6
rlabel metal1 11989 6970 11989 6970 0 Inst_RAM_IO_switch_matrix.W2BEG7
rlabel metal1 13892 7378 13892 7378 0 Inst_RAM_IO_switch_matrix.W2BEGb0
rlabel metal2 4370 7888 4370 7888 0 Inst_RAM_IO_switch_matrix.W2BEGb1
rlabel metal2 8418 8585 8418 8585 0 Inst_RAM_IO_switch_matrix.W2BEGb2
rlabel metal1 6026 8534 6026 8534 0 Inst_RAM_IO_switch_matrix.W2BEGb3
rlabel metal2 10074 9333 10074 9333 0 Inst_RAM_IO_switch_matrix.W2BEGb4
rlabel metal1 4462 9350 4462 9350 0 Inst_RAM_IO_switch_matrix.W2BEGb5
rlabel metal1 3450 4998 3450 4998 0 Inst_RAM_IO_switch_matrix.W2BEGb6
rlabel metal1 9246 9146 9246 9146 0 Inst_RAM_IO_switch_matrix.W2BEGb7
rlabel metal1 7590 16728 7590 16728 0 Inst_RAM_IO_switch_matrix.W6BEG0
rlabel metal1 5750 30294 5750 30294 0 Inst_RAM_IO_switch_matrix.W6BEG1
rlabel metal2 6026 17102 6026 17102 0 Inst_RAM_IO_switch_matrix.W6BEG10
rlabel via2 16054 16643 16054 16643 0 Inst_RAM_IO_switch_matrix.W6BEG11
rlabel metal2 5474 18173 5474 18173 0 Inst_RAM_IO_switch_matrix.W6BEG2
rlabel metal2 5474 14960 5474 14960 0 Inst_RAM_IO_switch_matrix.W6BEG3
rlabel metal2 9614 15351 9614 15351 0 Inst_RAM_IO_switch_matrix.W6BEG4
rlabel via2 4462 12053 4462 12053 0 Inst_RAM_IO_switch_matrix.W6BEG5
rlabel metal2 2254 14756 2254 14756 0 Inst_RAM_IO_switch_matrix.W6BEG6
rlabel metal2 15502 15521 15502 15521 0 Inst_RAM_IO_switch_matrix.W6BEG7
rlabel metal1 15594 16218 15594 16218 0 Inst_RAM_IO_switch_matrix.W6BEG8
rlabel metal1 5152 16218 5152 16218 0 Inst_RAM_IO_switch_matrix.W6BEG9
rlabel metal1 4600 10030 4600 10030 0 Inst_RAM_IO_switch_matrix.WW4BEG0
rlabel metal1 3726 11594 3726 11594 0 Inst_RAM_IO_switch_matrix.WW4BEG1
rlabel metal1 6578 12852 6578 12852 0 Inst_RAM_IO_switch_matrix.WW4BEG10
rlabel metal1 4738 13940 4738 13940 0 Inst_RAM_IO_switch_matrix.WW4BEG11
rlabel via2 15962 13243 15962 13243 0 Inst_RAM_IO_switch_matrix.WW4BEG12
rlabel metal2 4554 13770 4554 13770 0 Inst_RAM_IO_switch_matrix.WW4BEG13
rlabel metal2 6210 15776 6210 15776 0 Inst_RAM_IO_switch_matrix.WW4BEG14
rlabel metal1 7176 12818 7176 12818 0 Inst_RAM_IO_switch_matrix.WW4BEG15
rlabel metal1 4922 9452 4922 9452 0 Inst_RAM_IO_switch_matrix.WW4BEG2
rlabel metal2 11270 11305 11270 11305 0 Inst_RAM_IO_switch_matrix.WW4BEG3
rlabel metal1 13754 10778 13754 10778 0 Inst_RAM_IO_switch_matrix.WW4BEG4
rlabel metal1 1150 11254 1150 11254 0 Inst_RAM_IO_switch_matrix.WW4BEG5
rlabel metal2 8234 13600 8234 13600 0 Inst_RAM_IO_switch_matrix.WW4BEG6
rlabel metal1 7038 12308 7038 12308 0 Inst_RAM_IO_switch_matrix.WW4BEG7
rlabel via2 16146 12699 16146 12699 0 Inst_RAM_IO_switch_matrix.WW4BEG8
rlabel metal1 5198 11322 5198 11322 0 Inst_RAM_IO_switch_matrix.WW4BEG9
rlabel metal1 13294 23834 13294 23834 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0
rlabel metal1 13432 24378 13432 24378 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1
rlabel metal1 13294 24650 13294 24650 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 12880 24922 12880 24922 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal1 12512 25466 12512 25466 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_
rlabel metal2 12190 25568 12190 25568 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_
rlabel metal1 8602 34102 8602 34102 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0
rlabel metal1 10166 33524 10166 33524 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1
rlabel metal1 10442 34000 10442 34000 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 9384 33626 9384 33626 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 10120 34102 10120 34102 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_
rlabel metal1 8786 34170 8786 34170 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_
rlabel metal1 7130 29138 7130 29138 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0
rlabel metal1 7682 28526 7682 28526 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1
rlabel metal1 8050 28628 8050 28628 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal1 7866 28662 7866 28662 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal1 8786 30056 8786 30056 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_
rlabel metal2 8602 30362 8602 30362 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_
rlabel metal1 14306 31450 14306 31450 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0
rlabel metal1 15824 31994 15824 31994 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1
rlabel metal2 13846 32674 13846 32674 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 15824 33082 15824 33082 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal1 15640 33014 15640 33014 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_
rlabel metal1 14996 33286 14996 33286 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_
rlabel metal1 16008 21522 16008 21522 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0
rlabel metal1 16192 20434 16192 20434 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1
rlabel metal1 16698 20944 16698 20944 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 16514 20400 16514 20400 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal1 16238 20842 16238 20842 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_
rlabel metal1 16560 20570 16560 20570 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_
rlabel metal1 8602 23188 8602 23188 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0
rlabel metal1 9108 23102 9108 23102 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1
rlabel metal1 8878 21998 8878 21998 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 9384 22066 9384 22066 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 9338 22202 9338 22202 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_
rlabel metal1 9752 21930 9752 21930 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_
rlabel metal2 7130 25160 7130 25160 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0
rlabel metal1 7820 24786 7820 24786 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1
rlabel metal1 6946 25840 6946 25840 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal2 7958 25432 7958 25432 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal1 8050 25364 8050 25364 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_
rlabel metal1 8372 25262 8372 25262 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_
rlabel metal1 16100 30906 16100 30906 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0
rlabel metal1 16376 31314 16376 31314 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1
rlabel metal1 16330 32436 16330 32436 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 16882 31348 16882 31348 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal2 16422 31450 16422 31450 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_
rlabel metal1 16836 30702 16836 30702 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_
rlabel metal1 2070 43418 2070 43418 0 N1BEG[0]
rlabel metal2 2622 43428 2622 43428 0 N1BEG[1]
rlabel metal2 2806 43972 2806 43972 0 N1BEG[2]
rlabel metal2 2990 43598 2990 43598 0 N1BEG[3]
rlabel metal2 2438 670 2438 670 0 N1END[0]
rlabel metal2 2622 636 2622 636 0 N1END[1]
rlabel metal2 2806 976 2806 976 0 N1END[2]
rlabel metal2 2990 1214 2990 1214 0 N1END[3]
rlabel metal2 3174 43870 3174 43870 0 N2BEG[0]
rlabel metal1 3220 42670 3220 42670 0 N2BEG[1]
rlabel metal1 3220 43350 3220 43350 0 N2BEG[2]
rlabel metal1 3680 42738 3680 42738 0 N2BEG[3]
rlabel metal1 3174 42296 3174 42296 0 N2BEG[4]
rlabel metal1 3818 42330 3818 42330 0 N2BEG[5]
rlabel metal1 4232 42738 4232 42738 0 N2BEG[6]
rlabel metal2 4462 43564 4462 43564 0 N2BEG[7]
rlabel metal2 4646 43972 4646 43972 0 N2BEGb[0]
rlabel metal1 4508 42330 4508 42330 0 N2BEGb[1]
rlabel metal1 4876 42738 4876 42738 0 N2BEGb[2]
rlabel metal1 5152 42330 5152 42330 0 N2BEGb[3]
rlabel metal1 5336 42738 5336 42738 0 N2BEGb[4]
rlabel metal2 5566 43972 5566 43972 0 N2BEGb[5]
rlabel metal2 5750 43428 5750 43428 0 N2BEGb[6]
rlabel metal1 5704 43146 5704 43146 0 N2BEGb[7]
rlabel metal2 4646 976 4646 976 0 N2END[0]
rlabel metal2 4830 364 4830 364 0 N2END[1]
rlabel metal2 5014 755 5014 755 0 N2END[2]
rlabel metal2 5198 738 5198 738 0 N2END[3]
rlabel metal2 5435 68 5435 68 0 N2END[4]
rlabel metal2 5566 636 5566 636 0 N2END[5]
rlabel metal2 5750 1554 5750 1554 0 N2END[6]
rlabel metal2 5881 68 5881 68 0 N2END[7]
rlabel metal2 3227 68 3227 68 0 N2MID[0]
rlabel metal2 3358 364 3358 364 0 N2MID[1]
rlabel metal2 3542 670 3542 670 0 N2MID[2]
rlabel metal2 3726 704 3726 704 0 N2MID[3]
rlabel metal2 3963 68 3963 68 0 N2MID[4]
rlabel metal1 4646 2380 4646 2380 0 N2MID[5]
rlabel metal2 4331 68 4331 68 0 N2MID[6]
rlabel metal2 4462 670 4462 670 0 N2MID[7]
rlabel metal1 6072 42738 6072 42738 0 N4BEG[0]
rlabel metal2 7958 43632 7958 43632 0 N4BEG[10]
rlabel metal1 8280 42330 8280 42330 0 N4BEG[11]
rlabel metal2 8326 43785 8326 43785 0 N4BEG[12]
rlabel metal1 8142 43350 8142 43350 0 N4BEG[13]
rlabel metal1 8510 43418 8510 43418 0 N4BEG[14]
rlabel metal2 8878 43513 8878 43513 0 N4BEG[15]
rlabel metal2 4186 43639 4186 43639 0 N4BEG[1]
rlabel metal1 6440 42738 6440 42738 0 N4BEG[2]
rlabel metal1 6348 41786 6348 41786 0 N4BEG[3]
rlabel metal2 6854 43428 6854 43428 0 N4BEG[4]
rlabel metal2 7038 43564 7038 43564 0 N4BEG[5]
rlabel metal2 7222 44057 7222 44057 0 N4BEG[6]
rlabel metal1 7222 43418 7222 43418 0 N4BEG[7]
rlabel metal2 7590 43428 7590 43428 0 N4BEG[8]
rlabel metal1 7544 42058 7544 42058 0 N4BEG[9]
rlabel metal1 3082 42092 3082 42092 0 N4BEG_outbuf_0.A
rlabel metal1 5290 41208 5290 41208 0 N4BEG_outbuf_0.X
rlabel metal3 1955 18292 1955 18292 0 N4BEG_outbuf_1.A
rlabel metal1 4370 41616 4370 41616 0 N4BEG_outbuf_1.X
rlabel metal3 4669 18836 4669 18836 0 N4BEG_outbuf_10.A
rlabel metal1 9430 42160 9430 42160 0 N4BEG_outbuf_10.X
rlabel metal3 9292 28968 9292 28968 0 N4BEG_outbuf_11.A
rlabel metal1 8510 41616 8510 41616 0 N4BEG_outbuf_11.X
rlabel metal4 1196 36712 1196 36712 0 N4BEG_outbuf_2.A
rlabel metal2 5658 40596 5658 40596 0 N4BEG_outbuf_2.X
rlabel metal1 920 36142 920 36142 0 N4BEG_outbuf_3.A
rlabel metal1 4692 41582 4692 41582 0 N4BEG_outbuf_3.X
rlabel metal1 14214 38352 14214 38352 0 N4BEG_outbuf_4.A
rlabel metal1 6578 41174 6578 41174 0 N4BEG_outbuf_4.X
rlabel metal3 8441 35836 8441 35836 0 N4BEG_outbuf_5.A
rlabel metal1 7268 41718 7268 41718 0 N4BEG_outbuf_5.X
rlabel metal2 12834 40494 12834 40494 0 N4BEG_outbuf_6.A
rlabel metal1 7314 41242 7314 41242 0 N4BEG_outbuf_6.X
rlabel metal3 1104 18972 1104 18972 0 N4BEG_outbuf_7.A
rlabel metal1 7038 41072 7038 41072 0 N4BEG_outbuf_7.X
rlabel metal3 9085 20740 9085 20740 0 N4BEG_outbuf_8.A
rlabel metal1 7498 40902 7498 40902 0 N4BEG_outbuf_8.X
rlabel metal3 15548 38556 15548 38556 0 N4BEG_outbuf_9.A
rlabel metal1 8280 41582 8280 41582 0 N4BEG_outbuf_9.X
rlabel metal2 6118 398 6118 398 0 N4END[0]
rlabel metal1 7866 3026 7866 3026 0 N4END[10]
rlabel metal2 8142 687 8142 687 0 N4END[11]
rlabel metal2 8326 619 8326 619 0 N4END[12]
rlabel metal2 8510 755 8510 755 0 N4END[13]
rlabel metal2 8641 68 8641 68 0 N4END[14]
rlabel metal2 8878 823 8878 823 0 N4END[15]
rlabel metal2 6302 755 6302 755 0 N4END[1]
rlabel metal2 6486 704 6486 704 0 N4END[2]
rlabel metal2 6670 364 6670 364 0 N4END[3]
rlabel metal2 6854 551 6854 551 0 N4END[4]
rlabel metal2 7038 959 7038 959 0 N4END[5]
rlabel metal2 7360 3026 7360 3026 0 N4END[6]
rlabel metal1 7406 2924 7406 2924 0 N4END[7]
rlabel metal2 7590 143 7590 143 0 N4END[8]
rlabel metal2 7774 959 7774 959 0 N4END[9]
rlabel metal3 20283 7140 20283 7140 0 RAM2FAB_D0_I0
rlabel metal2 9890 4896 9890 4896 0 RAM2FAB_D0_I1
rlabel metal1 16514 8024 16514 8024 0 RAM2FAB_D0_I2
rlabel metal2 16054 9180 16054 9180 0 RAM2FAB_D0_I3
rlabel metal2 14858 5695 14858 5695 0 RAM2FAB_D1_I0
rlabel metal1 12374 5678 12374 5678 0 RAM2FAB_D1_I1
rlabel metal2 14582 5508 14582 5508 0 RAM2FAB_D1_I2
rlabel metal1 10350 4148 10350 4148 0 RAM2FAB_D1_I3
rlabel metal3 16514 3128 16514 3128 0 RAM2FAB_D2_I0
rlabel metal3 21594 3332 21594 3332 0 RAM2FAB_D2_I1
rlabel metal3 20306 3876 20306 3876 0 RAM2FAB_D2_I2
rlabel metal3 16836 4080 16836 4080 0 RAM2FAB_D2_I3
rlabel metal2 17618 2244 17618 2244 0 RAM2FAB_D3_I0
rlabel metal2 10396 2346 10396 2346 0 RAM2FAB_D3_I1
rlabel via2 14766 1275 14766 1275 0 RAM2FAB_D3_I2
rlabel metal3 13202 1768 13202 1768 0 RAM2FAB_D3_I3
rlabel metal2 9062 636 9062 636 0 S1BEG[0]
rlabel metal2 9246 823 9246 823 0 S1BEG[1]
rlabel metal2 9430 908 9430 908 0 S1BEG[2]
rlabel metal2 9614 908 9614 908 0 S1BEG[3]
rlabel metal2 9062 43904 9062 43904 0 S1END[0]
rlabel metal2 9246 43598 9246 43598 0 S1END[1]
rlabel metal2 9430 43904 9430 43904 0 S1END[2]
rlabel metal2 9614 43904 9614 43904 0 S1END[3]
rlabel metal1 10672 1190 10672 1190 0 S2BEG[0]
rlabel metal2 11638 1829 11638 1829 0 S2BEG[1]
rlabel metal2 11691 68 11691 68 0 S2BEG[2]
rlabel metal1 11408 1190 11408 1190 0 S2BEG[3]
rlabel metal1 11868 1462 11868 1462 0 S2BEG[4]
rlabel metal2 12190 636 12190 636 0 S2BEG[5]
rlabel metal2 12420 1530 12420 1530 0 S2BEG[6]
rlabel metal1 13248 1190 13248 1190 0 S2BEG[7]
rlabel metal2 9798 636 9798 636 0 S2BEGb[0]
rlabel metal1 9338 1292 9338 1292 0 S2BEGb[1]
rlabel metal2 10166 551 10166 551 0 S2BEGb[2]
rlabel metal1 10120 1462 10120 1462 0 S2BEGb[3]
rlabel metal2 10534 908 10534 908 0 S2BEGb[4]
rlabel metal2 9154 884 9154 884 0 S2BEGb[5]
rlabel metal1 10902 1734 10902 1734 0 S2BEGb[6]
rlabel metal2 11086 364 11086 364 0 S2BEGb[7]
rlabel metal2 9798 43394 9798 43394 0 S2END[0]
rlabel metal2 9982 43972 9982 43972 0 S2END[1]
rlabel metal2 10166 44176 10166 44176 0 S2END[2]
rlabel metal2 10350 44057 10350 44057 0 S2END[3]
rlabel metal2 10534 43598 10534 43598 0 S2END[4]
rlabel metal2 10718 44193 10718 44193 0 S2END[5]
rlabel metal2 10902 44125 10902 44125 0 S2END[6]
rlabel metal2 11086 44125 11086 44125 0 S2END[7]
rlabel metal2 11270 44193 11270 44193 0 S2MID[0]
rlabel metal2 11454 43598 11454 43598 0 S2MID[1]
rlabel metal2 11638 44193 11638 44193 0 S2MID[2]
rlabel metal2 11822 44261 11822 44261 0 S2MID[3]
rlabel metal2 12006 43904 12006 43904 0 S2MID[4]
rlabel metal2 12190 43904 12190 43904 0 S2MID[5]
rlabel metal2 12374 43904 12374 43904 0 S2MID[6]
rlabel metal2 12558 44057 12558 44057 0 S2MID[7]
rlabel metal1 13340 1870 13340 1870 0 S4BEG[0]
rlabel metal2 14582 432 14582 432 0 S4BEG[10]
rlabel metal2 14766 211 14766 211 0 S4BEG[11]
rlabel metal2 14950 160 14950 160 0 S4BEG[12]
rlabel metal2 15134 211 15134 211 0 S4BEG[13]
rlabel metal2 15318 126 15318 126 0 S4BEG[14]
rlabel metal2 15502 194 15502 194 0 S4BEG[15]
rlabel metal2 12979 68 12979 68 0 S4BEG[1]
rlabel metal1 13340 1734 13340 1734 0 S4BEG[2]
rlabel metal2 13340 1734 13340 1734 0 S4BEG[3]
rlabel metal1 13938 1734 13938 1734 0 S4BEG[4]
rlabel metal1 12420 1258 12420 1258 0 S4BEG[5]
rlabel metal2 13846 160 13846 160 0 S4BEG[6]
rlabel metal2 14030 262 14030 262 0 S4BEG[7]
rlabel metal2 14214 228 14214 228 0 S4BEG[8]
rlabel metal2 14398 262 14398 262 0 S4BEG[9]
rlabel metal1 13018 42228 13018 42228 0 S4BEG_outbuf_0.A
rlabel metal2 18906 25772 18906 25772 0 S4BEG_outbuf_0.X
rlabel metal1 13524 42194 13524 42194 0 S4BEG_outbuf_1.A
rlabel metal1 13064 36550 13064 36550 0 S4BEG_outbuf_1.X
rlabel metal1 15686 42296 15686 42296 0 S4BEG_outbuf_10.A
rlabel metal2 14996 38522 14996 38522 0 S4BEG_outbuf_10.X
rlabel metal1 15134 41616 15134 41616 0 S4BEG_outbuf_11.A
rlabel metal2 20516 38828 20516 38828 0 S4BEG_outbuf_11.X
rlabel metal1 13754 42228 13754 42228 0 S4BEG_outbuf_2.A
rlabel metal1 14628 37774 14628 37774 0 S4BEG_outbuf_2.X
rlabel metal1 14214 42160 14214 42160 0 S4BEG_outbuf_3.A
rlabel metal2 14306 40154 14306 40154 0 S4BEG_outbuf_3.X
rlabel metal2 14490 42636 14490 42636 0 S4BEG_outbuf_4.A
rlabel metal1 14536 41990 14536 41990 0 S4BEG_outbuf_4.X
rlabel viali 14214 41580 14214 41580 0 S4BEG_outbuf_5.A
rlabel metal3 18400 23596 18400 23596 0 S4BEG_outbuf_5.X
rlabel metal1 14858 42228 14858 42228 0 S4BEG_outbuf_6.A
rlabel metal2 14858 41769 14858 41769 0 S4BEG_outbuf_6.X
rlabel metal1 15088 42602 15088 42602 0 S4BEG_outbuf_7.A
rlabel metal3 17319 20604 17319 20604 0 S4BEG_outbuf_7.X
rlabel metal1 15502 42194 15502 42194 0 S4BEG_outbuf_8.A
rlabel metal4 19780 26996 19780 26996 0 S4BEG_outbuf_8.X
rlabel metal1 14858 41582 14858 41582 0 S4BEG_outbuf_9.A
rlabel metal3 14927 41140 14927 41140 0 S4BEG_outbuf_9.X
rlabel metal2 12742 43904 12742 43904 0 S4END[0]
rlabel metal1 14582 41208 14582 41208 0 S4END[10]
rlabel metal1 14812 41242 14812 41242 0 S4END[11]
rlabel metal2 14950 44261 14950 44261 0 S4END[12]
rlabel metal2 15134 43904 15134 43904 0 S4END[13]
rlabel metal2 15318 44125 15318 44125 0 S4END[14]
rlabel metal2 15502 44465 15502 44465 0 S4END[15]
rlabel metal2 12926 43938 12926 43938 0 S4END[1]
rlabel metal2 13110 43598 13110 43598 0 S4END[2]
rlabel metal2 13294 43972 13294 43972 0 S4END[3]
rlabel metal2 13478 44261 13478 44261 0 S4END[4]
rlabel metal2 13662 44074 13662 44074 0 S4END[5]
rlabel metal2 13846 44193 13846 44193 0 S4END[6]
rlabel metal2 14030 43649 14030 43649 0 S4END[7]
rlabel metal2 14214 44261 14214 44261 0 S4END[8]
rlabel metal2 14398 43989 14398 43989 0 S4END[9]
rlabel metal1 14628 38862 14628 38862 0 UserCLK
rlabel via2 16238 40715 16238 40715 0 UserCLKo
rlabel metal3 1096 4964 1096 4964 0 W1BEG[0]
rlabel metal3 728 5236 728 5236 0 W1BEG[1]
rlabel metal1 4347 4794 4347 4794 0 W1BEG[2]
rlabel metal3 774 5780 774 5780 0 W1BEG[3]
rlabel metal3 1648 6052 1648 6052 0 W2BEG[0]
rlabel metal3 1004 6324 1004 6324 0 W2BEG[1]
rlabel metal1 2300 4454 2300 4454 0 W2BEG[2]
rlabel metal2 4002 6375 4002 6375 0 W2BEG[3]
rlabel metal3 1556 7140 1556 7140 0 W2BEG[4]
rlabel metal1 3036 6970 3036 6970 0 W2BEG[5]
rlabel metal3 774 7684 774 7684 0 W2BEG[6]
rlabel metal3 2108 7956 2108 7956 0 W2BEG[7]
rlabel metal3 1648 8228 1648 8228 0 W2BEGb[0]
rlabel metal3 682 8500 682 8500 0 W2BEGb[1]
rlabel metal3 1234 8772 1234 8772 0 W2BEGb[2]
rlabel metal3 958 9044 958 9044 0 W2BEGb[3]
rlabel metal3 866 9316 866 9316 0 W2BEGb[4]
rlabel metal3 728 9588 728 9588 0 W2BEGb[5]
rlabel metal2 4278 9435 4278 9435 0 W2BEGb[6]
rlabel metal2 4462 7021 4462 7021 0 W2BEGb[7]
rlabel metal3 498 14756 498 14756 0 W6BEG[0]
rlabel metal3 866 17476 866 17476 0 W6BEG[10]
rlabel metal3 1418 17748 1418 17748 0 W6BEG[11]
rlabel metal3 1050 15028 1050 15028 0 W6BEG[1]
rlabel metal3 866 15300 866 15300 0 W6BEG[2]
rlabel metal3 1142 15572 1142 15572 0 W6BEG[3]
rlabel metal3 912 15844 912 15844 0 W6BEG[4]
rlabel metal3 498 16116 498 16116 0 W6BEG[5]
rlabel metal3 406 16388 406 16388 0 W6BEG[6]
rlabel metal3 958 16660 958 16660 0 W6BEG[7]
rlabel metal3 866 16932 866 16932 0 W6BEG[8]
rlabel metal3 1142 17204 1142 17204 0 W6BEG[9]
rlabel metal3 1234 10404 1234 10404 0 WW4BEG[0]
rlabel metal3 958 13124 958 13124 0 WW4BEG[10]
rlabel metal3 2062 13396 2062 13396 0 WW4BEG[11]
rlabel metal3 820 13668 820 13668 0 WW4BEG[12]
rlabel metal3 1096 13940 1096 13940 0 WW4BEG[13]
rlabel metal3 199 14212 199 14212 0 WW4BEG[14]
rlabel metal3 199 14484 199 14484 0 WW4BEG[15]
rlabel metal3 590 10676 590 10676 0 WW4BEG[1]
rlabel metal3 498 10948 498 10948 0 WW4BEG[2]
rlabel metal2 4186 10727 4186 10727 0 WW4BEG[3]
rlabel metal3 1050 11492 1050 11492 0 WW4BEG[4]
rlabel metal3 1004 11764 1004 11764 0 WW4BEG[5]
rlabel metal3 866 12036 866 12036 0 WW4BEG[6]
rlabel metal2 1702 11815 1702 11815 0 WW4BEG[7]
rlabel via2 5566 11883 5566 11883 0 WW4BEG[8]
rlabel metal2 4186 12631 4186 12631 0 WW4BEG[9]
rlabel metal1 18584 26486 18584 26486 0 data_inbuf_0.X
rlabel metal1 18860 27098 18860 27098 0 data_inbuf_1.X
rlabel metal2 17158 32963 17158 32963 0 data_inbuf_10.X
rlabel via2 19366 33269 19366 33269 0 data_inbuf_11.X
rlabel metal1 19642 34136 19642 34136 0 data_inbuf_12.X
rlabel metal1 18998 34170 18998 34170 0 data_inbuf_13.X
rlabel metal1 19136 35054 19136 35054 0 data_inbuf_14.X
rlabel metal1 18170 34170 18170 34170 0 data_inbuf_15.X
rlabel metal1 18630 35632 18630 35632 0 data_inbuf_16.X
rlabel metal1 17066 36142 17066 36142 0 data_inbuf_17.X
rlabel metal1 18952 36006 18952 36006 0 data_inbuf_18.X
rlabel metal1 19090 36550 19090 36550 0 data_inbuf_19.X
rlabel metal1 19320 27438 19320 27438 0 data_inbuf_2.X
rlabel metal1 18354 36890 18354 36890 0 data_inbuf_20.X
rlabel metal1 18906 37434 18906 37434 0 data_inbuf_21.X
rlabel metal1 18722 37944 18722 37944 0 data_inbuf_22.X
rlabel metal1 18906 38522 18906 38522 0 data_inbuf_23.X
rlabel metal1 18262 38420 18262 38420 0 data_inbuf_24.X
rlabel metal1 19136 38454 19136 38454 0 data_inbuf_25.X
rlabel metal1 19136 39610 19136 39610 0 data_inbuf_26.X
rlabel metal1 18538 40154 18538 40154 0 data_inbuf_27.X
rlabel metal1 19550 39610 19550 39610 0 data_inbuf_28.X
rlabel metal1 17986 38930 17986 38930 0 data_inbuf_29.X
rlabel metal1 19458 29172 19458 29172 0 data_inbuf_3.X
rlabel metal1 18584 39814 18584 39814 0 data_inbuf_30.X
rlabel metal1 15134 40528 15134 40528 0 data_inbuf_31.X
rlabel metal1 19320 29274 19320 29274 0 data_inbuf_4.X
rlabel metal1 19412 29750 19412 29750 0 data_inbuf_5.X
rlabel metal1 18860 29614 18860 29614 0 data_inbuf_6.X
rlabel metal1 18952 30362 18952 30362 0 data_inbuf_7.X
rlabel metal1 19389 30702 19389 30702 0 data_inbuf_8.X
rlabel metal1 18538 31824 18538 31824 0 data_inbuf_9.X
rlabel metal2 19182 27778 19182 27778 0 data_outbuf_0.X
rlabel metal1 19090 27472 19090 27472 0 data_outbuf_1.X
rlabel metal1 18262 33490 18262 33490 0 data_outbuf_10.X
rlabel metal1 20010 34714 20010 34714 0 data_outbuf_11.X
rlabel metal1 18676 33490 18676 33490 0 data_outbuf_12.X
rlabel metal1 18630 33966 18630 33966 0 data_outbuf_13.X
rlabel metal2 18906 35666 18906 35666 0 data_outbuf_14.X
rlabel metal1 17894 35700 17894 35700 0 data_outbuf_15.X
rlabel metal1 18906 35700 18906 35700 0 data_outbuf_16.X
rlabel metal1 18814 36176 18814 36176 0 data_outbuf_17.X
rlabel metal1 19734 37706 19734 37706 0 data_outbuf_18.X
rlabel metal2 19826 37502 19826 37502 0 data_outbuf_19.X
rlabel metal1 19274 27608 19274 27608 0 data_outbuf_2.X
rlabel metal1 18170 37264 18170 37264 0 data_outbuf_20.X
rlabel metal1 18998 37740 18998 37740 0 data_outbuf_21.X
rlabel metal1 19550 39066 19550 39066 0 data_outbuf_22.X
rlabel metal1 19090 38930 19090 38930 0 data_outbuf_23.X
rlabel metal1 19688 39270 19688 39270 0 data_outbuf_24.X
rlabel metal2 19550 39304 19550 39304 0 data_outbuf_25.X
rlabel metal1 16606 39372 16606 39372 0 data_outbuf_26.X
rlabel metal1 18860 40494 18860 40494 0 data_outbuf_27.X
rlabel metal1 17526 40460 17526 40460 0 data_outbuf_28.X
rlabel metal1 17986 39066 17986 39066 0 data_outbuf_29.X
rlabel metal1 19274 28968 19274 28968 0 data_outbuf_3.X
rlabel metal1 18078 39406 18078 39406 0 data_outbuf_30.X
rlabel via1 18450 38930 18450 38930 0 data_outbuf_31.X
rlabel metal1 19550 30362 19550 30362 0 data_outbuf_4.X
rlabel metal2 17710 30617 17710 30617 0 data_outbuf_5.X
rlabel metal1 18814 29818 18814 29818 0 data_outbuf_6.X
rlabel viali 19090 30703 19090 30703 0 data_outbuf_7.X
rlabel metal2 19274 30991 19274 30991 0 data_outbuf_8.X
rlabel metal1 18492 31994 18492 31994 0 data_outbuf_9.X
rlabel metal3 8188 19176 8188 19176 0 net1
rlabel metal1 2852 23698 2852 23698 0 net10
rlabel metal1 17066 38930 17066 38930 0 net100
rlabel metal1 11040 19414 11040 19414 0 net101
rlabel metal2 598 25772 598 25772 0 net102
rlabel metal1 5014 22678 5014 22678 0 net103
rlabel metal1 12052 8942 12052 8942 0 net104
rlabel via3 9453 29036 9453 29036 0 net105
rlabel metal3 7199 20740 7199 20740 0 net106
rlabel metal3 5796 11016 5796 11016 0 net107
rlabel metal2 17342 33881 17342 33881 0 net108
rlabel via3 10189 34612 10189 34612 0 net109
rlabel metal1 1610 30770 1610 30770 0 net11
rlabel metal2 6348 5236 6348 5236 0 net110
rlabel metal2 7406 4182 7406 4182 0 net111
rlabel metal3 8027 18156 8027 18156 0 net112
rlabel metal1 9890 29512 9890 29512 0 net113
rlabel metal2 782 23868 782 23868 0 net114
rlabel metal1 5796 11730 5796 11730 0 net115
rlabel metal2 10350 34340 10350 34340 0 net116
rlabel metal2 10534 35445 10534 35445 0 net117
rlabel metal1 4186 7820 4186 7820 0 net118
rlabel metal1 4830 4522 4830 4522 0 net119
rlabel metal2 1886 24395 1886 24395 0 net12
rlabel metal2 1380 19380 1380 19380 0 net120
rlabel metal3 4439 10948 4439 10948 0 net121
rlabel metal1 6854 1904 6854 1904 0 net122
rlabel metal1 7498 1360 7498 1360 0 net123
rlabel metal1 7084 1938 7084 1938 0 net124
rlabel metal1 7912 2006 7912 2006 0 net125
rlabel metal1 7866 1938 7866 1938 0 net126
rlabel metal1 8280 1938 8280 1938 0 net127
rlabel metal2 4462 33439 4462 33439 0 net128
rlabel metal1 5244 17646 5244 17646 0 net129
rlabel via1 11730 26282 11730 26282 0 net13
rlabel metal1 12650 12104 12650 12104 0 net130
rlabel metal1 5382 1802 5382 1802 0 net131
rlabel metal1 6026 1224 6026 1224 0 net132
rlabel metal1 6026 2040 6026 2040 0 net133
rlabel metal1 6854 1326 6854 1326 0 net134
rlabel metal1 6486 1972 6486 1972 0 net135
rlabel metal1 6532 1326 6532 1326 0 net136
rlabel metal1 16882 5712 16882 5712 0 net137
rlabel metal1 16422 7888 16422 7888 0 net138
rlabel metal1 15594 8466 15594 8466 0 net139
rlabel metal1 3128 18938 3128 18938 0 net14
rlabel metal1 16238 9520 16238 9520 0 net140
rlabel metal1 13570 5168 13570 5168 0 net141
rlabel metal1 12236 5202 12236 5202 0 net142
rlabel metal1 15134 4794 15134 4794 0 net143
rlabel metal1 18712 7378 18712 7378 0 net144
rlabel metal1 15180 5202 15180 5202 0 net145
rlabel metal1 14623 4182 14623 4182 0 net146
rlabel metal1 13156 3366 13156 3366 0 net147
rlabel metal1 13708 3910 13708 3910 0 net148
rlabel metal1 13248 4454 13248 4454 0 net149
rlabel metal1 3036 18598 3036 18598 0 net15
rlabel metal1 11086 2924 11086 2924 0 net150
rlabel metal1 13110 3468 13110 3468 0 net151
rlabel metal1 13386 4556 13386 4556 0 net152
rlabel metal2 9430 17442 9430 17442 0 net153
rlabel via2 3726 33541 3726 33541 0 net154
rlabel metal1 3772 18326 3772 18326 0 net155
rlabel metal1 12052 19482 12052 19482 0 net156
rlabel metal2 9568 41400 9568 41400 0 net157
rlabel metal3 8165 41684 8165 41684 0 net158
rlabel metal2 5796 41004 5796 41004 0 net159
rlabel via2 2070 18683 2070 18683 0 net16
rlabel metal1 9798 38182 9798 38182 0 net160
rlabel metal1 9936 35802 9936 35802 0 net161
rlabel metal3 9959 39644 9959 39644 0 net162
rlabel metal3 14329 18156 14329 18156 0 net163
rlabel metal2 10304 41400 10304 41400 0 net164
rlabel metal1 8694 29172 8694 29172 0 net165
rlabel metal2 11592 41400 11592 41400 0 net166
rlabel metal2 1334 42613 1334 42613 0 net167
rlabel metal2 11776 41400 11776 41400 0 net168
rlabel metal1 9430 35700 9430 35700 0 net169
rlabel via1 11086 20893 11086 20893 0 net17
rlabel metal2 11776 34068 11776 34068 0 net170
rlabel metal1 12926 43078 12926 43078 0 net171
rlabel metal1 13110 42568 13110 42568 0 net172
rlabel metal2 12512 19516 12512 19516 0 net173
rlabel metal1 14720 42194 14720 42194 0 net174
rlabel metal1 14996 41242 14996 41242 0 net175
rlabel metal2 15226 41327 15226 41327 0 net176
rlabel metal1 16790 42024 16790 42024 0 net177
rlabel metal1 16146 42160 16146 42160 0 net178
rlabel metal2 14444 41820 14444 41820 0 net179
rlabel metal1 8096 7310 8096 7310 0 net18
rlabel metal2 13570 43129 13570 43129 0 net180
rlabel metal2 2346 42579 2346 42579 0 net181
rlabel metal1 13616 42874 13616 42874 0 net182
rlabel metal1 13708 42670 13708 42670 0 net183
rlabel metal1 13938 43248 13938 43248 0 net184
rlabel metal1 14904 42670 14904 42670 0 net185
rlabel metal1 16468 42330 16468 42330 0 net186
rlabel metal1 14766 43282 14766 43282 0 net187
rlabel metal1 15778 42058 15778 42058 0 net188
rlabel metal2 18722 8687 18722 8687 0 net189
rlabel metal1 1794 30634 1794 30634 0 net19
rlabel metal1 11224 5338 11224 5338 0 net190
rlabel metal1 20056 7446 20056 7446 0 net191
rlabel metal2 19688 14892 19688 14892 0 net192
rlabel metal1 19320 15878 19320 15878 0 net193
rlabel metal1 20102 16490 20102 16490 0 net194
rlabel metal1 19872 17170 19872 17170 0 net195
rlabel metal1 20194 17272 20194 17272 0 net196
rlabel metal1 19642 13974 19642 13974 0 net197
rlabel metal1 19550 12954 19550 12954 0 net198
rlabel metal1 19826 15062 19826 15062 0 net199
rlabel metal2 1886 34561 1886 34561 0 net2
rlabel metal2 3634 21913 3634 21913 0 net20
rlabel metal1 20194 15368 20194 15368 0 net200
rlabel metal1 18952 12818 18952 12818 0 net201
rlabel metal1 20516 12750 20516 12750 0 net202
rlabel metal1 18446 12614 18446 12614 0 net203
rlabel metal1 20194 12852 20194 12852 0 net204
rlabel metal1 20010 24718 20010 24718 0 net205
rlabel metal1 19780 27030 19780 27030 0 net206
rlabel metal1 19642 26894 19642 26894 0 net207
rlabel viali 19817 26350 19817 26350 0 net208
rlabel metal1 20332 22678 20332 22678 0 net209
rlabel via2 3082 27931 3082 27931 0 net21
rlabel metal1 20884 23290 20884 23290 0 net210
rlabel metal1 20102 23766 20102 23766 0 net211
rlabel metal1 19826 25874 19826 25874 0 net212
rlabel metal1 20884 37366 20884 37366 0 net213
rlabel metal1 21850 37366 21850 37366 0 net214
rlabel metal1 20148 21522 20148 21522 0 net215
rlabel metal2 20286 21828 20286 21828 0 net216
rlabel metal1 19688 18326 19688 18326 0 net217
rlabel metal1 20654 18666 20654 18666 0 net218
rlabel metal1 19826 19448 19826 19448 0 net219
rlabel metal1 6440 20842 6440 20842 0 net22
rlabel metal2 20148 21964 20148 21964 0 net220
rlabel metal1 20102 27438 20102 27438 0 net221
rlabel metal1 20148 32878 20148 32878 0 net222
rlabel metal1 19734 32844 19734 32844 0 net223
rlabel metal1 20194 33592 20194 33592 0 net224
rlabel metal1 19366 33864 19366 33864 0 net225
rlabel metal1 19872 34646 19872 34646 0 net226
rlabel metal2 18170 35224 18170 35224 0 net227
rlabel metal1 19665 35054 19665 35054 0 net228
rlabel metal1 19412 36346 19412 36346 0 net229
rlabel via1 14042 30226 14042 30226 0 net23
rlabel metal1 19596 37162 19596 37162 0 net230
rlabel metal1 19665 37230 19665 37230 0 net231
rlabel metal1 19274 27370 19274 27370 0 net232
rlabel metal1 19090 37094 19090 37094 0 net233
rlabel metal1 20194 38420 20194 38420 0 net234
rlabel metal1 20148 38998 20148 38998 0 net235
rlabel metal1 18906 39066 18906 39066 0 net236
rlabel metal1 20194 40120 20194 40120 0 net237
rlabel metal1 19642 38760 19642 38760 0 net238
rlabel metal1 16514 39542 16514 39542 0 net239
rlabel metal1 2323 27302 2323 27302 0 net24
rlabel metal1 19044 40698 19044 40698 0 net240
rlabel metal1 17204 40630 17204 40630 0 net241
rlabel metal1 19366 39848 19366 39848 0 net242
rlabel metal1 20010 28118 20010 28118 0 net243
rlabel metal1 17756 39610 17756 39610 0 net244
rlabel metal1 19734 38964 19734 38964 0 net245
rlabel metal1 20148 28526 20148 28526 0 net246
rlabel metal2 20194 29784 20194 29784 0 net247
rlabel metal1 18998 29614 18998 29614 0 net248
rlabel metal1 20194 30260 20194 30260 0 net249
rlabel metal1 3871 22678 3871 22678 0 net25
rlabel metal1 19162 30702 19162 30702 0 net250
rlabel metal1 20194 31416 20194 31416 0 net251
rlabel metal1 18722 31892 18722 31892 0 net252
rlabel metal1 15732 41242 15732 41242 0 net253
rlabel metal1 12972 41718 12972 41718 0 net254
rlabel metal1 13110 42330 13110 42330 0 net255
rlabel metal1 14536 40902 14536 40902 0 net256
rlabel metal1 13662 41786 13662 41786 0 net257
rlabel metal1 17526 40358 17526 40358 0 net258
rlabel metal1 17158 39882 17158 39882 0 net259
rlabel via2 1702 29563 1702 29563 0 net26
rlabel metal1 18170 39610 18170 39610 0 net260
rlabel metal1 17250 40154 17250 40154 0 net261
rlabel metal1 18446 39066 18446 39066 0 net262
rlabel metal1 18170 39270 18170 39270 0 net263
rlabel metal1 18584 41242 18584 41242 0 net264
rlabel metal1 18538 42806 18538 42806 0 net265
rlabel metal2 12190 42109 12190 42109 0 net266
rlabel metal1 18630 42874 18630 42874 0 net267
rlabel metal2 15226 40919 15226 40919 0 net268
rlabel metal1 13800 41718 13800 41718 0 net269
rlabel via2 1702 28475 1702 28475 0 net27
rlabel metal1 17572 41242 17572 41242 0 net270
rlabel metal1 16606 41480 16606 41480 0 net271
rlabel metal1 17572 40154 17572 40154 0 net272
rlabel metal2 1518 43452 1518 43452 0 net273
rlabel metal1 1932 42262 1932 42262 0 net274
rlabel metal1 2990 41786 2990 41786 0 net275
rlabel metal1 2162 42568 2162 42568 0 net276
rlabel metal1 2392 41718 2392 41718 0 net277
rlabel metal1 2530 41786 2530 41786 0 net278
rlabel metal1 2254 42330 2254 42330 0 net279
rlabel metal1 1656 31314 1656 31314 0 net28
rlabel metal1 3772 41242 3772 41242 0 net280
rlabel metal1 3358 41786 3358 41786 0 net281
rlabel metal1 3404 41242 3404 41242 0 net282
rlabel metal2 3174 42160 3174 42160 0 net283
rlabel metal2 12650 42160 12650 42160 0 net284
rlabel metal1 1794 42772 1794 42772 0 net285
rlabel metal2 4002 41321 4002 41321 0 net286
rlabel metal1 4094 41718 4094 41718 0 net287
rlabel metal1 4600 41242 4600 41242 0 net288
rlabel metal1 5060 41242 5060 41242 0 net289
rlabel metal1 1748 30158 1748 30158 0 net29
rlabel metal1 5106 40970 5106 40970 0 net290
rlabel metal1 5152 41786 5152 41786 0 net291
rlabel metal2 3726 42466 3726 42466 0 net292
rlabel metal1 5704 42602 5704 42602 0 net293
rlabel metal1 9246 42296 9246 42296 0 net294
rlabel metal1 8280 41786 8280 41786 0 net295
rlabel metal1 9614 42704 9614 42704 0 net296
rlabel metal2 8970 42738 8970 42738 0 net297
rlabel metal1 8694 41718 8694 41718 0 net298
rlabel metal1 9890 42568 9890 42568 0 net299
rlabel metal1 2530 29750 2530 29750 0 net3
rlabel via2 2622 28611 2622 28611 0 net30
rlabel metal2 4186 42534 4186 42534 0 net300
rlabel metal1 6348 42602 6348 42602 0 net301
rlabel metal1 5842 41616 5842 41616 0 net302
rlabel metal1 5934 40970 5934 40970 0 net303
rlabel metal1 6302 42670 6302 42670 0 net304
rlabel metal1 7084 42670 7084 42670 0 net305
rlabel metal1 6808 41242 6808 41242 0 net306
rlabel metal1 6900 42262 6900 42262 0 net307
rlabel metal1 7544 41786 7544 41786 0 net308
rlabel metal2 7866 1564 7866 1564 0 net309
rlabel metal2 9200 28220 9200 28220 0 net31
rlabel metal1 8510 2380 8510 2380 0 net310
rlabel metal1 8786 2040 8786 2040 0 net311
rlabel metal2 11822 2091 11822 2091 0 net312
rlabel metal1 11224 2278 11224 2278 0 net313
rlabel metal2 11454 2516 11454 2516 0 net314
rlabel metal1 10534 1870 10534 1870 0 net315
rlabel metal1 11822 1870 11822 1870 0 net316
rlabel metal1 12834 2618 12834 2618 0 net317
rlabel metal1 11132 2550 11132 2550 0 net318
rlabel metal2 12926 935 12926 935 0 net319
rlabel via1 7843 38862 7843 38862 0 net32
rlabel metal1 14858 1836 14858 1836 0 net320
rlabel metal1 9384 2890 9384 2890 0 net321
rlabel metal1 8418 1394 8418 1394 0 net322
rlabel metal1 9752 1938 9752 1938 0 net323
rlabel metal1 9614 2448 9614 2448 0 net324
rlabel metal1 10442 1904 10442 1904 0 net325
rlabel metal1 9108 1326 9108 1326 0 net326
rlabel metal1 10166 2006 10166 2006 0 net327
rlabel metal1 9476 1258 9476 1258 0 net328
rlabel metal2 14122 1666 14122 1666 0 net329
rlabel metal1 8050 23800 8050 23800 0 net33
rlabel metal1 11868 2006 11868 2006 0 net330
rlabel metal1 15042 3026 15042 3026 0 net331
rlabel metal1 14904 4114 14904 4114 0 net332
rlabel metal1 15640 3094 15640 3094 0 net333
rlabel metal3 11132 4896 11132 4896 0 net334
rlabel via2 15870 3485 15870 3485 0 net335
rlabel metal1 13248 2006 13248 2006 0 net336
rlabel metal2 17802 1054 17802 1054 0 net337
rlabel metal1 13570 2448 13570 2448 0 net338
rlabel metal1 13837 2006 13837 2006 0 net339
rlabel metal2 4830 26758 4830 26758 0 net34
rlabel metal2 13938 646 13938 646 0 net340
rlabel metal1 14490 2006 14490 2006 0 net341
rlabel metal1 14029 3026 14029 3026 0 net342
rlabel metal1 19274 2346 19274 2346 0 net343
rlabel metal1 17204 2346 17204 2346 0 net344
rlabel metal1 16100 40494 16100 40494 0 net345
rlabel metal2 7314 4097 7314 4097 0 net346
rlabel metal2 6486 6086 6486 6086 0 net347
rlabel metal1 4554 3706 4554 3706 0 net348
rlabel metal2 6854 3961 6854 3961 0 net349
rlabel metal1 13616 28526 13616 28526 0 net35
rlabel metal1 5290 4726 5290 4726 0 net350
rlabel metal1 4370 4216 4370 4216 0 net351
rlabel metal2 4094 5066 4094 5066 0 net352
rlabel metal1 2944 5338 2944 5338 0 net353
rlabel metal2 3358 5372 3358 5372 0 net354
rlabel metal1 4370 6664 4370 6664 0 net355
rlabel metal1 4278 3944 4278 3944 0 net356
rlabel metal1 11546 7480 11546 7480 0 net357
rlabel metal2 13938 7327 13938 7327 0 net358
rlabel metal1 5290 6936 5290 6936 0 net359
rlabel metal1 5106 27098 5106 27098 0 net36
rlabel metal1 2024 4794 2024 4794 0 net360
rlabel metal2 4554 7854 4554 7854 0 net361
rlabel metal1 4462 6698 4462 6698 0 net362
rlabel metal2 1978 4862 1978 4862 0 net363
rlabel metal1 4462 8976 4462 8976 0 net364
rlabel metal2 4738 7786 4738 7786 0 net365
rlabel metal1 1748 11730 1748 11730 0 net366
rlabel metal1 2254 16218 2254 16218 0 net367
rlabel metal2 1518 16592 1518 16592 0 net368
rlabel metal4 1656 22080 1656 22080 0 net369
rlabel metal2 1886 32232 1886 32232 0 net37
rlabel metal1 1702 13226 1702 13226 0 net370
rlabel metal1 4002 15334 4002 15334 0 net371
rlabel metal1 4370 15368 4370 15368 0 net372
rlabel metal1 1656 12954 1656 12954 0 net373
rlabel metal1 1794 14314 1794 14314 0 net374
rlabel metal2 3082 15266 3082 15266 0 net375
rlabel metal1 1610 16150 1610 16150 0 net376
rlabel metal1 2576 17646 2576 17646 0 net377
rlabel metal2 4370 9418 4370 9418 0 net378
rlabel via2 6394 12699 6394 12699 0 net379
rlabel metal1 4048 25126 4048 25126 0 net38
rlabel metal2 4462 13464 4462 13464 0 net380
rlabel metal1 1564 10234 1564 10234 0 net381
rlabel metal2 4370 13056 4370 13056 0 net382
rlabel metal1 3174 12886 3174 12886 0 net383
rlabel metal1 4462 12920 4462 12920 0 net384
rlabel metal1 2070 8568 2070 8568 0 net385
rlabel metal1 1840 6358 1840 6358 0 net386
rlabel metal1 2024 7514 2024 7514 0 net387
rlabel metal2 4830 9435 4830 9435 0 net388
rlabel metal2 1518 7718 1518 7718 0 net389
rlabel metal3 14674 31756 14674 31756 0 net39
rlabel metal2 2070 9962 2070 9962 0 net390
rlabel metal1 4830 10506 4830 10506 0 net391
rlabel metal2 5382 10710 5382 10710 0 net392
rlabel metal1 4370 12104 4370 12104 0 net393
rlabel metal1 12466 19448 12466 19448 0 net394
rlabel metal1 13110 21114 13110 21114 0 net395
rlabel metal1 1886 20910 1886 20910 0 net396
rlabel metal2 8602 19652 8602 19652 0 net397
rlabel metal2 12374 35054 12374 35054 0 net398
rlabel via1 11831 20910 11831 20910 0 net399
rlabel metal2 13018 33116 13018 33116 0 net4
rlabel metal1 3588 24038 3588 24038 0 net40
rlabel metal1 9154 6358 9154 6358 0 net400
rlabel metal1 7498 27030 7498 27030 0 net401
rlabel metal2 13938 27030 13938 27030 0 net402
rlabel metal2 15870 18938 15870 18938 0 net403
rlabel metal2 8786 37196 8786 37196 0 net404
rlabel metal2 5014 22039 5014 22039 0 net405
rlabel metal1 10074 19448 10074 19448 0 net406
rlabel metal1 3358 37842 3358 37842 0 net407
rlabel metal1 4232 22202 4232 22202 0 net408
rlabel metal2 14858 19550 14858 19550 0 net409
rlabel metal1 5336 29614 5336 29614 0 net41
rlabel via2 2530 24667 2530 24667 0 net42
rlabel metal1 14306 23154 14306 23154 0 net43
rlabel metal1 1656 26010 1656 26010 0 net44
rlabel metal1 4462 25262 4462 25262 0 net45
rlabel metal1 14214 33354 14214 33354 0 net46
rlabel metal1 6026 26282 6026 26282 0 net47
rlabel metal2 6578 35173 6578 35173 0 net48
rlabel via1 1793 26350 1793 26350 0 net49
rlabel via2 12098 21539 12098 21539 0 net5
rlabel via1 5197 25874 5197 25874 0 net50
rlabel metal2 2346 35292 2346 35292 0 net51
rlabel metal1 20561 21998 20561 21998 0 net52
rlabel metal1 4967 13294 4967 13294 0 net53
rlabel via1 6761 35054 6761 35054 0 net54
rlabel metal1 16790 19482 16790 19482 0 net55
rlabel metal1 16145 14382 16145 14382 0 net56
rlabel viali 6660 21552 6660 21552 0 net57
rlabel via1 19549 25262 19549 25262 0 net58
rlabel via1 1885 20434 1885 20434 0 net59
rlabel metal1 2438 21454 2438 21454 0 net6
rlabel metal2 2254 31892 2254 31892 0 net60
rlabel metal2 18170 36703 18170 36703 0 net61
rlabel metal1 18906 37230 18906 37230 0 net62
rlabel metal2 17296 26962 17296 26962 0 net63
rlabel metal1 5290 38420 5290 38420 0 net64
rlabel via1 11821 6290 11821 6290 0 net65
rlabel metal1 9430 39406 9430 39406 0 net66
rlabel metal1 2115 21522 2115 21522 0 net67
rlabel metal2 782 18938 782 18938 0 net68
rlabel metal1 2162 40970 2162 40970 0 net69
rlabel metal1 7866 21658 7866 21658 0 net7
rlabel via2 2714 40443 2714 40443 0 net70
rlabel metal1 2530 18054 2530 18054 0 net71
rlabel metal2 12466 39644 12466 39644 0 net72
rlabel metal1 14075 11730 14075 11730 0 net73
rlabel metal1 644 21386 644 21386 0 net74
rlabel metal2 3864 25738 3864 25738 0 net75
rlabel metal1 1702 34102 1702 34102 0 net76
rlabel metal2 17618 29512 17618 29512 0 net77
rlabel via3 5221 23868 5221 23868 0 net78
rlabel metal2 2484 34612 2484 34612 0 net79
rlabel metal2 1702 20451 1702 20451 0 net8
rlabel metal1 6762 33864 6762 33864 0 net80
rlabel metal1 2530 38862 2530 38862 0 net81
rlabel metal1 19182 5746 19182 5746 0 net82
rlabel metal4 15548 2448 15548 2448 0 net83
rlabel metal1 16330 2516 16330 2516 0 net84
rlabel via2 16330 3077 16330 3077 0 net85
rlabel metal1 12144 2890 12144 2890 0 net86
rlabel metal1 17940 3026 17940 3026 0 net87
rlabel metal1 11546 2822 11546 2822 0 net88
rlabel metal1 12190 3706 12190 3706 0 net89
rlabel metal1 10764 20978 10764 20978 0 net9
rlabel metal1 11546 2890 11546 2890 0 net90
rlabel metal1 18262 6392 18262 6392 0 net91
rlabel metal3 16399 1292 16399 1292 0 net92
rlabel metal1 12466 40052 12466 40052 0 net93
rlabel metal2 5934 37536 5934 37536 0 net94
rlabel metal2 16928 39508 16928 39508 0 net95
rlabel metal1 15502 9078 15502 9078 0 net96
rlabel metal1 16698 40494 16698 40494 0 net97
rlabel metal2 8188 28390 8188 28390 0 net98
rlabel metal1 17434 13430 17434 13430 0 net99
rlabel metal1 15502 39610 15502 39610 0 strobe_inbuf_0.X
rlabel metal1 15732 40698 15732 40698 0 strobe_inbuf_1.X
rlabel metal1 17342 20774 17342 20774 0 strobe_inbuf_10.X
rlabel metal3 20401 20876 20401 20876 0 strobe_inbuf_11.X
rlabel via3 16997 40052 16997 40052 0 strobe_inbuf_12.X
rlabel via3 17181 38692 17181 38692 0 strobe_inbuf_13.X
rlabel metal3 18032 15028 18032 15028 0 strobe_inbuf_14.X
rlabel metal1 17710 21114 17710 21114 0 strobe_inbuf_15.X
rlabel metal1 20286 19686 20286 19686 0 strobe_inbuf_16.X
rlabel metal3 20539 18292 20539 18292 0 strobe_inbuf_17.X
rlabel metal3 18055 40052 18055 40052 0 strobe_inbuf_18.X
rlabel metal2 21252 33660 21252 33660 0 strobe_inbuf_19.X
rlabel metal1 15916 40970 15916 40970 0 strobe_inbuf_2.X
rlabel metal1 16284 41242 16284 41242 0 strobe_inbuf_3.X
rlabel metal1 16836 41242 16836 41242 0 strobe_inbuf_4.X
rlabel metal1 16468 15130 16468 15130 0 strobe_inbuf_5.X
rlabel metal1 16606 40698 16606 40698 0 strobe_inbuf_6.X
rlabel metal2 19044 39474 19044 39474 0 strobe_inbuf_7.X
rlabel metal1 17066 40698 17066 40698 0 strobe_inbuf_8.X
rlabel metal1 17250 39066 17250 39066 0 strobe_inbuf_9.X
rlabel metal2 15502 40868 15502 40868 0 strobe_outbuf_0.X
rlabel metal2 19090 41276 19090 41276 0 strobe_outbuf_1.X
rlabel metal1 16928 40902 16928 40902 0 strobe_outbuf_10.X
rlabel metal1 12926 42228 12926 42228 0 strobe_outbuf_11.X
rlabel metal1 16790 40154 16790 40154 0 strobe_outbuf_12.X
rlabel metal1 16376 39610 16376 39610 0 strobe_outbuf_13.X
rlabel metal2 17802 40732 17802 40732 0 strobe_outbuf_14.X
rlabel metal1 17296 39542 17296 39542 0 strobe_outbuf_15.X
rlabel metal1 20194 39542 20194 39542 0 strobe_outbuf_16.X
rlabel metal1 17342 40052 17342 40052 0 strobe_outbuf_17.X
rlabel metal1 18722 38964 18722 38964 0 strobe_outbuf_18.X
rlabel metal1 17710 39440 17710 39440 0 strobe_outbuf_19.X
rlabel metal1 19780 40562 19780 40562 0 strobe_outbuf_2.X
rlabel metal1 16238 41480 16238 41480 0 strobe_outbuf_3.X
rlabel metal2 16882 42058 16882 42058 0 strobe_outbuf_4.X
rlabel metal2 16468 41140 16468 41140 0 strobe_outbuf_5.X
rlabel metal1 13938 41650 13938 41650 0 strobe_outbuf_6.X
rlabel metal1 17802 41072 17802 41072 0 strobe_outbuf_7.X
rlabel metal1 17066 41208 17066 41208 0 strobe_outbuf_8.X
rlabel metal1 17434 39610 17434 39610 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 22000 44700
<< end >>
