* NGSPICE file created from DSP.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__dlxbp_1 abstract view
.subckt sky130_fd_sc_hd__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_2 abstract view
.subckt sky130_fd_sc_hd__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311ai_4 abstract view
.subckt sky130_fd_sc_hd__o311ai_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

.subckt DSP Tile_X0Y0_E1BEG[0] Tile_X0Y0_E1BEG[1] Tile_X0Y0_E1BEG[2] Tile_X0Y0_E1BEG[3]
+ Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2BEG[0]
+ Tile_X0Y0_E2BEG[1] Tile_X0Y0_E2BEG[2] Tile_X0Y0_E2BEG[3] Tile_X0Y0_E2BEG[4] Tile_X0Y0_E2BEG[5]
+ Tile_X0Y0_E2BEG[6] Tile_X0Y0_E2BEG[7] Tile_X0Y0_E2BEGb[0] Tile_X0Y0_E2BEGb[1] Tile_X0Y0_E2BEGb[2]
+ Tile_X0Y0_E2BEGb[3] Tile_X0Y0_E2BEGb[4] Tile_X0Y0_E2BEGb[5] Tile_X0Y0_E2BEGb[6]
+ Tile_X0Y0_E2BEGb[7] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6BEG[0] Tile_X0Y0_E6BEG[10] Tile_X0Y0_E6BEG[11]
+ Tile_X0Y0_E6BEG[1] Tile_X0Y0_E6BEG[2] Tile_X0Y0_E6BEG[3] Tile_X0Y0_E6BEG[4] Tile_X0Y0_E6BEG[5]
+ Tile_X0Y0_E6BEG[6] Tile_X0Y0_E6BEG[7] Tile_X0Y0_E6BEG[8] Tile_X0Y0_E6BEG[9] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4BEG[0] Tile_X0Y0_EE4BEG[10] Tile_X0Y0_EE4BEG[11]
+ Tile_X0Y0_EE4BEG[12] Tile_X0Y0_EE4BEG[13] Tile_X0Y0_EE4BEG[14] Tile_X0Y0_EE4BEG[15]
+ Tile_X0Y0_EE4BEG[1] Tile_X0Y0_EE4BEG[2] Tile_X0Y0_EE4BEG[3] Tile_X0Y0_EE4BEG[4]
+ Tile_X0Y0_EE4BEG[5] Tile_X0Y0_EE4BEG[6] Tile_X0Y0_EE4BEG[7] Tile_X0Y0_EE4BEG[8]
+ Tile_X0Y0_EE4BEG[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_NN4BEG[0] Tile_X0Y0_NN4BEG[10] Tile_X0Y0_NN4BEG[11]
+ Tile_X0Y0_NN4BEG[12] Tile_X0Y0_NN4BEG[13] Tile_X0Y0_NN4BEG[14] Tile_X0Y0_NN4BEG[15]
+ Tile_X0Y0_NN4BEG[1] Tile_X0Y0_NN4BEG[2] Tile_X0Y0_NN4BEG[3] Tile_X0Y0_NN4BEG[4]
+ Tile_X0Y0_NN4BEG[5] Tile_X0Y0_NN4BEG[6] Tile_X0Y0_NN4BEG[7] Tile_X0Y0_NN4BEG[8]
+ Tile_X0Y0_NN4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3]
+ Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4]
+ Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1]
+ Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6]
+ Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12]
+ Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7]
+ Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_SS4END[0] Tile_X0Y0_SS4END[10] Tile_X0Y0_SS4END[11]
+ Tile_X0Y0_SS4END[12] Tile_X0Y0_SS4END[13] Tile_X0Y0_SS4END[14] Tile_X0Y0_SS4END[15]
+ Tile_X0Y0_SS4END[1] Tile_X0Y0_SS4END[2] Tile_X0Y0_SS4END[3] Tile_X0Y0_SS4END[4]
+ Tile_X0Y0_SS4END[5] Tile_X0Y0_SS4END[6] Tile_X0Y0_SS4END[7] Tile_X0Y0_SS4END[8]
+ Tile_X0Y0_SS4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[1] Tile_X0Y0_W1END[2] Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4]
+ Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1]
+ Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5]
+ Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W2END[0] Tile_X0Y0_W2END[1] Tile_X0Y0_W2END[2]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W2END[4] Tile_X0Y0_W2END[5] Tile_X0Y0_W2END[6] Tile_X0Y0_W2END[7]
+ Tile_X0Y0_W2MID[0] Tile_X0Y0_W2MID[1] Tile_X0Y0_W2MID[2] Tile_X0Y0_W2MID[3] Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2MID[5] Tile_X0Y0_W2MID[6] Tile_X0Y0_W2MID[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_W6END[0] Tile_X0Y0_W6END[10] Tile_X0Y0_W6END[11] Tile_X0Y0_W6END[1] Tile_X0Y0_W6END[2]
+ Tile_X0Y0_W6END[3] Tile_X0Y0_W6END[4] Tile_X0Y0_W6END[5] Tile_X0Y0_W6END[6] Tile_X0Y0_W6END[7]
+ Tile_X0Y0_W6END[8] Tile_X0Y0_W6END[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11]
+ Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15]
+ Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4]
+ Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8]
+ Tile_X0Y0_WW4BEG[9] Tile_X0Y0_WW4END[0] Tile_X0Y0_WW4END[10] Tile_X0Y0_WW4END[11]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_WW4END[13] Tile_X0Y0_WW4END[14] Tile_X0Y0_WW4END[15]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_WW4END[2] Tile_X0Y0_WW4END[3] Tile_X0Y0_WW4END[4]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_WW4END[6] Tile_X0Y0_WW4END[7] Tile_X0Y0_WW4END[8]
+ Tile_X0Y0_WW4END[9] Tile_X0Y1_E1BEG[0] Tile_X0Y1_E1BEG[1] Tile_X0Y1_E1BEG[2] Tile_X0Y1_E1BEG[3]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2BEG[0]
+ Tile_X0Y1_E2BEG[1] Tile_X0Y1_E2BEG[2] Tile_X0Y1_E2BEG[3] Tile_X0Y1_E2BEG[4] Tile_X0Y1_E2BEG[5]
+ Tile_X0Y1_E2BEG[6] Tile_X0Y1_E2BEG[7] Tile_X0Y1_E2BEGb[0] Tile_X0Y1_E2BEGb[1] Tile_X0Y1_E2BEGb[2]
+ Tile_X0Y1_E2BEGb[3] Tile_X0Y1_E2BEGb[4] Tile_X0Y1_E2BEGb[5] Tile_X0Y1_E2BEGb[6]
+ Tile_X0Y1_E2BEGb[7] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6BEG[0] Tile_X0Y1_E6BEG[10] Tile_X0Y1_E6BEG[11]
+ Tile_X0Y1_E6BEG[1] Tile_X0Y1_E6BEG[2] Tile_X0Y1_E6BEG[3] Tile_X0Y1_E6BEG[4] Tile_X0Y1_E6BEG[5]
+ Tile_X0Y1_E6BEG[6] Tile_X0Y1_E6BEG[7] Tile_X0Y1_E6BEG[8] Tile_X0Y1_E6BEG[9] Tile_X0Y1_E6END[0]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3]
+ Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_EE4BEG[0] Tile_X0Y1_EE4BEG[10] Tile_X0Y1_EE4BEG[11]
+ Tile_X0Y1_EE4BEG[12] Tile_X0Y1_EE4BEG[13] Tile_X0Y1_EE4BEG[14] Tile_X0Y1_EE4BEG[15]
+ Tile_X0Y1_EE4BEG[1] Tile_X0Y1_EE4BEG[2] Tile_X0Y1_EE4BEG[3] Tile_X0Y1_EE4BEG[4]
+ Tile_X0Y1_EE4BEG[5] Tile_X0Y1_EE4BEG[6] Tile_X0Y1_EE4BEG[7] Tile_X0Y1_EE4BEG[8]
+ Tile_X0Y1_EE4BEG[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_NN4END[0]
+ Tile_X0Y1_NN4END[10] Tile_X0Y1_NN4END[11] Tile_X0Y1_NN4END[12] Tile_X0Y1_NN4END[13]
+ Tile_X0Y1_NN4END[14] Tile_X0Y1_NN4END[15] Tile_X0Y1_NN4END[1] Tile_X0Y1_NN4END[2]
+ Tile_X0Y1_NN4END[3] Tile_X0Y1_NN4END[4] Tile_X0Y1_NN4END[5] Tile_X0Y1_NN4END[6]
+ Tile_X0Y1_NN4END[7] Tile_X0Y1_NN4END[8] Tile_X0Y1_NN4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1]
+ Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2]
+ Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7]
+ Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_SS4BEG[0] Tile_X0Y1_SS4BEG[10] Tile_X0Y1_SS4BEG[11]
+ Tile_X0Y1_SS4BEG[12] Tile_X0Y1_SS4BEG[13] Tile_X0Y1_SS4BEG[14] Tile_X0Y1_SS4BEG[15]
+ Tile_X0Y1_SS4BEG[1] Tile_X0Y1_SS4BEG[2] Tile_X0Y1_SS4BEG[3] Tile_X0Y1_SS4BEG[4]
+ Tile_X0Y1_SS4BEG[5] Tile_X0Y1_SS4BEG[6] Tile_X0Y1_SS4BEG[7] Tile_X0Y1_SS4BEG[8]
+ Tile_X0Y1_SS4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[1] Tile_X0Y1_W1END[2] Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4]
+ Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1]
+ Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5]
+ Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W2END[0] Tile_X0Y1_W2END[1] Tile_X0Y1_W2END[2]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W2END[4] Tile_X0Y1_W2END[5] Tile_X0Y1_W2END[6] Tile_X0Y1_W2END[7]
+ Tile_X0Y1_W2MID[0] Tile_X0Y1_W2MID[1] Tile_X0Y1_W2MID[2] Tile_X0Y1_W2MID[3] Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2MID[5] Tile_X0Y1_W2MID[6] Tile_X0Y1_W2MID[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[10] Tile_X0Y1_W6END[11] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[2]
+ Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[4] Tile_X0Y1_W6END[5] Tile_X0Y1_W6END[6] Tile_X0Y1_W6END[7]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W6END[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11]
+ Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15]
+ Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4]
+ Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8]
+ Tile_X0Y1_WW4BEG[9] Tile_X0Y1_WW4END[0] Tile_X0Y1_WW4END[10] Tile_X0Y1_WW4END[11]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[15]
+ Tile_X0Y1_WW4END[1] Tile_X0Y1_WW4END[2] Tile_X0Y1_WW4END[3] Tile_X0Y1_WW4END[4]
+ Tile_X0Y1_WW4END[5] Tile_X0Y1_WW4END[6] Tile_X0Y1_WW4END[7] Tile_X0Y1_WW4END[8]
+ Tile_X0Y1_WW4END[9] VGND VPWR
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6 net257 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[198\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[379\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12 net232 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[364\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23 net244 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[375\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.S4END_inbuf_7._0_ Tile_X0Y0_DSP_top.S4BEG\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG_i\[7\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[96\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[107\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_32_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._27_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID3
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 sky130_fd_sc_hd__clkbuf_1
XANTENNA_224 Tile_X0Y0_DSP_top.S4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_202 Tile_X0Y1_DSP_bot.SS4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_213 net309 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_363_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 VGND VGND VPWR VPWR net737
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1590_ Tile_X0Y1_DSP_bot.Inst_MULADD._0733_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0754_ sky130_fd_sc_hd__inv_2
X_294_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb2 VGND VGND VPWR VPWR net677
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1024_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\] Tile_X0Y1_DSP_bot.Inst_MULADD._0191_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0196_ Tile_X0Y1_DSP_bot.Inst_MULADD._0070_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0197_ sky130_fd_sc_hd__o211a_2
XFILLER_0_155_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput401 net401 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_112_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput434 net434 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput412 net412 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput423 net423 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput467 net467 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[14] sky130_fd_sc_hd__clkbuf_4
Xoutput478 net478 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[6] sky130_fd_sc_hd__clkbuf_4
Xoutput445 net445 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[23] sky130_fd_sc_hd__clkbuf_4
Xoutput456 net456 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[4] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16 net236 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[272\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27 net248 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[283\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput489 net489 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._89_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q13
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 sky130_fd_sc_hd__buf_12
XFILLER_0_69_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_147_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[27\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_60_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[330\] Tile_X0Y0_DSP_top.ConfigBits\[331\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_130_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.strobe_inbuf_3._0_ Tile_X0Y0_DSP_top.FrameStrobe\[3\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7 net258 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[39\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1711_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0005_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_346_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb2 VGND VGND VPWR VPWR net729
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1642_ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0801_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0803_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_83_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_396 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1573_ Tile_X0Y1_DSP_bot.C13 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[13\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0738_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_277_ Tile_X0Y1_DSP_bot.FrameData_O\[29\] VGND VGND VPWR VPWR net652 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._12_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot8
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C10 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11 net231 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[395\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22 net243 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[406\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1007_ Tile_X0Y1_DSP_bot.Inst_MULADD._0179_ Tile_X0Y1_DSP_bot.Inst_MULADD._0180_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0181_ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[138\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_91_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[149\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_148_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[256\] Tile_X0Y0_DSP_top.ConfigBits\[257\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_129_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9 net260 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[297\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst0
+ net286 net308 net184 net186 Tile_X0Y1_DSP_bot.ConfigBits\[256\] Tile_X0Y1_DSP_bot.ConfigBits\[257\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[182\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.SS4END_inbuf_2._0_ Tile_X0Y0_DSP_top.SS4BEG\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_200_ Tile_X0Y1_DSP_bot.E1BEG\[0\] VGND VGND VPWR VPWR net583 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_131_ Tile_X0Y0_DSP_top.N4BEG\[11\] VGND VGND VPWR VPWR net504 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_inst0
+ net284 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3 net337 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[101\] Tile_X0Y1_DSP_bot.ConfigBits\[102\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_062_ Tile_X0Y0_DSP_top.FrameData_O\[14\] VGND VGND VPWR VPWR net435 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15 net235 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[303\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26 net247 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[314\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_126_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_329_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR net703
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1625_ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.ConfigBits\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0787_ sky130_fd_sc_hd__nand2_2
XFILLER_0_83_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1556_ Tile_X0Y1_DSP_bot.Inst_MULADD._0720_ Tile_X0Y1_DSP_bot.Inst_MULADD._0721_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1487_ Tile_X0Y1_DSP_bot.Inst_MULADD._0646_ Tile_X0Y1_DSP_bot.Inst_MULADD._0649_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0650_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0654_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID6
+ net19 net151 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 Tile_X0Y0_DSP_top.ConfigBits\[166\]
+ Tile_X0Y0_DSP_top.ConfigBits\[167\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[294\] Tile_X0Y0_DSP_top.ConfigBits\[295\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.data_outbuf_7._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[7\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.EE4END_inbuf_1._0_ net224 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_38_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[33\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_114_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 VGND VGND VPWR VPWR net496
+ sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top.strobe_inbuf_10._0_ Tile_X0Y0_DSP_top.FrameStrobe\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[10\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[278\] Tile_X0Y1_DSP_bot.ConfigBits\[279\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG5 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1410_ Tile_X0Y1_DSP_bot.Inst_MULADD._0575_ Tile_X0Y1_DSP_bot.Inst_MULADD._0576_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0578_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0579_
+ sky130_fd_sc_hd__o21bai_2
XFILLER_0_80_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_045_ Tile_X0Y0_DSP_top.EE4BEG\[13\] VGND VGND VPWR VPWR net418 sky130_fd_sc_hd__buf_1
XFILLER_0_123_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.WW4END_inbuf_9._0_ net169 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1341_ Tile_X0Y1_DSP_bot.Inst_MULADD._0504_ Tile_X0Y1_DSP_bot.Inst_MULADD._0510_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0511_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[180\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19 net239 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[211\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1272_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ Tile_X0Y1_DSP_bot.Inst_MULADD._0359_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0441_ Tile_X0Y1_DSP_bot.Inst_MULADD._0366_ Tile_X0Y1_DSP_bot.Inst_MULADD._0368_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0442_ sky130_fd_sc_hd__o32ai_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._0987_ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0138_ Tile_X0Y1_DSP_bot.Inst_MULADD._0146_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0161_ sky130_fd_sc_hd__a22o_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID3
+ net16 net96 net148 Tile_X0Y0_DSP_top.ConfigBits\[208\] Tile_X0Y0_DSP_top.ConfigBits\[209\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_112_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1608_ Tile_X0Y1_DSP_bot.Inst_MULADD._0765_ Tile_X0Y1_DSP_bot.Inst_MULADD._0771_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0428_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0772_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_141_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1539_ Tile_X0Y1_DSP_bot.Inst_MULADD._0137_ Tile_X0Y1_DSP_bot.Inst_MULADD._0351_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0704_ Tile_X0Y1_DSP_bot.Inst_MULADD._0656_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0705_ sky130_fd_sc_hd__o31a_1
XFILLER_0_141_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._60_ net149 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb4
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4 net255 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[100\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[281\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.data_outbuf_7._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[7\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.strobe_outbuf_12._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[12\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[12\] sky130_fd_sc_hd__buf_6
Xinput301 Tile_X0Y1_N4END[0] VGND VGND VPWR VPWR net301 sky130_fd_sc_hd__clkbuf_2
Xinput312 Tile_X0Y1_N4END[5] VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14 net234 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[334\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25 net246 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[345\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput345 Tile_X0Y1_W2END[7] VGND VGND VPWR VPWR net345 sky130_fd_sc_hd__clkbuf_4
Xinput334 Tile_X0Y1_W1END[0] VGND VGND VPWR VPWR net334 sky130_fd_sc_hd__buf_4
Xinput323 Tile_X0Y1_NN4END[15] VGND VGND VPWR VPWR net323 sky130_fd_sc_hd__clkbuf_1
Xinput367 Tile_X0Y1_WW4END[10] VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__clkbuf_1
Xinput378 Tile_X0Y1_WW4END[6] VGND VGND VPWR VPWR net378 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.ConfigBits\[316\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[317\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
Xinput356 Tile_X0Y1_W6END[11] VGND VGND VPWR VPWR net356 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0910_ Tile_X0Y1_DSP_bot.ConfigBits\[2\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.E6BEG_outbuf_5._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_5 Tile_X0Y0_DSP_top.FrameStrobe\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_028_ Tile_X0Y0_DSP_top.E6BEG\[8\] VGND VGND VPWR VPWR net412 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1324_ Tile_X0Y1_DSP_bot.Inst_MULADD._0436_ Tile_X0Y1_DSP_bot.Inst_MULADD._0492_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0493_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0494_
+ sky130_fd_sc_hd__nand3_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1255_ Tile_X0Y1_DSP_bot.Inst_MULADD._0341_ Tile_X0Y1_DSP_bot.Inst_MULADD._0425_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0426_ sky130_fd_sc_hd__xor2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_W1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG1 Tile_X0Y0_DSP_top.ConfigBits\[84\]
+ Tile_X0Y0_DSP_top.ConfigBits\[85\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1186_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.Inst_MULADD._0355_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0356_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0357_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.strobe_outbuf_8._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[8\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._43_ net96 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb3
+ sky130_fd_sc_hd__clkbuf_2
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29 net250 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[253\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18 net238 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[242\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_79_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[366\] Tile_X0Y0_DSP_top.ConfigBits\[367\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput120 Tile_X0Y0_SS4END[12] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1040_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ Tile_X0Y1_DSP_bot.Inst_MULADD._0211_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0212_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0213_
+ sky130_fd_sc_hd__o21ai_2
Xinput131 Tile_X0Y0_SS4END[8] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_1
Xinput153 Tile_X0Y0_W6END[0] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
Xinput142 Tile_X0Y0_W2END[5] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__clkbuf_2
Xinput164 Tile_X0Y0_W6END[9] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
Xinput175 Tile_X0Y0_WW4END[4] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.strobe_outbuf_1._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[1\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[1\] sky130_fd_sc_hd__buf_8
Xinput186 Tile_X0Y1_E2END[1] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_2
Xinput197 Tile_X0Y1_E2MID[4] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__buf_2
XFILLER_0_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_143_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
Xoutput627 net627 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput616 net616 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput605 net605 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput638 net638 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[16] sky130_fd_sc_hd__buf_2
Xoutput649 net649 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[26] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1307_ Tile_X0Y1_DSP_bot.Inst_MULADD._0461_ Tile_X0Y1_DSP_bot.Inst_MULADD._0467_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0476_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0477_
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y0_DSP_top.WW4BEG_outbuf_6._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[6\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1238_ Tile_X0Y1_DSP_bot.Inst_MULADD._0408_ Tile_X0Y1_DSP_bot.Inst_MULADD._0353_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0395_ Tile_X0Y1_DSP_bot.Inst_MULADD._0396_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0409_ sky130_fd_sc_hd__a22oi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1169_ Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ Tile_X0Y1_DSP_bot.Inst_MULADD._0339_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0340_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y0_DSP_top.E6END_inbuf_3._0_ net28 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_118_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[80\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2 sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7 net258 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[199\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[380\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13 net233 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[365\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24 net245 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[376\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_130_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[97\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[108\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_142_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30 net252 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[30\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_130_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_inst0
+ net282 net182 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.ConfigBits\[51\] Tile_X0Y1_DSP_bot.ConfigBits\[52\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._26_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID2
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb2 sky130_fd_sc_hd__clkbuf_1
XANTENNA_214 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_225 Tile_X0Y0_DSP_top.S4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_203 Tile_X0Y1_DSP_bot.SS4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.strobe_inbuf_16._0_ net268 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[16\]
+ sky130_fd_sc_hd__clkbuf_1
X_362_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net736
+ sky130_fd_sc_hd__buf_1
XFILLER_0_67_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_293_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb1 VGND VGND VPWR VPWR net676
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.E6BEG_outbuf_1._0_ Tile_X0Y0_DSP_top.E6BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1023_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.A3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0196_ sky130_fd_sc_hd__or2_1
XFILLER_0_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput402 net402 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_124_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput435 net435 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[14] sky130_fd_sc_hd__buf_2
Xoutput413 net413 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput424 net424 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput468 net468 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput446 net446 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[24] sky130_fd_sc_hd__buf_2
Xoutput457 net457 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._88_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q12
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 sky130_fd_sc_hd__buf_12
XFILLER_0_10_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17 net237 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[273\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput479 net479 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28 net249 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[284\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.E6END_inbuf_3._0_ net208 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_72_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[330\] Tile_X0Y0_DSP_top.ConfigBits\[331\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_60_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._09_ net14 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEGb\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1710_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0004_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8 net259 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[40\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_345_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb1 VGND VGND VPWR VPWR net728
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1641_ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.ConfigBits\[4\] Tile_X0Y1_DSP_bot.Inst_MULADD._0801_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0802_ sky130_fd_sc_hd__a221o_1
XFILLER_0_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1572_ Tile_X0Y1_DSP_bot.Inst_MULADD._0733_ Tile_X0Y1_DSP_bot.Inst_MULADD._0734_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0712_ Tile_X0Y1_DSP_bot.Inst_MULADD._0714_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0737_ sky130_fd_sc_hd__o211ai_2
X_276_ Tile_X0Y1_DSP_bot.FrameData_O\[28\] VGND VGND VPWR VPWR net651 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._11_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot7
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B7 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12 net232 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[396\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23 net244 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[407\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1006_ Tile_X0Y1_DSP_bot.Inst_MULADD._0176_ Tile_X0Y1_DSP_bot.Inst_MULADD._0178_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0175_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0180_
+ sky130_fd_sc_hd__or3_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[128\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[139\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_115_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst1
+ net204 Tile_X0Y0_DSP_top.SS4BEG\[1\] net339 net357 Tile_X0Y1_DSP_bot.ConfigBits\[256\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[257\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.N4BEG_outbuf_9._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4END\[9\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[86\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[183\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_130_ Tile_X0Y0_DSP_top.N4BEG\[10\] VGND VGND VPWR VPWR net503 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[101\] Tile_X0Y1_DSP_bot.ConfigBits\[102\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_33_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_061_ Tile_X0Y0_DSP_top.FrameData_O\[13\] VGND VGND VPWR VPWR net434 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16 net236 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[304\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27 net248 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[315\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1624_ Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ Tile_X0Y1_DSP_bot.Inst_MULADD._0785_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0786_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q15
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_153_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 net4 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[19\] Tile_X0Y0_DSP_top.ConfigBits\[20\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
X_328_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 VGND VGND VPWR VPWR net702
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1555_ Tile_X0Y1_DSP_bot.Inst_MULADD._0714_ Tile_X0Y1_DSP_bot.Inst_MULADD._0715_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0719_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0721_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_259_ Tile_X0Y1_DSP_bot.FrameData_O\[11\] VGND VGND VPWR VPWR net633 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1486_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0653_ sky130_fd_sc_hd__and4_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[296\] Tile_X0Y0_DSP_top.ConfigBits\[297\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG4 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID2
+ net15 net95 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG5 Tile_X0Y0_DSP_top.ConfigBits\[168\]
+ Tile_X0Y0_DSP_top.ConfigBits\[169\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst0
+ net282 net288 net310 net188 Tile_X0Y1_DSP_bot.ConfigBits\[296\] Tile_X0Y1_DSP_bot.ConfigBits\[297\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_117_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.W6BEG_outbuf_9._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_144_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top.N4END_inbuf_7._0_ Tile_X0Y0_DSP_top.N4END\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG_i\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_113_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 VGND VGND VPWR VPWR net495
+ sky130_fd_sc_hd__buf_1
XFILLER_0_108_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_044_ Tile_X0Y0_DSP_top.EE4BEG\[12\] VGND VGND VPWR VPWR net417 sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1340_ Tile_X0Y1_DSP_bot.Inst_MULADD._0341_ Tile_X0Y1_DSP_bot.Inst_MULADD._0508_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0509_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0510_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_150_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[181\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[170\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_131_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1271_ Tile_X0Y1_DSP_bot.Inst_MULADD._0265_ Tile_X0Y1_DSP_bot.Inst_MULADD._0267_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0441_
+ sky130_fd_sc_hd__o21ai_2
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END2
+ net7 net21 Tile_X0Y0_DSP_top.ConfigBits\[346\] Tile_X0Y0_DSP_top.ConfigBits\[347\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0986_ Tile_X0Y1_DSP_bot.Inst_MULADD._0145_ Tile_X0Y1_DSP_bot.Inst_MULADD._0138_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0149_ Tile_X0Y1_DSP_bot.Inst_MULADD._0114_ Tile_X0Y1_DSP_bot.Inst_MULADD._0147_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0160_ sky130_fd_sc_hd__a221oi_4
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1607_ Tile_X0Y1_DSP_bot.Inst_MULADD._0741_ Tile_X0Y1_DSP_bot.Inst_MULADD._0767_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0770_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0771_
+ sky130_fd_sc_hd__a21boi_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID5
+ net18 net98 net150 Tile_X0Y0_DSP_top.ConfigBits\[210\] Tile_X0Y0_DSP_top.ConfigBits\[211\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.NN4END_inbuf_2._0_ net329 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1538_ Tile_X0Y1_DSP_bot.Inst_MULADD._0154_ Tile_X0Y1_DSP_bot.Inst_MULADD._0646_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_ Tile_X0Y1_DSP_bot.Inst_MULADD._0655_ Tile_X0Y1_DSP_bot.Inst_MULADD._0651_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0704_ sky130_fd_sc_hd__o311a_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1469_ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0637_ sky130_fd_sc_hd__and2_1
XTile_X0Y0_DSP_top.N4BEG_outbuf_5._0_ Tile_X0Y0_DSP_top.N4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[5\] sky130_fd_sc_hd__buf_2
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5 net256 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[101\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_149_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[282\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.NN4BEG_outbuf_9._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_117_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput302 Tile_X0Y1_N4END[10] VGND VGND VPWR VPWR net302 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15 net235 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[335\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26 net247 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[346\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput335 Tile_X0Y1_W1END[1] VGND VGND VPWR VPWR net335 sky130_fd_sc_hd__buf_4
Xinput324 Tile_X0Y1_NN4END[1] VGND VGND VPWR VPWR net324 sky130_fd_sc_hd__buf_1
Xinput313 Tile_X0Y1_N4END[6] VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__clkbuf_1
Xinput346 Tile_X0Y1_W2MID[0] VGND VGND VPWR VPWR net346 sky130_fd_sc_hd__clkbuf_4
Xinput368 Tile_X0Y1_WW4END[11] VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__clkbuf_1
Xinput379 Tile_X0Y1_WW4END[7] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__clkbuf_1
Xinput357 Tile_X0Y1_W6END[1] VGND VGND VPWR VPWR net357 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[318\] Tile_X0Y1_DSP_bot.ConfigBits\[319\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG7 sky130_fd_sc_hd__mux4_1
XFILLER_0_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.data_outbuf_29._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[29\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[29\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.N4END_inbuf_7._0_ net303 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_6 Tile_X0Y0_DSP_top.FrameStrobe\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_027_ Tile_X0Y0_DSP_top.E6BEG\[7\] VGND VGND VPWR VPWR net411 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_2._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END2 sky130_fd_sc_hd__buf_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1323_ Tile_X0Y1_DSP_bot.Inst_MULADD._0483_ Tile_X0Y1_DSP_bot.Inst_MULADD._0490_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0491_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0493_
+ sky130_fd_sc_hd__nand3_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1254_ Tile_X0Y1_DSP_bot.Inst_MULADD._0421_ Tile_X0Y1_DSP_bot.Inst_MULADD._0424_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0425_ sky130_fd_sc_hd__xnor2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_W1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG2 Tile_X0Y0_DSP_top.ConfigBits\[86\]
+ Tile_X0Y0_DSP_top.ConfigBits\[87\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1
+ sky130_fd_sc_hd__mux4_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1185_ Tile_X0Y1_DSP_bot.Inst_MULADD._0026_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0356_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_119_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0969_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0143_ sky130_fd_sc_hd__and2_2
XFILLER_0_17_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_5._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.S4BEG_outbuf_9._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[9\] sky130_fd_sc_hd__buf_2
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.W6BEG_outbuf_5._0_ Tile_X0Y0_DSP_top.W6BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[5\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._42_ net95 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb2
+ sky130_fd_sc_hd__clkbuf_2
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[212\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19 net239 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[243\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[368\] Tile_X0Y0_DSP_top.ConfigBits\[369\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 sky130_fd_sc_hd__mux4_2
XFILLER_0_118_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst0
+ net3 net135 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.ConfigBits\[108\] Tile_X0Y0_DSP_top.ConfigBits\[109\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst0
+ net282 net290 net182 net190 Tile_X0Y1_DSP_bot.ConfigBits\[368\] Tile_X0Y1_DSP_bot.ConfigBits\[369\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput110 Tile_X0Y0_S4END[3] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_2
Xinput121 Tile_X0Y0_SS4END[13] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
Xinput132 Tile_X0Y0_SS4END[9] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
Xinput154 Tile_X0Y0_W6END[10] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
Xinput143 Tile_X0Y0_W2END[6] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput176 Tile_X0Y0_WW4END[5] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xinput165 Tile_X0Y0_WW4END[0] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_2
Xinput187 Tile_X0Y1_E2END[2] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__buf_2
Xinput198 Tile_X0Y1_E2MID[5] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__buf_2
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG0 net299
+ net199 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG6
+ Tile_X0Y1_DSP_bot.ConfigBits\[184\] Tile_X0Y1_DSP_bot.ConfigBits\[185\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END1 net4 net6 net24 Tile_X0Y0_DSP_top.ConfigBits\[310\]
+ Tile_X0Y0_DSP_top.ConfigBits\[311\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput617 net617 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput606 net606 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput628 net628 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput639 net639 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1306_ Tile_X0Y1_DSP_bot.Inst_MULADD._0474_ Tile_X0Y1_DSP_bot.Inst_MULADD._0475_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0476_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1237_ Tile_X0Y1_DSP_bot.Inst_MULADD._0345_ Tile_X0Y1_DSP_bot.Inst_MULADD._0397_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0408_ sky130_fd_sc_hd__or2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1168_ Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0340_ sky130_fd_sc_hd__nand2_1
XFILLER_0_118_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[80\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1099_ Tile_X0Y1_DSP_bot.Inst_MULADD._0269_ Tile_X0Y1_DSP_bot.Inst_MULADD._0270_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0070_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0271_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_159_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8 net259 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[200\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[381\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14 net234 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[366\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25 net246 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[377\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[98\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[109\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_130_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20 net241 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[20\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31 net253 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[31\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG0
+ Tile_X0Y1_DSP_bot.ConfigBits\[51\] Tile_X0Y1_DSP_bot.ConfigBits\[52\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.data_inbuf_4._0_ net255 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._25_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID1
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb1 sky130_fd_sc_hd__clkbuf_2
XANTENNA_204 Tile_X0Y1_DSP_bot.SS4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_215 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_226 Tile_X0Y1_DSP_bot.EE4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_361_ Tile_X0Y1_DSP_bot.W6BEG\[9\] VGND VGND VPWR VPWR net746 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG0 net310
+ net188 net341 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[400\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[401\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.data_outbuf_25._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[25\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[25\] sky130_fd_sc_hd__clkbuf_1
X_292_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb0 VGND VGND VPWR VPWR net675
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1022_ Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ Tile_X0Y1_DSP_bot.Inst_MULADD._0044_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0141_ Tile_X0Y1_DSP_bot.Inst_MULADD._0188_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0195_ sky130_fd_sc_hd__nand4_4
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.data_outbuf_16._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[16\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput403 net403 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[10] sky130_fd_sc_hd__buf_2
Xoutput425 net425 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput414 net414 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[0] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.S4BEG_outbuf_5._0_ Tile_X0Y0_DSP_top.S4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[5\] sky130_fd_sc_hd__clkbuf_1
Xoutput469 net469 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput447 net447 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[25] sky130_fd_sc_hd__clkbuf_4
Xoutput436 net436 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput458 net458 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[6] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._87_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q11
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 sky130_fd_sc_hd__buf_12
XFILLER_0_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18 net238 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[274\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29 net250 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[285\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[332\] Tile_X0Y0_DSP_top.ConfigBits\[333\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 sky130_fd_sc_hd__mux4_2
XFILLER_0_103_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END7
+ net41 net92 net144 Tile_X0Y0_DSP_top.ConfigBits\[230\] Tile_X0Y0_DSP_top.ConfigBits\[231\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_13_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst0
+ net289 net183 net189 net201 Tile_X0Y1_DSP_bot.ConfigBits\[332\] Tile_X0Y1_DSP_bot.ConfigBits\[333\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._08_ net13 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEGb\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9 net260 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[41\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_153_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_344_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb0 VGND VGND VPWR VPWR net727
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1640_ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ Tile_X0Y1_DSP_bot.Inst_MULADD._0800_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0801_ sky130_fd_sc_hd__and2b_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1571_ Tile_X0Y1_DSP_bot.Inst_MULADD._0711_ Tile_X0Y1_DSP_bot.Inst_MULADD._0725_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0735_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0736_
+ sky130_fd_sc_hd__o21ai_1
X_275_ Tile_X0Y1_DSP_bot.FrameData_O\[27\] VGND VGND VPWR VPWR net650 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._10_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot6
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B6 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13 net233 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[397\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24 net245 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[408\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1005_ Tile_X0Y1_DSP_bot.Inst_MULADD._0175_ Tile_X0Y1_DSP_bot.Inst_MULADD._0176_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0178_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0179_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[129\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[140\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30 net252 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[62\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_115_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst2
+ net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[256\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[257\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[86\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_156_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[184\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_060_ Tile_X0Y0_DSP_top.FrameData_O\[12\] VGND VGND VPWR VPWR net433 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.W6END_inbuf_1._0_ net158 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28 net249 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[316\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17 net237 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[305\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_327_ Tile_X0Y1_DSP_bot.SS4BEG\[11\] VGND VGND VPWR VPWR net701 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1623_ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0786_ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG1
+ Tile_X0Y0_DSP_top.ConfigBits\[19\] Tile_X0Y0_DSP_top.ConfigBits\[20\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0 net229 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[320\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_101_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1554_ Tile_X0Y1_DSP_bot.Inst_MULADD._0714_ Tile_X0Y1_DSP_bot.Inst_MULADD._0715_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0719_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0720_
+ sky130_fd_sc_hd__nand3_1
X_258_ Tile_X0Y1_DSP_bot.FrameData_O\[10\] VGND VGND VPWR VPWR net632 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_189_ Tile_X0Y0_DSP_top.WW4BEG\[5\] VGND VGND VPWR VPWR net578 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1485_ Tile_X0Y1_DSP_bot.Inst_MULADD._0192_ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0599_ Tile_X0Y1_DSP_bot.Inst_MULADD._0651_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0652_ sky130_fd_sc_hd__o211ai_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID4
+ net97 net149 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 Tile_X0Y0_DSP_top.ConfigBits\[170\]
+ Tile_X0Y0_DSP_top.ConfigBits\[171\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG2
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst1
+ net204 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb3 net341 net357 Tile_X0Y1_DSP_bot.ConfigBits\[296\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[297\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 net82 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[101\] Tile_X0Y0_DSP_top.ConfigBits\[102\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_5._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_112_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 VGND VGND VPWR VPWR net494
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_043_ Tile_X0Y0_DSP_top.EE4BEG\[11\] VGND VGND VPWR VPWR net416 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[160\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[171\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_131_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1270_ Tile_X0Y1_DSP_bot.Inst_MULADD._0070_ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0359_ Tile_X0Y1_DSP_bot.Inst_MULADD._0050_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0440_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.W6END_inbuf_1._0_ net359 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0985_ Tile_X0Y1_DSP_bot.Inst_MULADD._0148_ Tile_X0Y1_DSP_bot.Inst_MULADD._0150_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0153_ Tile_X0Y1_DSP_bot.Inst_MULADD._0157_ Tile_X0Y1_DSP_bot.Inst_MULADD._0158_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0159_ sky130_fd_sc_hd__o2111ai_4
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst1
+ net87 net109 net139 net153 Tile_X0Y0_DSP_top.ConfigBits\[346\] Tile_X0Y0_DSP_top.ConfigBits\[347\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1606_ Tile_X0Y1_DSP_bot.Inst_MULADD._0768_ Tile_X0Y1_DSP_bot.Inst_MULADD._0639_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0769_ Tile_X0Y1_DSP_bot.Inst_MULADD._0744_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0770_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_21_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID1
+ net14 net94 net146 Tile_X0Y0_DSP_top.ConfigBits\[212\] Tile_X0Y0_DSP_top.ConfigBits\[213\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1537_ Tile_X0Y1_DSP_bot.Inst_MULADD._0700_ Tile_X0Y1_DSP_bot.Inst_MULADD._0701_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0664_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0703_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1468_ Tile_X0Y1_DSP_bot.Inst_MULADD._0630_ Tile_X0Y1_DSP_bot.Inst_MULADD._0632_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0635_ Tile_X0Y1_DSP_bot.Inst_MULADD._0579_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0636_ sky130_fd_sc_hd__a22o_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1399_ Tile_X0Y1_DSP_bot.Inst_MULADD._0567_ Tile_X0Y1_DSP_bot.Inst_MULADD._0467_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0481_ Tile_X0Y1_DSP_bot.Inst_MULADD._0464_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0568_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_20_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6 net257 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[102\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_153_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[283\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput303 Tile_X0Y1_N4END[11] VGND VGND VPWR VPWR net303 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16 net236 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[336\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput336 Tile_X0Y1_W1END[2] VGND VGND VPWR VPWR net336 sky130_fd_sc_hd__buf_4
Xinput325 Tile_X0Y1_NN4END[2] VGND VGND VPWR VPWR net325 sky130_fd_sc_hd__clkbuf_2
Xinput314 Tile_X0Y1_N4END[7] VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.WW4END_inbuf_3._0_ net379 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27 net248 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[347\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput347 Tile_X0Y1_W2MID[1] VGND VGND VPWR VPWR net347 sky130_fd_sc_hd__clkbuf_4
Xinput358 Tile_X0Y1_W6END[2] VGND VGND VPWR VPWR net358 sky130_fd_sc_hd__clkbuf_1
Xinput369 Tile_X0Y1_WW4END[12] VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_123_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_7 Tile_X0Y0_DSP_top.FrameStrobe\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_026_ Tile_X0Y0_DSP_top.E6BEG\[6\] VGND VGND VPWR VPWR net410 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1322_ Tile_X0Y1_DSP_bot.Inst_MULADD._0483_ Tile_X0Y1_DSP_bot.Inst_MULADD._0490_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0491_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0492_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_158_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END0
+ net3 net9 Tile_X0Y0_DSP_top.ConfigBits\[258\] Tile_X0Y0_DSP_top.ConfigBits\[259\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_104_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1253_ Tile_X0Y1_DSP_bot.Inst_MULADD._0422_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0423_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0424_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_W1BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG3 Tile_X0Y0_DSP_top.ConfigBits\[88\]
+ Tile_X0Y0_DSP_top.ConfigBits\[89\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1184_ Tile_X0Y1_DSP_bot.A7 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0355_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_107_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0968_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.B2
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0142_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0899_ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_114_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.N4END_inbuf_11._0_ Tile_X0Y0_DSP_top.N4END\[15\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._41_ net94 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb1
+ sky130_fd_sc_hd__buf_2
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 net4 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[75\] Tile_X0Y0_DSP_top.ConfigBits\[76\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[202\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[213\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.inst_clk_buf Tile_X0Y0_DSP_top.UserCLK VGND VGND VPWR VPWR net534
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb5 net335 Tile_X0Y1_DSP_bot.ConfigBits\[368\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[369\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[108\] Tile_X0Y0_DSP_top.ConfigBits\[109\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_120_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput111 Tile_X0Y0_S4END[4] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
Xinput100 Tile_X0Y0_S2MID[7] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_4
Xinput122 Tile_X0Y0_SS4END[14] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
Xinput144 Tile_X0Y0_W2END[7] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_2
Xinput133 Tile_X0Y0_W1END[0] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__buf_4
Xinput155 Tile_X0Y0_W6END[11] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
Xinput177 Tile_X0Y0_WW4END[6] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xinput166 Tile_X0Y0_WW4END[10] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
Xinput199 Tile_X0Y1_E2MID[6] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__clkbuf_4
Xinput188 Tile_X0Y1_E2END[3] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG1 net295
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG2 net348 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG6
+ Tile_X0Y1_DSP_bot.ConfigBits\[186\] Tile_X0Y1_DSP_bot.ConfigBits\[187\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_85_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst1
+ net86 net108 net138 net156 Tile_X0Y0_DSP_top.ConfigBits\[310\] Tile_X0Y0_DSP_top.ConfigBits\[311\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_151_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput618 net618 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput607 net607 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[2] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG0 net8
+ net126 net173 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2 Tile_X0Y0_DSP_top.ConfigBits\[382\]
+ Tile_X0Y0_DSP_top.ConfigBits\[383\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG0
+ sky130_fd_sc_hd__mux4_1
X_009_ Tile_X0Y0_DSP_top.E2BEG\[5\] VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput629 net629 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[8] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1305_ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_ Tile_X0Y1_DSP_bot.Inst_MULADD._0472_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0347_ Tile_X0Y1_DSP_bot.Inst_MULADD._0473_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0475_ sky130_fd_sc_hd__nand4_1
XFILLER_0_94_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1236_ Tile_X0Y1_DSP_bot.Inst_MULADD._0404_ Tile_X0Y1_DSP_bot.Inst_MULADD._0405_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0406_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0407_
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1167_ Tile_X0Y1_DSP_bot.Inst_MULADD._0249_ Tile_X0Y1_DSP_bot.Inst_MULADD._0338_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0339_ sky130_fd_sc_hd__xor2_2
XFILLER_0_118_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.data_inbuf_30._0_ net72 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[30\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1098_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.A4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0270_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_134_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9 net260 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[201\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[382\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15 net235 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[367\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26 net247 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[378\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.SS4END_inbuf_11._0_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[99\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[110\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10 net230 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[10\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21 net242 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[21\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst0
+ net284 net292 net184 net192 Tile_X0Y1_DSP_bot.ConfigBits\[280\] Tile_X0Y1_DSP_bot.ConfigBits\[281\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.data_inbuf_21._0_ net62 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[21\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._24_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb0 sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[86\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_216 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_205 Tile_X0Y1_DSP_bot.SS4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_227 Tile_X0Y1_DSP_bot.EE4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_360_ Tile_X0Y1_DSP_bot.W6BEG\[8\] VGND VGND VPWR VPWR net745 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG1 net325
+ net187 Tile_X0Y0_DSP_top.S4BEG\[2\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[402\] Tile_X0Y1_DSP_bot.ConfigBits\[403\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_291_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG7 VGND VGND VPWR VPWR net674
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.strobe_inbuf_6._0_ Tile_X0Y0_DSP_top.FrameStrobe\[6\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1021_ Tile_X0Y1_DSP_bot.Inst_MULADD._0142_ Tile_X0Y1_DSP_bot.Inst_MULADD._0143_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ Tile_X0Y1_DSP_bot.Inst_MULADD._0138_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0194_ sky130_fd_sc_hd__o211ai_4
XTile_X0Y0_DSP_top.data_inbuf_12._0_ net52 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[12\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput404 net404 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput415 net415 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[10] sky130_fd_sc_hd__buf_2
Xoutput426 net426 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_0_22_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput448 net448 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[26] sky130_fd_sc_hd__clkbuf_4
Xoutput437 net437 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[16] sky130_fd_sc_hd__clkbuf_4
Xoutput459 net459 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[244\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_22_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._86_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q10
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 sky130_fd_sc_hd__buf_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19 net239 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[275\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1219_ Tile_X0Y1_DSP_bot.Inst_MULADD._0367_ Tile_X0Y1_DSP_bot.Inst_MULADD._0368_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0369_ Tile_X0Y1_DSP_bot.Inst_MULADD._0370_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0390_ sky130_fd_sc_hd__o211a_2
XFILLER_0_89_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.data_inbuf_30._0_ net252 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[30\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_159_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_147_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb4 Tile_X0Y0_DSP_top.S4BEG\[0\]
+ net342 net374 Tile_X0Y1_DSP_bot.ConfigBits\[332\] Tile_X0Y1_DSP_bot.ConfigBits\[333\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END3
+ net8 net88 net172 Tile_X0Y0_DSP_top.ConfigBits\[232\] Tile_X0Y0_DSP_top.ConfigBits\[233\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_95_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._07_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG7
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_157_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.SS4END_inbuf_5._0_ Tile_X0Y0_DSP_top.SS4BEG\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] sky130_fd_sc_hd__buf_2
XFILLER_0_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.data_inbuf_21._0_ net242 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[21\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_343_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG7 VGND VGND VPWR VPWR net726
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1570_ Tile_X0Y1_DSP_bot.Inst_MULADD._0733_ Tile_X0Y1_DSP_bot.Inst_MULADD._0734_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0735_ sky130_fd_sc_hd__nor2_1
X_274_ Tile_X0Y1_DSP_bot.FrameData_O\[26\] VGND VGND VPWR VPWR net649 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14 net234 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[398\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25 net246 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[409\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1004_ Tile_X0Y1_DSP_bot.Inst_MULADD._0127_ Tile_X0Y1_DSP_bot.Inst_MULADD._0177_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0125_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0178_
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[130\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_78_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[141\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31 net253 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[63\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20 net241 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[52\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.data_inbuf_12._0_ net232 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[12\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.ConfigBits\[256\] Tile_X0Y1_DSP_bot.ConfigBits\[257\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1699_ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ Tile_X0Y1_DSP_bot.Inst_MULADD._0785_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0015_ sky130_fd_sc_hd__nor2_1
XTile_X0Y0_DSP_top.S4END_inbuf_11._0_ net107 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[11\]
+ sky130_fd_sc_hd__buf_1
XFILLER_0_100_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._69_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG7
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[185\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_N1BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[6\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[7\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_92_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.EE4END_inbuf_4._0_ net227 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29 net250 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[317\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18 net238 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[306\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_83_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.strobe_inbuf_13._0_ Tile_X0Y0_DSP_top.FrameStrobe\[13\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[13\] sky130_fd_sc_hd__clkbuf_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_326_ Tile_X0Y1_DSP_bot.SS4BEG\[10\] VGND VGND VPWR VPWR net700 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1622_ Tile_X0Y1_DSP_bot.Inst_MULADD._0781_ Tile_X0Y1_DSP_bot.Inst_MULADD._0784_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0785_ sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1 net240 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[321\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_153_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1553_ Tile_X0Y1_DSP_bot.Inst_MULADD._0717_ Tile_X0Y1_DSP_bot.Inst_MULADD._0718_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0719_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_257_ Tile_X0Y1_DSP_bot.FrameData_O\[9\] VGND VGND VPWR VPWR net662 sky130_fd_sc_hd__clkbuf_1
X_188_ Tile_X0Y0_DSP_top.WW4BEG\[4\] VGND VGND VPWR VPWR net577 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1484_ Tile_X0Y1_DSP_bot.Inst_MULADD._0646_ Tile_X0Y1_DSP_bot.Inst_MULADD._0649_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0650_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0651_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG3 net13
+ net93 net145 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 Tile_X0Y0_DSP_top.ConfigBits\[172\]
+ Tile_X0Y0_DSP_top.ConfigBits\[173\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[296\] Tile_X0Y1_DSP_bot.ConfigBits\[297\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG2
+ Tile_X0Y0_DSP_top.ConfigBits\[101\] Tile_X0Y0_DSP_top.ConfigBits\[102\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.SS4END_inbuf_1._0_ net128 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[1\]
+ sky130_fd_sc_hd__buf_4
X_111_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG7 VGND VGND VPWR VPWR net493
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_042_ Tile_X0Y0_DSP_top.EE4BEG\[10\] VGND VGND VPWR VPWR net415 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[161\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[172\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30 net252 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[94\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.strobe_outbuf_15._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[15\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[15\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0984_ Tile_X0Y1_DSP_bot.Inst_MULADD._0145_ Tile_X0Y1_DSP_bot.Inst_MULADD._0138_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0149_ Tile_X0Y1_DSP_bot.Inst_MULADD._0114_ Tile_X0Y1_DSP_bot.Inst_MULADD._0147_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0158_ sky130_fd_sc_hd__a221o_2
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[346\] Tile_X0Y0_DSP_top.ConfigBits\[347\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.E6BEG_outbuf_8._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1605_ Tile_X0Y1_DSP_bot.Inst_MULADD._0722_ Tile_X0Y1_DSP_bot.Inst_MULADD._0683_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0769_ sky130_fd_sc_hd__nor2_1
X_309_ Tile_X0Y1_DSP_bot.S4BEG\[9\] VGND VGND VPWR VPWR net698 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1536_ Tile_X0Y1_DSP_bot.Inst_MULADD._0700_ Tile_X0Y1_DSP_bot.Inst_MULADD._0701_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0664_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0702_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_141_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_122_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1467_ Tile_X0Y1_DSP_bot.Inst_MULADD._0516_ Tile_X0Y1_DSP_bot.Inst_MULADD._0581_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0635_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1398_ Tile_X0Y1_DSP_bot.Inst_MULADD._0479_ Tile_X0Y1_DSP_bot.Inst_MULADD._0480_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0567_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7 net258 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[103\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_149_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[284\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.EE4END_inbuf_11._0_ net219 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17 net237 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[337\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28 net249 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[348\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput326 Tile_X0Y1_NN4END[3] VGND VGND VPWR VPWR net326 sky130_fd_sc_hd__clkbuf_2
Xinput315 Tile_X0Y1_N4END[8] VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_1
Xinput304 Tile_X0Y1_N4END[12] VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__clkbuf_1
Xinput348 Tile_X0Y1_W2MID[2] VGND VGND VPWR VPWR net348 sky130_fd_sc_hd__buf_2
Xinput337 Tile_X0Y1_W1END[3] VGND VGND VPWR VPWR net337 sky130_fd_sc_hd__clkbuf_8
Xinput359 Tile_X0Y1_W6END[3] VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.EE4END_inbuf_0._0_ net43 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 Tile_X0Y0_DSP_top.FrameStrobe\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_151_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_025_ Tile_X0Y0_DSP_top.E6BEG\[5\] VGND VGND VPWR VPWR net409 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1321_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0349_ Tile_X0Y1_DSP_bot.Inst_MULADD._0345_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0491_ sky130_fd_sc_hd__a31o_4
XFILLER_0_21_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst1
+ net21 net89 net141 net153 Tile_X0Y0_DSP_top.ConfigBits\[258\] Tile_X0Y0_DSP_top.ConfigBits\[259\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1252_ Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0423_ sky130_fd_sc_hd__clkbuf_4
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1183_ Tile_X0Y1_DSP_bot.Inst_MULADD._0353_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0354_ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.strobe_outbuf_4._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[4\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[4\] sky130_fd_sc_hd__buf_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_W1BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG0 Tile_X0Y0_DSP_top.ConfigBits\[90\]
+ Tile_X0Y0_DSP_top.ConfigBits\[91\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.NN4BEG_outbuf_10._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG\[10\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0967_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.Inst_MULADD._0139_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0140_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0141_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_8_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0898_ Tile_X0Y1_DSP_bot.Inst_MULADD._0073_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_84_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.WW4BEG_outbuf_9._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[9\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1519_ Tile_X0Y1_DSP_bot.Inst_MULADD._0638_ Tile_X0Y1_DSP_bot.Inst_MULADD._0639_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0683_ Tile_X0Y1_DSP_bot.Inst_MULADD._0684_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0686_ sky130_fd_sc_hd__o22a_1
XTile_X0Y0_DSP_top.E6END_inbuf_6._0_ net31 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._40_ net93 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb0
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_57_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG3
+ Tile_X0Y0_DSP_top.ConfigBits\[75\] Tile_X0Y0_DSP_top.ConfigBits\[76\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[192\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_79_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[203\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_152_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[368\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[369\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[108\] Tile_X0Y0_DSP_top.ConfigBits\[109\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput101 Tile_X0Y0_S4END[0] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__buf_2
Xinput112 Tile_X0Y0_S4END[5] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
Xinput123 Tile_X0Y0_SS4END[15] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput145 Tile_X0Y0_W2MID[0] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__buf_2
Xinput134 Tile_X0Y0_W1END[1] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_4
Xinput156 Tile_X0Y0_W6END[1] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_4
Xinput167 Tile_X0Y0_WW4END[11] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
Xinput178 Tile_X0Y0_WW4END[7] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_2._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.strobe_inbuf_19._0_ net271 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[19\]
+ sky130_fd_sc_hd__clkbuf_1
Xinput189 Tile_X0Y1_E2END[4] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END6
+ net3 net11 Tile_X0Y0_DSP_top.ConfigBits\[298\] Tile_X0Y0_DSP_top.ConfigBits\[299\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG2 net197
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG4 net350 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ Tile_X0Y1_DSP_bot.ConfigBits\[188\] Tile_X0Y1_DSP_bot.ConfigBits\[189\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_66_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.E6BEG_outbuf_4._0_ Tile_X0Y0_DSP_top.E6BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[310\] Tile_X0Y0_DSP_top.ConfigBits\[311\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput608 net608 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_008_ Tile_X0Y0_DSP_top.E2BEG\[4\] VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput619 net619 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[13] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1304_ Tile_X0Y1_DSP_bot.Inst_MULADD._0347_ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0472_ Tile_X0Y1_DSP_bot.Inst_MULADD._0473_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0474_ sky130_fd_sc_hd__a22o_1
XTile_X0Y0_DSP_top.strobe_outbuf_10._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[10\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[10\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END2
+ net7 net144 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG2 Tile_X0Y0_DSP_top.ConfigBits\[384\]
+ Tile_X0Y0_DSP_top.ConfigBits\[385\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG1
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1235_ Tile_X0Y1_DSP_bot.Inst_MULADD._0345_ Tile_X0Y1_DSP_bot.Inst_MULADD._0397_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0353_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0406_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1166_ Tile_X0Y1_DSP_bot.Inst_MULADD._0335_ Tile_X0Y1_DSP_bot.Inst_MULADD._0337_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0338_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1097_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0269_ sky130_fd_sc_hd__and2_2
XFILLER_0_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.data_inbuf_1._0_ net60 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[383\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16 net236 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[368\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27 net248 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[379\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[100\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[111\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22 net243 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[22\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11 net231 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[11\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._23_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG7 sky130_fd_sc_hd__clkbuf_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb7
+ net335 net337 Tile_X0Y1_DSP_bot.ConfigBits\[280\] Tile_X0Y1_DSP_bot.ConfigBits\[281\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_99_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[87\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.E6END_inbuf_6._0_ net211 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XANTENNA_206 Tile_X0Y1_DSP_bot.SS4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_217 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_228 Tile_X0Y1_DSP_bot.S4BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG2 net308
+ Tile_X0Y0_DSP_top.SS4BEG\[1\] net342 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[404\] Tile_X0Y1_DSP_bot.ConfigBits\[405\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG2 sky130_fd_sc_hd__mux4_2
X_290_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG6 VGND VGND VPWR VPWR net673
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1020_ Tile_X0Y1_DSP_bot.Inst_MULADD._0044_ Tile_X0Y1_DSP_bot.Inst_MULADD._0141_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0192_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0193_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_98_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput405 net405 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput416 net416 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput449 net449 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput438 net438 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput427 net427 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[245\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._85_ net353 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb7
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[234\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1218_ Tile_X0Y1_DSP_bot.Inst_MULADD._0365_ Tile_X0Y1_DSP_bot.Inst_MULADD._0377_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0389_ sky130_fd_sc_hd__nand2_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1149_ Tile_X0Y1_DSP_bot.Inst_MULADD._0199_ Tile_X0Y1_DSP_bot.Inst_MULADD._0235_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0306_ Tile_X0Y1_DSP_bot.Inst_MULADD._0291_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0321_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.SS4BEG_outbuf_2._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_60_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[332\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[333\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END5
+ net10 net124 net142 Tile_X0Y0_DSP_top.ConfigBits\[234\] Tile_X0Y0_DSP_top.ConfigBits\[235\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG2 sky130_fd_sc_hd__mux4_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._06_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_342_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG6 VGND VGND VPWR VPWR net725
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_273_ Tile_X0Y1_DSP_bot.FrameData_O\[25\] VGND VGND VPWR VPWR net648 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.data_outbuf_10._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15 net235 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[399\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1003_ Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ Tile_X0Y1_DSP_bot.Inst_MULADD._0097_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0123_ Tile_X0Y1_DSP_bot.Inst_MULADD._0124_ Tile_X0Y1_DSP_bot.Inst_MULADD._0098_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0177_ sky130_fd_sc_hd__o221a_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26 net247 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[410\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[131\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[142\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10 net230 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[42\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21 net242 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[53\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_138_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[258\] Tile_X0Y1_DSP_bot.ConfigBits\[259\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1698_ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ Tile_X0Y1_DSP_bot.Inst_MULADD._0783_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0773_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0014_
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_112_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END0
+ net1 net5 Tile_X0Y0_DSP_top.ConfigBits\[370\] Tile_X0Y0_DSP_top.ConfigBits\[371\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._68_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[186\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_N1BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[8\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[9\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_77_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0 net229 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[64\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[276\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19 net239 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[307\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_325_ Tile_X0Y1_DSP_bot.SS4BEG\[9\] VGND VGND VPWR VPWR net714 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1621_ Tile_X0Y1_DSP_bot.Inst_MULADD._0782_ Tile_X0Y1_DSP_bot.Inst_MULADD._0783_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0778_ Tile_X0Y1_DSP_bot.Inst_MULADD._0780_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0784_ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_138_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2 net251 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[322\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_153_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1552_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] Tile_X0Y1_DSP_bot.Inst_MULADD._0423_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0718_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_256_ Tile_X0Y1_DSP_bot.FrameData_O\[8\] VGND VGND VPWR VPWR net661 sky130_fd_sc_hd__clkbuf_1
X_187_ Tile_X0Y0_DSP_top.WW4BEG\[3\] VGND VGND VPWR VPWR net576 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1483_ Tile_X0Y1_DSP_bot.Inst_MULADD._0261_ Tile_X0Y1_DSP_bot.Inst_MULADD._0263_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0650_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_3_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[296\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[297\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.NN4END_inbuf_5._0_ net332 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_27_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.N4BEG_outbuf_8._0_ Tile_X0Y0_DSP_top.N4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[8\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_110_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG6 VGND VGND VPWR VPWR net492
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_041_ Tile_X0Y0_DSP_top.EE4BEG\[9\] VGND VGND VPWR VPWR net429 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[173\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[162\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31 net253 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[95\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20 net241 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[84\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0983_ Tile_X0Y1_DSP_bot.Inst_MULADD._0156_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0157_ sky130_fd_sc_hd__clkbuf_4
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[346\] Tile_X0Y0_DSP_top.ConfigBits\[347\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1604_ Tile_X0Y1_DSP_bot.Inst_MULADD._0632_ Tile_X0Y1_DSP_bot.Inst_MULADD._0689_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0768_ sky130_fd_sc_hd__nand2_1
X_308_ Tile_X0Y1_DSP_bot.S4BEG\[8\] VGND VGND VPWR VPWR net697 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1535_ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0698_ Tile_X0Y1_DSP_bot.Inst_MULADD._0699_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0701_ sky130_fd_sc_hd__nand4_4
X_239_ Tile_X0Y1_DSP_bot.EE4BEG\[7\] VGND VGND VPWR VPWR net628 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_5._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4END\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1466_ Tile_X0Y1_DSP_bot.Inst_MULADD._0516_ Tile_X0Y1_DSP_bot.Inst_MULADD._0581_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0633_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0634_
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1397_ Tile_X0Y1_DSP_bot.Inst_MULADD._0490_ Tile_X0Y1_DSP_bot.Inst_MULADD._0493_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0563_ Tile_X0Y1_DSP_bot.Inst_MULADD._0565_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0566_ sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END7
+ net4 net12 Tile_X0Y0_DSP_top.ConfigBits\[334\] Tile_X0Y0_DSP_top.ConfigBits\[335\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8 net259 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[104\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[285\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_8._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[8\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.W6BEG_outbuf_8._0_ Tile_X0Y0_DSP_top.W6BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput327 Tile_X0Y1_NN4END[4] VGND VGND VPWR VPWR net327 sky130_fd_sc_hd__clkbuf_1
Xinput305 Tile_X0Y1_N4END[13] VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
Xinput316 Tile_X0Y1_N4END[9] VGND VGND VPWR VPWR net316 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29 net250 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[349\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18 net238 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[338\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput338 Tile_X0Y1_W2END[0] VGND VGND VPWR VPWR net338 sky130_fd_sc_hd__buf_2
Xinput349 Tile_X0Y1_W2MID[3] VGND VGND VPWR VPWR net349 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_9 Tile_X0Y0_DSP_top.FrameStrobe\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_024_ Tile_X0Y0_DSP_top.E6BEG\[4\] VGND VGND VPWR VPWR net408 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1320_ Tile_X0Y1_DSP_bot.Inst_MULADD._0484_ Tile_X0Y1_DSP_bot.Inst_MULADD._0488_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0391_ Tile_X0Y1_DSP_bot.Inst_MULADD._0407_ Tile_X0Y1_DSP_bot.Inst_MULADD._0489_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0490_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[258\] Tile_X0Y0_DSP_top.ConfigBits\[259\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1251_ Tile_X0Y1_DSP_bot.C7 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[7\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0422_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1182_ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ Tile_X0Y1_DSP_bot.Inst_MULADD._0351_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0352_ Tile_X0Y1_DSP_bot.Inst_MULADD._0345_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0353_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_88_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID7
+ net20 net100 net152 Tile_X0Y0_DSP_top.ConfigBits\[182\] Tile_X0Y0_DSP_top.ConfigBits\[183\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0966_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0140_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0897_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.Inst_MULADD._0061_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0062_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0073_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.NN4END_inbuf_1._0_ Tile_X0Y0_DSP_top.NN4END\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1518_ Tile_X0Y1_DSP_bot.Inst_MULADD._0638_ Tile_X0Y1_DSP_bot.Inst_MULADD._0639_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0683_ Tile_X0Y1_DSP_bot.Inst_MULADD._0684_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0685_ sky130_fd_sc_hd__nor4_1
XFILLER_0_4_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1449_ Tile_X0Y1_DSP_bot.Inst_MULADD._0613_ Tile_X0Y1_DSP_bot.Inst_MULADD._0611_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0612_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0617_
+ sky130_fd_sc_hd__nand3b_2
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[193\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[204\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.EE4BEG_outbuf_2._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[2\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[368\] Tile_X0Y1_DSP_bot.ConfigBits\[369\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_160_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG2
+ Tile_X0Y0_DSP_top.ConfigBits\[108\] Tile_X0Y0_DSP_top.ConfigBits\[109\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput102 Tile_X0Y0_S4END[10] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.data_inbuf_7._0_ net258 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
Xinput113 Tile_X0Y0_S4END[6] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
Xinput124 Tile_X0Y0_SS4END[1] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__buf_2
Xinput135 Tile_X0Y0_W1END[2] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_4
Xinput157 Tile_X0Y0_W6END[2] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_1
Xinput168 Tile_X0Y0_WW4END[12] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
Xinput146 Tile_X0Y0_W2MID[1] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__buf_2
Xinput179 Tile_X0Y0_WW4END[8] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst1
+ net81 net83 net91 net135 Tile_X0Y0_DSP_top.ConfigBits\[298\] Tile_X0Y0_DSP_top.ConfigBits\[299\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.data_outbuf_28._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[28\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[28\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG3 net293
+ net193 net346 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 Tile_X0Y1_DSP_bot.ConfigBits\[190\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[191\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG3
+ sky130_fd_sc_hd__mux4_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[310\] Tile_X0Y0_DSP_top.ConfigBits\[311\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput609 net609 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[4] sky130_fd_sc_hd__clkbuf_4
X_007_ Tile_X0Y0_DSP_top.E2BEG\[3\] VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1303_ Tile_X0Y1_DSP_bot.Inst_MULADD._0063_ Tile_X0Y1_DSP_bot.Inst_MULADD._0299_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0380_ Tile_X0Y1_DSP_bot.Inst_MULADD._0382_ Tile_X0Y1_DSP_bot.Inst_MULADD._0372_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0473_ sky130_fd_sc_hd__o221ai_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END1
+ net40 net108 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 Tile_X0Y0_DSP_top.ConfigBits\[386\]
+ Tile_X0Y0_DSP_top.ConfigBits\[387\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1234_ Tile_X0Y1_DSP_bot.Inst_MULADD._0385_ Tile_X0Y1_DSP_bot.Inst_MULADD._0386_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0290_ Tile_X0Y1_DSP_bot.Inst_MULADD._0289_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0405_ sky130_fd_sc_hd__o22a_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1165_ Tile_X0Y1_DSP_bot.Inst_MULADD._0325_ Tile_X0Y1_DSP_bot.Inst_MULADD._0331_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0336_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0337_
+ sky130_fd_sc_hd__nand3_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1096_ Tile_X0Y1_DSP_bot.Inst_MULADD._0030_ Tile_X0Y1_DSP_bot.Inst_MULADD._0031_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0265_ Tile_X0Y1_DSP_bot.Inst_MULADD._0267_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0268_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.data_outbuf_19._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[19\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[19\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._0949_ Tile_X0Y1_DSP_bot.Inst_MULADD._0122_ Tile_X0Y1_DSP_bot.Inst_MULADD._0082_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0121_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0124_
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28 net249 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[380\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17 net237 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[369\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[101\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.S4BEG_outbuf_8._0_ Tile_X0Y0_DSP_top.S4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[112\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12 net232 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[12\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23 net244 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[23\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._22_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG6 sky130_fd_sc_hd__clkbuf_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[280\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[281\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XANTENNA_207 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[88\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_218 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_229 Tile_X0Y1_DSP_bot.S4BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG3 net222
+ Tile_X0Y0_DSP_top.S4BEG\[0\] net373 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[406\] Tile_X0Y1_DSP_bot.ConfigBits\[407\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_48_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0 net229 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[224\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput406 net406 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput417 net417 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput439 net439 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[18] sky130_fd_sc_hd__buf_2
Xoutput428 net428 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[8] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[224\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._84_ net352 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb6
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[235\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.S4END_inbuf_0._0_ net111 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1217_ Tile_X0Y1_DSP_bot.Inst_MULADD._0378_ Tile_X0Y1_DSP_bot.Inst_MULADD._0384_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0387_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0388_
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1148_ Tile_X0Y1_DSP_bot.Inst_MULADD._0310_ Tile_X0Y1_DSP_bot.Inst_MULADD._0311_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0317_ Tile_X0Y1_DSP_bot.Inst_MULADD._0303_ Tile_X0Y1_DSP_bot.Inst_MULADD._0307_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0320_ sky130_fd_sc_hd__a221oi_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1079_ Tile_X0Y1_DSP_bot.Inst_MULADD._0199_ Tile_X0Y1_DSP_bot.Inst_MULADD._0217_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0221_ Tile_X0Y1_DSP_bot.Inst_MULADD._0222_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0251_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_54_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[332\] Tile_X0Y1_DSP_bot.ConfigBits\[333\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END2
+ net6 net86 net138 Tile_X0Y0_DSP_top.ConfigBits\[236\] Tile_X0Y0_DSP_top.ConfigBits\[237\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG3 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.strobe_inbuf_0._0_ net261 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._05_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_341_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG5 VGND VGND VPWR VPWR net724
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_272_ Tile_X0Y1_DSP_bot.FrameData_O\[24\] VGND VGND VPWR VPWR net647 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.W6END_inbuf_4._0_ net161 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16 net236 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[400\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1002_ Tile_X0Y1_DSP_bot.Inst_MULADD._0168_ Tile_X0Y1_DSP_bot.Inst_MULADD._0171_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0173_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0176_
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27 net248 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[411\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[143\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[132\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11 net231 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[43\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22 net243 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[54\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_144_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1697_ Tile_X0Y1_DSP_bot.Inst_MULADD._0841_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._67_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb5 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst1
+ net81 net83 net85 net133 Tile_X0Y0_DSP_top.ConfigBits\[370\] Tile_X0Y0_DSP_top.ConfigBits\[371\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_57_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.S4END_inbuf_0._0_ Tile_X0Y0_DSP_top.S4BEG\[4\] VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.S4BEG_i\[0\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_8._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[187\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_N1BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[10\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[11\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1 net240 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[65\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_143_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_222 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[266\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[277\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG0 net292
+ net192 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb7 net366 Tile_X0Y1_DSP_bot.ConfigBits\[248\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[249\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_324_ Tile_X0Y1_DSP_bot.SS4BEG\[8\] VGND VGND VPWR VPWR net713 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1620_ Tile_X0Y1_DSP_bot.Inst_MULADD._0765_ Tile_X0Y1_DSP_bot.Inst_MULADD._0771_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0783_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1551_ Tile_X0Y1_DSP_bot.Inst_MULADD._0423_ Tile_X0Y1_DSP_bot.Inst_MULADD._0716_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0717_ sky130_fd_sc_hd__nor2_1
X_255_ Tile_X0Y1_DSP_bot.FrameData_O\[7\] VGND VGND VPWR VPWR net660 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3 net254 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[323\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_186_ Tile_X0Y0_DSP_top.WW4BEG\[2\] VGND VGND VPWR VPWR net575 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1482_ Tile_X0Y1_DSP_bot.Inst_MULADD._0101_ Tile_X0Y1_DSP_bot.Inst_MULADD._0132_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0647_ Tile_X0Y1_DSP_bot.Inst_MULADD._0648_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0649_ sky130_fd_sc_hd__o2bb2ai_1
XTile_X0Y1_DSP_bot.W6END_inbuf_4._0_ net362 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[298\] Tile_X0Y1_DSP_bot.ConfigBits\[299\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_99_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1749_ net333 Tile_X0Y1_DSP_bot.C7 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[22\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_040_ Tile_X0Y0_DSP_top.EE4BEG\[8\] VGND VGND VPWR VPWR net428 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[174\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_116_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[163\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10 net230 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[74\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21 net242 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[85\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.WW4END_inbuf_6._0_ net367 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[38\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG\[12\] sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0982_ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ Tile_X0Y1_DSP_bot.Inst_MULADD._0049_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0154_ Tile_X0Y1_DSP_bot.Inst_MULADD._0155_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0156_ sky130_fd_sc_hd__or4_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[348\] Tile_X0Y0_DSP_top.ConfigBits\[349\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1603_ Tile_X0Y1_DSP_bot.Inst_MULADD._0725_ Tile_X0Y1_DSP_bot.Inst_MULADD._0766_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0717_ Tile_X0Y1_DSP_bot.Inst_MULADD._0718_ Tile_X0Y1_DSP_bot.Inst_MULADD._0743_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0767_ sky130_fd_sc_hd__o41ai_2
X_307_ Tile_X0Y1_DSP_bot.S4BEG\[7\] VGND VGND VPWR VPWR net696 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1534_ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0698_ Tile_X0Y1_DSP_bot.Inst_MULADD._0699_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0700_ sky130_fd_sc_hd__a22o_1
X_238_ Tile_X0Y1_DSP_bot.EE4BEG\[6\] VGND VGND VPWR VPWR net627 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_169_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb5 VGND VGND VPWR VPWR net552
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1465_ Tile_X0Y1_DSP_bot.Inst_MULADD._0579_ Tile_X0Y1_DSP_bot.Inst_MULADD._0630_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0632_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0633_
+ sky130_fd_sc_hd__nand3_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1396_ Tile_X0Y1_DSP_bot.Inst_MULADD._0557_ Tile_X0Y1_DSP_bot.Inst_MULADD._0562_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0565_ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst1
+ net84 net92 net134 net136 Tile_X0Y0_DSP_top.ConfigBits\[334\] Tile_X0Y0_DSP_top.ConfigBits\[335\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9 net260 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[105\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[286\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[308\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput317 Tile_X0Y1_NN4END[0] VGND VGND VPWR VPWR net317 sky130_fd_sc_hd__buf_1
Xinput306 Tile_X0Y1_N4END[14] VGND VGND VPWR VPWR net306 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19 net239 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[339\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput339 Tile_X0Y1_W2END[1] VGND VGND VPWR VPWR net339 sky130_fd_sc_hd__buf_2
Xinput328 Tile_X0Y1_NN4END[5] VGND VGND VPWR VPWR net328 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_023_ Tile_X0Y0_DSP_top.E6BEG\[3\] VGND VGND VPWR VPWR net407 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[258\] Tile_X0Y0_DSP_top.ConfigBits\[259\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1250_ Tile_X0Y1_DSP_bot.Inst_MULADD._0342_ Tile_X0Y1_DSP_bot.Inst_MULADD._0417_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0420_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0421_
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1181_ Tile_X0Y1_DSP_bot.Inst_MULADD._0299_ Tile_X0Y1_DSP_bot.Inst_MULADD._0049_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0283_ Tile_X0Y1_DSP_bot.Inst_MULADD._0343_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0352_ sky130_fd_sc_hd__o211a_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID3
+ net16 net96 net148 Tile_X0Y0_DSP_top.ConfigBits\[184\] Tile_X0Y0_DSP_top.ConfigBits\[185\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_16_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0965_ Tile_X0Y1_DSP_bot.A4 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0139_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_inst0
+ net283 net183 net336 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.ConfigBits\[22\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[23\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_123_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0896_ Tile_X0Y1_DSP_bot.A0 Tile_X0Y1_DSP_bot.Inst_MULADD._0025_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0027_ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0072_ sky130_fd_sc_hd__o211a_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1517_ Tile_X0Y1_DSP_bot.Inst_MULADD._0677_ Tile_X0Y1_DSP_bot.Inst_MULADD._0679_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0682_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0684_
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot.NN4END_inbuf_11._0_ net323 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.data_outbuf_0._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[0\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1448_ Tile_X0Y1_DSP_bot.Inst_MULADD._0461_ Tile_X0Y1_DSP_bot.Inst_MULADD._0488_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0556_ Tile_X0Y1_DSP_bot.Inst_MULADD._0615_ Tile_X0Y1_DSP_bot.Inst_MULADD._0563_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0616_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_40_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1379_ Tile_X0Y1_DSP_bot.Inst_MULADD._0546_ Tile_X0Y1_DSP_bot.Inst_MULADD._0547_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0548_ sky130_fd_sc_hd__nand2_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[205\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[194\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_160_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[370\] Tile_X0Y1_DSP_bot.ConfigBits\[371\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG4 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[110\] Tile_X0Y0_DSP_top.ConfigBits\[111\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_3_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_11._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput114 Tile_X0Y0_S4END[7] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xinput125 Tile_X0Y0_SS4END[2] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_2
Xinput103 Tile_X0Y0_S4END[11] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.data_inbuf_24._0_ net65 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[24\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.WW4END_inbuf_2._0_ net177 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_1
Xinput136 Tile_X0Y0_W1END[3] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__buf_4
Xinput158 Tile_X0Y0_W6END[3] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_1
Xinput169 Tile_X0Y0_WW4END[13] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
Xinput147 Tile_X0Y0_W2MID[2] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[298\] Tile_X0Y0_DSP_top.ConfigBits\[299\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.strobe_inbuf_9._0_ Tile_X0Y0_DSP_top.FrameStrobe\[9\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[9\] sky130_fd_sc_hd__clkbuf_1
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[312\] Tile_X0Y0_DSP_top.ConfigBits\[313\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_006_ Tile_X0Y0_DSP_top.E2BEG\[2\] VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1302_ Tile_X0Y1_DSP_bot.Inst_MULADD._0468_ Tile_X0Y1_DSP_bot.Inst_MULADD._0470_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0471_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0472_
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END0
+ net117 net153 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 Tile_X0Y0_DSP_top.ConfigBits\[388\]
+ Tile_X0Y0_DSP_top.ConfigBits\[389\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1233_ Tile_X0Y1_DSP_bot.Inst_MULADD._0402_ Tile_X0Y1_DSP_bot.Inst_MULADD._0403_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0390_ Tile_X0Y1_DSP_bot.Inst_MULADD._0389_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0404_ sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1164_ Tile_X0Y1_DSP_bot.Inst_MULADD._0333_ Tile_X0Y1_DSP_bot.Inst_MULADD._0334_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0336_ sky130_fd_sc_hd__nor2_1
XTile_X0Y0_DSP_top.data_inbuf_15._0_ net55 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[15\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1095_ Tile_X0Y1_DSP_bot.Inst_MULADD._0266_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0267_ sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[44\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG\[12\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0948_ Tile_X0Y1_DSP_bot.Inst_MULADD._0121_ Tile_X0Y1_DSP_bot.Inst_MULADD._0122_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0082_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0123_
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29 net250 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[381\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18 net238 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[370\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0879_ Tile_X0Y1_DSP_bot.Inst_MULADD._0046_ Tile_X0Y1_DSP_bot.Inst_MULADD._0052_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0054_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0056_
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[113\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[102\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13 net233 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[13\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24 net245 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[24\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.data_outbuf_0._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[0\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._21_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG5 sky130_fd_sc_hd__clkbuf_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.ConfigBits\[280\] Tile_X0Y1_DSP_bot.ConfigBits\[281\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[89\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_208 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_219 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_118_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.SS4END_inbuf_8._0_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.data_inbuf_24._0_ net245 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[24\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_156_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1 net240 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[225\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_112_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput407 net407 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput418 net418 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput429 net429 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[9] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[225\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[236\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._83_ net351 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb5
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1216_ Tile_X0Y1_DSP_bot.Inst_MULADD._0385_ Tile_X0Y1_DSP_bot.Inst_MULADD._0386_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0290_ Tile_X0Y1_DSP_bot.Inst_MULADD._0289_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0387_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_129_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1147_ Tile_X0Y1_DSP_bot.Inst_MULADD._0223_ Tile_X0Y1_DSP_bot.Inst_MULADD._0250_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0307_ Tile_X0Y1_DSP_bot.Inst_MULADD._0318_ Tile_X0Y1_DSP_bot.Inst_MULADD._0313_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0319_ sky130_fd_sc_hd__o221ai_4
XTile_X0Y0_DSP_top.strobe_outbuf_1._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[1\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[1\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1078_ Tile_X0Y1_DSP_bot.Inst_MULADD._0224_ Tile_X0Y1_DSP_bot.Inst_MULADD._0225_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0157_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0250_
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y1_DSP_bot.data_inbuf_15._0_ net235 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[15\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_147_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[334\] Tile_X0Y1_DSP_bot.ConfigBits\[335\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[21\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 sky130_fd_sc_hd__o21ai_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._04_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG4
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_N4BEG0 net287 net308
+ net204 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[14\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[15\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.N4END\[12\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.inst_clk_buf net333 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.UserCLK
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_340_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG4 VGND VGND VPWR VPWR net723
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_271_ Tile_X0Y1_DSP_bot.FrameData_O\[23\] VGND VGND VPWR VPWR net646 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst0
+ net184 net337 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.ConfigBits\[110\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[111\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_121_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG0 net300
+ net200 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG7 net353 Tile_X0Y1_DSP_bot.ConfigBits\[200\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[201\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_121_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1001_ Tile_X0Y1_DSP_bot.Inst_MULADD._0174_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0175_ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28 net249 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[412\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.EE4END_inbuf_7._0_ net215 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17 net237 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[401\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[144\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[133\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12 net232 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[44\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23 net244 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[55\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.strobe_inbuf_16._0_ Tile_X0Y0_DSP_top.FrameStrobe\[16\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1696_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0746_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0841_ sky130_fd_sc_hd__and2b_1
XFILLER_0_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._66_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[370\] Tile_X0Y0_DSP_top.ConfigBits\[371\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[188\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_N1BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[12\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[13\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_81_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2 net251 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[66\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_128_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput760 net760 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.SS4END_inbuf_4._0_ net131 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[256\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[267\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG1 net288
+ net188 Tile_X0Y0_DSP_top.SS4BEG\[0\] net341 Tile_X0Y1_DSP_bot.ConfigBits\[250\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[251\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_83_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_323_ Tile_X0Y1_DSP_bot.SS4BEG\[7\] VGND VGND VPWR VPWR net712 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1550_ Tile_X0Y1_DSP_bot.C12 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[12\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0716_
+ sky130_fd_sc_hd__mux2_1
X_254_ Tile_X0Y1_DSP_bot.FrameData_O\[6\] VGND VGND VPWR VPWR net659 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4 net255 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[324\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_185_ Tile_X0Y0_DSP_top.WW4BEG\[1\] VGND VGND VPWR VPWR net574 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.strobe_outbuf_18._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[18\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[18\] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1481_ Tile_X0Y1_DSP_bot.Inst_MULADD._0025_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0648_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_142_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1748_ net333 Tile_X0Y1_DSP_bot.C6 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1679_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0181_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0833_ sky130_fd_sc_hd__and2b_1
XFILLER_0_2_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[23\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._49_ net296 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END3
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_148_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[164\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[175\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11 net231 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[75\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22 net243 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[86\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[27\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4END\[13\] sky130_fd_sc_hd__o21ai_1
Xoutput590 net590 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.EE4END_inbuf_3._0_ net46 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_88_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[38\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0981_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ Tile_X0Y1_DSP_bot.B4
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0152_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0155_
+ sky130_fd_sc_hd__o21ai_4
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1602_ Tile_X0Y1_DSP_bot.Inst_MULADD._0713_ Tile_X0Y1_DSP_bot.Inst_MULADD._0692_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0695_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0766_
+ sky130_fd_sc_hd__and3_1
X_306_ Tile_X0Y1_DSP_bot.S4BEG\[6\] VGND VGND VPWR VPWR net695 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1533_ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0696_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0697_ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0699_ sky130_fd_sc_hd__nand4_4
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_237_ Tile_X0Y1_DSP_bot.EE4BEG\[5\] VGND VGND VPWR VPWR net626 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_168_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb4 VGND VGND VPWR VPWR net551
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1464_ Tile_X0Y1_DSP_bot.Inst_MULADD._0624_ Tile_X0Y1_DSP_bot.Inst_MULADD._0626_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0631_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0632_
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_122_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_099_ Tile_X0Y0_DSP_top.FrameStrobe_O\[19\] VGND VGND VPWR VPWR net472 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1395_ Tile_X0Y1_DSP_bot.Inst_MULADD._0557_ Tile_X0Y1_DSP_bot.Inst_MULADD._0562_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0563_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0564_
+ sky130_fd_sc_hd__a21boi_4
XTile_X0Y1_DSP_bot.strobe_outbuf_7._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[7\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[7\] sky130_fd_sc_hd__clkbuf_16
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[334\] Tile_X0Y0_DSP_top.ConfigBits\[335\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.N4BEG_outbuf_2._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END2 sky130_fd_sc_hd__buf_2
XFILLER_0_1_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[287\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_62_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.E6END_inbuf_9._0_ net23 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[298\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[309\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_140_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput307 Tile_X0Y1_N4END[15] VGND VGND VPWR VPWR net307 sky130_fd_sc_hd__clkbuf_1
Xinput318 Tile_X0Y1_NN4END[10] VGND VGND VPWR VPWR net318 sky130_fd_sc_hd__clkbuf_1
Xinput329 Tile_X0Y1_NN4END[6] VGND VGND VPWR VPWR net329 sky130_fd_sc_hd__clkbuf_1
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_022_ Tile_X0Y0_DSP_top.E6BEG\[2\] VGND VGND VPWR VPWR net406 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[260\] Tile_X0Y0_DSP_top.ConfigBits\[261\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1180_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B7
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0346_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0351_
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_5._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[5\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst0
+ net287 net309 net181 net187 Tile_X0Y1_DSP_bot.ConfigBits\[260\] Tile_X0Y1_DSP_bot.ConfigBits\[261\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID5
+ net18 net98 net150 Tile_X0Y0_DSP_top.ConfigBits\[186\] Tile_X0Y0_DSP_top.ConfigBits\[187\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_69_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[22\] Tile_X0Y1_DSP_bot.ConfigBits\[23\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0964_ Tile_X0Y1_DSP_bot.Inst_MULADD._0044_ Tile_X0Y1_DSP_bot.Inst_MULADD._0112_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0137_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0138_ sky130_fd_sc_hd__o2bb2ai_4
XTile_X0Y0_DSP_top.E6BEG_outbuf_7._0_ Tile_X0Y0_DSP_top.E6BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0895_ Tile_X0Y1_DSP_bot.Inst_MULADD._0070_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ sky130_fd_sc_hd__buf_4
XFILLER_0_84_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[100\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1516_ Tile_X0Y1_DSP_bot.Inst_MULADD._0677_ Tile_X0Y1_DSP_bot.Inst_MULADD._0679_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0682_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0683_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_40_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.strobe_outbuf_13._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[13\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[13\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1447_ Tile_X0Y1_DSP_bot.Inst_MULADD._0552_ Tile_X0Y1_DSP_bot.Inst_MULADD._0554_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0535_ Tile_X0Y1_DSP_bot.Inst_MULADD._0539_ Tile_X0Y1_DSP_bot.Inst_MULADD._0559_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0615_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1378_ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ Tile_X0Y1_DSP_bot.Inst_MULADD._0543_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0545_ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0547_ sky130_fd_sc_hd__nand4_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.W6BEG_outbuf_2._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.data_inbuf_4._0_ net75 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_inst0
+ net281 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0 net334 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[104\] Tile_X0Y1_DSP_bot.ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[206\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[195\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net3 net83 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.ConfigBits\[36\] Tile_X0Y0_DSP_top.ConfigBits\[37\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_145_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.N4END_inbuf_0._0_ Tile_X0Y0_DSP_top.N4END\[4\] VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_i\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput126 Tile_X0Y0_SS4END[3] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_1
Xinput115 Tile_X0Y0_S4END[8] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
Xinput104 Tile_X0Y0_S4END[12] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.E6END_inbuf_9._0_ net203 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
Xinput159 Tile_X0Y0_W6END[4] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_1
Xinput137 Tile_X0Y0_W2END[0] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__buf_2
Xinput148 Tile_X0Y0_W2MID[3] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[298\] Tile_X0Y0_DSP_top.ConfigBits\[299\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_005_ Tile_X0Y0_DSP_top.E2BEG\[1\] VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1301_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B6
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ Tile_X0Y1_DSP_bot.Inst_MULADD._0293_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0471_ sky130_fd_sc_hd__o211a_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1232_ Tile_X0Y1_DSP_bot.Inst_MULADD._0365_ Tile_X0Y1_DSP_bot.Inst_MULADD._0371_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0403_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1163_ Tile_X0Y1_DSP_bot.Inst_MULADD._0325_ Tile_X0Y1_DSP_bot.Inst_MULADD._0331_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0333_ Tile_X0Y1_DSP_bot.Inst_MULADD._0334_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0335_ sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[44\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1094_ Tile_X0Y1_DSP_bot.Inst_MULADD._0026_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0266_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0947_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0120_ Tile_X0Y1_DSP_bot.Inst_MULADD._0117_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0122_ sky130_fd_sc_hd__a22o_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[340\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19 net239 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[371\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0878_ Tile_X0Y1_DSP_bot.Inst_MULADD._0046_ Tile_X0Y1_DSP_bot.Inst_MULADD._0052_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0054_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0055_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_127_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[114\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[103\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14 net234 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[14\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25 net246 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[25\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.data_outbuf_31._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[31\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[31\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.NN4BEG_outbuf_2._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._20_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG4 sky130_fd_sc_hd__clkbuf_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[282\] Tile_X0Y1_DSP_bot.ConfigBits\[283\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG6 sky130_fd_sc_hd__mux4_2
XFILLER_0_84_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[90\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_209 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.SS4BEG_outbuf_5._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.data_outbuf_22._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[22\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[22\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_133_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_121_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.N4END_inbuf_0._0_ net311 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[0\]
+ sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG0 net299
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG6 net352 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[160\] Tile_X0Y1_DSP_bot.ConfigBits\[161\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_156_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2 net251 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[226\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_81_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.data_outbuf_13._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[13\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput408 net408 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[4] sky130_fd_sc_hd__buf_2
XFILLER_0_112_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput419 net419 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[14] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[226\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[237\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._82_ net350 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb4
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1215_ Tile_X0Y1_DSP_bot.Inst_MULADD._0195_ Tile_X0Y1_DSP_bot.Inst_MULADD._0287_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0275_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0386_
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot.S4BEG_outbuf_2._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[2\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1146_ Tile_X0Y1_DSP_bot.Inst_MULADD._0303_ Tile_X0Y1_DSP_bot.Inst_MULADD._0317_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0298_ Tile_X0Y1_DSP_bot.Inst_MULADD._0301_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0318_ sky130_fd_sc_hd__o2bb2ai_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1077_ Tile_X0Y1_DSP_bot.Inst_MULADD._0183_ Tile_X0Y1_DSP_bot.Inst_MULADD._0245_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0244_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0249_
+ sky130_fd_sc_hd__o21bai_4
XFILLER_0_159_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[106\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_73 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[21\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_inst0
+ net283 net183 net336 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.ConfigBits\[78\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[79\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._03_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG3
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_N4BEG1 net288 net309
+ net201 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.ConfigBits\[16\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[17\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.N4END\[13\]
+ sky130_fd_sc_hd__mux4_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_270_ Tile_X0Y1_DSP_bot.FrameData_O\[22\] VGND VGND VPWR VPWR net645 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.ConfigBits\[110\] Tile_X0Y1_DSP_bot.ConfigBits\[111\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG1 net296
+ net196 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG3 net349 Tile_X0Y1_DSP_bot.ConfigBits\[202\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[203\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG1
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG0 Tile_X0Y0_DSP_top.ConfigBits\[112\]
+ Tile_X0Y0_DSP_top.ConfigBits\[113\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1000_ Tile_X0Y1_DSP_bot.Inst_MULADD._0168_ Tile_X0Y1_DSP_bot.Inst_MULADD._0171_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0173_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0174_
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29 net250 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[413\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18 net238 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[402\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[145\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[134\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13 net233 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[45\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24 net245 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[56\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1695_ Tile_X0Y1_DSP_bot.Inst_MULADD._0840_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._65_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb3 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[370\] Tile_X0Y0_DSP_top.ConfigBits\[371\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1129_ Tile_X0Y1_DSP_bot.Inst_MULADD._0205_ Tile_X0Y1_DSP_bot.Inst_MULADD._0215_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0301_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_156_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[189\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_81_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.NN4END_inbuf_8._0_ net320 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3 net254 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[67\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput750 net750 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput761 net761 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[8] sky130_fd_sc_hd__clkbuf_4
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[268\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[257\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG2 net324
+ net190 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb5 net343 Tile_X0Y1_DSP_bot.ConfigBits\[252\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[253\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG2
+ sky130_fd_sc_hd__mux4_2
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_322_ Tile_X0Y1_DSP_bot.SS4BEG\[6\] VGND VGND VPWR VPWR net711 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_253_ Tile_X0Y1_DSP_bot.FrameData_O\[5\] VGND VGND VPWR VPWR net658 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5 net256 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[325\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_184_ Tile_X0Y0_DSP_top.WW4BEG\[0\] VGND VGND VPWR VPWR net567 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1480_ Tile_X0Y1_DSP_bot.Inst_MULADD._0025_ Tile_X0Y1_DSP_bot.A7
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0647_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1747_ net333 Tile_X0Y1_DSP_bot.C5 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_8._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4END\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1678_ Tile_X0Y1_DSP_bot.Inst_MULADD._0832_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[24\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._48_ net295 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END2
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[176\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[165\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12 net232 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[76\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23 net244 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[87\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[27\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
Xoutput580 net580 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput591 net591 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[4] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_158_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0980_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ Tile_X0Y1_DSP_bot.Inst_MULADD._0100_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0101_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0154_
+ sky130_fd_sc_hd__o21a_2
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1601_ Tile_X0Y1_DSP_bot.Inst_MULADD._0763_ Tile_X0Y1_DSP_bot.Inst_MULADD._0764_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0765_ sky130_fd_sc_hd__nand2_1
X_305_ Tile_X0Y1_DSP_bot.S4BEG\[5\] VGND VGND VPWR VPWR net694 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1532_ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0696_ Tile_X0Y1_DSP_bot.Inst_MULADD._0697_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0698_ sky130_fd_sc_hd__a22o_1
X_236_ Tile_X0Y1_DSP_bot.EE4BEG\[4\] VGND VGND VPWR VPWR net625 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_167_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb3 VGND VGND VPWR VPWR net550
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1463_ Tile_X0Y1_DSP_bot.Inst_MULADD._0628_ Tile_X0Y1_DSP_bot.Inst_MULADD._0629_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0631_ sky130_fd_sc_hd__nor2_1
XFILLER_0_122_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_098_ Tile_X0Y0_DSP_top.FrameStrobe_O\[18\] VGND VGND VPWR VPWR net471 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1394_ Tile_X0Y1_DSP_bot.Inst_MULADD._0478_ Tile_X0Y1_DSP_bot.Inst_MULADD._0473_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0472_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0563_
+ sky130_fd_sc_hd__a21boi_4
XFILLER_0_20_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[334\] Tile_X0Y0_DSP_top.ConfigBits\[335\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END1 net40 Tile_X0Y0_DSP_top.ConfigBits\[278\]
+ Tile_X0Y0_DSP_top.ConfigBits\[279\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.NN4END_inbuf_4._0_ Tile_X0Y0_DSP_top.NN4END\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[299\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[288\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput308 Tile_X0Y1_N4END[1] VGND VGND VPWR VPWR net308 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput319 Tile_X0Y1_NN4END[11] VGND VGND VPWR VPWR net319 sky130_fd_sc_hd__clkbuf_1
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.EE4BEG_outbuf_5._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_021_ Tile_X0Y0_DSP_top.E6BEG\[1\] VGND VGND VPWR VPWR net405 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG0 net291
+ net191 Tile_X0Y0_DSP_top.SS4BEG\[3\] net344 Tile_X0Y1_DSP_bot.ConfigBits\[224\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[225\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst1
+ net201 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb2 net340 net354 Tile_X0Y1_DSP_bot.ConfigBits\[260\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[261\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID1
+ net14 net94 net146 Tile_X0Y0_DSP_top.ConfigBits\[188\] Tile_X0Y0_DSP_top.ConfigBits\[189\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0963_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.A4
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0136_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0137_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_29_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0 net229 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[128\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_139_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0894_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.Inst_MULADD._0068_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0069_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0070_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_154_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[100\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1515_ Tile_X0Y1_DSP_bot.Inst_MULADD._0680_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0682_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_219_ Tile_X0Y1_DSP_bot.E2BEGb\[7\] VGND VGND VPWR VPWR net602 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1446_ Tile_X0Y1_DSP_bot.Inst_MULADD._0611_ Tile_X0Y1_DSP_bot.Inst_MULADD._0612_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0613_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0614_
+ sky130_fd_sc_hd__a21boi_4
XFILLER_0_122_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1377_ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ Tile_X0Y1_DSP_bot.Inst_MULADD._0347_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0543_ Tile_X0Y1_DSP_bot.Inst_MULADD._0545_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0546_ sky130_fd_sc_hd__a22o_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[104\] Tile_X0Y1_DSP_bot.ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[207\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[196\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG0
+ Tile_X0Y0_DSP_top.ConfigBits\[36\] Tile_X0Y0_DSP_top.ConfigBits\[37\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput127 Tile_X0Y0_SS4END[4] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
Xinput116 Tile_X0Y0_S4END[9] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
Xinput105 Tile_X0Y0_S4END[13] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 net1 net133 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[22\] Tile_X0Y0_DSP_top.ConfigBits\[23\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
Xinput149 Tile_X0Y0_W2MID[4] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_2
Xinput138 Tile_X0Y0_W2END[1] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__buf_2
XFILLER_0_98_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[300\] Tile_X0Y0_DSP_top.ConfigBits\[301\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG5 sky130_fd_sc_hd__mux4_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst0
+ net283 net289 net301 net189 Tile_X0Y1_DSP_bot.ConfigBits\[300\] Tile_X0Y1_DSP_bot.ConfigBits\[301\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst0
+ net4 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.ConfigBits\[48\] Tile_X0Y0_DSP_top.ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_004_ Tile_X0Y0_DSP_top.E2BEG\[0\] VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1300_ Tile_X0Y1_DSP_bot.Inst_MULADD._0374_ Tile_X0Y1_DSP_bot.Inst_MULADD._0469_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0380_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0470_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0382_ Tile_X0Y1_DSP_bot.Inst_MULADD._0381_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0383_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0402_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1162_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] Tile_X0Y1_DSP_bot.Inst_MULADD._0085_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0334_ sky130_fd_sc_hd__and2b_1
XTile_X0Y1_DSP_bot.WW4END_inbuf_11._0_ net372 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1093_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.A6
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0265_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0946_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0117_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0120_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0121_ sky130_fd_sc_hd__nand4_4
XFILLER_0_84_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[341\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[330\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_127_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._0877_ Tile_X0Y1_DSP_bot.Inst_MULADD._0053_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[3\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0054_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[74\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG0 sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[104\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[115\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15 net235 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[15\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26 net247 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[26\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.S4END_inbuf_3._0_ net114 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1429_ Tile_X0Y1_DSP_bot.Inst_MULADD._0594_ Tile_X0Y1_DSP_bot.Inst_MULADD._0596_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0108_ Tile_X0Y1_DSP_bot.Inst_MULADD._0351_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0597_ sky130_fd_sc_hd__o2bb2ai_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[91\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END3
+ net8 net24 Tile_X0Y0_DSP_top.ConfigBits\[350\] Tile_X0Y0_DSP_top.ConfigBits\[351\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.strobe_inbuf_3._0_ net274 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[3\]
+ sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG1 net195
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG2 net348 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[162\] Tile_X0Y1_DSP_bot.ConfigBits\[163\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_156_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3 net254 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[227\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.W6END_inbuf_7._0_ net164 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._81_ net349 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb3
+ sky130_fd_sc_hd__clkbuf_1
Xoutput409 net409 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[227\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_10_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[238\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1214_ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0274_ Tile_X0Y1_DSP_bot.Inst_MULADD._0259_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0385_ sky130_fd_sc_hd__and4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1145_ Tile_X0Y1_DSP_bot.Inst_MULADD._0306_ Tile_X0Y1_DSP_bot.Inst_MULADD._0291_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0317_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1076_ Tile_X0Y1_DSP_bot.Inst_MULADD._0248_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 sky130_fd_sc_hd__buf_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[106\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._0929_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.S4END_inbuf_3._0_ Tile_X0Y0_DSP_top.S4BEG\[7\] VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.S4BEG_i\[3\] sky130_fd_sc_hd__clkbuf_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_inst1
+ net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[78\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[79\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._02_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEG\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_N4BEG2 net285 net310
+ net357 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.ConfigBits\[18\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[19\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.N4END\[14\]
+ sky130_fd_sc_hd__mux4_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[110\] Tile_X0Y1_DSP_bot.ConfigBits\[111\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.SS4END_inbuf_11._0_ net123 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG2 net298
+ net198 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG5 net351 Tile_X0Y1_DSP_bot.ConfigBits\[204\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[205\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG1 Tile_X0Y0_DSP_top.ConfigBits\[114\]
+ Tile_X0Y0_DSP_top.ConfigBits\[115\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[372\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19 net239 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[403\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[135\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[146\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_115_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14 net234 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[46\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25 net246 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[57\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1694_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0723_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0840_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_137_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.W6END_inbuf_7._0_ net365 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._64_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb2 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[372\] Tile_X0Y0_DSP_top.ConfigBits\[373\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG7 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1128_ Tile_X0Y1_DSP_bot.Inst_MULADD._0299_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0300_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst0
+ net283 net291 net183 net191 Tile_X0Y1_DSP_bot.ConfigBits\[372\] Tile_X0Y1_DSP_bot.ConfigBits\[373\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1059_ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0189_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0232_ sky130_fd_sc_hd__a41o_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[190\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_147_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[80\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG0 sky130_fd_sc_hd__o21ai_2
XFILLER_0_147_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4 net255 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[68\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput762 net762 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput751 net751 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput740 net740 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END2 net1 net41 net21 Tile_X0Y0_DSP_top.ConfigBits\[314\]
+ Tile_X0Y0_DSP_top.ConfigBits\[315\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[269\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[258\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_321_ Tile_X0Y1_DSP_bot.SS4BEG\[5\] VGND VGND VPWR VPWR net710 sky130_fd_sc_hd__clkbuf_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG3 net286
+ net222 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb1 net339 Tile_X0Y1_DSP_bot.ConfigBits\[254\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[255\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_76_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_252_ Tile_X0Y1_DSP_bot.FrameData_O\[4\] VGND VGND VPWR VPWR net657 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_183_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG1 VGND VGND VPWR VPWR net557
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6 net257 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[326\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_24_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.WW4END_inbuf_9._0_ net370 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1746_ net333 Tile_X0Y1_DSP_bot.C4 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1677_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0130_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0832_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[25\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_140_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._47_ net294 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END1
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_76_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_61_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[166\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_131_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[177\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13 net233 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[77\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24 net245 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[88\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_131_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput570 net570 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput581 net581 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput592 net592 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1600_ Tile_X0Y1_DSP_bot.Inst_MULADD._0755_ Tile_X0Y1_DSP_bot.Inst_MULADD._0760_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0762_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0764_
+ sky130_fd_sc_hd__nand3_2
X_304_ Tile_X0Y1_DSP_bot.S4BEG\[4\] VGND VGND VPWR VPWR net693 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1531_ Tile_X0Y1_DSP_bot.Inst_MULADD._0273_ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0660_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0697_
+ sky130_fd_sc_hd__o21ai_2
X_235_ Tile_X0Y1_DSP_bot.EE4BEG\[3\] VGND VGND VPWR VPWR net624 sky130_fd_sc_hd__clkbuf_1
X_166_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb2 VGND VGND VPWR VPWR net549
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1462_ Tile_X0Y1_DSP_bot.Inst_MULADD._0624_ Tile_X0Y1_DSP_bot.Inst_MULADD._0626_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0628_ Tile_X0Y1_DSP_bot.Inst_MULADD._0629_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0630_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_52_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ Tile_X0Y0_DSP_top.FrameStrobe_O\[17\] VGND VGND VPWR VPWR net470 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1393_ Tile_X0Y1_DSP_bot.Inst_MULADD._0484_ Tile_X0Y1_DSP_bot.Inst_MULADD._0558_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0560_ Tile_X0Y1_DSP_bot.Inst_MULADD._0561_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0562_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_122_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[336\] Tile_X0Y0_DSP_top.ConfigBits\[337\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 sky130_fd_sc_hd__mux4_2
XFILLER_0_137_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst1
+ net24 net86 net138 net156 Tile_X0Y0_DSP_top.ConfigBits\[278\] Tile_X0Y0_DSP_top.ConfigBits\[279\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst0
+ net282 net290 net182 net190 Tile_X0Y1_DSP_bot.ConfigBits\[336\] Tile_X0Y1_DSP_bot.ConfigBits\[337\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_190 Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1729_ net333 Tile_X0Y1_DSP_bot.A3 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_160_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.data_outbuf_3._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[3\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_140_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[300\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[289\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput309 Tile_X0Y1_N4END[2] VGND VGND VPWR VPWR net309 sky130_fd_sc_hd__buf_2
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_020_ Tile_X0Y0_DSP_top.E6BEG\[0\] VGND VGND VPWR VPWR net402 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.WW4END_inbuf_5._0_ net180 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG1 net317
+ net187 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb2 net340 Tile_X0Y1_DSP_bot.ConfigBits\[226\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[227\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG1
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.data_inbuf_27._0_ net68 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[27\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[260\] Tile_X0Y1_DSP_bot.ConfigBits\[261\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0962_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] Tile_X0Y1_DSP_bot.Inst_MULADD._0026_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0136_ sky130_fd_sc_hd__or2b_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1 net240 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[129\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[310\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0893_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0069_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_218_ Tile_X0Y1_DSP_bot.E2BEGb\[6\] VGND VGND VPWR VPWR net601 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1514_ Tile_X0Y1_DSP_bot.Inst_MULADD._0423_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ sky130_fd_sc_hd__clkbuf_4
X_149_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG1 VGND VGND VPWR VPWR net522
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1445_ Tile_X0Y1_DSP_bot.Inst_MULADD._0553_ Tile_X0Y1_DSP_bot.Inst_MULADD._0545_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0543_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0613_
+ sky130_fd_sc_hd__a21boi_2
XFILLER_0_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1376_ Tile_X0Y1_DSP_bot.Inst_MULADD._0108_ Tile_X0Y1_DSP_bot.Inst_MULADD._0299_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0445_ Tile_X0Y1_DSP_bot.Inst_MULADD._0544_ Tile_X0Y1_DSP_bot.Inst_MULADD._0452_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0545_ sky130_fd_sc_hd__o221ai_4
XTile_X0Y0_DSP_top.data_inbuf_18._0_ net58 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[18\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[208\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[197\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.data_outbuf_3._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[3\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[3\] sky130_fd_sc_hd__clkbuf_1
Xinput106 Tile_X0Y0_S4END[14] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
Xinput117 Tile_X0Y0_SS4END[0] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG1
+ Tile_X0Y0_DSP_top.ConfigBits\[22\] Tile_X0Y0_DSP_top.ConfigBits\[23\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
Xinput128 Tile_X0Y0_SS4END[5] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
Xinput139 Tile_X0Y0_W2END[2] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__buf_2
XFILLER_0_78_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.EE4END_inbuf_11._0_ net39 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst1
+ net201 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb4 net342 net354 Tile_X0Y1_DSP_bot.ConfigBits\[300\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[301\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[48\] Tile_X0Y0_DSP_top.ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_003_ Tile_X0Y0_DSP_top.E1BEG\[3\] VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_90 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.E6BEG_outbuf_1._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[1\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1230_ Tile_X0Y1_DSP_bot.Inst_MULADD._0392_ Tile_X0Y1_DSP_bot.Inst_MULADD._0399_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0400_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0401_
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1161_ Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ Tile_X0Y1_DSP_bot.Inst_MULADD._0332_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0333_ sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot.data_inbuf_27._0_ net248 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[27\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1092_ Tile_X0Y1_DSP_bot.Inst_MULADD._0261_ Tile_X0Y1_DSP_bot.Inst_MULADD._0263_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0264_
+ sky130_fd_sc_hd__o21ai_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0945_ Tile_X0Y1_DSP_bot.Inst_MULADD._0118_ Tile_X0Y1_DSP_bot.Inst_MULADD._0119_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0105_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0120_
+ sky130_fd_sc_hd__o21bai_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[331\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[320\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0876_ Tile_X0Y1_DSP_bot.C1 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[1\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[2\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0053_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[74\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[105\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16 net236 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[16\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_7_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27 net248 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[27\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1428_ Tile_X0Y1_DSP_bot.Inst_MULADD._0025_ Tile_X0Y1_DSP_bot.A4
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0136_ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_ Tile_X0Y1_DSP_bot.Inst_MULADD._0595_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0596_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1359_ Tile_X0Y1_DSP_bot.Inst_MULADD._0192_ Tile_X0Y1_DSP_bot.Inst_MULADD._0527_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0525_ Tile_X0Y1_DSP_bot.Inst_MULADD._0523_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0528_ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.strobe_outbuf_4._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[4\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[4\] sky130_fd_sc_hd__clkbuf_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.data_inbuf_18._0_ net238 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[18\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[92\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst1
+ net88 net110 net140 net156 Tile_X0Y0_DSP_top.ConfigBits\[350\] Tile_X0Y0_DSP_top.ConfigBits\[351\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG2 net297
+ net197 net350 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[164\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[165\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4 net255 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[228\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_81_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._80_ net348 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb2
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[228\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_10_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[239\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1213_ Tile_X0Y1_DSP_bot.Inst_MULADD._0381_ Tile_X0Y1_DSP_bot.Inst_MULADD._0382_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0383_ Tile_X0Y1_DSP_bot.Inst_MULADD._0365_ Tile_X0Y1_DSP_bot.Inst_MULADD._0371_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0384_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_129_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1144_ Tile_X0Y1_DSP_bot.Inst_MULADD._0254_ Tile_X0Y1_DSP_bot.Inst_MULADD._0315_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0316_ sky130_fd_sc_hd__nor2_1
XTile_X0Y0_DSP_top.WW4BEG_outbuf_2._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1075_ Tile_X0Y1_DSP_bot.Inst_MULADD._0247_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0248_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.strobe_inbuf_19._0_ Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[19\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG2.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0928_ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0859_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] Tile_X0Y1_DSP_bot.Inst_MULADD._0021_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0036_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0
+ sky130_fd_sc_hd__a21bo_4
XFILLER_0_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._01_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEG\[1\] sky130_fd_sc_hd__clkbuf_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_S1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG1 Tile_X0Y0_DSP_top.ConfigBits\[56\]
+ Tile_X0Y0_DSP_top.ConfigBits\[57\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux4_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_N4BEG3 net286 net301
+ net354 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.ConfigBits\[20\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[21\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.N4END\[15\]
+ sky130_fd_sc_hd__mux4_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END5
+ net2 net10 Tile_X0Y0_DSP_top.ConfigBits\[262\] Tile_X0Y0_DSP_top.ConfigBits\[263\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[110\] Tile_X0Y1_DSP_bot.ConfigBits\[111\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.strobe_inbuf_12._0_ net264 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[12\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_307 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG2 Tile_X0Y0_DSP_top.ConfigBits\[116\]
+ Tile_X0Y0_DSP_top.ConfigBits\[117\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG3 net294
+ net194 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG1 net347 Tile_X0Y1_DSP_bot.ConfigBits\[206\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[207\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG3
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[362\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[373\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.SS4END_inbuf_7._0_ net119 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[136\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[147\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26 net247 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[58\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15 net235 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[47\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_145_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 net1 net133 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[78\] Tile_X0Y0_DSP_top.ConfigBits\[79\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1693_ Tile_X0Y1_DSP_bot.Inst_MULADD._0839_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._63_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb1 sky130_fd_sc_hd__buf_1
XFILLER_0_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1127_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B6
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0293_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0299_
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb6 net336 Tile_X0Y1_DSP_bot.ConfigBits\[372\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[373\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1058_ Tile_X0Y1_DSP_bot.Inst_MULADD._0188_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[191\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[80\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5 net256 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[69\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput730 net730 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput752 net752 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput741 net741 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst1
+ net109 net125 net139 net153 Tile_X0Y0_DSP_top.ConfigBits\[314\] Tile_X0Y0_DSP_top.ConfigBits\[315\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_C0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[134\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[135\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C0 sky130_fd_sc_hd__mux4_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[270\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[259\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_320_ Tile_X0Y1_DSP_bot.SS4BEG\[4\] VGND VGND VPWR VPWR net709 sky130_fd_sc_hd__clkbuf_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot10 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG2 Tile_X0Y0_DSP_top.ConfigBits\[132\]
+ Tile_X0Y0_DSP_top.ConfigBits\[133\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot10
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_36_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_251_ Tile_X0Y1_DSP_bot.FrameData_O\[3\] VGND VGND VPWR VPWR net656 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_182_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 VGND VGND VPWR VPWR net556
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7 net258 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[327\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.EE4END_inbuf_6._0_ net34 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst0
+ net281 net285 net181 net213 Tile_X0Y1_DSP_bot.ConfigBits\[284\] Tile_X0Y1_DSP_bot.ConfigBits\[285\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1745_ net333 Tile_X0Y1_DSP_bot.C3 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1676_ Tile_X0Y1_DSP_bot.Inst_MULADD._0831_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._46_ net293 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END0
+ sky130_fd_sc_hd__buf_2
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[26\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.WW4BEG_outbuf_10._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG\[10\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.N4BEG_outbuf_5._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4END\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_148_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[404\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[167\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[178\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25 net246 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[89\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14 net234 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[78\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_131_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput560 net560 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput571 net571 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput582 net582 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput593 net593 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[6] sky130_fd_sc_hd__clkbuf_4
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_126_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_303_ Tile_X0Y1_DSP_bot.S4BEG\[3\] VGND VGND VPWR VPWR net692 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1530_ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_ Tile_X0Y1_DSP_bot.Inst_MULADD._0660_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0696_ sky130_fd_sc_hd__or2_2
X_234_ Tile_X0Y1_DSP_bot.EE4BEG\[2\] VGND VGND VPWR VPWR net623 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_165_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb1 VGND VGND VPWR VPWR net548
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1461_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] Tile_X0Y1_DSP_bot.Inst_MULADD._0423_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0629_ sky130_fd_sc_hd__and2b_1
X_096_ Tile_X0Y0_DSP_top.FrameStrobe_O\[16\] VGND VGND VPWR VPWR net469 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1392_ Tile_X0Y1_DSP_bot.Inst_MULADD._0552_ Tile_X0Y1_DSP_bot.Inst_MULADD._0554_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0551_ Tile_X0Y1_DSP_bot.Inst_MULADD._0534_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0561_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_122_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_8._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_137_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[278\] Tile_X0Y0_DSP_top.ConfigBits\[279\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb5
+ net335 net337 Tile_X0Y1_DSP_bot.ConfigBits\[336\] Tile_X0Y1_DSP_bot.ConfigBits\[337\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_180 Tile_X0Y0_DSP_top.S4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1728_ net333 Tile_X0Y1_DSP_bot.A2 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top.strobe_outbuf_16._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[16\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[16\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1659_ Tile_X0Y1_DSP_bot.Inst_MULADD._0813_ Tile_X0Y1_DSP_bot.Inst_MULADD._0814_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0818_ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0819_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_140_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[290\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.W6BEG_outbuf_5._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[5\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[301\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.data_inbuf_7._0_ net78 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._29_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG7
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.N4END_inbuf_3._0_ Tile_X0Y0_DSP_top.N4END\[7\] VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_i\[3\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG2 net289
+ net213 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb4 net342 Tile_X0Y1_DSP_bot.ConfigBits\[228\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[229\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG2
+ sky130_fd_sc_hd__mux4_2
Xoutput390 net390 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[260\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[261\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0961_ Tile_X0Y1_DSP_bot.Inst_MULADD._0133_ Tile_X0Y1_DSP_bot.Inst_MULADD._0134_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0117_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0135_
+ sky130_fd_sc_hd__o21ai_4
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2 net251 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[130\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[311\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0892_ Tile_X0Y1_DSP_bot.B2 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0068_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_84_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1513_ Tile_X0Y1_DSP_bot.C11 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[11\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0680_
+ sky130_fd_sc_hd__mux2_1
X_217_ Tile_X0Y1_DSP_bot.E2BEGb\[5\] VGND VGND VPWR VPWR net600 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_148_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 VGND VGND VPWR VPWR net521
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1444_ Tile_X0Y1_DSP_bot.Inst_MULADD._0549_ Tile_X0Y1_DSP_bot.Inst_MULADD._0607_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0610_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0612_
+ sky130_fd_sc_hd__nand3_4
X_079_ Tile_X0Y0_DSP_top.FrameData_O\[31\] VGND VGND VPWR VPWR net454 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1375_ Tile_X0Y1_DSP_bot.Inst_MULADD._0155_ Tile_X0Y1_DSP_bot.Inst_MULADD._0137_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0449_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0544_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[198\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.N4BEG_outbuf_1._0_ Tile_X0Y0_DSP_top.N4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[209\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.NN4BEG_outbuf_5._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[5\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput107 Tile_X0Y0_S4END[15] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xinput118 Tile_X0Y0_SS4END[10] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
Xinput129 Tile_X0Y0_SS4END[6] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.SS4BEG_outbuf_8._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[48\] Tile_X0Y0_DSP_top.ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[300\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[301\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.data_outbuf_25._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[25\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[25\] sky130_fd_sc_hd__clkbuf_1
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_002_ Tile_X0Y0_DSP_top.E1BEG\[2\] VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__clkbuf_1
XANTENNA_80 Tile_X0Y0_DSP_top.W6BEG\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.N4END_inbuf_3._0_ net314 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1160_ Tile_X0Y1_DSP_bot.C6 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[6\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0332_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1091_ Tile_X0Y1_DSP_bot.Inst_MULADD._0262_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0263_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0944_ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0109_ Tile_X0Y1_DSP_bot.Inst_MULADD._0114_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0119_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_69_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[332\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[321\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_57_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0875_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ Tile_X0Y1_DSP_bot.Inst_MULADD._0049_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0050_ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0052_ sky130_fd_sc_hd__or4_2
XFILLER_0_115_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.data_outbuf_16._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[16\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17 net237 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[17\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_80_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28 net249 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[28\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1427_ Tile_X0Y1_DSP_bot.Inst_MULADD._0525_ Tile_X0Y1_DSP_bot.Inst_MULADD._0523_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0192_ Tile_X0Y1_DSP_bot.Inst_MULADD._0527_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0595_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_1._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.S4BEG_outbuf_5._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[5\] sky130_fd_sc_hd__buf_2
XFILLER_0_110_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1358_ Tile_X0Y1_DSP_bot.Inst_MULADD._0265_ Tile_X0Y1_DSP_bot.Inst_MULADD._0267_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0527_ sky130_fd_sc_hd__o211ai_4
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.W6BEG_outbuf_1._0_ Tile_X0Y0_DSP_top.W6BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1289_ Tile_X0Y1_DSP_bot.Inst_MULADD._0369_ Tile_X0Y1_DSP_bot.Inst_MULADD._0370_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0459_ sky130_fd_sc_hd__nand2_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[93\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[350\] Tile_X0Y0_DSP_top.ConfigBits\[351\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG3 net293
+ net193 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[166\] Tile_X0Y1_DSP_bot.ConfigBits\[167\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_98_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5 net256 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[229\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[240\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_120_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[229\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1212_ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0375_ Tile_X0Y1_DSP_bot.Inst_MULADD._0372_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0383_ sky130_fd_sc_hd__a22o_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1143_ Tile_X0Y1_DSP_bot.Inst_MULADD._0305_ Tile_X0Y1_DSP_bot.Inst_MULADD._0313_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0314_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0315_
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1074_ Tile_X0Y1_DSP_bot.Inst_MULADD._0183_ Tile_X0Y1_DSP_bot.Inst_MULADD._0246_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0247_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_159_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0927_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ Tile_X0Y1_DSP_bot.Inst_MULADD._0100_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0101_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0102_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_155_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_115_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0858_ Tile_X0Y1_DSP_bot.ConfigBits\[5\] Tile_X0Y1_DSP_bot.Inst_MULADD._0034_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0035_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0036_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_5_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.data_outbuf_30._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[30\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[30\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._00_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEG\[0\] sky130_fd_sc_hd__clkbuf_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_S1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG2 Tile_X0Y0_DSP_top.ConfigBits\[58\]
+ Tile_X0Y0_DSP_top.ConfigBits\[59\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__mux4_2
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst1
+ net82 net90 net134 net136 Tile_X0Y0_DSP_top.ConfigBits\[262\] Tile_X0Y0_DSP_top.ConfigBits\[263\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_inbuf_0._0_ net229 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[112\] Tile_X0Y1_DSP_bot.ConfigBits\[113\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.data_outbuf_21._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[21\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[21\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG3 Tile_X0Y0_DSP_top.ConfigBits\[118\]
+ Tile_X0Y0_DSP_top.ConfigBits\[119\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_12_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[363\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[352\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[137\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16 net236 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[48\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27 net248 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[59\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1761_ net333 Tile_X0Y1_DSP_bot.C19 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1692_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0687_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0839_ sky130_fd_sc_hd__and2b_1
XFILLER_0_54_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG3
+ Tile_X0Y0_DSP_top.ConfigBits\[78\] Tile_X0Y0_DSP_top.ConfigBits\[79\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.data_outbuf_12._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[12\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._62_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb0 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.S4BEG_outbuf_1._0_ Tile_X0Y0_DSP_top.S4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1126_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0297_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0298_
+ sky130_fd_sc_hd__and3_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[372\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[373\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1057_ Tile_X0Y1_DSP_bot.Inst_MULADD._0141_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ sky130_fd_sc_hd__buf_4
Xinput290 Tile_X0Y1_N2END[5] VGND VGND VPWR VPWR net290 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[146\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG0.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_81_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6 net257 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[70\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_81_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END7
+ net4 net12 Tile_X0Y0_DSP_top.ConfigBits\[302\] Tile_X0Y0_DSP_top.ConfigBits\[303\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput720 net720 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput731 net731 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput753 net753 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput742 net742 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[314\] Tile_X0Y0_DSP_top.ConfigBits\[315\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_C1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[136\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[137\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C1 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_B0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[126\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[127\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B0 sky130_fd_sc_hd__mux4_2
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[271\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[260\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot11 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG3 Tile_X0Y0_DSP_top.ConfigBits\[134\]
+ Tile_X0Y0_DSP_top.ConfigBits\[135\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot11
+ sky130_fd_sc_hd__mux4_1
X_250_ Tile_X0Y1_DSP_bot.FrameData_O\[2\] VGND VGND VPWR VPWR net653 sky130_fd_sc_hd__clkbuf_1
X_181_ Tile_X0Y0_DSP_top.W6BEG\[9\] VGND VGND VPWR VPWR net566 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8 net259 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[328\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_134_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_129_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1744_ net333 Tile_X0Y1_DSP_bot.C2 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb0
+ net334 net336 Tile_X0Y1_DSP_bot.ConfigBits\[284\] Tile_X0Y1_DSP_bot.ConfigBits\[285\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
X_379_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR net753
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1675_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0093_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_152_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._45_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG7
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID7 sky130_fd_sc_hd__buf_2
XFILLER_0_50_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[27\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1109_ Tile_X0Y1_DSP_bot.Inst_MULADD._0255_ Tile_X0Y1_DSP_bot.Inst_MULADD._0277_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0280_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0281_
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_148_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.NN4END_inbuf_7._0_ Tile_X0Y0_DSP_top.NN4END\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[405\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[394\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[168\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15 net235 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[79\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[179\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26 net247 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[90\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput561 net561 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput572 net572 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput550 net550 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[3] sky130_fd_sc_hd__clkbuf_4
Xoutput583 net583 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput594 net594 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.EE4BEG_outbuf_8._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_302_ Tile_X0Y1_DSP_bot.S4BEG\[2\] VGND VGND VPWR VPWR net691 sky130_fd_sc_hd__clkbuf_1
X_233_ Tile_X0Y1_DSP_bot.EE4BEG\[1\] VGND VGND VPWR VPWR net622 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_164_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb0 VGND VGND VPWR VPWR net547
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1460_ Tile_X0Y1_DSP_bot.Inst_MULADD._0423_ Tile_X0Y1_DSP_bot.Inst_MULADD._0627_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0628_ sky130_fd_sc_hd__nor2_1
X_095_ Tile_X0Y0_DSP_top.FrameStrobe_O\[15\] VGND VGND VPWR VPWR net468 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1391_ Tile_X0Y1_DSP_bot.Inst_MULADD._0535_ Tile_X0Y1_DSP_bot.Inst_MULADD._0539_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0555_ Tile_X0Y1_DSP_bot.Inst_MULADD._0559_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0560_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_20_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[278\] Tile_X0Y0_DSP_top.ConfigBits\[279\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[336\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[337\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_157_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_170 Tile_X0Y0_DSP_top.FrameStrobe\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_181 Tile_X0Y0_DSP_top.S4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_145_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1727_ net333 Tile_X0Y1_DSP_bot.A1 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_1._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1658_ Tile_X0Y1_DSP_bot.Inst_MULADD._0816_ Tile_X0Y1_DSP_bot.Inst_MULADD._0817_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0818_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1589_ Tile_X0Y1_DSP_bot.Inst_MULADD._0752_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0753_ sky130_fd_sc_hd__inv_2
XFILLER_0_70_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[291\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[302\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._28_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.N4END_inbuf_11._0_ net307 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID6
+ net19 net99 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 Tile_X0Y0_DSP_top.ConfigBits\[174\]
+ Tile_X0Y0_DSP_top.ConfigBits\[175\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG3 net285
+ net185 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb0 net375 Tile_X0Y1_DSP_bot.ConfigBits\[230\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[231\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG3
+ sky130_fd_sc_hd__mux4_2
Xoutput391 net391 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[262\] Tile_X0Y1_DSP_bot.ConfigBits\[263\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG1 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0960_ Tile_X0Y1_DSP_bot.Inst_MULADD._0115_ Tile_X0Y1_DSP_bot.Inst_MULADD._0116_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0105_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0134_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3 net254 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[131\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0891_ Tile_X0Y1_DSP_bot.ConfigBits\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[312\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1512_ Tile_X0Y1_DSP_bot.Inst_MULADD._0614_ Tile_X0Y1_DSP_bot.Inst_MULADD._0618_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0623_ Tile_X0Y1_DSP_bot.Inst_MULADD._0625_ Tile_X0Y1_DSP_bot.Inst_MULADD._0678_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0679_ sky130_fd_sc_hd__o221ai_4
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_216_ Tile_X0Y1_DSP_bot.E2BEGb\[4\] VGND VGND VPWR VPWR net599 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_147_ Tile_X0Y0_DSP_top.NN4BEG\[11\] VGND VGND VPWR VPWR net520 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1443_ Tile_X0Y1_DSP_bot.Inst_MULADD._0607_ Tile_X0Y1_DSP_bot.Inst_MULADD._0610_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0549_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0611_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_078_ Tile_X0Y0_DSP_top.FrameData_O\[30\] VGND VGND VPWR VPWR net453 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1374_ Tile_X0Y1_DSP_bot.Inst_MULADD._0540_ Tile_X0Y1_DSP_bot.Inst_MULADD._0541_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0542_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0543_
+ sky130_fd_sc_hd__o21ai_2
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[199\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[210\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.S4END_inbuf_6._0_ net102 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[6\]
+ sky130_fd_sc_hd__buf_4
XFILLER_0_160_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 VGND VGND VPWR VPWR net763
+ sky130_fd_sc_hd__buf_8
XFILLER_0_101_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput108 Tile_X0Y0_S4END[1] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_4
Xinput119 Tile_X0Y0_SS4END[11] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.ConfigBits\[300\] Tile_X0Y1_DSP_bot.ConfigBits\[301\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1
+ Tile_X0Y0_DSP_top.ConfigBits\[48\] Tile_X0Y0_DSP_top.ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_70 Tile_X0Y0_DSP_top.S4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_001_ Tile_X0Y0_DSP_top.E1BEG\[1\] VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__clkbuf_1
XANTENNA_81 Tile_X0Y1_DSP_bot.E6BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_22_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.strobe_inbuf_6._0_ net277 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1090_ Tile_X0Y1_DSP_bot.Inst_MULADD._0026_ Tile_X0Y1_DSP_bot.A5
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0262_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0943_ Tile_X0Y1_DSP_bot.Inst_MULADD._0064_ Tile_X0Y1_DSP_bot.Inst_MULADD._0065_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ Tile_X0Y1_DSP_bot.Inst_MULADD._0109_ Tile_X0Y1_DSP_bot.Inst_MULADD._0114_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0118_ sky130_fd_sc_hd__o2111a_1
XTile_X0Y0_DSP_top.SS4BEG_outbuf_10._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG\[10\] sky130_fd_sc_hd__clkbuf_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[333\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[322\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0874_ Tile_X0Y1_DSP_bot.A0 Tile_X0Y1_DSP_bot.Inst_MULADD._0037_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0027_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0051_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_127_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18 net238 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[18\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29 net250 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[29\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1426_ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0523_ Tile_X0Y1_DSP_bot.Inst_MULADD._0525_ Tile_X0Y1_DSP_bot.Inst_MULADD._0593_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0594_ sky130_fd_sc_hd__a221o_2
XFILLER_0_7_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1357_ Tile_X0Y1_DSP_bot.Inst_MULADD._0523_ Tile_X0Y1_DSP_bot.Inst_MULADD._0524_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0525_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0526_
+ sky130_fd_sc_hd__a21oi_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1288_ Tile_X0Y1_DSP_bot.Inst_MULADD._0451_ Tile_X0Y1_DSP_bot.Inst_MULADD._0453_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0455_ Tile_X0Y1_DSP_bot.Inst_MULADD._0457_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0458_ sky130_fd_sc_hd__a22o_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[94\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_95_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.NN4END_inbuf_11._0_ Tile_X0Y0_DSP_top.NN4END\[15\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_1
Xinput90 Tile_X0Y0_S2END[5] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.S4END_inbuf_6._0_ Tile_X0Y0_DSP_top.S4BEG\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[350\] Tile_X0Y0_DSP_top.ConfigBits\[351\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_149_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6 net257 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[230\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END0
+ net1 net5 Tile_X0Y0_DSP_top.ConfigBits\[338\] Tile_X0Y0_DSP_top.ConfigBits\[339\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[230\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[241\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1211_ Tile_X0Y1_DSP_bot.Inst_MULADD._0108_ Tile_X0Y1_DSP_bot.Inst_MULADD._0155_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0137_ Tile_X0Y1_DSP_bot.Inst_MULADD._0154_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0382_ sky130_fd_sc_hd__o22a_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1142_ Tile_X0Y1_DSP_bot.Inst_MULADD._0157_ Tile_X0Y1_DSP_bot.Inst_MULADD._0237_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0251_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0314_
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1073_ Tile_X0Y1_DSP_bot.Inst_MULADD._0244_ Tile_X0Y1_DSP_bot.Inst_MULADD._0245_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0926_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0101_ sky130_fd_sc_hd__nand2_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0857_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0023_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0035_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1409_ Tile_X0Y1_DSP_bot.Inst_MULADD._0577_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0423_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0578_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot.S4END_inbuf_11._0_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.S4BEG_i\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_S1BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG3 Tile_X0Y0_DSP_top.ConfigBits\[60\]
+ Tile_X0Y0_DSP_top.ConfigBits\[61\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2
+ sky130_fd_sc_hd__mux4_2
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[262\] Tile_X0Y0_DSP_top.ConfigBits\[263\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_88_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[152\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C8 sky130_fd_sc_hd__o21ai_1
XTile_X0Y0_DSP_top.strobe_inbuf_2._0_ Tile_X0Y0_DSP_top.FrameStrobe\[2\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[2\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG0 Tile_X0Y0_DSP_top.ConfigBits\[120\]
+ Tile_X0Y0_DSP_top.ConfigBits\[121\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot4
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[353\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[364\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._59_ net148 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb3
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17 net237 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[49\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28 net249 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[60\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1760_ net333 Tile_X0Y1_DSP_bot.C18 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_156_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1691_ Tile_X0Y1_DSP_bot.Inst_MULADD._0838_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._61_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG7 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1125_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ Tile_X0Y1_DSP_bot.Inst_MULADD._0206_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_ Tile_X0Y1_DSP_bot.Inst_MULADD._0296_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0297_ sky130_fd_sc_hd__a31oi_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.ConfigBits\[372\] Tile_X0Y1_DSP_bot.ConfigBits\[373\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1056_ Tile_X0Y1_DSP_bot.Inst_MULADD._0050_ Tile_X0Y1_DSP_bot.Inst_MULADD._0137_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0192_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0229_ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput280 Tile_X0Y1_FrameStrobe[9] VGND VGND VPWR VPWR net280 sky130_fd_sc_hd__clkbuf_16
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[146\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
Xinput291 Tile_X0Y1_N2END[6] VGND VGND VPWR VPWR net291 sky130_fd_sc_hd__buf_2
XFILLER_0_18_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7 net258 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[71\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0909_ Tile_X0Y1_DSP_bot.ConfigBits\[3\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst1
+ net82 net84 net92 net136 Tile_X0Y0_DSP_top.ConfigBits\[302\] Tile_X0Y0_DSP_top.ConfigBits\[303\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_53_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput721 net721 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput710 net710 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput754 net754 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput732 net732 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput743 net743 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_W1BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[90\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[91\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[314\] Tile_X0Y0_DSP_top.ConfigBits\[315\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_C2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[138\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[139\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C2 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_B1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[128\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[129\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B1 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_A0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[118\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[119\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A0 sky130_fd_sc_hd__mux4_2
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[261\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[272\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.SS4END_inbuf_1._0_ Tile_X0Y0_DSP_top.SS4BEG\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot12 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG0 Tile_X0Y0_DSP_top.ConfigBits\[136\]
+ Tile_X0Y0_DSP_top.ConfigBits\[137\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot12
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_134_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_180_ Tile_X0Y0_DSP_top.W6BEG\[8\] VGND VGND VPWR VPWR net565 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9 net260 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[329\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_126_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[214\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1743_ net333 Tile_X0Y1_DSP_bot.C1 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_378_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net752
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[284\] Tile_X0Y1_DSP_bot.ConfigBits\[285\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_55_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1674_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._44_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID6 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[28\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1108_ Tile_X0Y1_DSP_bot.Inst_MULADD._0274_ Tile_X0Y1_DSP_bot.Inst_MULADD._0259_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0278_ Tile_X0Y1_DSP_bot.Inst_MULADD._0279_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0280_ sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1039_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0212_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.data_outbuf_6._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[6\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[6\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[384\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[395\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_131_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[169\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16 net236 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[80\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27 net248 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[91\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput562 net562 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput551 net551 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput540 net540 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput573 net573 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput584 net584 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput595 net595 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[0] sky130_fd_sc_hd__buf_2
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.EE4END_inbuf_0._0_ net223 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_301_ Tile_X0Y1_DSP_bot.S4BEG\[1\] VGND VGND VPWR VPWR net690 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_11._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.NN4END\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_232_ Tile_X0Y1_DSP_bot.EE4BEG\[0\] VGND VGND VPWR VPWR net615 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_163_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG7 VGND VGND VPWR VPWR net546
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_094_ Tile_X0Y0_DSP_top.FrameStrobe_O\[14\] VGND VGND VPWR VPWR net467 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1390_ Tile_X0Y1_DSP_bot.Inst_MULADD._0463_ Tile_X0Y1_DSP_bot.Inst_MULADD._0457_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0529_ Tile_X0Y1_DSP_bot.Inst_MULADD._0533_ Tile_X0Y1_DSP_bot.Inst_MULADD._0443_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0559_ sky130_fd_sc_hd__a221o_2
XTile_X0Y0_DSP_top.WW4END_inbuf_8._0_ net168 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[280\] Tile_X0Y0_DSP_top.ConfigBits\[281\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.ConfigBits\[336\] Tile_X0Y1_DSP_bot.ConfigBits\[337\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_160 Tile_X0Y0_DSP_top.FrameStrobe\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_193 Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 Tile_X0Y0_DSP_top.S4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_171 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_157_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1726_ net333 Tile_X0Y1_DSP_bot.A0 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1657_ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.Inst_MULADD._0810_
+ Tile_X0Y1_DSP_bot.ConfigBits\[4\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0817_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_140_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1588_ Tile_X0Y1_DSP_bot.Inst_MULADD._0711_ Tile_X0Y1_DSP_bot.Inst_MULADD._0734_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0752_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[303\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_121_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[292\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._27_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID2
+ net95 net147 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG6 Tile_X0Y0_DSP_top.ConfigBits\[176\]
+ Tile_X0Y0_DSP_top.ConfigBits\[177\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_outbuf_6._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[6\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput392 net392 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[6] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.strobe_outbuf_11._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[11\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[11\] sky130_fd_sc_hd__buf_8
XFILLER_0_69_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0890_ Tile_X0Y1_DSP_bot.Inst_MULADD._0064_ Tile_X0Y1_DSP_bot.Inst_MULADD._0065_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0066_
+ sky130_fd_sc_hd__o21ai_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4 net255 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[132\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[313\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_113_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1511_ Tile_X0Y1_DSP_bot.Inst_MULADD._0676_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0678_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_215_ Tile_X0Y1_DSP_bot.E2BEGb\[3\] VGND VGND VPWR VPWR net598 sky130_fd_sc_hd__clkbuf_1
X_146_ Tile_X0Y0_DSP_top.NN4BEG\[10\] VGND VGND VPWR VPWR net519 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1442_ Tile_X0Y1_DSP_bot.Inst_MULADD._0597_ Tile_X0Y1_DSP_bot.Inst_MULADD._0598_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0608_ Tile_X0Y1_DSP_bot.Inst_MULADD._0609_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0610_ sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot.E6BEG_outbuf_4._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_077_ Tile_X0Y0_DSP_top.FrameData_O\[29\] VGND VGND VPWR VPWR net451 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1373_ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_ Tile_X0Y1_DSP_bot.Inst_MULADD._0107_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0196_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0542_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_20_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[200\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[211\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1709_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0003_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 VGND VGND VPWR VPWR net764
+ sky130_fd_sc_hd__clkbuf_8
XTile_X0Y0_DSP_top.strobe_outbuf_7._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[7\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[7\] sky130_fd_sc_hd__clkbuf_1
Xinput109 Tile_X0Y0_S4END[2] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_2
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[302\] Tile_X0Y1_DSP_bot.ConfigBits\[303\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG3 sky130_fd_sc_hd__mux4_2
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[50\] Tile_X0Y0_DSP_top.ConfigBits\[51\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.E6BEG\[10\] sky130_fd_sc_hd__mux4_1
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_151_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_71 Tile_X0Y0_DSP_top.S4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_000_ Tile_X0Y0_DSP_top.E1BEG\[0\] VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_60 Tile_X0Y0_DSP_top.N4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_82 Tile_X0Y1_DSP_bot.E6BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.strobe_outbuf_0._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[0\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[0\] sky130_fd_sc_hd__buf_8
XFILLER_0_134_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0942_ Tile_X0Y1_DSP_bot.Inst_MULADD._0105_ Tile_X0Y1_DSP_bot.Inst_MULADD._0115_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0116_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0117_
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_69_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[334\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[323\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0873_ Tile_X0Y1_DSP_bot.Inst_MULADD._0047_ Tile_X0Y1_DSP_bot.B1
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0043_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0050_
+ sky130_fd_sc_hd__a21boi_4
XFILLER_0_127_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[20\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_159_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19 net239 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[19\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_129_ Tile_X0Y0_DSP_top.N4BEG\[9\] VGND VGND VPWR VPWR net517 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1425_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0593_ sky130_fd_sc_hd__and4_1
XFILLER_0_110_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1356_ Tile_X0Y1_DSP_bot.Inst_MULADD._0025_ Tile_X0Y1_DSP_bot.A4
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0136_ Tile_X0Y1_DSP_bot.Inst_MULADD._0213_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0525_ sky130_fd_sc_hd__o211a_1
XTile_X0Y0_DSP_top.WW4BEG_outbuf_5._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[5\] sky130_fd_sc_hd__clkbuf_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1287_ Tile_X0Y1_DSP_bot.Inst_MULADD._0368_ Tile_X0Y1_DSP_bot.Inst_MULADD._0366_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0358_ Tile_X0Y1_DSP_bot.Inst_MULADD._0456_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0457_ sky130_fd_sc_hd__o211ai_4
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.E6END_inbuf_2._0_ net27 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[95\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput91 Tile_X0Y0_S2END[6] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__buf_2
Xinput80 Tile_X0Y0_FrameData[9] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[352\] Tile_X0Y0_DSP_top.ConfigBits\[353\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_149_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_S4BEG0 net24 net87
+ net108 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.ConfigBits\[64\]
+ Tile_X0Y0_DSP_top.ConfigBits\[65\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst0
+ net284 net286 net186 net204 Tile_X0Y1_DSP_bot.ConfigBits\[352\] Tile_X0Y1_DSP_bot.ConfigBits\[353\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.strobe_inbuf_15._0_ net267 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[15\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7 net258 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[231\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst1
+ net81 net85 net133 net135 Tile_X0Y0_DSP_top.ConfigBits\[338\] Tile_X0Y0_DSP_top.ConfigBits\[339\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[231\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.E6BEG_outbuf_0._0_ Tile_X0Y0_DSP_top.E6BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[0\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[242\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1210_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ Tile_X0Y1_DSP_bot.Inst_MULADD._0380_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0381_ sky130_fd_sc_hd__a41o_1
XFILLER_0_120_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1141_ Tile_X0Y1_DSP_bot.Inst_MULADD._0307_ Tile_X0Y1_DSP_bot.Inst_MULADD._0309_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0312_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0313_
+ sky130_fd_sc_hd__o21bai_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1072_ Tile_X0Y1_DSP_bot.Inst_MULADD._0243_ Tile_X0Y1_DSP_bot.Inst_MULADD._0241_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0240_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0245_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_97_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0925_ Tile_X0Y1_DSP_bot.B3 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0100_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_155_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0856_ Tile_X0Y1_DSP_bot.Inst_MULADD._0023_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0034_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_38_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1408_ Tile_X0Y1_DSP_bot.C9 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[9\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0577_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1339_ Tile_X0Y1_DSP_bot.Inst_MULADD._0421_ Tile_X0Y1_DSP_bot.Inst_MULADD._0424_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0509_ sky130_fd_sc_hd__nand2_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_S1BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG0 Tile_X0Y0_DSP_top.ConfigBits\[62\]
+ Tile_X0Y0_DSP_top.ConfigBits\[63\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3
+ sky130_fd_sc_hd__mux4_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[262\] Tile_X0Y0_DSP_top.ConfigBits\[263\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.E6END_inbuf_2._0_ net207 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[152\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG1 Tile_X0Y0_DSP_top.ConfigBits\[122\]
+ Tile_X0Y0_DSP_top.ConfigBits\[123\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot5
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_inst0
+ net284 net184 net337 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[25\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[26\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[354\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[365\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._58_ net147 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb2
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18 net238 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[50\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29 net250 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[61\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1690_ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ Tile_X0Y1_DSP_bot.Inst_MULADD._0634_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0636_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0838_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_82_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._60_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG6 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.EE4END_inbuf_9._0_ net37 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1124_ Tile_X0Y1_DSP_bot.Inst_MULADD._0040_ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0296_ sky130_fd_sc_hd__and4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[374\] Tile_X0Y1_DSP_bot.ConfigBits\[375\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1055_ Tile_X0Y1_DSP_bot.Inst_MULADD._0146_ Tile_X0Y1_DSP_bot.Inst_MULADD._0194_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0198_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0228_
+ sky130_fd_sc_hd__a21o_1
Xinput270 Tile_X0Y1_FrameStrobe[18] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__clkbuf_1
Xinput281 Tile_X0Y1_N1END[0] VGND VGND VPWR VPWR net281 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
Xinput292 Tile_X0Y1_N2END[7] VGND VGND VPWR VPWR net292 sky130_fd_sc_hd__buf_2
XFILLER_0_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0908_ Tile_X0Y1_DSP_bot.Inst_MULADD._0082_ Tile_X0Y1_DSP_bot.Inst_MULADD._0083_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0084_ sky130_fd_sc_hd__or2b_1
XFILLER_0_128_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8 net259 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[72\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[302\] Tile_X0Y0_DSP_top.ConfigBits\[303\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput711 net711 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput700 net700 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput733 net733 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput722 net722 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput744 net744 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput755 net755 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_W1BEG1 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[92\] Tile_X0Y1_DSP_bot.ConfigBits\[93\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.N4BEG_outbuf_8._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4END\[8\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[316\] Tile_X0Y0_DSP_top.ConfigBits\[317\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_B2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[130\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[131\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B2 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_C3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[140\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[141\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C3 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_A1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[120\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[121\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A1 sky130_fd_sc_hd__mux4_2
XFILLER_0_146_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[262\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[273\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_138_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot13 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG1 Tile_X0Y0_DSP_top.ConfigBits\[138\]
+ Tile_X0Y0_DSP_top.ConfigBits\[139\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot13
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[215\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_143_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1742_ net333 Tile_X0Y1_DSP_bot.C0 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_129_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_377_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR net751
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[284\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[285\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1673_ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ Tile_X0Y1_DSP_bot.Inst_MULADD._0058_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0001_ sky130_fd_sc_hd__nor2_1
XFILLER_0_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._43_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID5 sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[29\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1107_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B2
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0279_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1038_ Tile_X0Y1_DSP_bot.B5 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0211_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.strobe_outbuf_19._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[19\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[19\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[385\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[396\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.W6BEG_outbuf_8._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_14_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28 net249 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[92\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17 net237 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[81\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput530 net530 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput563 net563 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput552 net552 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput541 net541 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput574 net574 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput585 net585 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput596 net596 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_300_ Tile_X0Y1_DSP_bot.S4BEG\[0\] VGND VGND VPWR VPWR net683 sky130_fd_sc_hd__clkbuf_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_154_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_231_ Tile_X0Y1_DSP_bot.E6BEG\[11\] VGND VGND VPWR VPWR net605 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_162_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG6 VGND VGND VPWR VPWR net545
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.N4END_inbuf_6._0_ Tile_X0Y0_DSP_top.N4END\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_093_ Tile_X0Y0_DSP_top.FrameStrobe_O\[13\] VGND VGND VPWR VPWR net466 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[338\] Tile_X0Y1_DSP_bot.ConfigBits\[339\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 sky130_fd_sc_hd__mux4_2
XFILLER_0_157_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_161 Tile_X0Y0_DSP_top.FrameStrobe\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_150 net291 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_194 Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_183 Tile_X0Y0_DSP_top.W6BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1725_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0019_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1656_ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.ConfigBits\[4\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0810_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0816_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_125_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1587_ Tile_X0Y1_DSP_bot.Inst_MULADD._0748_ Tile_X0Y1_DSP_bot.Inst_MULADD._0749_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0751_ sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot.NN4END_inbuf_1._0_ net328 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._26_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[304\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[293\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst0
+ net183 net336 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.ConfigBits\[114\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[115\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
Xinput1 Tile_X0Y0_E1END[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.N4BEG_outbuf_4._0_ Tile_X0Y0_DSP_top.N4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[4\] sky130_fd_sc_hd__clkbuf_2
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.NN4BEG_outbuf_8._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG2 net17
+ net97 net149 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6 Tile_X0Y0_DSP_top.ConfigBits\[178\]
+ Tile_X0Y0_DSP_top.ConfigBits\[179\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG2
+ sky130_fd_sc_hd__mux4_2
Xoutput393 net393 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput382 net382 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[0] sky130_fd_sc_hd__buf_2
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5 net256 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[133\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_127_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[314\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.data_outbuf_28._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[28\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[28\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1510_ Tile_X0Y1_DSP_bot.Inst_MULADD._0642_ Tile_X0Y1_DSP_bot.Inst_MULADD._0676_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0677_ sky130_fd_sc_hd__nand2_2
XFILLER_0_25_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_214_ Tile_X0Y1_DSP_bot.E2BEGb\[2\] VGND VGND VPWR VPWR net597 sky130_fd_sc_hd__clkbuf_1
X_145_ Tile_X0Y0_DSP_top.NN4BEG\[9\] VGND VGND VPWR VPWR net533 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1441_ Tile_X0Y1_DSP_bot.Inst_MULADD._0605_ Tile_X0Y1_DSP_bot.Inst_MULADD._0533_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0603_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0609_
+ sky130_fd_sc_hd__a21oi_2
X_076_ Tile_X0Y0_DSP_top.FrameData_O\[28\] VGND VGND VPWR VPWR net450 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1372_ Tile_X0Y1_DSP_bot.Inst_MULADD._0448_ Tile_X0Y1_DSP_bot.Inst_MULADD._0449_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0445_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0541_
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot.N4END_inbuf_6._0_ net302 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_1._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END1 sky130_fd_sc_hd__buf_1
XFILLER_0_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[201\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame6_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.data_outbuf_19._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[19\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[19\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1708_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0002_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_4._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1639_ Tile_X0Y1_DSP_bot.C17 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[17\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0800_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot.S4BEG_outbuf_8._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.W6BEG_outbuf_4._0_ Tile_X0Y0_DSP_top.W6BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[4\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._09_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot5
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B5 sky130_fd_sc_hd__buf_2
XFILLER_0_138_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_50 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_61 Tile_X0Y0_DSP_top.N4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 Tile_X0Y0_DSP_top.S4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 Tile_X0Y1_DSP_bot.E6BEG_i\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_94 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0941_ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0109_ Tile_X0Y1_DSP_bot.Inst_MULADD._0114_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0116_ sky130_fd_sc_hd__a22o_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[324\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0872_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.Inst_MULADD._0038_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0039_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0049_
+ sky130_fd_sc_hd__o21a_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[335\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_150_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[21\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[10\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_128_ Tile_X0Y0_DSP_top.N4BEG\[8\] VGND VGND VPWR VPWR net516 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1424_ Tile_X0Y1_DSP_bot.Inst_MULADD._0573_ Tile_X0Y1_DSP_bot.Inst_MULADD._0591_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_059_ Tile_X0Y0_DSP_top.FrameData_O\[11\] VGND VGND VPWR VPWR net432 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1355_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0524_ sky130_fd_sc_hd__nand4_2
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1286_ Tile_X0Y1_DSP_bot.Inst_MULADD._0359_ Tile_X0Y1_DSP_bot.Inst_MULADD._0439_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0440_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0456_
+ sky130_fd_sc_hd__o21ai_2
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput81 Tile_X0Y0_S1END[0] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_4
Xinput70 Tile_X0Y0_FrameData[29] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_6
XFILLER_0_141_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput92 Tile_X0Y0_S2END[7] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_S4BEG1 net21 net88
+ net109 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.ConfigBits\[66\]
+ Tile_X0Y0_DSP_top.ConfigBits\[67\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb1 Tile_X0Y0_DSP_top.S4BEG\[1\]
+ net339 net357 Tile_X0Y1_DSP_bot.ConfigBits\[352\] Tile_X0Y1_DSP_bot.ConfigBits\[353\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_inbuf_3._0_ net254 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[47\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG\[15\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8 net259 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[232\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.data_outbuf_24._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[24\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[24\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[338\] Tile_X0Y0_DSP_top.ConfigBits\[339\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_109_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[232\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[243\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1140_ Tile_X0Y1_DSP_bot.Inst_MULADD._0310_ Tile_X0Y1_DSP_bot.Inst_MULADD._0311_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0312_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1071_ Tile_X0Y1_DSP_bot.Inst_MULADD._0240_ Tile_X0Y1_DSP_bot.Inst_MULADD._0241_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0243_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0244_
+ sky130_fd_sc_hd__a21boi_1
XFILLER_0_89_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0924_ Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ Tile_X0Y1_DSP_bot.Inst_MULADD._0097_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0098_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0099_
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0855_ Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top.data_outbuf_15._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[15\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1407_ Tile_X0Y1_DSP_bot.Inst_MULADD._0494_ Tile_X0Y1_DSP_bot.Inst_MULADD._0520_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0574_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0576_
+ sky130_fd_sc_hd__and3_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.S4BEG_outbuf_4._0_ Tile_X0Y0_DSP_top.S4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1338_ Tile_X0Y1_DSP_bot.Inst_MULADD._0420_ Tile_X0Y1_DSP_bot.Inst_MULADD._0507_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0424_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0508_
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y0_DSP_top.WW4END_inbuf_11._0_ net171 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1269_ Tile_X0Y1_DSP_bot.Inst_MULADD._0265_ Tile_X0Y1_DSP_bot.Inst_MULADD._0267_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_ Tile_X0Y1_DSP_bot.Inst_MULADD._0070_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0439_ sky130_fd_sc_hd__o211ai_4
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[264\] Tile_X0Y0_DSP_top.ConfigBits\[265\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 sky130_fd_sc_hd__mux4_2
XFILLER_0_158_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst0
+ net288 net310 net182 net188 Tile_X0Y1_DSP_bot.ConfigBits\[264\] Tile_X0Y1_DSP_bot.ConfigBits\[265\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_114_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG2 Tile_X0Y0_DSP_top.ConfigBits\[124\]
+ Tile_X0Y0_DSP_top.ConfigBits\[125\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot6
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[25\] Tile_X0Y1_DSP_bot.ConfigBits\[26\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[366\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[355\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[52\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._57_ net146 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb1
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19 net239 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[51\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_86_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG0 net310
+ net213 Tile_X0Y0_DSP_top.S4BEG\[3\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG4
+ Tile_X0Y1_DSP_bot.ConfigBits\[408\] Tile_X0Y1_DSP_bot.ConfigBits\[409\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_156_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_inst0
+ net282 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 net335 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.ConfigBits\[107\] Tile_X0Y1_DSP_bot.ConfigBits\[108\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 net4 net84 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[39\] Tile_X0Y0_DSP_top.ConfigBits\[40\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1123_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0295_ sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1054_ Tile_X0Y1_DSP_bot.Inst_MULADD._0197_ Tile_X0Y1_DSP_bot.Inst_MULADD._0193_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0195_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0227_
+ sky130_fd_sc_hd__and3_1
Xinput271 Tile_X0Y1_FrameStrobe[19] VGND VGND VPWR VPWR net271 sky130_fd_sc_hd__clkbuf_1
Xinput260 Tile_X0Y1_FrameData[9] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__buf_6
Xinput293 Tile_X0Y1_N2MID[0] VGND VGND VPWR VPWR net293 sky130_fd_sc_hd__clkbuf_4
Xinput282 Tile_X0Y1_N1END[1] VGND VGND VPWR VPWR net282 sky130_fd_sc_hd__buf_4
XFILLER_0_58_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0907_ Tile_X0Y1_DSP_bot.Inst_MULADD._0077_ Tile_X0Y1_DSP_bot.Inst_MULADD._0081_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0052_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0083_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9 net260 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[73\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[302\] Tile_X0Y0_DSP_top.ConfigBits\[303\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput712 net712 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput701 net701 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput734 net734 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput723 net723 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput745 net745 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput756 net756 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_W1BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[94\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[95\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_B3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[132\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[133\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B3 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_A2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[122\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[123\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A2 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_C4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[142\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[143\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C4 sky130_fd_sc_hd__mux4_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[274\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[263\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_91_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot14 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG2 Tile_X0Y0_DSP_top.ConfigBits\[140\]
+ Tile_X0Y0_DSP_top.ConfigBits\[141\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot14
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END7
+ net12 net92 net165 Tile_X0Y0_DSP_top.ConfigBits\[238\] Tile_X0Y0_DSP_top.ConfigBits\[239\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.W6END_inbuf_0._0_ net157 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[53\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG\[15\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_99_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[216\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1741_ net333 Tile_X0Y1_DSP_bot.B7 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_376_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net750
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[286\] Tile_X0Y1_DSP_bot.ConfigBits\[287\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG7 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1672_ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ Tile_X0Y1_DSP_bot.Inst_MULADD._0034_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0035_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0000_
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_82_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._42_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG4
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID4 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[30\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1106_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\] Tile_X0Y1_DSP_bot.Inst_MULADD._0047_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0278_ sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1037_ Tile_X0Y1_DSP_bot.Inst_MULADD._0205_ Tile_X0Y1_DSP_bot.Inst_MULADD._0206_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0209_ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0210_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[397\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[386\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_4._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0 net229 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[352\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput520 net520 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29 net250 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[93\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18 net238 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[82\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput531 net531 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput553 net553 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[6] sky130_fd_sc_hd__clkbuf_4
Xoutput542 net542 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput564 net564 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput575 net575 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput586 net586 VGND VGND VPWR VPWR Tile_X0Y1_E1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput597 net597 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[2] sky130_fd_sc_hd__buf_2
XFILLER_0_139_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_230_ Tile_X0Y1_DSP_bot.E6BEG\[10\] VGND VGND VPWR VPWR net604 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_161_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG5 VGND VGND VPWR VPWR net544
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_092_ Tile_X0Y0_DSP_top.FrameStrobe_O\[12\] VGND VGND VPWR VPWR net465 sky130_fd_sc_hd__buf_1
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.W6END_inbuf_0._0_ net358 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_140 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 net291 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 Tile_X0Y0_DSP_top.WW4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 Tile_X0Y0_DSP_top.FrameStrobe\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_inst0
+ net284 net184 net337 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[81\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[82\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XANTENNA_173 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG0 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_195 Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1724_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0018_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_359_ Tile_X0Y1_DSP_bot.W6BEG\[7\] VGND VGND VPWR VPWR net744 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1655_ Tile_X0Y1_DSP_bot.Inst_MULADD._0811_ Tile_X0Y1_DSP_bot.Inst_MULADD._0812_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0813_ Tile_X0Y1_DSP_bot.Inst_MULADD._0814_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0815_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_102_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1586_ Tile_X0Y1_DSP_bot.Inst_MULADD._0748_ Tile_X0Y1_DSP_bot.Inst_MULADD._0749_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0750_ sky130_fd_sc_hd__and2_1
XFILLER_0_113_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._25_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[305\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[294\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_121_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.ConfigBits\[114\] Tile_X0Y1_DSP_bot.ConfigBits\[115\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
Xinput2 Tile_X0Y0_E1END[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_127_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.S4END_inbuf_9._0_ net105 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[9\]
+ sky130_fd_sc_hd__buf_1
XFILLER_0_156_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_GHa_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID0
+ net13 net145 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 Tile_X0Y0_DSP_top.ConfigBits\[180\]
+ Tile_X0Y0_DSP_top.ConfigBits\[181\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput394 net394 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput383 net383 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[1] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.WW4END_inbuf_2._0_ net378 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6 net257 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[134\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[315\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_213_ Tile_X0Y1_DSP_bot.E2BEGb\[1\] VGND VGND VPWR VPWR net596 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_144_ Tile_X0Y0_DSP_top.NN4BEG\[8\] VGND VGND VPWR VPWR net532 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1440_ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_ Tile_X0Y1_DSP_bot.Inst_MULADD._0439_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0533_ Tile_X0Y1_DSP_bot.Inst_MULADD._0603_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0608_ sky130_fd_sc_hd__o211a_1
XTile_X0Y1_DSP_bot.strobe_inbuf_9._0_ net280 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
X_075_ Tile_X0Y0_DSP_top.FrameData_O\[27\] VGND VGND VPWR VPWR net449 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1371_ Tile_X0Y1_DSP_bot.Inst_MULADD._0448_ Tile_X0Y1_DSP_bot.Inst_MULADD._0449_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0540_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[94\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1707_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0001_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_113_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1638_ Tile_X0Y1_DSP_bot.Inst_MULADD._0795_ Tile_X0Y1_DSP_bot.Inst_MULADD._0790_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0799_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1569_ Tile_X0Y1_DSP_bot.Inst_MULADD._0702_ Tile_X0Y1_DSP_bot.Inst_MULADD._0707_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0730_ Tile_X0Y1_DSP_bot.Inst_MULADD._0732_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0734_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._08_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.B4 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.N4END_inbuf_10._0_ Tile_X0Y0_DSP_top.N4END\[14\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_40 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_62 Tile_X0Y0_DSP_top.N4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 Tile_X0Y0_DSP_top.S4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.S4END_inbuf_9._0_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG1
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.S4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_84 Tile_X0Y1_DSP_bot.E6BEG_i\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_95 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_104_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0940_ Tile_X0Y1_DSP_bot.Inst_MULADD._0064_ Tile_X0Y1_DSP_bot.Inst_MULADD._0065_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ Tile_X0Y1_DSP_bot.Inst_MULADD._0109_ Tile_X0Y1_DSP_bot.Inst_MULADD._0114_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0115_ sky130_fd_sc_hd__o2111ai_4
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[325\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0871_ Tile_X0Y1_DSP_bot.Inst_MULADD._0047_ Tile_X0Y1_DSP_bot.B0
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0030_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0048_
+ sky130_fd_sc_hd__a21boi_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[336\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[0\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[11\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_127_ Tile_X0Y0_DSP_top.N4BEG\[7\] VGND VGND VPWR VPWR net515 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1423_ Tile_X0Y1_DSP_bot.Inst_MULADD._0572_ Tile_X0Y1_DSP_bot.Inst_MULADD._0590_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0494_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0591_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_159_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_058_ Tile_X0Y0_DSP_top.FrameData_O\[10\] VGND VGND VPWR VPWR net431 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1354_ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_ Tile_X0Y1_DSP_bot.Inst_MULADD._0188_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0273_ Tile_X0Y1_DSP_bot.Inst_MULADD._0154_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0523_ sky130_fd_sc_hd__o2bb2ai_4
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1285_ Tile_X0Y1_DSP_bot.Inst_MULADD._0442_ Tile_X0Y1_DSP_bot.Inst_MULADD._0444_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0455_ sky130_fd_sc_hd__nand2_4
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.SS4END_inbuf_10._0_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG2
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput82 Tile_X0Y0_S1END[1] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__clkbuf_4
Xinput71 Tile_X0Y0_FrameData[2] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_8
Xinput60 Tile_X0Y0_FrameData[1] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_8
Xinput93 Tile_X0Y0_S2MID[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_S4BEG2 net85 net110
+ net156 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.ConfigBits\[68\]
+ Tile_X0Y0_DSP_top.ConfigBits\[69\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst2
+ net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[352\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[353\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.data_inbuf_20._0_ net61 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[20\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[47\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9 net260 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[233\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[338\] Tile_X0Y0_DSP_top.ConfigBits\[339\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END2 net7 Tile_X0Y0_DSP_top.ConfigBits\[282\]
+ Tile_X0Y0_DSP_top.ConfigBits\[283\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.strobe_inbuf_5._0_ Tile_X0Y0_DSP_top.FrameStrobe\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[233\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1070_ Tile_X0Y1_DSP_bot.Inst_MULADD._0242_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[5\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0243_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.data_inbuf_11._0_ net51 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[118\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_97_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0923_ Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0098_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0854_ Tile_X0Y1_DSP_bot.Inst_MULADD._0030_ Tile_X0Y1_DSP_bot.Inst_MULADD._0031_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ sky130_fd_sc_hd__nand2_8
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END3
+ net8 net140 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.ConfigBits\[390\]
+ Tile_X0Y0_DSP_top.ConfigBits\[391\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[100\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG0 sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1406_ Tile_X0Y1_DSP_bot.Inst_MULADD._0494_ Tile_X0Y1_DSP_bot.Inst_MULADD._0520_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0574_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0575_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1337_ Tile_X0Y1_DSP_bot.Inst_MULADD._0319_ Tile_X0Y1_DSP_bot.Inst_MULADD._0506_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0342_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0507_
+ sky130_fd_sc_hd__a21o_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1268_ Tile_X0Y1_DSP_bot.Inst_MULADD._0359_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0438_ sky130_fd_sc_hd__buf_4
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1199_ Tile_X0Y1_DSP_bot.Inst_MULADD._0070_ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0358_ Tile_X0Y1_DSP_bot.Inst_MULADD._0360_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0370_ sky130_fd_sc_hd__a22o_2
XFILLER_0_88_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst1
+ net204 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb3 net341 net373 Tile_X0Y1_DSP_bot.ConfigBits\[264\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[265\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_146_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG3 Tile_X0Y0_DSP_top.ConfigBits\[126\]
+ Tile_X0Y0_DSP_top.ConfigBits\[127\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot7
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[367\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[356\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[53\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[42\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._56_ net145 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb0
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG1 net309
+ Tile_X0Y0_DSP_top.SS4BEG\[2\] net340 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG4
+ Tile_X0Y1_DSP_bot.ConfigBits\[410\] Tile_X0Y1_DSP_bot.ConfigBits\[411\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.SS4END_inbuf_4._0_ Tile_X0Y0_DSP_top.SS4BEG\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[4\] sky130_fd_sc_hd__buf_2
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.data_inbuf_20._0_ net241 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[20\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[107\] Tile_X0Y1_DSP_bot.ConfigBits\[108\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG0
+ Tile_X0Y0_DSP_top.ConfigBits\[39\] Tile_X0Y0_DSP_top.ConfigBits\[40\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_105_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1122_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ Tile_X0Y1_DSP_bot.B6
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0293_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0294_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_156_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1053_ Tile_X0Y1_DSP_bot.Inst_MULADD._0224_ Tile_X0Y1_DSP_bot.Inst_MULADD._0225_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0157_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0226_
+ sky130_fd_sc_hd__a21o_1
Xinput261 Tile_X0Y1_FrameStrobe[0] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__buf_8
Xinput272 Tile_X0Y1_FrameStrobe[1] VGND VGND VPWR VPWR net272 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput250 Tile_X0Y1_FrameData[29] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__clkbuf_8
Xinput294 Tile_X0Y1_N2MID[1] VGND VGND VPWR VPWR net294 sky130_fd_sc_hd__buf_2
Xinput283 Tile_X0Y1_N1END[2] VGND VGND VPWR VPWR net283 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 net2 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[25\] Tile_X0Y0_DSP_top.ConfigBits\[26\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.data_inbuf_11._0_ net231 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0906_ Tile_X0Y1_DSP_bot.Inst_MULADD._0077_ Tile_X0Y1_DSP_bot.Inst_MULADD._0081_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0052_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0082_
+ sky130_fd_sc_hd__nor3_2
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[304\] Tile_X0Y0_DSP_top.ConfigBits\[305\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG6 sky130_fd_sc_hd__mux4_2
XFILLER_0_41_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput702 net702 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput724 net724 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput713 net713 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput735 net735 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[0] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.S4END_inbuf_10._0_ net106 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[10\]
+ sky130_fd_sc_hd__dlymetal6s2s_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst0
+ net3 net135 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.ConfigBits\[52\] Tile_X0Y0_DSP_top.ConfigBits\[53\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput757 net757 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput746 net746 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[9] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst0
+ net282 net290 net182 net190 Tile_X0Y1_DSP_bot.ConfigBits\[304\] Tile_X0Y1_DSP_bot.ConfigBits\[305\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_W1BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[96\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[97\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_146_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_A3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[124\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[125\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A3 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_C5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[144\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[145\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C5 sky130_fd_sc_hd__mux4_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[264\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.data_outbuf_9._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[9\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[9\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[275\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot15 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG3 Tile_X0Y0_DSP_top.ConfigBits\[142\]
+ Tile_X0Y0_DSP_top.ConfigBits\[143\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot15
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_91_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END3
+ net8 net117 net140 Tile_X0Y0_DSP_top.ConfigBits\[240\] Tile_X0Y0_DSP_top.ConfigBits\[241\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG1 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[53\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.EE4END_inbuf_3._0_ net226 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._39_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[217\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1740_ net333 Tile_X0Y1_DSP_bot.B6 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XTile_X0Y0_DSP_top.strobe_inbuf_12._0_ Tile_X0Y0_DSP_top.FrameStrobe\[12\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_375_ Tile_X0Y1_DSP_bot.WW4BEG\[11\] VGND VGND VPWR VPWR net749 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1671_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._41_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG3
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID3 sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[31\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1105_ Tile_X0Y1_DSP_bot.Inst_MULADD._0264_ Tile_X0Y1_DSP_bot.Inst_MULADD._0268_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0272_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0277_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_92_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1036_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B5
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0208_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0209_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_116_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END4
+ net9 net21 Tile_X0Y0_DSP_top.ConfigBits\[354\] Tile_X0Y0_DSP_top.ConfigBits\[355\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[387\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[398\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[84\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1 net240 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[353\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_73_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput510 net510 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19 net239 net262 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[83\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame10_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput521 net521 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput532 net532 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[8] sky130_fd_sc_hd__buf_2
Xoutput554 net554 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput543 net543 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput565 net565 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput576 net576 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput587 net587 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput598 net598 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.SS4END_inbuf_0._0_ net127 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_160_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG4 VGND VGND VPWR VPWR net543
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.data_outbuf_9._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[9\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[9\] sky130_fd_sc_hd__clkbuf_1
X_091_ Tile_X0Y0_DSP_top.FrameStrobe_O\[11\] VGND VGND VPWR VPWR net464 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.strobe_outbuf_14._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[14\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[14\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_157_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_130 Tile_X0Y1_DSP_bot.SS4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 net291 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_174 Tile_X0Y0_DSP_top.N4BEG\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 Tile_X0Y0_DSP_top.FrameStrobe\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[81\] Tile_X0Y1_DSP_bot.ConfigBits\[82\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XANTENNA_185 Tile_X0Y1_DSP_bot.EE4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1723_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0017_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_358_ Tile_X0Y1_DSP_bot.W6BEG\[6\] VGND VGND VPWR VPWR net743 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.E6BEG_outbuf_7._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1654_ Tile_X0Y1_DSP_bot.Inst_MULADD._0787_ Tile_X0Y1_DSP_bot.Inst_MULADD._0803_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0798_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0814_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_125_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1585_ Tile_X0Y1_DSP_bot.Inst_MULADD._0701_ Tile_X0Y1_DSP_bot.Inst_MULADD._0728_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0730_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0749_
+ sky130_fd_sc_hd__o21ai_1
X_289_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG5 VGND VGND VPWR VPWR net672
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._24_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEG\[2\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[306\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[295\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[114\] Tile_X0Y1_DSP_bot.ConfigBits\[115\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 Tile_X0Y0_E1END[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1019_ Tile_X0Y1_DSP_bot.Inst_MULADD._0191_ Tile_X0Y1_DSP_bot.A5
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0187_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0192_
+ sky130_fd_sc_hd__a21boi_4
XFILLER_0_36_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_143_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.EE4END_inbuf_10._0_ net218 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput395 net395 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput384 net384 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7 net258 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[135\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[316\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_212_ Tile_X0Y1_DSP_bot.E2BEGb\[0\] VGND VGND VPWR VPWR net595 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst0
+ net284 net292 net184 net192 Tile_X0Y1_DSP_bot.ConfigBits\[376\] Tile_X0Y1_DSP_bot.ConfigBits\[377\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_143_ Tile_X0Y0_DSP_top.NN4BEG\[7\] VGND VGND VPWR VPWR net531 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_074_ Tile_X0Y0_DSP_top.FrameData_O\[26\] VGND VGND VPWR VPWR net448 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1370_ Tile_X0Y1_DSP_bot.Inst_MULADD._0455_ Tile_X0Y1_DSP_bot.Inst_MULADD._0454_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0537_ Tile_X0Y1_DSP_bot.Inst_MULADD._0538_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0539_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[94\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.strobe_outbuf_3._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[3\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[3\] sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END3 net2 net8 net24 Tile_X0Y0_DSP_top.ConfigBits\[318\]
+ Tile_X0Y0_DSP_top.ConfigBits\[319\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_7_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1706_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0000_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1637_ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.Inst_MULADD._0789_
+ Tile_X0Y1_DSP_bot.ConfigBits\[4\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0798_
+ sky130_fd_sc_hd__nand3_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1568_ Tile_X0Y1_DSP_bot.Inst_MULADD._0730_ Tile_X0Y1_DSP_bot.Inst_MULADD._0732_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0702_ Tile_X0Y1_DSP_bot.Inst_MULADD._0707_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0733_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_141_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.WW4BEG_outbuf_8._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[8\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1499_ Tile_X0Y1_DSP_bot.Inst_MULADD._0597_ Tile_X0Y1_DSP_bot.Inst_MULADD._0598_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0604_ Tile_X0Y1_DSP_bot.Inst_MULADD._0609_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0666_ sky130_fd_sc_hd__a31oi_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._07_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_138_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.E6END_inbuf_5._0_ net30 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_41 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_30 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG2 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 Tile_X0Y0_DSP_top.N4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_74 Tile_X0Y0_DSP_top.S4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_96 Tile_X0Y1_DSP_bot.N4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 Tile_X0Y1_DSP_bot.EE4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_132_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_1._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_159_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.strobe_inbuf_18._0_ net270 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[18\]
+ sky130_fd_sc_hd__clkbuf_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._0870_ Tile_X0Y1_DSP_bot.ConfigBits\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0047_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[337\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[326\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[12\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[1\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_126_ Tile_X0Y0_DSP_top.N4BEG\[6\] VGND VGND VPWR VPWR net514 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.E6BEG_outbuf_3._0_ Tile_X0Y0_DSP_top.E6BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1422_ Tile_X0Y1_DSP_bot.Inst_MULADD._0588_ Tile_X0Y1_DSP_bot.Inst_MULADD._0589_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0590_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_150_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_123_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_057_ Tile_X0Y0_DSP_top.FrameData_O\[9\] VGND VGND VPWR VPWR net461 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1353_ Tile_X0Y1_DSP_bot.Inst_MULADD._0050_ Tile_X0Y1_DSP_bot.Inst_MULADD._0273_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0522_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_21_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1284_ Tile_X0Y1_DSP_bot.Inst_MULADD._0444_ Tile_X0Y1_DSP_bot.Inst_MULADD._0442_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0451_ Tile_X0Y1_DSP_bot.Inst_MULADD._0453_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0454_ sky130_fd_sc_hd__o211ai_4
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.data_inbuf_0._0_ net49 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._0999_ Tile_X0Y1_DSP_bot.Inst_MULADD._0172_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0173_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_140_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput72 Tile_X0Y0_FrameData[30] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_8
Xinput61 Tile_X0Y0_FrameData[20] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_6
Xinput50 Tile_X0Y0_FrameData[10] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput94 Tile_X0Y0_S2MID[1] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_4
Xinput83 Tile_X0Y0_S1END[2] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_S4BEG3 net86 net101
+ net153 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.ConfigBits\[70\]
+ Tile_X0Y0_DSP_top.ConfigBits\[71\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[352\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[353\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID7
+ net20 net100 net152 Tile_X0Y0_DSP_top.ConfigBits\[190\] Tile_X0Y0_DSP_top.ConfigBits\[191\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.E6END_inbuf_5._0_ net210 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_94_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[340\] Tile_X0Y0_DSP_top.ConfigBits\[341\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7 sky130_fd_sc_hd__mux4_2
XFILLER_0_124_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst1
+ net21 net87 net139 net174 Tile_X0Y0_DSP_top.ConfigBits\[282\] Tile_X0Y0_DSP_top.ConfigBits\[283\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_120_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst0
+ net283 net291 net183 net191 Tile_X0Y1_DSP_bot.ConfigBits\[340\] Tile_X0Y1_DSP_bot.ConfigBits\[341\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_132_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[119\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0922_ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ Tile_X0Y1_DSP_bot.C3
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0096_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0097_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0853_ Tile_X0Y1_DSP_bot.ConfigBits\[1\] Tile_X0Y1_DSP_bot.B0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0031_ sky130_fd_sc_hd__or2b_4
XFILLER_0_57_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END2
+ net7 net109 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG3 Tile_X0Y0_DSP_top.ConfigBits\[392\]
+ Tile_X0Y0_DSP_top.ConfigBits\[393\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[100\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
X_109_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG5 VGND VGND VPWR VPWR net491
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1405_ Tile_X0Y1_DSP_bot.Inst_MULADD._0564_ Tile_X0Y1_DSP_bot.Inst_MULADD._0566_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0573_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0574_
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1336_ Tile_X0Y1_DSP_bot.Inst_MULADD._0410_ Tile_X0Y1_DSP_bot.Inst_MULADD._0505_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0411_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0506_
+ sky130_fd_sc_hd__o21ai_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1267_ Tile_X0Y1_DSP_bot.Inst_MULADD._0395_ Tile_X0Y1_DSP_bot.Inst_MULADD._0398_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0391_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0437_
+ sky130_fd_sc_hd__a21oi_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1198_ Tile_X0Y1_DSP_bot.Inst_MULADD._0271_ Tile_X0Y1_DSP_bot.Inst_MULADD._0363_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0259_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0369_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_135_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[264\] Tile_X0Y1_DSP_bot.ConfigBits\[265\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.SS4BEG_outbuf_1._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[1\] sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG0 Tile_X0Y0_DSP_top.ConfigBits\[128\]
+ Tile_X0Y0_DSP_top.ConfigBits\[129\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot8
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_5_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[368\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[357\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[43\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[32\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._55_ net144 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG7
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG2 net204
+ Tile_X0Y0_DSP_top.S4BEG\[1\] net375 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.ConfigBits\[412\] Tile_X0Y1_DSP_bot.ConfigBits\[413\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_0_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_137_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1121_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[6\] Tile_X0Y1_DSP_bot.Inst_MULADD._0079_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0293_ sky130_fd_sc_hd__or2b_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1052_ Tile_X0Y1_DSP_bot.Inst_MULADD._0164_ Tile_X0Y1_DSP_bot.Inst_MULADD._0163_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0158_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0225_
+ sky130_fd_sc_hd__o21a_1
Xinput262 Tile_X0Y1_FrameStrobe[10] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__buf_8
Xinput240 Tile_X0Y1_FrameData[1] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_8
Xinput251 Tile_X0Y1_FrameData[2] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__buf_6
Xinput295 Tile_X0Y1_N2MID[2] VGND VGND VPWR VPWR net295 sky130_fd_sc_hd__clkbuf_4
Xinput284 Tile_X0Y1_N1END[3] VGND VGND VPWR VPWR net284 sky130_fd_sc_hd__buf_4
Xinput273 Tile_X0Y1_FrameStrobe[2] VGND VGND VPWR VPWR net273 sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._0905_ Tile_X0Y1_DSP_bot.Inst_MULADD._0076_ Tile_X0Y1_DSP_bot.Inst_MULADD._0078_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ Tile_X0Y1_DSP_bot.Inst_MULADD._0080_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0081_ sky130_fd_sc_hd__o2bb2a_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG1
+ Tile_X0Y0_DSP_top.ConfigBits\[25\] Tile_X0Y0_DSP_top.ConfigBits\[26\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput703 net703 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput725 net725 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput714 net714 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput736 net736 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput758 net758 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput747 net747 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[0] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb5 net335 Tile_X0Y1_DSP_bot.ConfigBits\[304\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[305\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[52\] Tile_X0Y0_DSP_top.ConfigBits\[53\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1319_ Tile_X0Y1_DSP_bot.Inst_MULADD._0474_ Tile_X0Y1_DSP_bot.Inst_MULADD._0475_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0461_ Tile_X0Y1_DSP_bot.Inst_MULADD._0467_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0489_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_146_52 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_C6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[146\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[147\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C6 sky130_fd_sc_hd__mux4_2
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[265\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_119_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END1
+ net10 net90 net142 Tile_X0Y0_DSP_top.ConfigBits\[242\] Tile_X0Y0_DSP_top.ConfigBits\[243\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_142_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst3_765
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst3_765/HI
+ net765 sky130_fd_sc_hd__conb_1
XFILLER_0_99_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG3.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._38_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[218\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.N4END_inbuf_9._0_ Tile_X0Y0_DSP_top.N4END\[13\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_374_ Tile_X0Y1_DSP_bot.WW4BEG\[10\] VGND VGND VPWR VPWR net748 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1670_ Tile_X0Y1_DSP_bot.Inst_MULADD._0428_ Tile_X0Y1_DSP_bot.Inst_MULADD._0820_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0828_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q19
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[83\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG3 sky130_fd_sc_hd__o21ai_1
XFILLER_0_133_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._40_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID2 sky130_fd_sc_hd__buf_2
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1104_ Tile_X0Y1_DSP_bot.Inst_MULADD._0259_ Tile_X0Y1_DSP_bot.Inst_MULADD._0272_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0275_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0276_
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1035_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\] Tile_X0Y1_DSP_bot.Inst_MULADD._0047_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0208_ sky130_fd_sc_hd__or2_2
XFILLER_0_92_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst1
+ net89 net101 net141 net153 Tile_X0Y0_DSP_top.ConfigBits\[354\] Tile_X0Y0_DSP_top.ConfigBits\[355\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[388\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[399\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_128_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[74\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[85\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2 net251 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[354\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.NN4END_inbuf_4._0_ net331 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput511 net511 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput500 net500 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput533 net533 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput522 net522 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput544 net544 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput566 net566 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput555 net555 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput577 net577 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput588 net588 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput599 net599 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[4] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.N4BEG_outbuf_7._0_ Tile_X0Y0_DSP_top.N4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[7\] sky130_fd_sc_hd__clkbuf_2
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_090_ Tile_X0Y0_DSP_top.FrameStrobe_O\[10\] VGND VGND VPWR VPWR net463 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG0 net326
+ Tile_X0Y0_DSP_top.S4BEG\[3\] net366 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[384\] Tile_X0Y1_DSP_bot.ConfigBits\[385\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_131 Tile_X0Y1_DSP_bot.SS4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 net140 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_120 Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_175 Tile_X0Y0_DSP_top.NN4BEG\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 Tile_X0Y0_DSP_top.FrameStrobe\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 net310 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_197 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1722_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0016_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_186 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_127_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_357_ Tile_X0Y1_DSP_bot.W6BEG\[5\] VGND VGND VPWR VPWR net742 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1653_ Tile_X0Y1_DSP_bot.Inst_MULADD._0795_ Tile_X0Y1_DSP_bot.Inst_MULADD._0790_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0802_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0813_
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_153_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.N4END_inbuf_9._0_ net305 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_125_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1584_ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_ Tile_X0Y1_DSP_bot.Inst_MULADD._0351_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0748_ sky130_fd_sc_hd__a211o_1
X_288_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG4 VGND VGND VPWR VPWR net671
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END6
+ net3 net11 Tile_X0Y0_DSP_top.ConfigBits\[266\] Tile_X0Y0_DSP_top.ConfigBits\[267\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_4._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4END\[4\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._23_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEG\[1\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[296\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[307\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[114\] Tile_X0Y1_DSP_bot.ConfigBits\[115\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
Xinput4 Tile_X0Y0_E1END[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1018_ Tile_X0Y1_DSP_bot.ConfigBits\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0191_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_7._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.W6BEG_outbuf_7._0_ Tile_X0Y0_DSP_top.W6BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[7\] sky130_fd_sc_hd__clkbuf_2
Xoutput396 net396 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[2] sky130_fd_sc_hd__buf_2
Xoutput385 net385 VGND VGND VPWR VPWR Tile_X0Y0_E1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_77_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 net2 net134 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[81\] Tile_X0Y0_DSP_top.ConfigBits\[82\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.S4BEG_outbuf_11._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[11\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END6
+ net11 net126 net143 Tile_X0Y0_DSP_top.ConfigBits\[214\] Tile_X0Y0_DSP_top.ConfigBits\[215\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8 net259 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[136\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[317\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_211_ Tile_X0Y1_DSP_bot.E2BEG\[7\] VGND VGND VPWR VPWR net594 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb7 net337 Tile_X0Y1_DSP_bot.ConfigBits\[376\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[377\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
X_142_ Tile_X0Y0_DSP_top.NN4BEG\[6\] VGND VGND VPWR VPWR net530 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_073_ Tile_X0Y0_DSP_top.FrameData_O\[25\] VGND VGND VPWR VPWR net447 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[89\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 sky130_fd_sc_hd__o21ai_2
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst1
+ net88 net110 net140 net156 Tile_X0Y0_DSP_top.ConfigBits\[318\] Tile_X0Y0_DSP_top.ConfigBits\[319\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1705_ Tile_X0Y1_DSP_bot.Inst_MULADD._0825_ Tile_X0Y1_DSP_bot.Inst_MULADD._0827_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0019_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1636_ Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0796_ Tile_X0Y1_DSP_bot.Inst_MULADD._0797_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q16 sky130_fd_sc_hd__a22o_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1567_ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0697_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_ Tile_X0Y1_DSP_bot.Inst_MULADD._0731_ Tile_X0Y1_DSP_bot.Inst_MULADD._0729_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0732_ sky130_fd_sc_hd__a311o_1
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.NN4END_inbuf_0._0_ Tile_X0Y0_DSP_top.NN4END\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1498_ Tile_X0Y1_DSP_bot.Inst_MULADD._0657_ Tile_X0Y1_DSP_bot.Inst_MULADD._0658_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0660_ Tile_X0Y1_DSP_bot.Inst_MULADD._0661_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0665_ sky130_fd_sc_hd__a22oi_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._06_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot2
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A6 sky130_fd_sc_hd__buf_2
XFILLER_0_138_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_154_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID6
+ net99 net151 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3 Tile_X0Y0_DSP_top.ConfigBits\[150\]
+ Tile_X0Y0_DSP_top.ConfigBits\[151\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_129_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_31 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG2 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 Tile_X0Y0_DSP_top.FrameStrobe\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 Tile_X0Y0_DSP_top.NN4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 Tile_X0Y0_DSP_top.S4BEG_i\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top.EE4BEG_outbuf_1._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[1\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_42 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_6_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_53 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_97 Tile_X0Y1_DSP_bot.NN4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_86 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.data_inbuf_6._0_ net257 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.data_outbuf_27._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[27\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[27\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[338\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[327\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[13\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[2\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_125_ Tile_X0Y0_DSP_top.N4BEG\[5\] VGND VGND VPWR VPWR net513 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1421_ Tile_X0Y1_DSP_bot.Inst_MULADD._0563_ Tile_X0Y1_DSP_bot.Inst_MULADD._0557_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0562_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0589_
+ sky130_fd_sc_hd__nand3b_1
X_056_ Tile_X0Y0_DSP_top.FrameData_O\[8\] VGND VGND VPWR VPWR net460 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1352_ Tile_X0Y1_DSP_bot.Inst_MULADD._0357_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0521_ sky130_fd_sc_hd__buf_4
XFILLER_0_150_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1283_ Tile_X0Y1_DSP_bot.Inst_MULADD._0196_ Tile_X0Y1_DSP_bot.Inst_MULADD._0107_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_ Tile_X0Y1_DSP_bot.Inst_MULADD._0450_ Tile_X0Y1_DSP_bot.Inst_MULADD._0452_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0453_ sky130_fd_sc_hd__a32o_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.data_outbuf_18._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[18\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[18\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0998_ Tile_X0Y1_DSP_bot.C4 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[4\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0172_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput40 Tile_X0Y0_EE4END[1] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1619_ Tile_X0Y1_DSP_bot.Inst_MULADD._0764_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0782_ sky130_fd_sc_hd__inv_2
Xinput73 Tile_X0Y0_FrameData[31] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_8
Xinput62 Tile_X0Y0_FrameData[21] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_6
Xinput51 Tile_X0Y0_FrameData[11] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_8
XTile_X0Y0_DSP_top.S4BEG_outbuf_7._0_ Tile_X0Y0_DSP_top.S4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[7\] sky130_fd_sc_hd__clkbuf_1
Xinput95 Tile_X0Y0_S2MID[2] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_4
Xinput84 Tile_X0Y0_S1END[3] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[354\] Tile_X0Y1_DSP_bot.ConfigBits\[355\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG0 sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID3
+ net16 net96 net148 Tile_X0Y0_DSP_top.ConfigBits\[192\] Tile_X0Y0_DSP_top.ConfigBits\[193\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_94_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[282\] Tile_X0Y0_DSP_top.ConfigBits\[283\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_62_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb6
+ net334 net336 Tile_X0Y1_DSP_bot.ConfigBits\[340\] Tile_X0Y1_DSP_bot.ConfigBits\[341\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_120_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[120\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0921_ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[3\] Tile_X0Y1_DSP_bot.Inst_MULADD._0086_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0096_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._0852_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\] Tile_X0Y1_DSP_bot.ConfigBits\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0030_ sky130_fd_sc_hd__nand2_4
XFILLER_0_155_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_123_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END1
+ net124 net141 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 Tile_X0Y0_DSP_top.ConfigBits\[394\]
+ Tile_X0Y0_DSP_top.ConfigBits\[395\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_53_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_108_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG4 VGND VGND VPWR VPWR net490
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1404_ Tile_X0Y1_DSP_bot.Inst_MULADD._0564_ Tile_X0Y1_DSP_bot.Inst_MULADD._0571_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0572_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0573_
+ sky130_fd_sc_hd__o21ai_4
X_039_ Tile_X0Y0_DSP_top.EE4BEG\[7\] VGND VGND VPWR VPWR net427 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1335_ Tile_X0Y1_DSP_bot.Inst_MULADD._0307_ Tile_X0Y1_DSP_bot.Inst_MULADD._0413_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0415_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0505_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1266_ Tile_X0Y1_DSP_bot.Inst_MULADD._0431_ Tile_X0Y1_DSP_bot.Inst_MULADD._0409_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0430_ Tile_X0Y1_DSP_bot.Inst_MULADD._0429_ Tile_X0Y1_DSP_bot.Inst_MULADD._0401_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0436_ sky130_fd_sc_hd__o32ai_4
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1197_ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0357_ Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0368_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_28_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.ConfigBits\[264\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[265\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_158_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0 net229 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[256\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_top2bot9 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG1 Tile_X0Y0_DSP_top.ConfigBits\[130\]
+ Tile_X0Y0_DSP_top.ConfigBits\[131\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot9
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[369\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[358\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[44\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[33\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._54_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG6 sky130_fd_sc_hd__clkbuf_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG3 net317
+ net201 net338 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG4 Tile_X0Y1_DSP_bot.ConfigBits\[414\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[415\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_145_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.W6END_inbuf_3._0_ net160 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1120_ Tile_X0Y1_DSP_bot.Inst_MULADD._0199_ Tile_X0Y1_DSP_bot.Inst_MULADD._0235_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0291_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0292_
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1051_ Tile_X0Y1_DSP_bot.Inst_MULADD._0199_ Tile_X0Y1_DSP_bot.Inst_MULADD._0217_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0221_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0224_
+ sky130_fd_sc_hd__o21ai_2
Xinput263 Tile_X0Y1_FrameStrobe[11] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__buf_8
Xinput241 Tile_X0Y1_FrameData[20] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_8
Xinput230 Tile_X0Y1_FrameData[10] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__buf_6
Xinput252 Tile_X0Y1_FrameData[30] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__buf_6
Xinput285 Tile_X0Y1_N2END[0] VGND VGND VPWR VPWR net285 sky130_fd_sc_hd__buf_2
Xinput296 Tile_X0Y1_N2MID[3] VGND VGND VPWR VPWR net296 sky130_fd_sc_hd__clkbuf_4
Xinput274 Tile_X0Y1_FrameStrobe[3] VGND VGND VPWR VPWR net274 sky130_fd_sc_hd__clkbuf_16
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst0
+ net299 net193 net199 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[156\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[157\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_81_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0904_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ Tile_X0Y1_DSP_bot.Inst_MULADD._0068_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0069_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0080_
+ sky130_fd_sc_hd__o21a_2
XFILLER_0_85_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput726 net726 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput715 net715 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput704 net704 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_111_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput759 net759 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput748 net748 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput737 net737 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[11] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[304\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[305\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[52\] Tile_X0Y0_DSP_top.ConfigBits\[53\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1318_ Tile_X0Y1_DSP_bot.Inst_MULADD._0487_ Tile_X0Y1_DSP_bot.Inst_MULADD._0466_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0476_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0488_
+ sky130_fd_sc_hd__a21o_2
XFILLER_0_39_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1249_ Tile_X0Y1_DSP_bot.Inst_MULADD._0417_ Tile_X0Y1_DSP_bot.Inst_MULADD._0419_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0342_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0420_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_C7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[148\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[149\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C7 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG6
+ Tile_X0Y0_DSP_top.ConfigBits\[144\] Tile_X0Y0_DSP_top.ConfigBits\[145\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_7._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_GH_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END1
+ net42 net86 net138 Tile_X0Y0_DSP_top.ConfigBits\[244\] Tile_X0Y0_DSP_top.ConfigBits\[245\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_32_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst3_766
+ VGND VGND VPWR VPWR net766 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst3_766/LO
+ sky130_fd_sc_hd__conb_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._37_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG5 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[219\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_373_ Tile_X0Y1_DSP_bot.WW4BEG\[9\] VGND VGND VPWR VPWR net762 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[83\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_137_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.W6END_inbuf_3._0_ net361 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0274_ Tile_X0Y1_DSP_bot.Inst_MULADD._0259_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0275_ sky130_fd_sc_hd__a22oi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1034_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[354\] Tile_X0Y0_DSP_top.ConfigBits\[355\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_148_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[389\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[400\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10 net50 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[64\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21 net62 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[75\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3 net254 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[355\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG0 net300
+ net200 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG7 net353 Tile_X0Y1_DSP_bot.ConfigBits\[208\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[209\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput501 net501 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput534 net534 VGND VGND VPWR VPWR Tile_X0Y0_UserCLKo sky130_fd_sc_hd__buf_2
Xoutput523 net523 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput512 net512 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput545 net545 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput556 net556 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput578 net578 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput567 net567 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput589 net589 VGND VGND VPWR VPWR Tile_X0Y1_E2BEG[2] sky130_fd_sc_hd__buf_2
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG1 net221
+ Tile_X0Y0_DSP_top.S4BEG\[2\] net345 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[386\] Tile_X0Y1_DSP_bot.ConfigBits\[387\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG1 sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[54\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.WW4END_inbuf_5._0_ net381 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_143 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 Tile_X0Y1_DSP_bot.SS4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_110 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 Tile_X0Y0_DSP_top.FrameStrobe\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 Tile_X0Y0_DSP_top.S4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 net310 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_198 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1721_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0015_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\] sky130_fd_sc_hd__dfxtp_1
X_356_ Tile_X0Y1_DSP_bot.W6BEG\[4\] VGND VGND VPWR VPWR net741 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1652_ Tile_X0Y1_DSP_bot.Inst_MULADD._0809_ Tile_X0Y1_DSP_bot.Inst_MULADD._0787_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0812_ sky130_fd_sc_hd__or2_1
XFILLER_0_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_113_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1583_ Tile_X0Y1_DSP_bot.Inst_MULADD._0747_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q13 sky130_fd_sc_hd__buf_1
X_287_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG3 VGND VGND VPWR VPWR net670
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst1
+ net83 net91 net133 net135 Tile_X0Y0_DSP_top.ConfigBits\[266\] Tile_X0Y0_DSP_top.ConfigBits\[267\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_140_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._22_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEG\[0\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[297\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_W6BEG1.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[116\] Tile_X0Y1_DSP_bot.ConfigBits\[117\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W6BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_127_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput5 Tile_X0Y0_E2END[0] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1017_ Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0141_ Tile_X0Y1_DSP_bot.Inst_MULADD._0188_ Tile_X0Y1_DSP_bot.Inst_MULADD._0189_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0190_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput386 net386 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput397 net397 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG3
+ Tile_X0Y0_DSP_top.ConfigBits\[81\] Tile_X0Y0_DSP_top.ConfigBits\[82\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END0
+ net7 net87 net139 Tile_X0Y0_DSP_top.ConfigBits\[216\] Tile_X0Y0_DSP_top.ConfigBits\[217\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG1 sky130_fd_sc_hd__mux4_2
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9 net260 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[137\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[318\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_210_ Tile_X0Y1_DSP_bot.E2BEG\[6\] VGND VGND VPWR VPWR net593 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[376\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[377\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
X_141_ Tile_X0Y0_DSP_top.NN4BEG\[5\] VGND VGND VPWR VPWR net529 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_072_ Tile_X0Y0_DSP_top.FrameData_O\[24\] VGND VGND VPWR VPWR net446 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END0
+ net1 net5 Tile_X0Y0_DSP_top.ConfigBits\[306\] Tile_X0Y0_DSP_top.ConfigBits\[307\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[89\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[318\] Tile_X0Y0_DSP_top.ConfigBits\[319\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1704_ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ Tile_X0Y1_DSP_bot.Inst_MULADD._0020_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0815_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0018_
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_83_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_339_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG3 VGND VGND VPWR VPWR net722
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1635_ Tile_X0Y1_DSP_bot.Inst_MULADD._0795_ Tile_X0Y1_DSP_bot.Inst_MULADD._0790_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0797_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1566_ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_ Tile_X0Y1_DSP_bot.Inst_MULADD._0660_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.NN4END_inbuf_10._0_ net322 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_51_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._05_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot1
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A5 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1497_ Tile_X0Y1_DSP_bot.Inst_MULADD._0644_ Tile_X0Y1_DSP_bot.Inst_MULADD._0645_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0657_ Tile_X0Y1_DSP_bot.Inst_MULADD._0658_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0664_ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG1 net15
+ net95 net147 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG3 Tile_X0Y0_DSP_top.ConfigBits\[152\]
+ Tile_X0Y0_DSP_top.ConfigBits\[153\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_19_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_21 Tile_X0Y0_DSP_top.FrameStrobe\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 Tile_X0Y0_DSP_top.FrameStrobe\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_32 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_65 Tile_X0Y0_DSP_top.NN4BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_54 Tile_X0Y0_DSP_top.N4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_76 Tile_X0Y0_DSP_top.S4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 Tile_X0Y1_DSP_bot.NN4BEG_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_112_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_10._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG\[10\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.data_inbuf_23._0_ net64 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[23\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.WW4END_inbuf_1._0_ net176 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[339\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[328\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[3\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[14\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_124_ Tile_X0Y0_DSP_top.N4BEG\[4\] VGND VGND VPWR VPWR net512 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.strobe_inbuf_8._0_ Tile_X0Y0_DSP_top.FrameStrobe\[8\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[8\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1420_ Tile_X0Y1_DSP_bot.Inst_MULADD._0569_ Tile_X0Y1_DSP_bot.Inst_MULADD._0570_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0563_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0588_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_150_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_055_ Tile_X0Y0_DSP_top.FrameData_O\[7\] VGND VGND VPWR VPWR net459 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1351_ Tile_X0Y1_DSP_bot.Inst_MULADD._0435_ Tile_X0Y1_DSP_bot.Inst_MULADD._0519_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_150_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1282_ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0141_ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0452_ sky130_fd_sc_hd__nand4_4
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.data_inbuf_14._0_ net54 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[14\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0997_ Tile_X0Y1_DSP_bot.Inst_MULADD._0135_ Tile_X0Y1_DSP_bot.Inst_MULADD._0159_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0165_ Tile_X0Y1_DSP_bot.Inst_MULADD._0169_ Tile_X0Y1_DSP_bot.Inst_MULADD._0170_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0171_ sky130_fd_sc_hd__a311o_1
XFILLER_0_158_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput30 Tile_X0Y0_E6END[7] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1618_ Tile_X0Y1_DSP_bot.Inst_MULADD._0765_ Tile_X0Y1_DSP_bot.Inst_MULADD._0771_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0778_ Tile_X0Y1_DSP_bot.Inst_MULADD._0780_ Tile_X0Y1_DSP_bot.Inst_MULADD._0764_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0781_ sky130_fd_sc_hd__o2111a_1
Xinput63 Tile_X0Y0_FrameData[22] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_8
Xinput52 Tile_X0Y0_FrameData[12] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_8
Xinput41 Tile_X0Y0_EE4END[2] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_2
Xinput96 Tile_X0Y0_S2MID[3] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__buf_4
Xinput85 Tile_X0Y0_S2END[0] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_2
Xinput74 Tile_X0Y0_FrameData[3] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1549_ Tile_X0Y1_DSP_bot.Inst_MULADD._0713_ Tile_X0Y1_DSP_bot.Inst_MULADD._0692_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0695_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0715_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID5
+ net18 net98 net150 Tile_X0Y0_DSP_top.ConfigBits\[194\] Tile_X0Y0_DSP_top.ConfigBits\[195\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_149_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[282\] Tile_X0Y0_DSP_top.ConfigBits\[283\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[340\] Tile_X0Y1_DSP_bot.ConfigBits\[341\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[121\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.SS4END_inbuf_7._0_ Tile_X0Y0_DSP_top.SS4BEG\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[7\] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.data_inbuf_23._0_ net244 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[23\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0920_ Tile_X0Y1_DSP_bot.Inst_MULADD._0095_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 sky130_fd_sc_hd__buf_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0851_ Tile_X0Y1_DSP_bot.Inst_MULADD._0028_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ sky130_fd_sc_hd__buf_4
XFILLER_0_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_107_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG3 VGND VGND VPWR VPWR net489
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_EF_BEG3 net42
+ net101 net172 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG3 Tile_X0Y0_DSP_top.ConfigBits\[396\]
+ Tile_X0Y0_DSP_top.ConfigBits\[397\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1403_ Tile_X0Y1_DSP_bot.Inst_MULADD._0483_ Tile_X0Y1_DSP_bot.Inst_MULADD._0491_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0490_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0572_
+ sky130_fd_sc_hd__a21boi_4
XFILLER_0_79_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_038_ Tile_X0Y0_DSP_top.EE4BEG\[6\] VGND VGND VPWR VPWR net426 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1334_ Tile_X0Y1_DSP_bot.Inst_MULADD._0502_ Tile_X0Y1_DSP_bot.Inst_MULADD._0503_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0504_ sky130_fd_sc_hd__nand2_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1265_ Tile_X0Y1_DSP_bot.Inst_MULADD._0434_ Tile_X0Y1_DSP_bot.Inst_MULADD._0416_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0342_ Tile_X0Y1_DSP_bot.Inst_MULADD._0417_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0435_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_95_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1196_ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_ Tile_X0Y1_DSP_bot.Inst_MULADD._0357_ Tile_X0Y1_DSP_bot.Inst_MULADD._0366_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0367_ sky130_fd_sc_hd__a41o_1
XFILLER_0_28_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.strobe_outbuf_0._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[0\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[0\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.data_inbuf_14._0_ net234 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[14\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[266\] Tile_X0Y1_DSP_bot.ConfigBits\[267\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_151_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1 net240 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[257\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[359\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[370\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[34\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[45\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._53_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG5 sky130_fd_sc_hd__clkbuf_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput220 Tile_X0Y1_EE4END[1] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1050_ Tile_X0Y1_DSP_bot.Inst_MULADD._0199_ Tile_X0Y1_DSP_bot.Inst_MULADD._0217_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0221_ Tile_X0Y1_DSP_bot.Inst_MULADD._0222_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0223_ sky130_fd_sc_hd__o211a_4
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_11._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG\[11\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.EE4END_inbuf_6._0_ net214 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
Xinput231 Tile_X0Y1_FrameData[11] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__buf_6
Xinput242 Tile_X0Y1_FrameData[21] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_8
Xinput253 Tile_X0Y1_FrameData[31] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__buf_6
Xinput286 Tile_X0Y1_N2END[1] VGND VGND VPWR VPWR net286 sky130_fd_sc_hd__clkbuf_2
Xinput297 Tile_X0Y1_N2MID[4] VGND VGND VPWR VPWR net297 sky130_fd_sc_hd__buf_2
Xinput275 Tile_X0Y1_FrameStrobe[4] VGND VGND VPWR VPWR net275 sky130_fd_sc_hd__buf_8
Xinput264 Tile_X0Y1_FrameStrobe[12] VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__clkbuf_16
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst1
+ net346 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[156\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[157\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_85_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.strobe_inbuf_15._0_ Tile_X0Y0_DSP_top.FrameStrobe\[15\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0903_ Tile_X0Y1_DSP_bot.ConfigBits\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ sky130_fd_sc_hd__buf_4
XFILLER_0_155_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_136_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput727 net727 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput716 net716 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput705 net705 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput749 net749 VGND VGND VPWR VPWR Tile_X0Y1_WW4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput738 net738 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[1] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG0 net199
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG6 net352 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG4
+ Tile_X0Y1_DSP_bot.ConfigBits\[168\] Tile_X0Y1_DSP_bot.ConfigBits\[169\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG0 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[304\] Tile_X0Y1_DSP_bot.ConfigBits\[305\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1317_ Tile_X0Y1_DSP_bot.Inst_MULADD._0485_ Tile_X0Y1_DSP_bot.Inst_MULADD._0486_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0454_ Tile_X0Y1_DSP_bot.Inst_MULADD._0443_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0487_ sky130_fd_sc_hd__o2bb2ai_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG2
+ Tile_X0Y0_DSP_top.ConfigBits\[52\] Tile_X0Y0_DSP_top.ConfigBits\[53\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1248_ Tile_X0Y1_DSP_bot.Inst_MULADD._0411_ Tile_X0Y1_DSP_bot.Inst_MULADD._0416_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0418_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0419_
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1179_ Tile_X0Y1_DSP_bot.Inst_MULADD._0345_ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0349_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0350_ sky130_fd_sc_hd__and4b_1
XFILLER_0_146_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6
+ Tile_X0Y0_DSP_top.ConfigBits\[144\] Tile_X0Y0_DSP_top.ConfigBits\[145\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_71_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._36_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG4 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.SS4END_inbuf_3._0_ net130 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[220\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_372_ Tile_X0Y1_DSP_bot.WW4BEG\[8\] VGND VGND VPWR VPWR net761 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_140_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.strobe_outbuf_17._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[17\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[17\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1102_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_ Tile_X0Y1_DSP_bot.Inst_MULADD._0188_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0273_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0274_ sky130_fd_sc_hd__o2bb2ai_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1033_ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0155_ Tile_X0Y1_DSP_bot.Inst_MULADD._0049_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0206_ sky130_fd_sc_hd__o2bb2ai_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[354\] Tile_X0Y0_DSP_top.ConfigBits\[355\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[390\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_128_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[401\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11 net51 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[65\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22 net63 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[76\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4 net255 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[356\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG1 net296
+ net196 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG3 net349 Tile_X0Y1_DSP_bot.ConfigBits\[210\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[211\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_143_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput502 net502 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[0] sky130_fd_sc_hd__buf_2
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput524 net524 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput513 net513 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[5] sky130_fd_sc_hd__buf_2
Xoutput535 net535 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput557 net557 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput568 net568 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput546 net546 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput579 net579 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[6] sky130_fd_sc_hd__clkbuf_4
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG2 net308
+ net204 net357 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[388\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[389\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[55\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._19_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG3 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.EE4END_inbuf_2._0_ net45 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_100 Tile_X0Y1_DSP_bot.NN4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 Tile_X0Y1_DSP_bot.SS4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 Tile_X0Y0_DSP_top.FrameStrobe\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 net151 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 net310 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1720_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0014_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_177 Tile_X0Y0_DSP_top.S4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 Tile_X0Y1_DSP_bot.SS4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_153_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_355_ Tile_X0Y1_DSP_bot.W6BEG\[3\] VGND VGND VPWR VPWR net740 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1651_ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.ConfigBits\[4\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0810_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0811_
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1582_ Tile_X0Y1_DSP_bot.Inst_MULADD._0746_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0747_
+ sky130_fd_sc_hd__mux2_1
X_286_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG2 VGND VGND VPWR VPWR net669
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_inst0
+ net283 net183 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.ConfigBits\[42\] Tile_X0Y1_DSP_bot.ConfigBits\[43\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[266\] Tile_X0Y0_DSP_top.ConfigBits\[267\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_23_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._21_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.strobe_outbuf_6._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[6\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[6\] sky130_fd_sc_hd__buf_8
XFILLER_0_127_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput6 Tile_X0Y0_E2END[1] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1016_ Tile_X0Y1_DSP_bot.Inst_MULADD._0142_ Tile_X0Y1_DSP_bot.Inst_MULADD._0143_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0112_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0189_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_160_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.N4BEG_outbuf_1._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END1 sky130_fd_sc_hd__buf_2
XFILLER_0_129_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.E6END_inbuf_8._0_ net22 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
Xoutput387 net387 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput398 net398 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[4] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END4
+ net33 net89 net141 Tile_X0Y0_DSP_top.ConfigBits\[218\] Tile_X0Y0_DSP_top.ConfigBits\[219\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_0_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[319\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_140_ Tile_X0Y0_DSP_top.NN4BEG\[4\] VGND VGND VPWR VPWR net528 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[376\] Tile_X0Y1_DSP_bot.ConfigBits\[377\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_135_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_071_ Tile_X0Y0_DSP_top.FrameData_O\[23\] VGND VGND VPWR VPWR net445 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_364 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_4._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[4\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst1
+ net81 net83 net117 net165 Tile_X0Y0_DSP_top.ConfigBits\[306\] Tile_X0Y0_DSP_top.ConfigBits\[307\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[318\] Tile_X0Y0_DSP_top.ConfigBits\[319\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_113_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1703_ Tile_X0Y1_DSP_bot.Inst_MULADD._0813_ Tile_X0Y1_DSP_bot.Inst_MULADD._0814_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0818_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0020_
+ sky130_fd_sc_hd__and3_1
XTile_X0Y0_DSP_top.E6BEG_outbuf_6._0_ Tile_X0Y0_DSP_top.E6BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[6\] sky130_fd_sc_hd__clkbuf_1
X_338_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG2 VGND VGND VPWR VPWR net721
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1634_ Tile_X0Y1_DSP_bot.Inst_MULADD._0790_ Tile_X0Y1_DSP_bot.Inst_MULADD._0795_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0796_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_153_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1565_ Tile_X0Y1_DSP_bot.Inst_MULADD._0696_ Tile_X0Y1_DSP_bot.Inst_MULADD._0699_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0729_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0730_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_269_ Tile_X0Y1_DSP_bot.FrameData_O\[21\] VGND VGND VPWR VPWR net644 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1496_ Tile_X0Y1_DSP_bot.Inst_MULADD._0643_ Tile_X0Y1_DSP_bot.Inst_MULADD._0659_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0662_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0663_
+ sky130_fd_sc_hd__nand3_2
XFILLER_0_3_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.strobe_outbuf_12._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[12\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[12\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._04_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.A4 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.W6BEG_outbuf_1._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.data_inbuf_3._0_ net74 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID4
+ net17 net149 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 Tile_X0Y0_DSP_top.ConfigBits\[154\]
+ Tile_X0Y0_DSP_top.ConfigBits\[155\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_59_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_22 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 Tile_X0Y0_DSP_top.FrameStrobe\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 Tile_X0Y0_DSP_top.N4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_66 Tile_X0Y0_DSP_top.S4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_99 Tile_X0Y1_DSP_bot.NN4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 Tile_X0Y0_DSP_top.S4BEG_i\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.E6END_inbuf_8._0_ net202 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[329\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame2_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[15\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[4\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_123_ Tile_X0Y0_DSP_top.N4BEG\[3\] VGND VGND VPWR VPWR net511 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_054_ Tile_X0Y0_DSP_top.FrameData_O\[6\] VGND VGND VPWR VPWR net458 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1350_ Tile_X0Y1_DSP_bot.Inst_MULADD._0517_ Tile_X0Y1_DSP_bot.Inst_MULADD._0492_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0518_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0519_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_150_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1281_ Tile_X0Y1_DSP_bot.Inst_MULADD._0446_ Tile_X0Y1_DSP_bot.Inst_MULADD._0450_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0451_ sky130_fd_sc_hd__nand2_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0996_ Tile_X0Y1_DSP_bot.Inst_MULADD._0159_ Tile_X0Y1_DSP_bot.Inst_MULADD._0165_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0135_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0170_
+ sky130_fd_sc_hd__a21oi_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_140_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput31 Tile_X0Y0_E6END[8] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput20 Tile_X0Y0_E2MID[7] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1617_ Tile_X0Y1_DSP_bot.Inst_MULADD._0351_ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0774_ Tile_X0Y1_DSP_bot.Inst_MULADD._0779_ Tile_X0Y1_DSP_bot.Inst_MULADD._0755_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0780_ sky130_fd_sc_hd__o311ai_4
Xinput64 Tile_X0Y0_FrameData[23] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_6
Xinput53 Tile_X0Y0_FrameData[13] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_8
Xinput42 Tile_X0Y0_EE4END[3] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1548_ Tile_X0Y1_DSP_bot.Inst_MULADD._0692_ Tile_X0Y1_DSP_bot.Inst_MULADD._0695_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0713_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0714_
+ sky130_fd_sc_hd__a21o_1
Xinput86 Tile_X0Y0_S2END[1] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__clkbuf_4
Xinput97 Tile_X0Y0_S2MID[4] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_4
Xinput75 Tile_X0Y0_FrameData[4] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_6
XTile_X0Y1_DSP_bot.data_outbuf_30._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[30\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[30\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1479_ Tile_X0Y1_DSP_bot.Inst_MULADD._0265_ Tile_X0Y1_DSP_bot.Inst_MULADD._0267_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0646_
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y0_DSP_top.NN4BEG_outbuf_1._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_149_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_CDb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID1
+ net14 net94 net146 Tile_X0Y0_DSP_top.ConfigBits\[196\] Tile_X0Y0_DSP_top.ConfigBits\[197\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_79_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_149_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[284\] Tile_X0Y0_DSP_top.ConfigBits\[285\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG1 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.SS4BEG_outbuf_4._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[340\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[341\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_outbuf_21._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[21\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[21\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[122\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0850_ Tile_X0Y1_DSP_bot.A0 Tile_X0Y1_DSP_bot.Inst_MULADD._0025_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0027_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0028_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0 net229 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[0\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_106_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG2 VGND VGND VPWR VPWR net488
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1402_ Tile_X0Y1_DSP_bot.Inst_MULADD._0563_ Tile_X0Y1_DSP_bot.Inst_MULADD._0569_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0570_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0571_
+ sky130_fd_sc_hd__nor3_1
XTile_X0Y1_DSP_bot.data_outbuf_12._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[12\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[12\] sky130_fd_sc_hd__clkbuf_1
X_037_ Tile_X0Y0_DSP_top.EE4BEG\[5\] VGND VGND VPWR VPWR net425 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1333_ Tile_X0Y1_DSP_bot.Inst_MULADD._0501_ Tile_X0Y1_DSP_bot.Inst_MULADD._0497_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0496_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0503_
+ sky130_fd_sc_hd__or3_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1264_ Tile_X0Y1_DSP_bot.Inst_MULADD._0429_ Tile_X0Y1_DSP_bot.Inst_MULADD._0433_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0319_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0434_
+ sky130_fd_sc_hd__a21oi_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.S4BEG_outbuf_1._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[1\] sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1195_ Tile_X0Y1_DSP_bot.Inst_MULADD._0261_ Tile_X0Y1_DSP_bot.Inst_MULADD._0263_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0070_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0366_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_88_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0979_ Tile_X0Y1_DSP_bot.Inst_MULADD._0028_ Tile_X0Y1_DSP_bot.Inst_MULADD._0151_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0152_ Tile_X0Y1_DSP_bot.Inst_MULADD._0040_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0153_ sky130_fd_sc_hd__a32o_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2 net251 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[258\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_114_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[360\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[371\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[35\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[46\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._52_ net141 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG4
+ sky130_fd_sc_hd__clkbuf_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput210 Tile_X0Y1_E6END[7] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
Xinput221 Tile_X0Y1_EE4END[2] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_2
Xinput254 Tile_X0Y1_FrameData[3] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__buf_6
Xinput232 Tile_X0Y1_FrameData[12] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_8
Xinput243 Tile_X0Y1_FrameData[22] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_8
Xinput287 Tile_X0Y1_N2END[2] VGND VGND VPWR VPWR net287 sky130_fd_sc_hd__clkbuf_2
Xinput276 Tile_X0Y1_FrameStrobe[5] VGND VGND VPWR VPWR net276 sky130_fd_sc_hd__clkbuf_16
Xinput265 Tile_X0Y1_FrameStrobe[13] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[156\] Tile_X0Y1_DSP_bot.ConfigBits\[157\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
Xinput298 Tile_X0Y1_N2MID[5] VGND VGND VPWR VPWR net298 sky130_fd_sc_hd__buf_2
XFILLER_0_58_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0902_ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0078_ sky130_fd_sc_hd__nand4_1
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput717 net717 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput706 net706 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput728 net728 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput739 net739 VGND VGND VPWR VPWR Tile_X0Y1_W6BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG1 net295
+ net195 net348 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG4 Tile_X0Y1_DSP_bot.ConfigBits\[170\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[171\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[306\] Tile_X0Y1_DSP_bot.ConfigBits\[307\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG4 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1316_ Tile_X0Y1_DSP_bot.Inst_MULADD._0455_ Tile_X0Y1_DSP_bot.Inst_MULADD._0457_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0486_ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[54\] Tile_X0Y0_DSP_top.ConfigBits\[55\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.E6BEG\[11\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1247_ Tile_X0Y1_DSP_bot.Inst_MULADD._0223_ Tile_X0Y1_DSP_bot.Inst_MULADD._0250_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0307_ Tile_X0Y1_DSP_bot.Inst_MULADD._0318_ Tile_X0Y1_DSP_bot.Inst_MULADD._0313_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0418_ sky130_fd_sc_hd__o221a_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1178_ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_ Tile_X0Y1_DSP_bot.Inst_MULADD._0049_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0283_ Tile_X0Y1_DSP_bot.Inst_MULADD._0343_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0349_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_55_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.NN4END_inbuf_7._0_ net319 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._35_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG3 sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[221\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_371_ Tile_X0Y1_DSP_bot.WW4BEG\[7\] VGND VGND VPWR VPWR net760 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1101_ Tile_X0Y1_DSP_bot.Inst_MULADD._0191_ Tile_X0Y1_DSP_bot.A6
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0257_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0273_
+ sky130_fd_sc_hd__a21boi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1032_ Tile_X0Y1_DSP_bot.Inst_MULADD._0040_ Tile_X0Y1_DSP_bot.Inst_MULADD._0073_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0205_ sky130_fd_sc_hd__nand4_4
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[356\] Tile_X0Y0_DSP_top.ConfigBits\[357\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_156_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst0
+ net281 net287 net187 net201 Tile_X0Y1_DSP_bot.ConfigBits\[356\] Tile_X0Y1_DSP_bot.ConfigBits\[357\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[391\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_132_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[402\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12 net52 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[66\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23 net64 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[77\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG2 net298
+ net198 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG5 net351 Tile_X0Y1_DSP_bot.ConfigBits\[212\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[213\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_7._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4END\[7\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5 net256 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[357\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput525 net525 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput503 net503 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput514 net514 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput536 net536 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput558 net558 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput569 net569 VGND VGND VPWR VPWR Tile_X0Y0_WW4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput547 net547 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_159_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG3 net301
+ net201 Tile_X0Y0_DSP_top.S4BEG\[0\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[390\] Tile_X0Y1_DSP_bot.ConfigBits\[391\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_130_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[56\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._18_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_112 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 Tile_X0Y1_DSP_bot.S4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 Tile_X0Y1_DSP_bot.SS4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_167 Tile_X0Y0_DSP_top.FrameStrobe\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 net345 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 net184 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_189 Tile_X0Y1_DSP_bot.SS4BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_178 Tile_X0Y0_DSP_top.S4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_354_ Tile_X0Y1_DSP_bot.W6BEG\[2\] VGND VGND VPWR VPWR net739 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1650_ Tile_X0Y1_DSP_bot.Inst_MULADD._0809_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0810_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1581_ Tile_X0Y1_DSP_bot.Inst_MULADD._0744_ Tile_X0Y1_DSP_bot.Inst_MULADD._0745_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0746_ sky130_fd_sc_hd__xor2_1
X_285_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG1 VGND VGND VPWR VPWR net668
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_inst1
+ net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[42\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[43\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[266\] Tile_X0Y0_DSP_top.ConfigBits\[267\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._20_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot16.X
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1015_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.Inst_MULADD._0186_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0187_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0188_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_127_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput7 Tile_X0Y0_E2END[2] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
XFILLER_0_36_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_inst0
+ net281 net181 net334 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[28\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[29\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.NN4END_inbuf_3._0_ Tile_X0Y0_DSP_top.NN4END\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst0
+ net184 net337 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.ConfigBits\[54\] Tile_X0Y1_DSP_bot.ConfigBits\[55\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput399 net399 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput388 net388 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[2] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_AB_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END0
+ net5 net85 net174 Tile_X0Y0_DSP_top.ConfigBits\[220\] Tile_X0Y0_DSP_top.ConfigBits\[221\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_93_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.EE4BEG_outbuf_4._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_11._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.SS4BEG\[11\] sky130_fd_sc_hd__buf_2
XFILLER_0_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[378\] Tile_X0Y1_DSP_bot.ConfigBits\[379\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6 sky130_fd_sc_hd__mux4_2
X_070_ Tile_X0Y0_DSP_top.FrameData_O\[22\] VGND VGND VPWR VPWR net444 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.data_inbuf_9._0_ net260 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[306\] Tile_X0Y0_DSP_top.ConfigBits\[307\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[320\] Tile_X0Y0_DSP_top.ConfigBits\[321\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2 sky130_fd_sc_hd__mux4_2
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1702_ Tile_X0Y1_DSP_bot.Inst_MULADD._0805_ Tile_X0Y1_DSP_bot.Inst_MULADD._0806_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0017_
+ sky130_fd_sc_hd__a21oi_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1633_ Tile_X0Y1_DSP_bot.Inst_MULADD._0780_ Tile_X0Y1_DSP_bot.Inst_MULADD._0793_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0794_ Tile_X0Y1_DSP_bot.Inst_MULADD._0770_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0795_ sky130_fd_sc_hd__o2bb2ai_2
X_337_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG1 VGND VGND VPWR VPWR net720
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst0
+ net324 net184 net186 net204 Tile_X0Y1_DSP_bot.ConfigBits\[320\] Tile_X0Y1_DSP_bot.ConfigBits\[321\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_141_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1564_ Tile_X0Y1_DSP_bot.Inst_MULADD._0701_ Tile_X0Y1_DSP_bot.Inst_MULADD._0728_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0729_ sky130_fd_sc_hd__xor2_1
XFILLER_0_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_268_ Tile_X0Y1_DSP_bot.FrameData_O\[20\] VGND VGND VPWR VPWR net643 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_199_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 VGND VGND VPWR VPWR net573
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1495_ Tile_X0Y1_DSP_bot.Inst_MULADD._0657_ Tile_X0Y1_DSP_bot.Inst_MULADD._0658_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0660_ Tile_X0Y1_DSP_bot.Inst_MULADD._0661_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_138_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_ABa_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID0
+ net13 net93 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG3 Tile_X0Y0_DSP_top.ConfigBits\[156\]
+ Tile_X0Y0_DSP_top.ConfigBits\[157\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0 net229 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[160\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_23 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 Tile_X0Y0_DSP_top.FrameStrobe\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 Tile_X0Y0_DSP_top.N4BEG\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_45 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_144_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_89 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 Tile_X0Y0_DSP_top.S4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 Tile_X0Y0_DSP_top.SS4BEG\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[5\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[16\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_25_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_122_ Tile_X0Y0_DSP_top.N4BEG\[2\] VGND VGND VPWR VPWR net510 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_053_ Tile_X0Y0_DSP_top.FrameData_O\[5\] VGND VGND VPWR VPWR net457 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG0 net326
+ net191 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb6 net344 Tile_X0Y1_DSP_bot.ConfigBits\[232\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[233\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1280_ Tile_X0Y1_DSP_bot.Inst_MULADD._0448_ Tile_X0Y1_DSP_bot.Inst_MULADD._0449_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0450_ sky130_fd_sc_hd__nand2_4
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.WW4END_inbuf_10._0_ net371 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0995_ Tile_X0Y1_DSP_bot.Inst_MULADD._0122_ Tile_X0Y1_DSP_bot.Inst_MULADD._0082_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0121_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0169_
+ sky130_fd_sc_hd__nand3_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput21 Tile_X0Y0_E6END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__buf_4
Xinput10 Tile_X0Y0_E2END[5] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1616_ Tile_X0Y1_DSP_bot.Inst_MULADD._0777_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0779_ sky130_fd_sc_hd__inv_2
Xinput54 Tile_X0Y0_FrameData[14] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_8
Xinput32 Tile_X0Y0_E6END[9] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput43 Tile_X0Y0_EE4END[4] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1547_ Tile_X0Y1_DSP_bot.Inst_MULADD._0710_ Tile_X0Y1_DSP_bot.Inst_MULADD._0712_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0713_ sky130_fd_sc_hd__nand2_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput98 Tile_X0Y0_S2MID[5] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_4
Xinput87 Tile_X0Y0_S2END[2] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_2
Xinput65 Tile_X0Y0_FrameData[24] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput76 Tile_X0Y0_FrameData[5] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__clkbuf_8
XTile_X0Y0_DSP_top.S4END_inbuf_2._0_ net113 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1478_ Tile_X0Y1_DSP_bot.Inst_MULADD._0155_ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0645_ sky130_fd_sc_hd__o211a_1
XFILLER_0_149_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.N4BEG_outbuf_11._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4END\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[342\] Tile_X0Y1_DSP_bot.ConfigBits\[343\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net83 net135 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.ConfigBits\[92\] Tile_X0Y0_DSP_top.ConfigBits\[93\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.strobe_inbuf_2._0_ net273 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[2\]
+ sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[123\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_85_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1 net240 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[1\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_155_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.W6END_inbuf_6._0_ net163 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_105_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG1 VGND VGND VPWR VPWR net487
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1401_ Tile_X0Y1_DSP_bot.Inst_MULADD._0484_ Tile_X0Y1_DSP_bot.Inst_MULADD._0558_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0560_ Tile_X0Y1_DSP_bot.Inst_MULADD._0561_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0570_ sky130_fd_sc_hd__o211a_2
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_036_ Tile_X0Y0_DSP_top.EE4BEG\[4\] VGND VGND VPWR VPWR net424 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1332_ Tile_X0Y1_DSP_bot.Inst_MULADD._0496_ Tile_X0Y1_DSP_bot.Inst_MULADD._0497_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0501_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0502_
+ sky130_fd_sc_hd__o21ai_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1263_ Tile_X0Y1_DSP_bot.Inst_MULADD._0432_ Tile_X0Y1_DSP_bot.Inst_MULADD._0414_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0433_ sky130_fd_sc_hd__nand2_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1194_ Tile_X0Y1_DSP_bot.Inst_MULADD._0361_ Tile_X0Y1_DSP_bot.Inst_MULADD._0362_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0364_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0365_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_88_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._0978_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\] Tile_X0Y1_DSP_bot.Inst_MULADD._0067_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0152_ sky130_fd_sc_hd__or2b_2
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3 net254 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[259\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[361\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.S4END_inbuf_2._0_ Tile_X0Y0_DSP_top.S4BEG\[6\] VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.S4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[36\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[47\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._51_ net140 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG3
+ sky130_fd_sc_hd__clkbuf_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.SS4END_inbuf_10._0_ net122 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_145_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput200 Tile_X0Y1_E2MID[7] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__clkbuf_4
Xinput211 Tile_X0Y1_E6END[8] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
Xinput222 Tile_X0Y1_EE4END[3] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__buf_1
Xinput233 Tile_X0Y1_FrameData[13] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_8
Xinput244 Tile_X0Y1_FrameData[23] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__buf_4
Xinput288 Tile_X0Y1_N2END[3] VGND VGND VPWR VPWR net288 sky130_fd_sc_hd__clkbuf_4
Xinput277 Tile_X0Y1_FrameStrobe[6] VGND VGND VPWR VPWR net277 sky130_fd_sc_hd__clkbuf_16
Xinput266 Tile_X0Y1_FrameStrobe[14] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ net765 net766 Tile_X0Y1_DSP_bot.ConfigBits\[156\] Tile_X0Y1_DSP_bot.ConfigBits\[157\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
Xinput255 Tile_X0Y1_FrameData[4] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_8
Xinput299 Tile_X0Y1_N2MID[6] VGND VGND VPWR VPWR net299 sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0901_ Tile_X0Y1_DSP_bot.Inst_MULADD._0050_ Tile_X0Y1_DSP_bot.Inst_MULADD._0063_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0066_ Tile_X0Y1_DSP_bot.Inst_MULADD._0072_ Tile_X0Y1_DSP_bot.Inst_MULADD._0076_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0077_ sky130_fd_sc_hd__o311a_1
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput718 net718 VGND VGND VPWR VPWR Tile_X0Y1_W1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput707 net707 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.W6END_inbuf_6._0_ net364 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
X_019_ Tile_X0Y0_DSP_top.E2BEGb\[7\] VGND VGND VPWR VPWR net401 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1315_ Tile_X0Y1_DSP_bot.Inst_MULADD._0450_ Tile_X0Y1_DSP_bot.Inst_MULADD._0446_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0462_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0485_
+ sky130_fd_sc_hd__a21o_1
Xoutput729 net729 VGND VGND VPWR VPWR Tile_X0Y1_W2BEGb[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG2 net297
+ net197 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ Tile_X0Y1_DSP_bot.ConfigBits\[172\] Tile_X0Y1_DSP_bot.ConfigBits\[173\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG2 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1246_ Tile_X0Y1_DSP_bot.Inst_MULADD._0305_ Tile_X0Y1_DSP_bot.Inst_MULADD._0329_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0411_ Tile_X0Y1_DSP_bot.Inst_MULADD._0416_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0417_ sky130_fd_sc_hd__a22oi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1177_ Tile_X0Y1_DSP_bot.Inst_MULADD._0347_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0348_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_127_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END1
+ net4 net6 Tile_X0Y0_DSP_top.ConfigBits\[246\] Tile_X0Y0_DSP_top.ConfigBits\[247\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._34_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG2 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[222\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
X_370_ Tile_X0Y1_DSP_bot.WW4BEG\[6\] VGND VGND VPWR VPWR net759 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_118_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.WW4END_inbuf_8._0_ net369 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1100_ Tile_X0Y1_DSP_bot.Inst_MULADD._0264_ Tile_X0Y1_DSP_bot.Inst_MULADD._0268_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0271_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0272_
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1031_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.Inst_MULADD._0202_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0203_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0204_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_116_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb2 Tile_X0Y0_DSP_top.S4BEG\[2\]
+ net340 net354 Tile_X0Y1_DSP_bot.ConfigBits\[356\] Tile_X0Y1_DSP_bot.ConfigBits\[357\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[392\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[403\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13 net53 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[67\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24 net65 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[78\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG3 net294
+ net194 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG1 net347 Tile_X0Y1_DSP_bot.ConfigBits\[214\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[215\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6 net257 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[358\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput526 net526 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput504 net504 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[11] sky130_fd_sc_hd__clkbuf_4
Xoutput515 net515 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput559 net559 VGND VGND VPWR VPWR Tile_X0Y0_W6BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput548 net548 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput537 net537 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1229_ Tile_X0Y1_DSP_bot.Inst_MULADD._0327_ Tile_X0Y1_DSP_bot.Inst_MULADD._0309_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0321_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0400_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_66_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_119_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[57\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_99_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._17_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_124 Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_102 Tile_X0Y1_DSP_bot.S4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_113 Tile_X0Y1_DSP_bot.SS4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 Tile_X0Y1_DSP_bot.SS4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 net198 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 net373 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_179 Tile_X0Y0_DSP_top.S4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_168 Tile_X0Y0_DSP_top.FrameStrobe\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_353_ Tile_X0Y1_DSP_bot.W6BEG\[1\] VGND VGND VPWR VPWR net738 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1580_ Tile_X0Y1_DSP_bot.Inst_MULADD._0690_ Tile_X0Y1_DSP_bot.Inst_MULADD._0721_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0720_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0745_
+ sky130_fd_sc_hd__a21bo_1
X_284_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG0 VGND VGND VPWR VPWR net667
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[268\] Tile_X0Y0_DSP_top.ConfigBits\[269\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 sky130_fd_sc_hd__mux4_2
XFILLER_0_121_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_121_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst0
+ net289 net301 net183 net189 Tile_X0Y1_DSP_bot.ConfigBits\[268\] Tile_X0Y1_DSP_bot.ConfigBits\[269\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1014_ Tile_X0Y1_DSP_bot.Inst_MULADD._0026_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0187_ sky130_fd_sc_hd__nand2_1
Xinput8 Tile_X0Y0_E2END[3] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_127_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[28\] Tile_X0Y1_DSP_bot.ConfigBits\[29\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_143_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.data_outbuf_2._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[2\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.ConfigBits\[54\] Tile_X0Y1_DSP_bot.ConfigBits\[55\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput389 net389 VGND VGND VPWR VPWR Tile_X0Y0_E2BEG[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._79_ net347 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb1
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 net1 net81 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[42\] Tile_X0Y0_DSP_top.ConfigBits\[43\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.data_inbuf_26._0_ net67 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[26\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.WW4END_inbuf_4._0_ net179 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[306\] Tile_X0Y0_DSP_top.ConfigBits\[307\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_S1BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[62\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[63\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0
+ sky130_fd_sc_hd__mux4_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1701_ Tile_X0Y1_DSP_bot.Inst_MULADD._0842_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0016_ sky130_fd_sc_hd__clkbuf_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1632_ Tile_X0Y1_DSP_bot.Inst_MULADD._0763_ Tile_X0Y1_DSP_bot.Inst_MULADD._0764_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0778_ Tile_X0Y1_DSP_bot.Inst_MULADD._0780_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0794_ sky130_fd_sc_hd__nand4_1
X_336_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG0 VGND VGND VPWR VPWR net719
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb1 Tile_X0Y0_DSP_top.S4BEG\[1\]
+ net339 net357 Tile_X0Y1_DSP_bot.ConfigBits\[320\] Tile_X0Y1_DSP_bot.ConfigBits\[321\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_141_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1563_ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_ Tile_X0Y1_DSP_bot.Inst_MULADD._0726_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0727_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0728_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_267_ Tile_X0Y1_DSP_bot.FrameData_O\[19\] VGND VGND VPWR VPWR net641 sky130_fd_sc_hd__clkbuf_1
X_198_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG2 VGND VGND VPWR VPWR net572
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1494_ Tile_X0Y1_DSP_bot.Inst_MULADD._0151_ Tile_X0Y1_DSP_bot.Inst_MULADD._0152_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0661_ sky130_fd_sc_hd__a32o_1
XTile_X0Y0_DSP_top.data_inbuf_17._0_ net57 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[17\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_154_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1 net240 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[161\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[342\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_13 Tile_X0Y0_DSP_top.FrameStrobe\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_57 Tile_X0Y0_DSP_top.N4BEG\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID3 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_35 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_24 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_68 Tile_X0Y0_DSP_top.S4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 Tile_X0Y0_DSP_top.SS4BEG\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.data_outbuf_2._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[2\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.EE4END_inbuf_10._0_ net38 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[6\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_92_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_121_ Tile_X0Y0_DSP_top.N4BEG\[1\] VGND VGND VPWR VPWR net509 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[17\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_052_ Tile_X0Y0_DSP_top.FrameData_O\[4\] VGND VGND VPWR VPWR net456 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG1 net287
+ net187 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb2 net374 Tile_X0Y1_DSP_bot.ConfigBits\[234\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[235\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.E6BEG_outbuf_0._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[0\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.data_inbuf_26._0_ net247 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[26\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0994_ Tile_X0Y1_DSP_bot.Inst_MULADD._0082_ Tile_X0Y1_DSP_bot.Inst_MULADD._0121_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0122_ Tile_X0Y1_DSP_bot.Inst_MULADD._0166_ Tile_X0Y1_DSP_bot.Inst_MULADD._0167_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0168_ sky130_fd_sc_hd__a32o_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_130_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 Tile_X0Y0_E6END[10] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 Tile_X0Y0_E2END[6] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1615_ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.Inst_MULADD._0777_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0778_ sky130_fd_sc_hd__nand2_1
X_319_ Tile_X0Y1_DSP_bot.SS4BEG\[3\] VGND VGND VPWR VPWR net708 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput55 Tile_X0Y0_FrameData[15] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_141_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput44 Tile_X0Y0_EE4END[5] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput33 Tile_X0Y0_EE4END[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1546_ Tile_X0Y1_DSP_bot.Inst_MULADD._0711_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0712_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput88 Tile_X0Y0_S2END[3] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__clkbuf_2
Xinput66 Tile_X0Y0_FrameData[25] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_8
Xinput77 Tile_X0Y0_FrameData[6] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput99 Tile_X0Y0_S2MID[6] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1477_ Tile_X0Y1_DSP_bot.Inst_MULADD._0209_ Tile_X0Y1_DSP_bot.Inst_MULADD._0273_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0644_ sky130_fd_sc_hd__o211a_1
XTile_X0Y0_DSP_top.strobe_outbuf_3._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[3\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[3\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.data_inbuf_17._0_ net237 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[17\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[41\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG\[13\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_inst0
+ net281 net181 net334 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[84\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[85\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG2
+ Tile_X0Y0_DSP_top.ConfigBits\[92\] Tile_X0Y0_DSP_top.ConfigBits\[93\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[124\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_85_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2 net251 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[2\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_104_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG0 VGND VGND VPWR VPWR net486
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1400_ Tile_X0Y1_DSP_bot.Inst_MULADD._0560_ Tile_X0Y1_DSP_bot.Inst_MULADD._0561_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0568_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0569_
+ sky130_fd_sc_hd__a21oi_1
X_035_ Tile_X0Y0_DSP_top.EE4BEG\[3\] VGND VGND VPWR VPWR net423 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1331_ Tile_X0Y1_DSP_bot.Inst_MULADD._0423_ Tile_X0Y1_DSP_bot.Inst_MULADD._0499_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0500_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0501_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1262_ Tile_X0Y1_DSP_bot.Inst_MULADD._0409_ Tile_X0Y1_DSP_bot.Inst_MULADD._0430_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0431_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0432_
+ sky130_fd_sc_hd__o21ai_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.EE4END_inbuf_9._0_ net217 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1193_ Tile_X0Y1_DSP_bot.Inst_MULADD._0050_ Tile_X0Y1_DSP_bot.Inst_MULADD._0192_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0268_ Tile_X0Y1_DSP_bot.Inst_MULADD._0271_ Tile_X0Y1_DSP_bot.Inst_MULADD._0363_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0364_ sky130_fd_sc_hd__o32a_1
XTile_X0Y0_DSP_top.WW4BEG_outbuf_1._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[1\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.strobe_inbuf_18._0_ Tile_X0Y0_DSP_top.FrameStrobe\[18\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._0977_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ Tile_X0Y1_DSP_bot.B4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0151_ sky130_fd_sc_hd__or2_2
XFILLER_0_29_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4 net255 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[260\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1529_ Tile_X0Y1_DSP_bot.Inst_MULADD._0691_ Tile_X0Y1_DSP_bot.Inst_MULADD._0591_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0573_ Tile_X0Y1_DSP_bot.Inst_MULADD._0694_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0695_ sky130_fd_sc_hd__a31oi_4
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[48\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[37\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._50_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG2 sky130_fd_sc_hd__clkbuf_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.strobe_inbuf_11._0_ net263 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[11\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_7_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput201 Tile_X0Y1_E6END[0] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_4
Xinput223 Tile_X0Y1_EE4END[4] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_1
Xinput212 Tile_X0Y1_E6END[9] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
Xinput234 Tile_X0Y1_FrameData[14] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_8
Xinput245 Tile_X0Y1_FrameData[24] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__clkbuf_8
Xinput278 Tile_X0Y1_FrameStrobe[7] VGND VGND VPWR VPWR net278 sky130_fd_sc_hd__buf_8
Xinput267 Tile_X0Y1_FrameStrobe[15] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_clr.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[158\] Tile_X0Y1_DSP_bot.ConfigBits\[159\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.clr sky130_fd_sc_hd__mux4_2
Xinput256 Tile_X0Y1_FrameData[5] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__clkbuf_8
Xinput289 Tile_X0Y1_N2END[4] VGND VGND VPWR VPWR net289 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.SS4END_inbuf_6._0_ net118 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0900_ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_155_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput708 net708 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[3] sky130_fd_sc_hd__clkbuf_4
X_018_ Tile_X0Y0_DSP_top.E2BEGb\[6\] VGND VGND VPWR VPWR net400 sky130_fd_sc_hd__clkbuf_1
Xoutput719 net719 VGND VGND VPWR VPWR Tile_X0Y1_W2BEG[0] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG3 net293
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG0 net346 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG4
+ Tile_X0Y1_DSP_bot.ConfigBits\[174\] Tile_X0Y1_DSP_bot.ConfigBits\[175\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG3 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1314_ Tile_X0Y1_DSP_bot.Inst_MULADD._0443_ Tile_X0Y1_DSP_bot.Inst_MULADD._0454_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0458_ Tile_X0Y1_DSP_bot.Inst_MULADD._0460_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0484_ sky130_fd_sc_hd__o211a_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1245_ Tile_X0Y1_DSP_bot.Inst_MULADD._0307_ Tile_X0Y1_DSP_bot.Inst_MULADD._0413_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0414_ Tile_X0Y1_DSP_bot.Inst_MULADD._0415_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0416_ sky130_fd_sc_hd__o211ai_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1176_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B7
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0346_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0347_
+ sky130_fd_sc_hd__o21a_4
XFILLER_0_71_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst1
+ net24 net124 net138 net156 Tile_X0Y0_DSP_top.ConfigBits\[246\] Tile_X0Y0_DSP_top.ConfigBits\[247\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_154_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._33_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG1 sky130_fd_sc_hd__clkbuf_2
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[223\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame5_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_67_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[47\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG\[13\] sky130_fd_sc_hd__o21ai_2
XFILLER_0_137_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1030_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0203_ sky130_fd_sc_hd__nand2_2
XTile_X0Y0_DSP_top.EE4END_inbuf_5._0_ net48 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_116_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[356\] Tile_X0Y1_DSP_bot.ConfigBits\[357\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_156_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[393\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14 net54 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[68\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_109_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25 net66 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[79\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7 net258 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[359\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput505 net505 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput527 net527 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput516 net516 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.strobe_outbuf_9._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[9\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[9\] sky130_fd_sc_hd__buf_8
Xoutput549 net549 VGND VGND VPWR VPWR Tile_X0Y0_W2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput538 net538 VGND VGND VPWR VPWR Tile_X0Y0_W1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._95_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q19
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 sky130_fd_sc_hd__buf_8
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1228_ Tile_X0Y1_DSP_bot.Inst_MULADD._0395_ Tile_X0Y1_DSP_bot.Inst_MULADD._0396_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0398_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0399_
+ sky130_fd_sc_hd__nand3_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END3 net8 Tile_X0Y0_DSP_top.ConfigBits\[286\]
+ Tile_X0Y0_DSP_top.ConfigBits\[287\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1159_ Tile_X0Y1_DSP_bot.Inst_MULADD._0185_ Tile_X0Y1_DSP_bot.Inst_MULADD._0326_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0330_ Tile_X0Y1_DSP_bot.Inst_MULADD._0166_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0331_ sky130_fd_sc_hd__nand4_4
XTile_X0Y1_DSP_bot.N4BEG_outbuf_4._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4END\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[58\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._16_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEG0 sky130_fd_sc_hd__clkbuf_1
XANTENNA_103 Tile_X0Y1_DSP_bot.S4BEG\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 Tile_X0Y1_DSP_bot.SS4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_136 Tile_X0Y1_DSP_bot.SS4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 net374 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 Tile_X0Y0_DSP_top.FrameStrobe\[18\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_352_ Tile_X0Y1_DSP_bot.W6BEG\[0\] VGND VGND VPWR VPWR net735 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_283_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3 VGND VGND VPWR VPWR net666
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst1
+ net201 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb4 net342 net354 Tile_X0Y1_DSP_bot.ConfigBits\[268\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[269\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_7._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[7\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1013_ Tile_X0Y1_DSP_bot.A5 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0186_
+ sky130_fd_sc_hd__inv_2
Xinput9 Tile_X0Y0_E2END[4] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[24\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.E6BEG_outbuf_9._0_ Tile_X0Y0_DSP_top.E6BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_156_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.strobe_outbuf_15._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[15\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[15\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_E1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG1 Tile_X0Y0_DSP_top.ConfigBits\[28\]
+ Tile_X0Y0_DSP_top.ConfigBits\[29\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E1BEG\[0\]
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst2
+ net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[54\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[55\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._78_ net346 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb0
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.data_inbuf_6._0_ net77 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.W6BEG_outbuf_4._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[4\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG0
+ Tile_X0Y0_DSP_top.ConfigBits\[42\] Tile_X0Y0_DSP_top.ConfigBits\[43\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.N4END_inbuf_2._0_ Tile_X0Y0_DSP_top.N4END\[6\] VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[308\] Tile_X0Y0_DSP_top.ConfigBits\[309\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG7 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_S1BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[64\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[65\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_87_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst0
+ net283 net291 net183 net191 Tile_X0Y1_DSP_bot.ConfigBits\[308\] Tile_X0Y1_DSP_bot.ConfigBits\[309\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1700_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0799_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0796_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0842_
+ sky130_fd_sc_hd__and3b_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1631_ Tile_X0Y1_DSP_bot.Inst_MULADD._0791_ Tile_X0Y1_DSP_bot.Inst_MULADD._0792_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0793_ sky130_fd_sc_hd__nand2_1
X_335_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net718
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_153_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1562_ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0727_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_266_ Tile_X0Y1_DSP_bot.FrameData_O\[18\] VGND VGND VPWR VPWR net640 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst2
+ net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[320\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[321\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_3_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_197_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 VGND VGND VPWR VPWR net571
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1493_ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0660_ sky130_fd_sc_hd__nand4_4
XFILLER_0_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.N4BEG_outbuf_0._0_ Tile_X0Y0_DSP_top.N4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2 net251 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[162\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[343\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_14 Tile_X0Y0_DSP_top.FrameStrobe\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_117_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_36 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_25 Tile_X0Y0_DSP_top.FrameStrobe\[19\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 Tile_X0Y0_DSP_top.N4BEG\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 Tile_X0Y0_DSP_top.S4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.NN4BEG_outbuf_4._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[4\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_120_ Tile_X0Y0_DSP_top.N4BEG\[0\] VGND VGND VPWR VPWR net502 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.SS4BEG_outbuf_7._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[18\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[7\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_135_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.data_outbuf_24._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[24\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[24\] sky130_fd_sc_hd__clkbuf_1
X_051_ Tile_X0Y0_DSP_top.FrameData_O\[3\] VGND VGND VPWR VPWR net455 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END5
+ net2 net10 Tile_X0Y0_DSP_top.ConfigBits\[358\] Tile_X0Y0_DSP_top.ConfigBits\[359\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_123_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG2 net289
+ net189 Tile_X0Y0_DSP_top.SS4BEG\[2\] net342 Tile_X0Y1_DSP_bot.ConfigBits\[236\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[237\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.N4END_inbuf_2._0_ net313 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.S4BEG_outbuf_11._0_ Tile_X0Y0_DSP_top.S4BEG_i\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_158_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0993_ Tile_X0Y1_DSP_bot.Inst_MULADD._0159_ Tile_X0Y1_DSP_bot.Inst_MULADD._0165_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0135_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0167_
+ sky130_fd_sc_hd__a21o_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_140_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput12 Tile_X0Y0_E2END[7] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_2
XFILLER_0_114_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1614_ Tile_X0Y1_DSP_bot.Inst_MULADD._0776_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[15\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0423_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0777_
+ sky130_fd_sc_hd__mux2_1
X_318_ Tile_X0Y1_DSP_bot.SS4BEG\[2\] VGND VGND VPWR VPWR net707 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.data_outbuf_15._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[15\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[15\] sky130_fd_sc_hd__clkbuf_1
Xinput23 Tile_X0Y0_E6END[11] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput34 Tile_X0Y0_EE4END[10] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 Tile_X0Y0_EE4END[6] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1545_ Tile_X0Y1_DSP_bot.Inst_MULADD._0709_ Tile_X0Y1_DSP_bot.Inst_MULADD._0706_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0707_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0711_
+ sky130_fd_sc_hd__nor3_1
X_249_ Tile_X0Y1_DSP_bot.FrameData_O\[1\] VGND VGND VPWR VPWR net642 sky130_fd_sc_hd__clkbuf_1
Xinput89 Tile_X0Y0_S2END[4] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_2
Xinput67 Tile_X0Y0_FrameData[26] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_8
Xinput56 Tile_X0Y0_FrameData[16] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_8
Xinput78 Tile_X0Y0_FrameData[7] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__clkbuf_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1476_ Tile_X0Y1_DSP_bot.Inst_MULADD._0597_ Tile_X0Y1_DSP_bot.Inst_MULADD._0598_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0604_ Tile_X0Y1_DSP_bot.Inst_MULADD._0609_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0643_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_0._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.S4BEG_outbuf_4._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[4\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.W6BEG_outbuf_0._0_ Tile_X0Y0_DSP_top.W6BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[30\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4END\[14\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[41\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[84\] Tile_X0Y1_DSP_bot.ConfigBits\[85\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[125\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_93_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3 net254 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[3\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_108_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_103_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3 VGND VGND VPWR VPWR net485
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_034_ Tile_X0Y0_DSP_top.EE4BEG\[2\] VGND VGND VPWR VPWR net422 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1330_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] Tile_X0Y1_DSP_bot.Inst_MULADD._0423_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0500_ sky130_fd_sc_hd__or2b_1
XFILLER_0_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1261_ Tile_X0Y1_DSP_bot.Inst_MULADD._0286_ Tile_X0Y1_DSP_bot.Inst_MULADD._0292_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0327_ Tile_X0Y1_DSP_bot.Inst_MULADD._0309_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0431_ sky130_fd_sc_hd__o22a_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1192_ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_ Tile_X0Y1_DSP_bot.Inst_MULADD._0188_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_ Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0363_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_119_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_158_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0976_ Tile_X0Y1_DSP_bot.Inst_MULADD._0114_ Tile_X0Y1_DSP_bot.Inst_MULADD._0149_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0150_ sky130_fd_sc_hd__nand2_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5 net256 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[261\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1528_ Tile_X0Y1_DSP_bot.Inst_MULADD._0670_ Tile_X0Y1_DSP_bot.Inst_MULADD._0673_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0693_ Tile_X0Y1_DSP_bot.Inst_MULADD._0641_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0694_ sky130_fd_sc_hd__o22ai_2
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1459_ Tile_X0Y1_DSP_bot.C10 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[10\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0627_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst0
+ net281 net285 net181 net185 Tile_X0Y1_DSP_bot.ConfigBits\[380\] Tile_X0Y1_DSP_bot.ConfigBits\[381\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[49\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[38\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.data_outbuf_20._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[20\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[20\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END4 net3 net9 net21 Tile_X0Y0_DSP_top.ConfigBits\[322\]
+ Tile_X0Y0_DSP_top.ConfigBits\[323\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[103\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG3 sky130_fd_sc_hd__o21ai_1
Xinput202 Tile_X0Y1_E6END[10] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_1
Xinput213 Tile_X0Y1_EE4END[0] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_2
Xinput224 Tile_X0Y1_EE4END[5] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_1
Xinput235 Tile_X0Y1_FrameData[15] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__clkbuf_8
Xinput279 Tile_X0Y1_FrameStrobe[8] VGND VGND VPWR VPWR net279 sky130_fd_sc_hd__clkbuf_16
Xinput268 Tile_X0Y1_FrameStrobe[16] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__clkbuf_1
Xinput257 Tile_X0Y1_FrameData[6] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_8
Xinput246 Tile_X0Y1_FrameData[25] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.data_outbuf_11._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput709 net709 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[4] sky130_fd_sc_hd__buf_2
X_017_ Tile_X0Y0_DSP_top.E2BEGb\[5\] VGND VGND VPWR VPWR net399 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1313_ Tile_X0Y1_DSP_bot.Inst_MULADD._0437_ Tile_X0Y1_DSP_bot.Inst_MULADD._0477_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0482_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0483_
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_104_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1244_ Tile_X0Y1_DSP_bot.Inst_MULADD._0205_ Tile_X0Y1_DSP_bot.Inst_MULADD._0215_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0415_ sky130_fd_sc_hd__a211oi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1175_ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[7\] Tile_X0Y1_DSP_bot.Inst_MULADD._0047_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0346_ sky130_fd_sc_hd__or2_2
XTile_X0Y0_DSP_top.S4BEG_outbuf_0._0_ Tile_X0Y0_DSP_top.S4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[0\] sky130_fd_sc_hd__buf_2
XFILLER_0_146_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0959_ Tile_X0Y1_DSP_bot.Inst_MULADD._0101_ Tile_X0Y1_DSP_bot.Inst_MULADD._0132_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0133_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[246\] Tile_X0Y0_DSP_top.ConfigBits\[247\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._32_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG0 sky130_fd_sc_hd__buf_2
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[47\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.ConfigBits\[356\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[357\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_39_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15 net55 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[69\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26 net67 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[80\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_109_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8 net259 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[360\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput506 net506 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[13] sky130_fd_sc_hd__clkbuf_4
Xoutput517 net517 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_0_124_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput528 net528 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[4] sky130_fd_sc_hd__buf_2
Xoutput539 net539 VGND VGND VPWR VPWR Tile_X0Y0_W2BEG[0] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._94_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q18
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 sky130_fd_sc_hd__buf_8
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1227_ Tile_X0Y1_DSP_bot.Inst_MULADD._0345_ Tile_X0Y1_DSP_bot.Inst_MULADD._0397_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0353_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0398_
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst1
+ net24 net88 net140 net156 Tile_X0Y0_DSP_top.ConfigBits\[286\] Tile_X0Y0_DSP_top.ConfigBits\[287\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1158_ Tile_X0Y1_DSP_bot.Inst_MULADD._0305_ Tile_X0Y1_DSP_bot.Inst_MULADD._0329_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0315_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0330_
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst0
+ net284 net292 net184 net192 Tile_X0Y1_DSP_bot.ConfigBits\[344\] Tile_X0Y1_DSP_bot.ConfigBits\[345\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1089_ Tile_X0Y1_DSP_bot.Inst_MULADD._0260_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0261_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_159_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.NN4END_inbuf_6._0_ Tile_X0Y0_DSP_top.NN4END\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_115_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[59\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._15_ net20 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEGb\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_104 Tile_X0Y1_DSP_bot.S4BEG\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 Tile_X0Y1_DSP_bot.SS4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 Tile_X0Y1_DSP_bot.SS4BEG_i\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top.EE4BEG_outbuf_7._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_148 net220 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 Tile_X0Y1_DSP_bot.SS4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_159 Tile_X0Y0_DSP_top.FrameStrobe\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_351_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb7 VGND VGND VPWR VPWR net734
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_282_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 VGND VGND VPWR VPWR net665
+ sky130_fd_sc_hd__buf_1
XFILLER_0_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[109\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG3 sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[268\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[269\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1012_ Tile_X0Y1_DSP_bot.Inst_MULADD._0121_ Tile_X0Y1_DSP_bot.Inst_MULADD._0122_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0167_ Tile_X0Y1_DSP_bot.Inst_MULADD._0082_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0185_ sky130_fd_sc_hd__and4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[24\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_E1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG2 Tile_X0Y0_DSP_top.ConfigBits\[30\]
+ Tile_X0Y0_DSP_top.ConfigBits\[31\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E1BEG\[1\]
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_0._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[0\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[54\] Tile_X0Y1_DSP_bot.ConfigBits\[55\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_124_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._77_ net345 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG7
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.N4END_inbuf_10._0_ net306 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30 net252 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[126\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_135_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_S1BEG2 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[66\] Tile_X0Y1_DSP_bot.ConfigBits\[67\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG2 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb6 net336 Tile_X0Y1_DSP_bot.ConfigBits\[308\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[309\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1630_ Tile_X0Y1_DSP_bot.Inst_MULADD._0755_ Tile_X0Y1_DSP_bot.Inst_MULADD._0760_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0762_ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.Inst_MULADD._0777_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0792_ sky130_fd_sc_hd__a32oi_1
X_334_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG2 VGND VGND VPWR VPWR net717
+ sky130_fd_sc_hd__clkbuf_1
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1561_ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0726_
+ sky130_fd_sc_hd__and3_1
X_265_ Tile_X0Y1_DSP_bot.FrameData_O\[17\] VGND VGND VPWR VPWR net639 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.ConfigBits\[320\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[321\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
X_196_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG0 VGND VGND VPWR VPWR net570
+ sky130_fd_sc_hd__buf_1
XFILLER_0_106_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1492_ Tile_X0Y1_DSP_bot.Inst_MULADD._0644_ Tile_X0Y1_DSP_bot.Inst_MULADD._0645_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0657_ Tile_X0Y1_DSP_bot.Inst_MULADD._0658_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0659_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3 net254 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[163\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[344\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_117_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_37 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_15 Tile_X0Y0_DSP_top.FrameStrobe\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID6 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_26 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG2 VGND VGND VPWR
+ VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_59 Tile_X0Y0_DSP_top.N4BEG\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_144_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1759_ net333 Tile_X0Y1_DSP_bot.C17 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[17\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.S4END_inbuf_5._0_ net116 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[5\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[19\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[8\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_150_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_050_ Tile_X0Y0_DSP_top.FrameData_O\[2\] VGND VGND VPWR VPWR net452 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst1
+ net82 net84 net90 net134 Tile_X0Y0_DSP_top.ConfigBits\[358\] Tile_X0Y0_DSP_top.ConfigBits\[359\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_103_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG3 net285
+ net220 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb0 net338 Tile_X0Y1_DSP_bot.ConfigBits\[238\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[239\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG3
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.strobe_inbuf_5._0_ net276 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0992_ Tile_X0Y1_DSP_bot.Inst_MULADD._0135_ Tile_X0Y1_DSP_bot.Inst_MULADD._0159_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0165_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0166_
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_158_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.W6END_inbuf_9._0_ net155 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1613_ Tile_X0Y1_DSP_bot.C15 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[15\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0776_
+ sky130_fd_sc_hd__mux2_1
X_317_ Tile_X0Y1_DSP_bot.SS4BEG\[1\] VGND VGND VPWR VPWR net706 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 Tile_X0Y0_E2MID[0] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
XFILLER_0_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput35 Tile_X0Y0_EE4END[11] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
Xinput24 Tile_X0Y0_E6END[1] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_4
Xinput46 Tile_X0Y0_EE4END[7] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_114_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1544_ Tile_X0Y1_DSP_bot.Inst_MULADD._0706_ Tile_X0Y1_DSP_bot.Inst_MULADD._0707_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0709_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0710_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_248_ Tile_X0Y1_DSP_bot.FrameData_O\[0\] VGND VGND VPWR VPWR net631 sky130_fd_sc_hd__clkbuf_1
Xinput68 Tile_X0Y0_FrameData[27] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_8
Xinput57 Tile_X0Y0_FrameData[17] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_8
Xinput79 Tile_X0Y0_FrameData[8] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_4
X_179_ Tile_X0Y0_DSP_top.W6BEG\[7\] VGND VGND VPWR VPWR net564 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1475_ Tile_X0Y1_DSP_bot.Inst_MULADD._0623_ Tile_X0Y1_DSP_bot.Inst_MULADD._0625_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0641_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0642_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[30\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.NN4END_inbuf_10._0_ Tile_X0Y0_DSP_top.NN4END\[14\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.S4END_inbuf_5._0_ Tile_X0Y0_DSP_top.S4BEG\[9\] VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.S4BEG_i\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END7
+ net4 net12 Tile_X0Y0_DSP_top.ConfigBits\[270\] Tile_X0Y0_DSP_top.ConfigBits\[271\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[126\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4 net255 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[4\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_102_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 VGND VGND VPWR VPWR net484
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_033_ Tile_X0Y0_DSP_top.EE4BEG\[1\] VGND VGND VPWR VPWR net421 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1260_ Tile_X0Y1_DSP_bot.Inst_MULADD._0405_ Tile_X0Y1_DSP_bot.Inst_MULADD._0393_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0394_ Tile_X0Y1_DSP_bot.Inst_MULADD._0398_ Tile_X0Y1_DSP_bot.Inst_MULADD._0395_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0430_ sky130_fd_sc_hd__o311a_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1191_ Tile_X0Y1_DSP_bot.Inst_MULADD._0142_ Tile_X0Y1_DSP_bot.Inst_MULADD._0143_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0188_ Tile_X0Y1_DSP_bot.Inst_MULADD._0358_ Tile_X0Y1_DSP_bot.Inst_MULADD._0360_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0362_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_135_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0975_ Tile_X0Y1_DSP_bot.Inst_MULADD._0064_ Tile_X0Y1_DSP_bot.Inst_MULADD._0065_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0070_ Tile_X0Y1_DSP_bot.Inst_MULADD._0109_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0149_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_139_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6 net257 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[262\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.W6END_inbuf_9._0_ net356 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1527_ Tile_X0Y1_DSP_bot.Inst_MULADD._0674_ Tile_X0Y1_DSP_bot.Inst_MULADD._0672_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0671_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0693_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1458_ Tile_X0Y1_DSP_bot.Inst_MULADD._0625_ Tile_X0Y1_DSP_bot.Inst_MULADD._0623_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0626_ sky130_fd_sc_hd__nand2_2
XTile_X0Y1_DSP_bot.S4END_inbuf_10._0_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG2
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.S4BEG_i\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb0 net334 Tile_X0Y1_DSP_bot.ConfigBits\[380\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[381\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1389_ Tile_X0Y1_DSP_bot.Inst_MULADD._0487_ Tile_X0Y1_DSP_bot.Inst_MULADD._0466_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0476_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0558_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[50\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[39\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_141_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst1
+ net89 net101 net141 net173 Tile_X0Y0_DSP_top.ConfigBits\[322\] Tile_X0Y0_DSP_top.ConfigBits\[323\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[103\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.strobe_inbuf_1._0_ Tile_X0Y0_DSP_top.FrameStrobe\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[1\] sky130_fd_sc_hd__clkbuf_1
Xinput214 Tile_X0Y1_EE4END[10] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
Xinput225 Tile_X0Y1_EE4END[6] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
Xinput203 Tile_X0Y1_E6END[11] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
Xinput236 Tile_X0Y1_FrameData[16] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__buf_4
Xinput269 Tile_X0Y1_FrameStrobe[17] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__clkbuf_1
Xinput258 Tile_X0Y1_FrameData[7] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__buf_6
Xinput247 Tile_X0Y1_FrameData[26] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_155_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_121_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_016_ Tile_X0Y0_DSP_top.E2BEGb\[4\] VGND VGND VPWR VPWR net398 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1312_ Tile_X0Y1_DSP_bot.Inst_MULADD._0479_ Tile_X0Y1_DSP_bot.Inst_MULADD._0480_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0464_ Tile_X0Y1_DSP_bot.Inst_MULADD._0481_ Tile_X0Y1_DSP_bot.Inst_MULADD._0467_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0482_ sky130_fd_sc_hd__o221ai_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1243_ Tile_X0Y1_DSP_bot.Inst_MULADD._0400_ Tile_X0Y1_DSP_bot.Inst_MULADD._0392_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0399_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0414_
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1174_ Tile_X0Y1_DSP_bot.Inst_MULADD._0283_ Tile_X0Y1_DSP_bot.Inst_MULADD._0343_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0344_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0345_
+ sky130_fd_sc_hd__a21oi_4
XFILLER_0_159_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0958_ Tile_X0Y1_DSP_bot.Inst_MULADD._0067_ Tile_X0Y1_DSP_bot.B3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0132_ sky130_fd_sc_hd__or2b_2
XFILLER_0_146_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0889_ Tile_X0Y1_DSP_bot.Inst_MULADD._0025_ Tile_X0Y1_DSP_bot.Inst_MULADD._0038_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0065_ sky130_fd_sc_hd__nor2_4
XFILLER_0_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[246\] Tile_X0Y0_DSP_top.ConfigBits\[247\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._31_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID7
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 sky130_fd_sc_hd__clkbuf_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.SS4END_inbuf_0._0_ Tile_X0Y0_DSP_top.SS4BEG\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[0\] sky130_fd_sc_hd__buf_4
XFILLER_0_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[77\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1 sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_156_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_156_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG1.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[358\] Tile_X0Y1_DSP_bot.ConfigBits\[359\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_73_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27 net68 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[81\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16 net56 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[70\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9 net260 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[361\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_81_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput518 net518 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput507 net507 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_0_1_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput529 net529 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[5] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._93_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q17
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 sky130_fd_sc_hd__buf_12
XFILLER_0_157_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1226_ Tile_X0Y1_DSP_bot.A0 Tile_X0Y1_DSP_bot.Inst_MULADD._0025_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0027_ Tile_X0Y1_DSP_bot.Inst_MULADD._0347_ Tile_X0Y1_DSP_bot.Inst_MULADD._0349_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0397_ sky130_fd_sc_hd__o2111ai_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[286\] Tile_X0Y0_DSP_top.ConfigBits\[287\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1157_ Tile_X0Y1_DSP_bot.Inst_MULADD._0223_ Tile_X0Y1_DSP_bot.Inst_MULADD._0250_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0327_ Tile_X0Y1_DSP_bot.Inst_MULADD._0328_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0329_ sky130_fd_sc_hd__a2bb2oi_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb7
+ net335 net337 Tile_X0Y1_DSP_bot.ConfigBits\[344\] Tile_X0Y1_DSP_bot.ConfigBits\[345\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1088_ Tile_X0Y1_DSP_bot.Inst_MULADD._0026_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0260_ sky130_fd_sc_hd__and2_1
XFILLER_0_106_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_159_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[246\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.data_outbuf_5._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[60\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._14_ net19 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEGb\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA_116 Tile_X0Y1_DSP_bot.SS4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 Tile_X0Y1_DSP_bot.S4BEG\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_127 Tile_X0Y1_DSP_bot.SS4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_149 net291 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_350_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb6 VGND VGND VPWR VPWR net733
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_281_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG1 VGND VGND VPWR VPWR net664
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_10._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.NN4END\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[109\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top.data_inbuf_29._0_ net70 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[29\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.WW4END_inbuf_7._0_ net167 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[268\] Tile_X0Y1_DSP_bot.ConfigBits\[269\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_S4BEG0 net204 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb2
+ Tile_X0Y0_DSP_top.S4BEG\[1\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.ConfigBits\[70\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[71\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1011_ Tile_X0Y1_DSP_bot.Inst_MULADD._0135_ Tile_X0Y1_DSP_bot.Inst_MULADD._0159_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0165_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0184_
+ sky130_fd_sc_hd__and3_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_156_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_E1BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG3 Tile_X0Y0_DSP_top.ConfigBits\[32\]
+ Tile_X0Y0_DSP_top.ConfigBits\[33\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E1BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG0.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[56\] Tile_X0Y1_DSP_bot.ConfigBits\[57\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG\[10\] sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._76_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG6 sky130_fd_sc_hd__buf_1
XFILLER_0_77_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1209_ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0380_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20 net241 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[116\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31 net253 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[127\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_130_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.data_outbuf_5._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[5\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.strobe_outbuf_10._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[10\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[10\] sky130_fd_sc_hd__buf_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_S1BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG0 Tile_X0Y1_DSP_bot.ConfigBits\[68\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[69\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[308\] Tile_X0Y1_DSP_bot.ConfigBits\[309\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_333_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net716
+ sky130_fd_sc_hd__clkbuf_1
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_153_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1560_ Tile_X0Y1_DSP_bot.Inst_MULADD._0692_ Tile_X0Y1_DSP_bot.Inst_MULADD._0695_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0713_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0725_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_264_ Tile_X0Y1_DSP_bot.FrameData_O\[16\] VGND VGND VPWR VPWR net638 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG0.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[322\] Tile_X0Y1_DSP_bot.ConfigBits\[323\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_24_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_195_ Tile_X0Y0_DSP_top.WW4BEG\[11\] VGND VGND VPWR VPWR net569 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1491_ Tile_X0Y1_DSP_bot.Inst_MULADD._0656_ Tile_X0Y1_DSP_bot.Inst_MULADD._0652_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0137_ Tile_X0Y1_DSP_bot.Inst_MULADD._0351_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0658_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG7
+ Tile_X0Y0_DSP_top.ConfigBits\[147\] Tile_X0Y0_DSP_top.ConfigBits\[148\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[83\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG1 sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot.E6BEG_outbuf_3._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.data_inbuf_29._0_ net250 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[29\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_129_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4 net255 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[164\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[345\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_117_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_38 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA_16 Tile_X0Y0_DSP_top.FrameStrobe\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1758_ net333 Tile_X0Y1_DSP_bot.C16 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[16\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_49 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1689_ Tile_X0Y1_DSP_bot.Inst_MULADD._0837_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0009_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.strobe_outbuf_6._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[6\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._59_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[12\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[9\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame12_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[358\] Tile_X0Y0_DSP_top.ConfigBits\[359\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_5_191 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput690 net690 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0991_ Tile_X0Y1_DSP_bot.Inst_MULADD._0160_ Tile_X0Y1_DSP_bot.Inst_MULADD._0163_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0164_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0165_
+ sky130_fd_sc_hd__o21ai_4
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1612_ Tile_X0Y1_DSP_bot.Inst_MULADD._0351_ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0774_ Tile_X0Y1_DSP_bot.Inst_MULADD._0755_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ sky130_fd_sc_hd__o31ai_4
X_316_ Tile_X0Y1_DSP_bot.SS4BEG\[0\] VGND VGND VPWR VPWR net699 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_141_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput25 Tile_X0Y0_E6END[2] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput36 Tile_X0Y0_EE4END[12] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput14 Tile_X0Y0_E2MID[1] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1543_ Tile_X0Y1_DSP_bot.Inst_MULADD._0669_ Tile_X0Y1_DSP_bot.Inst_MULADD._0708_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0663_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0709_
+ sky130_fd_sc_hd__o21a_1
X_247_ Tile_X0Y1_DSP_bot.EE4BEG\[15\] VGND VGND VPWR VPWR net621 sky130_fd_sc_hd__clkbuf_1
Xinput69 Tile_X0Y0_FrameData[28] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_8
Xinput58 Tile_X0Y0_FrameData[18] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_8
XTile_X0Y0_DSP_top.EE4BEG_outbuf_11._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG\[11\] sky130_fd_sc_hd__clkbuf_1
Xinput47 Tile_X0Y0_EE4END[8] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_1
X_178_ Tile_X0Y0_DSP_top.W6BEG\[6\] VGND VGND VPWR VPWR net563 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1474_ Tile_X0Y1_DSP_bot.Inst_MULADD._0570_ Tile_X0Y1_DSP_bot.Inst_MULADD._0616_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0617_ Tile_X0Y1_DSP_bot.Inst_MULADD._0640_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0641_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_12_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30 net252 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[158\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.WW4BEG_outbuf_4._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[4\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[4\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG2.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_74_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.E6END_inbuf_1._0_ net26 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_59_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_130_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst1
+ net84 net92 net134 net136 Tile_X0Y0_DSP_top.ConfigBits\[270\] Tile_X0Y0_DSP_top.ConfigBits\[271\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[127\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5 net256 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[5\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.strobe_inbuf_14._0_ net266 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[14\]
+ sky130_fd_sc_hd__clkbuf_1
X_101_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1 VGND VGND VPWR VPWR net483
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.cus_mux41_buf_inst0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG6
+ Tile_X0Y1_DSP_bot.ConfigBits\[150\] Tile_X0Y1_DSP_bot.ConfigBits\[151\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_46_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_032_ Tile_X0Y0_DSP_top.EE4BEG\[0\] VGND VGND VPWR VPWR net414 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1190_ Tile_X0Y1_DSP_bot.Inst_MULADD._0080_ Tile_X0Y1_DSP_bot.Inst_MULADD._0192_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0358_ Tile_X0Y1_DSP_bot.Inst_MULADD._0360_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0361_ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.SS4END_inbuf_9._0_ net121 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0974_ Tile_X0Y1_DSP_bot.Inst_MULADD._0138_ Tile_X0Y1_DSP_bot.Inst_MULADD._0145_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0147_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0148_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7 net258 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[263\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_44_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1526_ Tile_X0Y1_DSP_bot.Inst_MULADD._0435_ Tile_X0Y1_DSP_bot.Inst_MULADD._0519_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0586_ Tile_X0Y1_DSP_bot.Inst_MULADD._0691_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0692_ sky130_fd_sc_hd__nand4_4
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1457_ Tile_X0Y1_DSP_bot.Inst_MULADD._0435_ Tile_X0Y1_DSP_bot.Inst_MULADD._0519_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0586_ Tile_X0Y1_DSP_bot.Inst_MULADD._0591_ Tile_X0Y1_DSP_bot.Inst_MULADD._0573_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0625_ sky130_fd_sc_hd__a32oi_4
XFILLER_0_12_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1388_ Tile_X0Y1_DSP_bot.Inst_MULADD._0534_ Tile_X0Y1_DSP_bot.Inst_MULADD._0549_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0556_ Tile_X0Y1_DSP_bot.Inst_MULADD._0461_ Tile_X0Y1_DSP_bot.Inst_MULADD._0488_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0557_ sky130_fd_sc_hd__o2111ai_4
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[380\] Tile_X0Y1_DSP_bot.ConfigBits\[381\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[40\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[51\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.E6END_inbuf_1._0_ net206 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_90_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[322\] Tile_X0Y0_DSP_top.ConfigBits\[323\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput226 Tile_X0Y1_EE4END[7] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
Xinput215 Tile_X0Y1_EE4END[11] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
Xinput204 Tile_X0Y1_E6END[1] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__buf_4
Xinput259 Tile_X0Y1_FrameData[8] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__buf_6
Xinput237 Tile_X0Y1_FrameData[17] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_4
Xinput248 Tile_X0Y1_FrameData[27] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_128_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_015_ Tile_X0Y0_DSP_top.E2BEGb\[3\] VGND VGND VPWR VPWR net397 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1311_ Tile_X0Y1_DSP_bot.Inst_MULADD._0443_ Tile_X0Y1_DSP_bot.Inst_MULADD._0454_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0460_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0481_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_39_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1242_ Tile_X0Y1_DSP_bot.Inst_MULADD._0407_ Tile_X0Y1_DSP_bot.Inst_MULADD._0396_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0406_ Tile_X0Y1_DSP_bot.Inst_MULADD._0412_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0413_ sky130_fd_sc_hd__a22oi_4
XTile_X0Y0_DSP_top.EE4END_inbuf_8._0_ net36 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1173_ Tile_X0Y1_DSP_bot.Inst_MULADD._0064_ Tile_X0Y1_DSP_bot.Inst_MULADD._0065_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0344_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_76_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0957_ Tile_X0Y1_DSP_bot.Inst_MULADD._0131_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 sky130_fd_sc_hd__buf_12
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0888_ Tile_X0Y1_DSP_bot.Inst_MULADD._0025_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0064_ sky130_fd_sc_hd__and2_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG0.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[248\] Tile_X0Y0_DSP_top.ConfigBits\[249\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG0 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1509_ Tile_X0Y1_DSP_bot.Inst_MULADD._0670_ Tile_X0Y1_DSP_bot.Inst_MULADD._0673_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0675_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0676_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._30_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID6
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 sky130_fd_sc_hd__clkbuf_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.N4BEG_outbuf_7._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4END\[7\] sky130_fd_sc_hd__clkbuf_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_145_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[77\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28 net69 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[82\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17 net57 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[71\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput508 net508 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[15] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._92_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q16
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 sky130_fd_sc_hd__buf_12
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput519 net519 VGND VGND VPWR VPWR Tile_X0Y0_NN4BEG[10] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1225_ Tile_X0Y1_DSP_bot.Inst_MULADD._0390_ Tile_X0Y1_DSP_bot.Inst_MULADD._0389_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0378_ Tile_X0Y1_DSP_bot.Inst_MULADD._0387_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0396_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_157_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[286\] Tile_X0Y0_DSP_top.ConfigBits\[287\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1156_ Tile_X0Y1_DSP_bot.Inst_MULADD._0286_ Tile_X0Y1_DSP_bot.Inst_MULADD._0292_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0304_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0328_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[344\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[345\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1087_ Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0188_ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0259_ sky130_fd_sc_hd__nand4_4
XFILLER_0_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[247\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.strobe_outbuf_18._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[18\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.data_inbuf_9._0_ net80 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.W6BEG_outbuf_7._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[7\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[61\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._13_ net18 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEGb\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 Tile_X0Y1_DSP_bot.S4BEG\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 Tile_X0Y1_DSP_bot.SS4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 Tile_X0Y1_DSP_bot.SS4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S1BEG0 VGND VGND VPWR VPWR net663
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.N4END_inbuf_5._0_ Tile_X0Y0_DSP_top.N4END\[9\] VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_i\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG3.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_121_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG3.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[270\] Tile_X0Y1_DSP_bot.ConfigBits\[271\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG3 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_S4BEG1 net201 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb3
+ Tile_X0Y0_DSP_top.S4BEG\[2\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1 Tile_X0Y1_DSP_bot.ConfigBits\[72\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[73\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1010_ Tile_X0Y1_DSP_bot.Inst_MULADD._0178_ Tile_X0Y1_DSP_bot.Inst_MULADD._0174_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0176_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0183_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_E1BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG0 Tile_X0Y0_DSP_top.ConfigBits\[34\]
+ Tile_X0Y0_DSP_top.ConfigBits\[35\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E1BEG\[3\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_124_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.NN4END_inbuf_0._0_ net327 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[0\]
+ sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._75_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG5 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1208_ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0379_ sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1139_ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0215_ Tile_X0Y1_DSP_bot.Inst_MULADD._0205_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0311_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10 net230 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[106\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.N4BEG_outbuf_3._0_ Tile_X0Y0_DSP_top.N4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21 net242 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[117\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.NN4BEG_outbuf_7._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[7\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_130_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_158_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.ConfigBits\[308\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[309\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_332_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net715
+ sky130_fd_sc_hd__clkbuf_1
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.data_outbuf_27._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[27\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[27\] sky130_fd_sc_hd__clkbuf_1
X_263_ Tile_X0Y1_DSP_bot.FrameData_O\[15\] VGND VGND VPWR VPWR net637 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1490_ Tile_X0Y1_DSP_bot.Inst_MULADD._0269_ Tile_X0Y1_DSP_bot.Inst_MULADD._0270_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0652_ Tile_X0Y1_DSP_bot.Inst_MULADD._0347_ Tile_X0Y1_DSP_bot.Inst_MULADD._0656_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0657_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_24_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_194_ Tile_X0Y0_DSP_top.WW4BEG\[10\] VGND VGND VPWR VPWR net568 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[83\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG7
+ Tile_X0Y0_DSP_top.ConfigBits\[147\] Tile_X0Y0_DSP_top.ConfigBits\[148\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.N4END_inbuf_5._0_ net316 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_121_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_0._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END0 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5 net256 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[165\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[346\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_86_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.data_outbuf_18._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[18\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[18\] sky130_fd_sc_hd__clkbuf_1
XANTENNA_17 Tile_X0Y0_DSP_top.FrameStrobe\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_117_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_39 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1757_ net333 Tile_X0Y1_DSP_bot.C15 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[15\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1688_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0584_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0837_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_3._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.S4BEG_outbuf_7._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[7\] sky130_fd_sc_hd__buf_2
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.W6BEG_outbuf_3._0_ Tile_X0Y0_DSP_top.W6BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._58_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_135_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_116_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[358\] Tile_X0Y0_DSP_top.ConfigBits\[359\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_21_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput680 net680 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput691 net691 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0990_ Tile_X0Y1_DSP_bot.Inst_MULADD._0157_ Tile_X0Y1_DSP_bot.Inst_MULADD._0153_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0164_ sky130_fd_sc_hd__nand2_2
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1611_ Tile_X0Y1_DSP_bot.Inst_MULADD._0273_ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0701_ Tile_X0Y1_DSP_bot.Inst_MULADD._0728_ Tile_X0Y1_DSP_bot.Inst_MULADD._0730_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0774_ sky130_fd_sc_hd__o221a_2
X_315_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 VGND VGND VPWR VPWR net689
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_141_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput26 Tile_X0Y0_E6END[3] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput37 Tile_X0Y0_EE4END[13] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput15 Tile_X0Y0_E2MID[2] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1542_ Tile_X0Y1_DSP_bot.Inst_MULADD._0664_ Tile_X0Y1_DSP_bot.Inst_MULADD._0665_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0666_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0708_
+ sky130_fd_sc_hd__o21a_1
X_246_ Tile_X0Y1_DSP_bot.EE4BEG\[14\] VGND VGND VPWR VPWR net620 sky130_fd_sc_hd__clkbuf_1
Xinput59 Tile_X0Y0_FrameData[19] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_6
Xinput48 Tile_X0Y0_EE4END[9] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_177_ Tile_X0Y0_DSP_top.W6BEG\[5\] VGND VGND VPWR VPWR net562 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1473_ Tile_X0Y1_DSP_bot.Inst_MULADD._0611_ Tile_X0Y1_DSP_bot.Inst_MULADD._0612_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0613_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0640_
+ sky130_fd_sc_hd__a21bo_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31 net253 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[159\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20 net241 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[148\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_149_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_319 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_inst0
+ net284 net184 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[45\] Tile_X0Y1_DSP_bot.ConfigBits\[46\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[270\] Tile_X0Y0_DSP_top.ConfigBits\[271\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_inbuf_2._0_ net251 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6 net257 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[6\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_100_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0 VGND VGND VPWR VPWR net482
+ sky130_fd_sc_hd__buf_1
XFILLER_0_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG6
+ Tile_X0Y1_DSP_bot.ConfigBits\[150\] Tile_X0Y1_DSP_bot.ConfigBits\[151\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C8.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.data_outbuf_23._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[23\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[23\] sky130_fd_sc_hd__clkbuf_1
X_031_ Tile_X0Y0_DSP_top.E6BEG\[11\] VGND VGND VPWR VPWR net404 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0973_ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0138_ Tile_X0Y1_DSP_bot.Inst_MULADD._0146_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0147_ sky130_fd_sc_hd__a22oi_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8 net259 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[264\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.data_outbuf_14._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[14\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1525_ Tile_X0Y1_DSP_bot.Inst_MULADD._0670_ Tile_X0Y1_DSP_bot.Inst_MULADD._0673_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0675_ Tile_X0Y1_DSP_bot.Inst_MULADD._0641_ Tile_X0Y1_DSP_bot.Inst_MULADD._0622_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0691_ sky130_fd_sc_hd__o2111a_2
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_229_ Tile_X0Y1_DSP_bot.E6BEG\[9\] VGND VGND VPWR VPWR net614 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1456_ Tile_X0Y1_DSP_bot.Inst_MULADD._0587_ Tile_X0Y1_DSP_bot.Inst_MULADD._0592_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0623_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0624_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_69_79 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1387_ Tile_X0Y1_DSP_bot.Inst_MULADD._0551_ Tile_X0Y1_DSP_bot.Inst_MULADD._0534_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0555_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0556_
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y0_DSP_top.S4BEG_outbuf_3._0_ Tile_X0Y0_DSP_top.S4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.ConfigBits\[380\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[381\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[11\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[41\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame11_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.WW4END_inbuf_10._0_ net170 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[10\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[322\] Tile_X0Y0_DSP_top.ConfigBits\[323\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.N4BEG_outbuf_11._0_ Tile_X0Y0_DSP_top.N4BEG_i\[11\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[11\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput227 Tile_X0Y1_EE4END[8] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
Xinput216 Tile_X0Y1_EE4END[12] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
Xinput205 Tile_X0Y1_E6END[2] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__clkbuf_1
Xinput238 Tile_X0Y1_FrameData[18] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_8
Xinput249 Tile_X0Y1_FrameData[28] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__buf_6
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30 net252 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[190\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_014_ Tile_X0Y0_DSP_top.E2BEGb\[2\] VGND VGND VPWR VPWR net396 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1310_ Tile_X0Y1_DSP_bot.Inst_MULADD._0472_ Tile_X0Y1_DSP_bot.Inst_MULADD._0478_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0473_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0480_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_151_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1241_ Tile_X0Y1_DSP_bot.Inst_MULADD._0395_ Tile_X0Y1_DSP_bot.Inst_MULADD._0396_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0412_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1172_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B5
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_ Tile_X0Y1_DSP_bot.Inst_MULADD._0208_ Tile_X0Y1_DSP_bot.Inst_MULADD._0282_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0343_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_159_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0956_ Tile_X0Y1_DSP_bot.Inst_MULADD._0130_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[3\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0131_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0887_ Tile_X0Y1_DSP_bot.Inst_MULADD._0025_ Tile_X0Y1_DSP_bot.Inst_MULADD._0061_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0062_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0063_
+ sky130_fd_sc_hd__o21a_2
XFILLER_0_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1508_ Tile_X0Y1_DSP_bot.Inst_MULADD._0674_ Tile_X0Y1_DSP_bot.Inst_MULADD._0672_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0671_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0675_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1439_ Tile_X0Y1_DSP_bot.Inst_MULADD._0597_ Tile_X0Y1_DSP_bot.Inst_MULADD._0598_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0604_ Tile_X0Y1_DSP_bot.Inst_MULADD._0606_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0607_ sky130_fd_sc_hd__nand4_4
XFILLER_0_110_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.NN4END_inbuf_9._0_ Tile_X0Y0_DSP_top.NN4END\[13\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_118_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_39_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18 net58 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[72\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29 net70 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[83\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput509 net509 VGND VGND VPWR VPWR Tile_X0Y0_N4BEG[1] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._91_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q15
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 sky130_fd_sc_hd__buf_12
XFILLER_0_34_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_151_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1224_ Tile_X0Y1_DSP_bot.Inst_MULADD._0393_ Tile_X0Y1_DSP_bot.Inst_MULADD._0394_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0387_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0395_
+ sky130_fd_sc_hd__o21bai_4
XFILLER_0_157_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG2.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[288\] Tile_X0Y0_DSP_top.ConfigBits\[289\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG2 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1155_ Tile_X0Y1_DSP_bot.Inst_MULADD._0298_ Tile_X0Y1_DSP_bot.Inst_MULADD._0301_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0327_ sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.ConfigBits\[344\] Tile_X0Y1_DSP_bot.ConfigBits\[345\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1086_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.Inst_MULADD._0256_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0257_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0258_
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst0
+ net284 net286 net308 net220 Tile_X0Y1_DSP_bot.ConfigBits\[288\] Tile_X0Y1_DSP_bot.ConfigBits\[289\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[248\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0939_ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0114_ sky130_fd_sc_hd__nand4_4
XFILLER_0_122_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_3._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[62\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._12_ net17 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEGb\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 Tile_X0Y1_DSP_bot.SS4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 Tile_X0Y1_DSP_bot.SS4BEG_i\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 Tile_X0Y1_DSP_bot.SS4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0 net229 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[384\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_S4BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb0
+ Tile_X0Y0_DSP_top.S4BEG\[3\] net357 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.ConfigBits\[74\] Tile_X0Y1_DSP_bot.ConfigBits\[75\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_124_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_124_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._74_ net342 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG4
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1207_ Tile_X0Y1_DSP_bot.Inst_MULADD._0365_ Tile_X0Y1_DSP_bot.Inst_MULADD._0371_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0377_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0378_
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1138_ Tile_X0Y1_DSP_bot.Inst_MULADD._0298_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0310_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1069_ Tile_X0Y1_DSP_bot.C5 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[5\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0242_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11 net231 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[107\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22 net243 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[118\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_89_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.S4END_inbuf_8._0_ net104 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.WW4END_inbuf_1._0_ net377 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG5.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[310\] Tile_X0Y1_DSP_bot.ConfigBits\[311\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG5 sky130_fd_sc_hd__mux4_2
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_331_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG3 VGND VGND VPWR VPWR net705
+ sky130_fd_sc_hd__clkbuf_1
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_262_ Tile_X0Y1_DSP_bot.FrameData_O\[14\] VGND VGND VPWR VPWR net636 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[149\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.X
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_134_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_193_ Tile_X0Y0_DSP_top.WW4BEG\[9\] VGND VGND VPWR VPWR net582 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG1.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.strobe_inbuf_8._0_ net279 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[8\]
+ sky130_fd_sc_hd__buf_1
XFILLER_0_121_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6 net257 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[166\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XANTENNA_29 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2 VGND VGND
+ VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[347\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1756_ net333 Tile_X0Y1_DSP_bot.C14 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[14\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_18 Tile_X0Y0_DSP_top.FrameStrobe\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1687_ Tile_X0Y1_DSP_bot.Inst_MULADD._0836_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0008_ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._57_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG3
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG4.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[360\] Tile_X0Y0_DSP_top.ConfigBits\[361\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG4 sky130_fd_sc_hd__mux4_2
XFILLER_0_131_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.S4END_inbuf_8._0_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S4BEG0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.S4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst0
+ net282 net288 net188 net204 Tile_X0Y1_DSP_bot.ConfigBits\[360\] Tile_X0Y1_DSP_bot.ConfigBits\[361\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
Xoutput681 net681 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput670 net670 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[3] sky130_fd_sc_hd__buf_2
Xoutput692 net692 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[3] sky130_fd_sc_hd__clkbuf_4
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG2 VGND VGND VPWR VPWR net688
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1610_ Tile_X0Y1_DSP_bot.Inst_MULADD._0772_ Tile_X0Y1_DSP_bot.Inst_MULADD._0773_
+ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\] Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q14 sky130_fd_sc_hd__a2bb2o_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1541_ Tile_X0Y1_DSP_bot.Inst_MULADD._0705_ Tile_X0Y1_DSP_bot.Inst_MULADD._0702_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0703_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0707_
+ sky130_fd_sc_hd__nor3_2
X_245_ Tile_X0Y1_DSP_bot.EE4BEG\[13\] VGND VGND VPWR VPWR net619 sky130_fd_sc_hd__clkbuf_1
Xinput27 Tile_X0Y0_E6END[4] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput16 Tile_X0Y0_E2MID[3] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_0_116_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput49 Tile_X0Y0_FrameData[0] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_8
Xinput38 Tile_X0Y0_EE4END[14] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
X_176_ Tile_X0Y0_DSP_top.W6BEG\[4\] VGND VGND VPWR VPWR net561 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1472_ Tile_X0Y1_DSP_bot.Inst_MULADD._0516_ Tile_X0Y1_DSP_bot.Inst_MULADD._0581_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0633_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0639_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10 net230 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[138\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21 net242 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[149\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1739_ net333 Tile_X0Y1_DSP_bot.B5 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_132_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_140_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG0
+ Tile_X0Y1_DSP_bot.ConfigBits\[45\] Tile_X0Y1_DSP_bot.ConfigBits\[46\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[270\] Tile_X0Y0_DSP_top.ConfigBits\[271\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_155_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7 net258 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[7\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_148_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_030_ Tile_X0Y0_DSP_top.E6BEG\[10\] VGND VGND VPWR VPWR net403 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_inst0
+ net282 net182 net335 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.ConfigBits\[31\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[32\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_73_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.strobe_inbuf_4._0_ Tile_X0Y0_DSP_top.FrameStrobe\[4\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst0
+ net183 net336 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.ConfigBits\[58\] Tile_X0Y1_DSP_bot.ConfigBits\[59\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.data_inbuf_10._0_ net50 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[10\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0972_ Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_ Tile_X0Y1_DSP_bot.Inst_MULADD._0141_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0146_ sky130_fd_sc_hd__nand4_4
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9 net260 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[265\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_154_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_154_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1524_ Tile_X0Y1_DSP_bot.Inst_MULADD._0632_ Tile_X0Y1_DSP_bot.Inst_MULADD._0634_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0689_ Tile_X0Y1_DSP_bot.Inst_MULADD._0683_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0690_ sky130_fd_sc_hd__a31oi_2
X_228_ Tile_X0Y1_DSP_bot.E6BEG\[8\] VGND VGND VPWR VPWR net613 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_159_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG3 VGND VGND VPWR VPWR net542
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1455_ Tile_X0Y1_DSP_bot.Inst_MULADD._0614_ Tile_X0Y1_DSP_bot.Inst_MULADD._0618_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0622_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0623_
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1386_ Tile_X0Y1_DSP_bot.Inst_MULADD._0552_ Tile_X0Y1_DSP_bot.Inst_MULADD._0554_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0555_ sky130_fd_sc_hd__nor2_2
XFILLER_0_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG7.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[382\] Tile_X0Y1_DSP_bot.ConfigBits\[383\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG7 sky130_fd_sc_hd__mux4_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_149_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_125_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[150\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_113_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG3.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[324\] Tile_X0Y0_DSP_top.ConfigBits\[325\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_11_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst0
+ net325 net181 net221 net201 Tile_X0Y1_DSP_bot.ConfigBits\[324\] Tile_X0Y1_DSP_bot.ConfigBits\[325\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
Xinput206 Tile_X0Y1_E6END[3] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__clkbuf_1
Xinput217 Tile_X0Y1_EE4END[13] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
Xinput228 Tile_X0Y1_EE4END[9] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
Xinput239 Tile_X0Y1_FrameData[19] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_8
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20 net241 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[180\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31 net253 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[191\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.SS4END_inbuf_3._0_ Tile_X0Y0_DSP_top.SS4BEG\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[3\] sky130_fd_sc_hd__clkbuf_4
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_013_ Tile_X0Y0_DSP_top.E2BEGb\[1\] VGND VGND VPWR VPWR net395 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1240_ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0297_ Tile_X0Y1_DSP_bot.Inst_MULADD._0401_ Tile_X0Y1_DSP_bot.Inst_MULADD._0410_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0411_ sky130_fd_sc_hd__o32ai_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID7
+ net20 net100 net152 Tile_X0Y0_DSP_top.ConfigBits\[198\] Tile_X0Y0_DSP_top.ConfigBits\[199\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG0
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1171_ Tile_X0Y1_DSP_bot.Inst_MULADD._0184_ Tile_X0Y1_DSP_bot.Inst_MULADD._0185_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0326_ Tile_X0Y1_DSP_bot.Inst_MULADD._0330_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0342_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_57_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.data_inbuf_10._0_ net230 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[10\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0955_ Tile_X0Y1_DSP_bot.Inst_MULADD._0128_ Tile_X0Y1_DSP_bot.Inst_MULADD._0129_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0130_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0886_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[2\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0062_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END3
+ net33 net110 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.ConfigBits\[398\]
+ Tile_X0Y0_DSP_top.ConfigBits\[399\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1507_ Tile_X0Y1_DSP_bot.Inst_MULADD._0663_ Tile_X0Y1_DSP_bot.Inst_MULADD._0667_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0669_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0674_
+ sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1438_ Tile_X0Y1_DSP_bot.Inst_MULADD._0605_ Tile_X0Y1_DSP_bot.Inst_MULADD._0533_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0603_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0606_
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1369_ Tile_X0Y1_DSP_bot.Inst_MULADD._0530_ Tile_X0Y1_DSP_bot.Inst_MULADD._0531_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0538_ sky130_fd_sc_hd__nand2_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.data_outbuf_8._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[8\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_133_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.EE4END_inbuf_2._0_ net225 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_156_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_136_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.strobe_inbuf_11._0_ Tile_X0Y0_DSP_top.FrameStrobe\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[11\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19 net59 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[73\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_151_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._90_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q14
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 sky130_fd_sc_hd__buf_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1223_ Tile_X0Y1_DSP_bot.Inst_MULADD._0381_ Tile_X0Y1_DSP_bot.Inst_MULADD._0382_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0383_ Tile_X0Y1_DSP_bot.Inst_MULADD._0365_ Tile_X0Y1_DSP_bot.Inst_MULADD._0371_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0394_ sky130_fd_sc_hd__o2111a_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1154_ Tile_X0Y1_DSP_bot.Inst_MULADD._0239_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0326_ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG6.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[346\] Tile_X0Y1_DSP_bot.ConfigBits\[347\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG6 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1085_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0257_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst1
+ net204 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb1 net339 net357 Tile_X0Y1_DSP_bot.ConfigBits\[288\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[289\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_159_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_159_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[249\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 net84 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[95\] Tile_X0Y0_DSP_top.ConfigBits\[96\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0938_ Tile_X0Y1_DSP_bot.Inst_MULADD._0112_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0113_ sky130_fd_sc_hd__buf_6
XFILLER_0_122_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_122_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._0869_ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0029_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0046_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_142_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30 net252 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[222\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[10\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[63\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame10_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._11_ net16 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEGb\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_119 Tile_X0Y1_DSP_bot.SS4BEG_i\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_108 Tile_X0Y1_DSP_bot.SS4BEG\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.data_outbuf_8._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[8\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1 net240 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[385\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_133_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_121_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.strobe_outbuf_13._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[13\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[13\] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_S4BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb1
+ Tile_X0Y0_DSP_top.S4BEG\[0\] net354 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[76\] Tile_X0Y1_DSP_bot.ConfigBits\[77\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_129_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_124_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.E6BEG_outbuf_6._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._73_ net341 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG3
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1206_ Tile_X0Y1_DSP_bot.Inst_MULADD._0373_ Tile_X0Y1_DSP_bot.Inst_MULADD._0375_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0376_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0377_
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1137_ Tile_X0Y1_DSP_bot.Inst_MULADD._0306_ Tile_X0Y1_DSP_bot.Inst_MULADD._0291_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0308_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0309_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[155\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C9 sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1068_ Tile_X0Y1_DSP_bot.Inst_MULADD._0223_ Tile_X0Y1_DSP_bot.Inst_MULADD._0226_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0238_ Tile_X0Y1_DSP_bot.Inst_MULADD._0171_ Tile_X0Y1_DSP_bot.Inst_MULADD._0166_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0241_ sky130_fd_sc_hd__o2111ai_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12 net232 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[108\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23 net244 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[119\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_77_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_147_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.strobe_outbuf_9._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[9\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_330_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.SS4BEG2 VGND VGND VPWR VPWR net704
+ sky130_fd_sc_hd__clkbuf_1
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_261_ Tile_X0Y1_DSP_bot.FrameData_O\[13\] VGND VGND VPWR VPWR net635 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[149\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
X_192_ Tile_X0Y0_DSP_top.WW4BEG\[8\] VGND VGND VPWR VPWR net581 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END2
+ net1 net7 Tile_X0Y0_DSP_top.ConfigBits\[250\] Tile_X0Y0_DSP_top.ConfigBits\[251\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.strobe_outbuf_2._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[2\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[2\] sky130_fd_sc_hd__buf_8
XFILLER_0_154_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7 net258 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[167\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[348\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1755_ net333 Tile_X0Y1_DSP_bot.C13 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[13\] sky130_fd_sc_hd__dfxtp_1
XANTENNA_19 Tile_X0Y0_DSP_top.FrameStrobe\[16\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1686_ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ Tile_X0Y1_DSP_bot.Inst_MULADD._0511_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0512_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0836_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_140_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_112_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.WW4BEG_outbuf_7._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[7\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[7\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._56_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG2 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.E6END_inbuf_4._0_ net29 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_131_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb3 Tile_X0Y0_DSP_top.S4BEG\[3\]
+ net341 net357 Tile_X0Y1_DSP_bot.ConfigBits\[360\] Tile_X0Y1_DSP_bot.ConfigBits\[361\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput671 net671 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput660 net660 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[7] sky130_fd_sc_hd__clkbuf_4
Xoutput682 net682 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[7] sky130_fd_sc_hd__buf_2
Xoutput693 net693 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_0._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.strobe_inbuf_17._0_ net269 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[17\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_313_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG1 VGND VGND VPWR VPWR net687
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1540_ Tile_X0Y1_DSP_bot.Inst_MULADD._0702_ Tile_X0Y1_DSP_bot.Inst_MULADD._0703_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0705_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0706_
+ sky130_fd_sc_hd__o21a_1
X_244_ Tile_X0Y1_DSP_bot.EE4BEG\[12\] VGND VGND VPWR VPWR net618 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput28 Tile_X0Y0_E6END[5] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 Tile_X0Y0_E2MID[4] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_134_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput39 Tile_X0Y0_EE4END[15] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_175_ Tile_X0Y0_DSP_top.W6BEG\[3\] VGND VGND VPWR VPWR net560 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1471_ Tile_X0Y1_DSP_bot.Inst_MULADD._0624_ Tile_X0Y1_DSP_bot.Inst_MULADD._0626_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0631_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0638_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.E6BEG_outbuf_2._0_ Tile_X0Y0_DSP_top.E6BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11 net231 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[139\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22 net243 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[150\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_114_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_114_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_114_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1738_ net333 Tile_X0Y1_DSP_bot.B4 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1669_ Tile_X0Y1_DSP_bot.Inst_MULADD._0825_ Tile_X0Y1_DSP_bot.Inst_MULADD._0827_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0828_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._39_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID1 sky130_fd_sc_hd__buf_1
XFILLER_0_48_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG6.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[272\] Tile_X0Y0_DSP_top.ConfigBits\[273\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG6 sky130_fd_sc_hd__mux4_2
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.E6END_inbuf_4._0_ net209 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst0
+ net282 net290 net182 net190 Tile_X0Y1_DSP_bot.ConfigBits\[272\] Tile_X0Y1_DSP_bot.ConfigBits\[273\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8 net259 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[8\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG1
+ Tile_X0Y1_DSP_bot.ConfigBits\[31\] Tile_X0Y1_DSP_bot.ConfigBits\[32\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_116_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput490 net490 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG0 net19
+ net99 net151 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG4 Tile_X0Y0_DSP_top.ConfigBits\[158\]
+ Tile_X0Y0_DSP_top.ConfigBits\[159\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.ConfigBits\[58\] Tile_X0Y1_DSP_bot.ConfigBits\[59\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0971_ Tile_X0Y1_DSP_bot.Inst_MULADD._0033_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_ Tile_X0Y1_DSP_bot.Inst_MULADD._0141_ Tile_X0Y1_DSP_bot.Inst_MULADD._0144_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0145_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_158_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 net2 net82 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[45\] Tile_X0Y0_DSP_top.ConfigBits\[46\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1523_ Tile_X0Y1_DSP_bot.Inst_MULADD._0677_ Tile_X0Y1_DSP_bot.Inst_MULADD._0679_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0682_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0689_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_227_ Tile_X0Y1_DSP_bot.E6BEG\[7\] VGND VGND VPWR VPWR net612 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_158_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG2 VGND VGND VPWR VPWR net541
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1454_ Tile_X0Y1_DSP_bot.Inst_MULADD._0614_ Tile_X0Y1_DSP_bot.Inst_MULADD._0620_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0621_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0622_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_089_ Tile_X0Y0_DSP_top.FrameStrobe_O\[9\] VGND VGND VPWR VPWR net481 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1385_ Tile_X0Y1_DSP_bot.Inst_MULADD._0543_ Tile_X0Y1_DSP_bot.Inst_MULADD._0545_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0553_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0554_
+ sky130_fd_sc_hd__and3_2
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[151\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_157_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.SS4BEG_outbuf_0._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[0\] sky130_fd_sc_hd__clkbuf_2
Xinput218 Tile_X0Y1_EE4END[14] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__clkbuf_1
Xinput207 Tile_X0Y1_E6END[4] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.S4BEG\[2\] Tile_X0Y0_DSP_top.SS4BEG\[2\] net340 net354 Tile_X0Y1_DSP_bot.ConfigBits\[324\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[325\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
Xinput229 Tile_X0Y1_FrameData[0] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21 net242 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[181\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10 net230 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[170\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_151_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_012_ Tile_X0Y0_DSP_top.E2BEGb\[0\] VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID3
+ net16 net96 net148 Tile_X0Y0_DSP_top.ConfigBits\[200\] Tile_X0Y0_DSP_top.ConfigBits\[201\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG1
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1170_ Tile_X0Y1_DSP_bot.Inst_MULADD._0325_ Tile_X0Y1_DSP_bot.Inst_MULADD._0336_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0331_ Tile_X0Y1_DSP_bot.Inst_MULADD._0249_ Tile_X0Y1_DSP_bot.Inst_MULADD._0335_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0341_ sky130_fd_sc_hd__a32oi_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0954_ Tile_X0Y1_DSP_bot.Inst_MULADD._0125_ Tile_X0Y1_DSP_bot.Inst_MULADD._0126_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0127_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0129_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_127_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0885_ Tile_X0Y1_DSP_bot.A2 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0061_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_84_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END2
+ net125 net139 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG4 Tile_X0Y0_DSP_top.ConfigBits\[400\]
+ Tile_X0Y0_DSP_top.ConfigBits\[401\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_142_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1506_ Tile_X0Y1_DSP_bot.Inst_MULADD._0671_ Tile_X0Y1_DSP_bot.Inst_MULADD._0672_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1437_ Tile_X0Y1_DSP_bot.Inst_MULADD._0050_ Tile_X0Y1_DSP_bot.Inst_MULADD._0080_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0273_ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0605_ sky130_fd_sc_hd__or4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1368_ Tile_X0Y1_DSP_bot.Inst_MULADD._0045_ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_ Tile_X0Y1_DSP_bot.Inst_MULADD._0080_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0537_ sky130_fd_sc_hd__a211o_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1299_ Tile_X0Y1_DSP_bot.Inst_MULADD._0196_ Tile_X0Y1_DSP_bot.Inst_MULADD._0107_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0151_ Tile_X0Y1_DSP_bot.Inst_MULADD._0152_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0469_ sky130_fd_sc_hd__nand4_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_137_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_160_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_156_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.N4END_inbuf_8._0_ Tile_X0Y0_DSP_top.N4END\[12\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_136_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1222_ Tile_X0Y1_DSP_bot.Inst_MULADD._0365_ Tile_X0Y1_DSP_bot.Inst_MULADD._0371_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0377_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0393_
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1153_ Tile_X0Y1_DSP_bot.Inst_MULADD._0252_ Tile_X0Y1_DSP_bot.Inst_MULADD._0253_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0316_ Tile_X0Y1_DSP_bot.Inst_MULADD._0324_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0325_ sky130_fd_sc_hd__o22ai_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1084_ Tile_X0Y1_DSP_bot.A6 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0256_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst2
+ net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[288\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[289\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_inst0
+ net282 net182 net335 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.ConfigBits\[87\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[88\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[250\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_159_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_EF_BEG2
+ Tile_X0Y0_DSP_top.ConfigBits\[95\] Tile_X0Y0_DSP_top.ConfigBits\[96\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0937_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ Tile_X0Y1_DSP_bot.Inst_MULADD._0110_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0111_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0112_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_57_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_115_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0868_ Tile_X0Y1_DSP_bot.Inst_MULADD._0044_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0045_ sky130_fd_sc_hd__buf_4
XTile_X0Y1_DSP_bot.NN4END_inbuf_3._0_ net330 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[3\]
+ sky130_fd_sc_hd__buf_2
XFILLER_0_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_130_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20 net241 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[212\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31 net253 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[223\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._10_ net15 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E2BEGb\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.N4BEG_outbuf_6._0_ Tile_X0Y0_DSP_top.N4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[6\] sky130_fd_sc_hd__buf_2
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2 net251 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[386\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_98_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_129_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.N4END_inbuf_8._0_ net304 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_3._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END3 sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._72_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG2 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1205_ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0375_ Tile_X0Y1_DSP_bot.Inst_MULADD._0372_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0376_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_93_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1136_ Tile_X0Y1_DSP_bot.Inst_MULADD._0227_ Tile_X0Y1_DSP_bot.Inst_MULADD._0228_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0217_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0308_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[155\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1067_ Tile_X0Y1_DSP_bot.Inst_MULADD._0184_ Tile_X0Y1_DSP_bot.Inst_MULADD._0185_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0239_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0240_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13 net233 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[109\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24 net245 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[120\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_6._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_115_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.W6BEG_outbuf_6._0_ Tile_X0Y0_DSP_top.W6BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[6\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.S4BEG_outbuf_10._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[10\] sky130_fd_sc_hd__clkbuf_4
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG0 net300
+ net200 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG7 net353 Tile_X0Y1_DSP_bot.ConfigBits\[216\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[217\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_top2bot17.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_36_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_260_ Tile_X0Y1_DSP_bot.FrameData_O\[12\] VGND VGND VPWR VPWR net634 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_191_ Tile_X0Y0_DSP_top.WW4BEG\[7\] VGND VGND VPWR VPWR net580 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG0 net188
+ Tile_X0Y0_DSP_top.SS4BEG\[3\] net374 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[392\] Tile_X0Y1_DSP_bot.ConfigBits\[393\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG0 sky130_fd_sc_hd__mux4_1
XFILLER_0_121_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst1
+ net21 net87 net139 net153 Tile_X0Y0_DSP_top.ConfigBits\[250\] Tile_X0Y0_DSP_top.ConfigBits\[251\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30 net252 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[254\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8 net259 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[168\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[349\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1754_ net333 Tile_X0Y1_DSP_bot.C12 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1685_ Tile_X0Y1_DSP_bot.Inst_MULADD._0835_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_152_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._55_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1119_ Tile_X0Y1_DSP_bot.Inst_MULADD._0288_ Tile_X0Y1_DSP_bot.Inst_MULADD._0289_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0290_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0291_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_53_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_116_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_143_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.EE4BEG_outbuf_0._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[360\] Tile_X0Y1_DSP_bot.ConfigBits\[361\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput672 net672 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput661 net661 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[8] sky130_fd_sc_hd__buf_2
Xoutput650 net650 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[27] sky130_fd_sc_hd__clkbuf_4
Xoutput683 net683 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[0] sky130_fd_sc_hd__buf_2
Xoutput694 net694 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[5] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END3
+ net11 net91 net143 Tile_X0Y0_DSP_top.ConfigBits\[222\] Tile_X0Y0_DSP_top.ConfigBits\[223\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG0 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_inbuf_5._0_ net256 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[5\]
+ sky130_fd_sc_hd__buf_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.data_outbuf_26._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[26\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[26\] sky130_fd_sc_hd__clkbuf_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END0 net9 Tile_X0Y0_DSP_top.ConfigBits\[290\]
+ Tile_X0Y0_DSP_top.ConfigBits\[291\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
X_312_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S4BEG0 VGND VGND VPWR VPWR net686
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_119_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_243_ Tile_X0Y1_DSP_bot.EE4BEG\[11\] VGND VGND VPWR VPWR net617 sky130_fd_sc_hd__clkbuf_1
Xinput18 Tile_X0Y0_E2MID[5] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 Tile_X0Y0_E6END[6] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_122_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_174_ Tile_X0Y0_DSP_top.W6BEG\[2\] VGND VGND VPWR VPWR net559 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1470_ Tile_X0Y1_DSP_bot.Inst_MULADD._0428_ Tile_X0Y1_DSP_bot.Inst_MULADD._0634_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0636_ Tile_X0Y1_DSP_bot.Inst_MULADD._0637_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q10 sky130_fd_sc_hd__a31o_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12 net232 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[140\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23 net244 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[151\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.data_outbuf_17._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[17\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1737_ net333 Tile_X0Y1_DSP_bot.B3 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1668_ Tile_X0Y1_DSP_bot.Inst_MULADD._0787_ Tile_X0Y1_DSP_bot.Inst_MULADD._0810_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0824_ Tile_X0Y1_DSP_bot.Inst_MULADD._0826_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0827_ sky130_fd_sc_hd__o211ai_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1599_ Tile_X0Y1_DSP_bot.Inst_MULADD._0755_ Tile_X0Y1_DSP_bot.Inst_MULADD._0760_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0762_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0763_
+ sky130_fd_sc_hd__a21o_1
XTile_X0Y0_DSP_top.S4BEG_outbuf_6._0_ Tile_X0Y0_DSP_top.S4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._38_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID0 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_48_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb5
+ net335 net337 Tile_X0Y1_DSP_bot.ConfigBits\[272\] Tile_X0Y1_DSP_bot.ConfigBits\[273\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_93_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9 net260 net264 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[9\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame12_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_148_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput480 net480 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[8] sky130_fd_sc_hd__clkbuf_4
Xoutput491 net491 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[5] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID2
+ net15 net147 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG4 Tile_X0Y0_DSP_top.ConfigBits\[160\]
+ Tile_X0Y0_DSP_top.ConfigBits\[161\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst2
+ net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[58\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[59\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0970_ Tile_X0Y1_DSP_bot.Inst_MULADD._0142_ Tile_X0Y1_DSP_bot.Inst_MULADD._0143_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0144_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_AB_BEG0
+ Tile_X0Y0_DSP_top.ConfigBits\[45\] Tile_X0Y0_DSP_top.ConfigBits\[46\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1522_ Tile_X0Y1_DSP_bot.Inst_MULADD._0688_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q11 sky130_fd_sc_hd__buf_1
X_226_ Tile_X0Y1_DSP_bot.E6BEG\[6\] VGND VGND VPWR VPWR net611 sky130_fd_sc_hd__clkbuf_1
X_157_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG1 VGND VGND VPWR VPWR net540
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1453_ Tile_X0Y1_DSP_bot.Inst_MULADD._0563_ Tile_X0Y1_DSP_bot.Inst_MULADD._0569_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0562_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0621_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_088_ Tile_X0Y0_DSP_top.FrameStrobe_O\[8\] VGND VGND VPWR VPWR net480 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1384_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B7
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0075_ Tile_X0Y1_DSP_bot.Inst_MULADD._0346_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0553_ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[152\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_157_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst0
+ net284 net292 net184 net192 Tile_X0Y1_DSP_bot.ConfigBits\[312\] Tile_X0Y1_DSP_bot.ConfigBits\[313\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_101_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput208 Tile_X0Y1_E6END[5] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[324\] Tile_X0Y1_DSP_bot.ConfigBits\[325\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
Xinput219 Tile_X0Y1_EE4END[15] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11 net231 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[171\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22 net243 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[182\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0 net229 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[288\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_151_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_011_ Tile_X0Y0_DSP_top.E2BEG\[7\] VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__buf_1
XFILLER_0_104_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.W6END_inbuf_2._0_ net159 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_276 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID5
+ net18 net98 net150 Tile_X0Y0_DSP_top.ConfigBits\[202\] Tile_X0Y0_DSP_top.ConfigBits\[203\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0953_ Tile_X0Y1_DSP_bot.Inst_MULADD._0125_ Tile_X0Y1_DSP_bot.Inst_MULADD._0126_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0127_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0128_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_29_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0884_ Tile_X0Y1_DSP_bot.Inst_MULADD._0046_ Tile_X0Y1_DSP_bot.Inst_MULADD._0052_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0054_ Tile_X0Y1_DSP_bot.Inst_MULADD._0057_ Tile_X0Y1_DSP_bot.Inst_MULADD._0034_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0060_ sky130_fd_sc_hd__a32o_1
XFILLER_0_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG2 net24
+ net108 net174 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y0_DSP_top.ConfigBits\[402\]
+ Tile_X0Y0_DSP_top.ConfigBits\[403\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1505_ Tile_X0Y1_DSP_bot.Inst_MULADD._0669_ Tile_X0Y1_DSP_bot.Inst_MULADD._0663_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0667_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0672_
+ sky130_fd_sc_hd__nand3b_1
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_209_ Tile_X0Y1_DSP_bot.E2BEG\[5\] VGND VGND VPWR VPWR net592 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1436_ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_ Tile_X0Y1_DSP_bot.Inst_MULADD._0439_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0533_ Tile_X0Y1_DSP_bot.Inst_MULADD._0603_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0604_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_96_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1367_ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0536_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1298_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0468_ sky130_fd_sc_hd__and4_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END6
+ net3 net11 Tile_X0Y0_DSP_top.ConfigBits\[362\] Tile_X0Y0_DSP_top.ConfigBits\[363\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_6._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_152_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1221_ Tile_X0Y1_DSP_bot.Inst_MULADD._0350_ Tile_X0Y1_DSP_bot.Inst_MULADD._0354_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0388_ Tile_X0Y1_DSP_bot.Inst_MULADD._0391_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0392_ sky130_fd_sc_hd__o22ai_4
XTile_X0Y1_DSP_bot.W6END_inbuf_2._0_ net360 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1152_ Tile_X0Y1_DSP_bot.Inst_MULADD._0166_ Tile_X0Y1_DSP_bot.Inst_MULADD._0239_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0319_ Tile_X0Y1_DSP_bot.Inst_MULADD._0323_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0324_ sky130_fd_sc_hd__a2bb2oi_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1083_ Tile_X0Y1_DSP_bot.Inst_MULADD._0189_ Tile_X0Y1_DSP_bot.Inst_MULADD._0229_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0195_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0255_
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[288\] Tile_X0Y1_DSP_bot.ConfigBits\[289\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_AB_BEG3
+ Tile_X0Y1_DSP_bot.ConfigBits\[87\] Tile_X0Y1_DSP_bot.ConfigBits\[88\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_SS4BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_159_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[251\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0936_ Tile_X0Y1_DSP_bot.Inst_MULADD._0026_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0111_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0867_ Tile_X0Y1_DSP_bot.ConfigBits\[1\] Tile_X0Y1_DSP_bot.Inst_MULADD._0042_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0043_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0044_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_57_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_123_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1419_ Tile_X0Y1_DSP_bot.Inst_MULADD._0435_ Tile_X0Y1_DSP_bot.Inst_MULADD._0519_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0586_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0587_
+ sky130_fd_sc_hd__nand3_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21 net242 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[213\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10 net230 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[202\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_138_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_133_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3 net254 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[387\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG0 net299
+ net199 net352 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG5 Tile_X0Y1_DSP_bot.ConfigBits\[176\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[177\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.WW4END_inbuf_4._0_ net380 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[18\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG0 sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._71_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG1 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1204_ Tile_X0Y1_DSP_bot.Inst_MULADD._0108_ Tile_X0Y1_DSP_bot.Inst_MULADD._0155_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0374_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0375_
+ sky130_fd_sc_hd__o21ai_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END3
+ net110 net165 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 Tile_X0Y0_DSP_top.ConfigBits\[374\]
+ Tile_X0Y0_DSP_top.ConfigBits\[375\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG0
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1135_ Tile_X0Y1_DSP_bot.Inst_MULADD._0199_ Tile_X0Y1_DSP_bot.Inst_MULADD._0235_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0306_ Tile_X0Y1_DSP_bot.Inst_MULADD._0291_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0307_ sky130_fd_sc_hd__o211a_4
XFILLER_0_93_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1066_ Tile_X0Y1_DSP_bot.Inst_MULADD._0223_ Tile_X0Y1_DSP_bot.Inst_MULADD._0226_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0238_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0239_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput380 Tile_X0Y1_WW4END[8] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25 net246 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[121\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14 net234 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[110\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END5
+ net2 net10 Tile_X0Y0_DSP_top.ConfigBits\[326\] Tile_X0Y0_DSP_top.ConfigBits\[327\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0919_ Tile_X0Y1_DSP_bot.Inst_MULADD._0093_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0095_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_115_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_130_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG1 net296
+ net196 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG3 net349 Tile_X0Y1_DSP_bot.ConfigBits\[218\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[219\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_76_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_146_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_190_ Tile_X0Y0_DSP_top.WW4BEG\[6\] VGND VGND VPWR VPWR net579 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG1 net309
+ net187 net345 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[394\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[395\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_91_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[250\] Tile_X0Y0_DSP_top.ConfigBits\[251\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20 net241 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[244\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31 net253 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[255\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9 net260 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[169\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[350\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1753_ net333 Tile_X0Y1_DSP_bot.C11 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1684_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0426_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0835_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_420 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._54_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEG0 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1118_ Tile_X0Y1_DSP_bot.Inst_MULADD._0284_ Tile_X0Y1_DSP_bot.Inst_MULADD._0285_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0290_ sky130_fd_sc_hd__nand2_2
XTile_X0Y0_DSP_top.data_inbuf_31._0_ net73 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[31\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1049_ Tile_X0Y1_DSP_bot.Inst_MULADD._0164_ Tile_X0Y1_DSP_bot.Inst_MULADD._0163_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0158_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0222_
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_58_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_143_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[360\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[361\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
Xoutput662 net662 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput640 net640 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput651 net651 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[28] sky130_fd_sc_hd__clkbuf_4
Xoutput673 net673 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput695 net695 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput684 net684 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[10] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END2
+ net7 net87 net173 Tile_X0Y0_DSP_top.ConfigBits\[224\] Tile_X0Y0_DSP_top.ConfigBits\[225\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG1 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.data_inbuf_22._0_ net63 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[22\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.WW4END_inbuf_0._0_ net175 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst1
+ net21 net89 net141 net153 Tile_X0Y0_DSP_top.ConfigBits\[290\] Tile_X0Y0_DSP_top.ConfigBits\[291\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
X_311_ Tile_X0Y1_DSP_bot.S4BEG\[11\] VGND VGND VPWR VPWR net685 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst0
+ net281 net285 net181 net185 Tile_X0Y1_DSP_bot.ConfigBits\[348\] Tile_X0Y1_DSP_bot.ConfigBits\[349\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
X_242_ Tile_X0Y1_DSP_bot.EE4BEG\[10\] VGND VGND VPWR VPWR net616 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput19 Tile_X0Y0_E2MID[6] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__buf_2
XFILLER_0_119_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_173_ Tile_X0Y0_DSP_top.W6BEG\[1\] VGND VGND VPWR VPWR net558 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.strobe_inbuf_7._0_ Tile_X0Y0_DSP_top.FrameStrobe\[7\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[7\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13 net233 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[141\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24 net245 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[152\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.data_inbuf_13._0_ net53 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[13\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[24\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4END\[12\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1736_ net333 Tile_X0Y1_DSP_bot.B2 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_130_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1667_ Tile_X0Y1_DSP_bot.Inst_MULADD._0814_ Tile_X0Y1_DSP_bot.Inst_MULADD._0813_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0817_ Tile_X0Y1_DSP_bot.Inst_MULADD._0816_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0826_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_125_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1598_ Tile_X0Y1_DSP_bot.Inst_MULADD._0761_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[14\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0762_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._37_ net200 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEGb\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[272\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[273\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_inbuf_31._0_ net253 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[31\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_148_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput470 net470 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[17] sky130_fd_sc_hd__clkbuf_4
Xoutput492 net492 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput481 net481 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[9] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30 net252 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[286\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID4
+ net17 net97 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 Tile_X0Y0_DSP_top.ConfigBits\[162\]
+ Tile_X0Y0_DSP_top.ConfigBits\[163\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG2
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDa_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHa_BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[58\] Tile_X0Y1_DSP_bot.ConfigBits\[59\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.SS4END_inbuf_6._0_ Tile_X0Y0_DSP_top.SS4BEG\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[6\] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.data_inbuf_22._0_ net243 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[22\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1521_ Tile_X0Y1_DSP_bot.Inst_MULADD._0687_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0688_
+ sky130_fd_sc_hd__mux2_1
X_225_ Tile_X0Y1_DSP_bot.E6BEG\[5\] VGND VGND VPWR VPWR net610 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1452_ Tile_X0Y1_DSP_bot.Inst_MULADD._0613_ Tile_X0Y1_DSP_bot.Inst_MULADD._0619_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0612_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0620_
+ sky130_fd_sc_hd__nor3b_1
X_156_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG0 VGND VGND VPWR VPWR net539
+ sky130_fd_sc_hd__clkbuf_1
X_087_ Tile_X0Y0_DSP_top.FrameStrobe_O\[7\] VGND VGND VPWR VPWR net479 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1383_ Tile_X0Y1_DSP_bot.Inst_MULADD._0543_ Tile_X0Y1_DSP_bot.Inst_MULADD._0545_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0063_ Tile_X0Y1_DSP_bot.Inst_MULADD._0351_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0552_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_122_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_125_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[153\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.data_inbuf_13._0_ net233 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[13\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_157_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_145_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1719_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0013_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb7 net337 Tile_X0Y1_DSP_bot.ConfigBits\[312\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[313\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput209 Tile_X0Y1_E6END[6] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[324\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[325\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[97\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.WW4BEG1 sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12 net232 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[172\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23 net244 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[183\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_66_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1 net240 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[289\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_151_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_010_ Tile_X0Y0_DSP_top.E2BEG\[6\] VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_EFb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID1
+ net14 net94 net146 Tile_X0Y0_DSP_top.ConfigBits\[204\] Tile_X0Y0_DSP_top.ConfigBits\[205\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_10._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG\[10\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.EE4END_inbuf_5._0_ net228 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0952_ Tile_X0Y1_DSP_bot.Inst_MULADD._0060_ Tile_X0Y1_DSP_bot.Inst_MULADD._0091_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0090_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0127_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_139_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.strobe_inbuf_14._0_ Tile_X0Y0_DSP_top.FrameStrobe\[14\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[14\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0883_ Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ Tile_X0Y1_DSP_bot.Inst_MULADD._0058_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0059_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_142_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_GH_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4END0
+ net21 net137 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG4 Tile_X0Y0_DSP_top.ConfigBits\[404\]
+ Tile_X0Y0_DSP_top.ConfigBits\[405\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG3
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1504_ Tile_X0Y1_DSP_bot.Inst_MULADD._0613_ Tile_X0Y1_DSP_bot.Inst_MULADD._0619_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0612_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0671_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_208_ Tile_X0Y1_DSP_bot.E2BEG\[4\] VGND VGND VPWR VPWR net591 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_139_ Tile_X0Y0_DSP_top.NN4BEG\[3\] VGND VGND VPWR VPWR net527 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1435_ Tile_X0Y1_DSP_bot.Inst_MULADD._0601_ Tile_X0Y1_DSP_bot.Inst_MULADD._0602_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0603_ sky130_fd_sc_hd__nand2_2
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1366_ Tile_X0Y1_DSP_bot.Inst_MULADD._0080_ Tile_X0Y1_DSP_bot.Inst_MULADD._0522_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0526_ Tile_X0Y1_DSP_bot.Inst_MULADD._0528_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0535_ sky130_fd_sc_hd__o22a_4
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1297_ Tile_X0Y1_DSP_bot.Inst_MULADD._0464_ Tile_X0Y1_DSP_bot.Inst_MULADD._0465_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0466_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0467_
+ sky130_fd_sc_hd__o21ai_4
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst1
+ net81 net83 net91 net135 Tile_X0Y0_DSP_top.ConfigBits\[362\] Tile_X0Y0_DSP_top.ConfigBits\[363\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_30 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_156_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.SS4END_inbuf_2._0_ net129 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[2\]
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.strobe_outbuf_16._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[16\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[16\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1220_ Tile_X0Y1_DSP_bot.Inst_MULADD._0389_ Tile_X0Y1_DSP_bot.Inst_MULADD._0390_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0387_ Tile_X0Y1_DSP_bot.Inst_MULADD._0378_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0391_ sky130_fd_sc_hd__o211a_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1151_ Tile_X0Y1_DSP_bot.Inst_MULADD._0320_ Tile_X0Y1_DSP_bot.Inst_MULADD._0322_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0314_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0323_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_66_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1082_ Tile_X0Y1_DSP_bot.Inst_MULADD._0223_ Tile_X0Y1_DSP_bot.Inst_MULADD._0226_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0184_ Tile_X0Y1_DSP_bot.Inst_MULADD._0238_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0254_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_89_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG0.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[290\] Tile_X0Y1_DSP_bot.ConfigBits\[291\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_106_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[252\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0935_ Tile_X0Y1_DSP_bot.A3 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0110_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_155_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.E6BEG_outbuf_9._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[9\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0866_ Tile_X0Y1_DSP_bot.ConfigBits\[1\] Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0043_ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END0
+ net1 net33 Tile_X0Y0_DSP_top.ConfigBits\[274\] Tile_X0Y0_DSP_top.ConfigBits\[275\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_127_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1418_ Tile_X0Y1_DSP_bot.Inst_MULADD._0564_ Tile_X0Y1_DSP_bot.Inst_MULADD._0566_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0573_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0586_
+ sky130_fd_sc_hd__o21a_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11 net231 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[203\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_40_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22 net243 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[214\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_147_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1349_ Tile_X0Y1_DSP_bot.Inst_MULADD._0492_ Tile_X0Y1_DSP_bot.Inst_MULADD._0493_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0436_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0518_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_158_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_133_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4 net255 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[388\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG1 net295
+ net195 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG5
+ Tile_X0Y1_DSP_bot.ConfigBits\[178\] Tile_X0Y1_DSP_bot.ConfigBits\[179\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_133_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[103\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.WW4BEG1 sky130_fd_sc_hd__o21ai_1
XTile_X0Y0_DSP_top.EE4END_inbuf_1._0_ net44 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_152_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[18\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_109_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_152_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._70_ net338 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEG0
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1203_ Tile_X0Y1_DSP_bot.Inst_MULADD._0269_ Tile_X0Y1_DSP_bot.Inst_MULADD._0270_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0374_
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y1_DSP_bot.strobe_outbuf_5._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[5\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[5\] sky130_fd_sc_hd__buf_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG1 net41
+ net109 net144 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG1 Tile_X0Y0_DSP_top.ConfigBits\[376\]
+ Tile_X0Y0_DSP_top.ConfigBits\[377\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1134_ Tile_X0Y1_DSP_bot.Inst_MULADD._0255_ Tile_X0Y1_DSP_bot.Inst_MULADD._0276_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0281_ Tile_X0Y1_DSP_bot.Inst_MULADD._0284_ Tile_X0Y1_DSP_bot.Inst_MULADD._0285_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0306_ sky130_fd_sc_hd__o2111ai_4
XFILLER_0_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1065_ Tile_X0Y1_DSP_bot.Inst_MULADD._0223_ Tile_X0Y1_DSP_bot.Inst_MULADD._0237_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0157_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0238_
+ sky130_fd_sc_hd__o21ai_4
Xinput381 Tile_X0Y1_WW4END[9] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__clkbuf_1
Xinput370 Tile_X0Y1_WW4END[13] VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26 net247 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[122\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15 net235 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[111\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_158_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst1
+ net82 net90 net134 net136 Tile_X0Y0_DSP_top.ConfigBits\[326\] Tile_X0Y0_DSP_top.ConfigBits\[327\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_117_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_N1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_CD_BEG1 Tile_X0Y0_DSP_top.ConfigBits\[0\]
+ Tile_X0Y0_DSP_top.ConfigBits\[1\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG0
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_77_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.N4BEG_outbuf_0._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END0 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.NN4BEG_outbuf_11._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.NN4BEG\[11\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0918_ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._0849_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[0\] Tile_X0Y1_DSP_bot.Inst_MULADD._0026_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0027_ sky130_fd_sc_hd__or2b_2
XFILLER_0_143_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.E6END_inbuf_7._0_ net32 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG2 net298
+ net198 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG5 net351 Tile_X0Y1_DSP_bot.ConfigBits\[220\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[221\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG2
+ sky130_fd_sc_hd__mux4_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_134_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG2 net324
+ net220 Tile_X0Y0_DSP_top.S4BEG\[1\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[396\] Tile_X0Y1_DSP_bot.ConfigBits\[397\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_0_32_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[250\] Tile_X0Y0_DSP_top.ConfigBits\[251\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_3._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_129_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10 net230 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[234\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21 net242 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[245\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_144_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[351\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame1_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1752_ net333 Tile_X0Y1_DSP_bot.C10 VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1683_ Tile_X0Y1_DSP_bot.Inst_MULADD._0829_ Tile_X0Y1_DSP_bot.Inst_MULADD._0339_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0006_ sky130_fd_sc_hd__nor2_1
XTile_X0Y0_DSP_top.E6BEG_outbuf_5._0_ Tile_X0Y0_DSP_top.E6BEG_i\[5\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_112_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._53_ net300 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END7
+ sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.strobe_outbuf_11._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[11\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1117_ Tile_X0Y1_DSP_bot.Inst_MULADD._0277_ Tile_X0Y1_DSP_bot.Inst_MULADD._0280_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0255_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0289_
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y1_DSP_bot.W6BEG_outbuf_0._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.data_inbuf_2._0_ net71 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1048_ Tile_X0Y1_DSP_bot.Inst_MULADD._0199_ Tile_X0Y1_DSP_bot.Inst_MULADD._0220_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0216_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0221_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_143_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG2.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[362\] Tile_X0Y1_DSP_bot.ConfigBits\[363\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2 sky130_fd_sc_hd__mux4_2
Xoutput663 net663 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput630 net630 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput641 net641 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput652 net652 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[29] sky130_fd_sc_hd__clkbuf_4
Xoutput674 net674 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput696 net696 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput685 net685 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[11] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END4
+ net9 net125 net141 Tile_X0Y0_DSP_top.ConfigBits\[226\] Tile_X0Y0_DSP_top.ConfigBits\[227\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG2 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.E6END_inbuf_7._0_ net212 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_310_ Tile_X0Y1_DSP_bot.S4BEG\[10\] VGND VGND VPWR VPWR net684 sky130_fd_sc_hd__clkbuf_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[290\] Tile_X0Y0_DSP_top.ConfigBits\[291\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb0
+ net334 net336 Tile_X0Y1_DSP_bot.ConfigBits\[348\] Tile_X0Y1_DSP_bot.ConfigBits\[349\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
X_241_ Tile_X0Y1_DSP_bot.EE4BEG\[9\] VGND VGND VPWR VPWR net630 sky130_fd_sc_hd__clkbuf_1
X_172_ Tile_X0Y0_DSP_top.W6BEG\[0\] VGND VGND VPWR VPWR net555 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25 net246 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[153\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14 net234 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[142\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[24\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_157_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_117_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1735_ net333 Tile_X0Y1_DSP_bot.B1 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1666_ Tile_X0Y1_DSP_bot.Inst_MULADD._0821_ Tile_X0Y1_DSP_bot.Inst_MULADD._0815_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0824_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0825_
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_82_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1597_ Tile_X0Y1_DSP_bot.C14 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[14\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0761_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._36_ net199 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEGb\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.NN4BEG_outbuf_0._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[0\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.ConfigBits\[272\] Tile_X0Y1_DSP_bot.ConfigBits\[273\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_78_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_148_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.SS4BEG_outbuf_3._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[3\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.data_outbuf_20._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[20\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[20\] sky130_fd_sc_hd__clkbuf_1
Xoutput471 net471 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[18] sky130_fd_sc_hd__clkbuf_4
Xoutput460 net460 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[8] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20 net241 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[276\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput482 net482 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[0] sky130_fd_sc_hd__buf_2
Xoutput493 net493 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[7] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31 net253 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[287\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_CDa_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID0
+ net93 net145 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG4 Tile_X0Y0_DSP_top.ConfigBits\[164\]
+ Tile_X0Y0_DSP_top.ConfigBits\[165\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDa_BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_E6BEG1.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[60\] Tile_X0Y1_DSP_bot.ConfigBits\[61\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG\[11\] sky130_fd_sc_hd__mux4_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1520_ Tile_X0Y1_DSP_bot.Inst_MULADD._0685_ Tile_X0Y1_DSP_bot.Inst_MULADD._0686_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0687_ sky130_fd_sc_hd__or2_1
X_224_ Tile_X0Y1_DSP_bot.E6BEG\[4\] VGND VGND VPWR VPWR net609 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1451_ Tile_X0Y1_DSP_bot.Inst_MULADD._0607_ Tile_X0Y1_DSP_bot.Inst_MULADD._0610_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0549_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0619_
+ sky130_fd_sc_hd__a21oi_1
X_155_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG3 VGND VGND VPWR VPWR net538
+ sky130_fd_sc_hd__clkbuf_1
X_086_ Tile_X0Y0_DSP_top.FrameStrobe_O\[6\] VGND VGND VPWR VPWR net478 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1382_ Tile_X0Y1_DSP_bot.Inst_MULADD._0455_ Tile_X0Y1_DSP_bot.Inst_MULADD._0454_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0550_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0551_
+ sky130_fd_sc_hd__a21oi_4
XTile_X0Y1_DSP_bot.data_outbuf_11._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[11\] sky130_fd_sc_hd__clkbuf_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.S4BEG_outbuf_0._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[0\] sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[154\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0 net229 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[32\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_145_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_145_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1718_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0012_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[312\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[313\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1649_ Tile_X0Y1_DSP_bot.Inst_MULADD._0808_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0809_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_113_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_113_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._19_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot15
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C17 sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG1.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[326\] Tile_X0Y1_DSP_bot.ConfigBits\[327\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[97\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13 net233 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[173\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24 net245 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[184\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_136_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2 net251 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[290\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_144_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._0951_ Tile_X0Y1_DSP_bot.Inst_MULADD._0124_ Tile_X0Y1_DSP_bot.Inst_MULADD._0123_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0099_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0126_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0882_ Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0059_ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1503_ Tile_X0Y1_DSP_bot.Inst_MULADD._0663_ Tile_X0Y1_DSP_bot.Inst_MULADD._0667_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0669_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0670_
+ sky130_fd_sc_hd__a21boi_2
XFILLER_0_92_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_207_ Tile_X0Y1_DSP_bot.E2BEG\[3\] VGND VGND VPWR VPWR net590 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_138_ Tile_X0Y0_DSP_top.NN4BEG\[2\] VGND VGND VPWR VPWR net526 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1434_ Tile_X0Y1_DSP_bot.Inst_MULADD._0261_ Tile_X0Y1_DSP_bot.Inst_MULADD._0263_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_ Tile_X0Y1_DSP_bot.Inst_MULADD._0599_ Tile_X0Y1_DSP_bot.Inst_MULADD._0600_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0602_ sky130_fd_sc_hd__o2111ai_1
X_069_ Tile_X0Y0_DSP_top.FrameData_O\[21\] VGND VGND VPWR VPWR net443 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1365_ Tile_X0Y1_DSP_bot.Inst_MULADD._0463_ Tile_X0Y1_DSP_bot.Inst_MULADD._0457_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0529_ Tile_X0Y1_DSP_bot.Inst_MULADD._0533_ Tile_X0Y1_DSP_bot.Inst_MULADD._0443_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0534_ sky130_fd_sc_hd__a221oi_4
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1296_ Tile_X0Y1_DSP_bot.Inst_MULADD._0365_ Tile_X0Y1_DSP_bot.Inst_MULADD._0377_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0390_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0466_
+ sky130_fd_sc_hd__a21oi_2
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[362\] Tile_X0Y0_DSP_top.ConfigBits\[363\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_118_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.NN4END_inbuf_6._0_ net318 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30 net252 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[318\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_133_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.N4BEG_outbuf_9._0_ Tile_X0Y0_DSP_top.N4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[9\] sky130_fd_sc_hd__buf_2
XFILLER_0_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_136_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1150_ Tile_X0Y1_DSP_bot.Inst_MULADD._0321_ Tile_X0Y1_DSP_bot.Inst_MULADD._0304_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0312_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0322_
+ sky130_fd_sc_hd__a21oi_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1081_ Tile_X0Y1_DSP_bot.Inst_MULADD._0238_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0253_ sky130_fd_sc_hd__inv_2
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_159_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[253\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_97_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0934_ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_ Tile_X0Y1_DSP_bot.Inst_MULADD._0073_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0108_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0109_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_155_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0865_ Tile_X0Y1_DSP_bot.B1 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0042_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst1
+ net81 net85 net133 net135 Tile_X0Y0_DSP_top.ConfigBits\[274\] Tile_X0Y0_DSP_top.ConfigBits\[275\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_142_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_6._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4END\[6\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12 net232 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[204\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1417_ Tile_X0Y1_DSP_bot.Inst_MULADD._0585_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 sky130_fd_sc_hd__buf_8
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23 net244 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[215\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1348_ Tile_X0Y1_DSP_bot.Inst_MULADD._0483_ Tile_X0Y1_DSP_bot.Inst_MULADD._0490_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0491_ Tile_X0Y1_DSP_bot.Inst_MULADD._0505_ Tile_X0Y1_DSP_bot.Inst_MULADD._0414_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0517_ sky130_fd_sc_hd__a32oi_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.cus_mux41_buf_inst0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG7
+ Tile_X0Y1_DSP_bot.ConfigBits\[153\] Tile_X0Y1_DSP_bot.ConfigBits\[154\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_147_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1279_ Tile_X0Y1_DSP_bot.Inst_MULADD._0101_ Tile_X0Y1_DSP_bot.Inst_MULADD._0132_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0261_ Tile_X0Y1_DSP_bot.Inst_MULADD._0263_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0449_ sky130_fd_sc_hd__o2bb2ai_4
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_9._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.W6BEG_outbuf_9._0_ Tile_X0Y0_DSP_top.W6BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[9\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5 net256 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[389\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG2 net297
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG4 net350 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5
+ Tile_X0Y1_DSP_bot.ConfigBits\[180\] Tile_X0Y1_DSP_bot.ConfigBits\[181\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_114_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[103\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_149_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_105_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1202_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B5
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ Tile_X0Y1_DSP_bot.Inst_MULADD._0208_ Tile_X0Y1_DSP_bot.Inst_MULADD._0372_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0373_ sky130_fd_sc_hd__o2111a_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END1
+ net24 net156 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG1 Tile_X0Y0_DSP_top.ConfigBits\[378\]
+ Tile_X0Y0_DSP_top.ConfigBits\[379\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1133_ Tile_X0Y1_DSP_bot.Inst_MULADD._0286_ Tile_X0Y1_DSP_bot.Inst_MULADD._0292_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0298_ Tile_X0Y1_DSP_bot.Inst_MULADD._0301_ Tile_X0Y1_DSP_bot.Inst_MULADD._0304_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0305_ sky130_fd_sc_hd__o221ai_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1064_ Tile_X0Y1_DSP_bot.Inst_MULADD._0236_ Tile_X0Y1_DSP_bot.Inst_MULADD._0221_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0222_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0237_
+ sky130_fd_sc_hd__a21oi_2
Xinput371 Tile_X0Y1_WW4END[14] VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__clkbuf_1
Xinput360 Tile_X0Y1_W6END[4] VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16 net236 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[112\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[326\] Tile_X0Y0_DSP_top.ConfigBits\[327\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27 net248 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[123\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_N1BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_EF_BEG2 Tile_X0Y0_DSP_top.ConfigBits\[2\]
+ Tile_X0Y0_DSP_top.ConfigBits\[3\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_128_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0917_ Tile_X0Y1_DSP_bot.Inst_MULADD._0060_ Tile_X0Y1_DSP_bot.Inst_MULADD._0092_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0093_ sky130_fd_sc_hd__xnor2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0848_ Tile_X0Y1_DSP_bot.ConfigBits\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0026_ sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.NN4END_inbuf_2._0_ Tile_X0Y0_DSP_top.NN4END\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG3 net294
+ net194 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG1 net347 Tile_X0Y1_DSP_bot.ConfigBits\[222\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[223\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_119_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.EE4BEG_outbuf_3._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_10._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.SS4BEG\[10\] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J_l_CD_BEG3 net301
+ Tile_X0Y0_DSP_top.SS4BEG\[0\] net354 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[398\] Tile_X0Y1_DSP_bot.ConfigBits\[399\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_114_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.data_inbuf_8._0_ net259 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG1.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[252\] Tile_X0Y0_DSP_top.ConfigBits\[253\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG1 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.data_outbuf_29._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[29\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[29\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11 net231 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[235\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22 net243 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[246\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1751_ net333 Tile_X0Y1_DSP_bot.C9 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1682_ Tile_X0Y1_DSP_bot.Inst_MULADD._0834_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0005_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_140_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_112_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._52_ net299 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END6
+ sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1116_ Tile_X0Y1_DSP_bot.Inst_MULADD._0272_ Tile_X0Y1_DSP_bot.Inst_MULADD._0259_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0287_ Tile_X0Y1_DSP_bot.Inst_MULADD._0195_ Tile_X0Y1_DSP_bot.Inst_MULADD._0275_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0288_ sky130_fd_sc_hd__a221oi_4
Xinput190 Tile_X0Y1_E2END[5] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1047_ Tile_X0Y1_DSP_bot.Inst_MULADD._0218_ Tile_X0Y1_DSP_bot.Inst_MULADD._0219_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0200_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0220_
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_inst0
+ net283 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2 net336 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.ConfigBits\[98\] Tile_X0Y1_DSP_bot.ConfigBits\[99\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_77_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.S4BEG_outbuf_9._0_ Tile_X0Y0_DSP_top.S4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput620 net620 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[14] sky130_fd_sc_hd__buf_2
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput631 net631 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[0] sky130_fd_sc_hd__buf_2
Xoutput642 net642 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput653 net653 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput664 net664 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[1] sky130_fd_sc_hd__buf_2
Xoutput675 net675 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput686 net686 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[12] sky130_fd_sc_hd__clkbuf_4
Xoutput697 net697 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[8] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2END_CD_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END0
+ net40 net85 net137 Tile_X0Y0_DSP_top.ConfigBits\[228\] Tile_X0Y0_DSP_top.ConfigBits\[229\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0 net229 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[192\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[290\] Tile_X0Y0_DSP_top.ConfigBits\[291\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[348\] Tile_X0Y1_DSP_bot.ConfigBits\[349\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
X_240_ Tile_X0Y1_DSP_bot.EE4BEG\[8\] VGND VGND VPWR VPWR net629 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_171_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb7 VGND VGND VPWR VPWR net554
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_134_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26 net247 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[154\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15 net235 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[143\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_99_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG0.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_74_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1734_ net333 Tile_X0Y1_DSP_bot.B0 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.B_reg\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_67_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_125_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_369_ Tile_X0Y1_DSP_bot.WW4BEG\[5\] VGND VGND VPWR VPWR net758 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1665_ Tile_X0Y1_DSP_bot.Inst_MULADD._0787_ Tile_X0Y1_DSP_bot.Inst_MULADD._0823_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0824_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1596_ Tile_X0Y1_DSP_bot.Inst_MULADD._0733_ Tile_X0Y1_DSP_bot.Inst_MULADD._0752_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0758_ Tile_X0Y1_DSP_bot.Inst_MULADD._0759_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0760_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.S4END_inbuf_1._0_ net112 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._35_ net198 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEGb\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.N4BEG_outbuf_10._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4END\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG4.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[274\] Tile_X0Y1_DSP_bot.ConfigBits\[275\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG4 sky130_fd_sc_hd__mux4_2
XFILLER_0_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput450 net450 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[28] sky130_fd_sc_hd__buf_2
Xoutput461 net461 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[9] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10 net230 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[266\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput472 net472 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[19] sky130_fd_sc_hd__clkbuf_4
Xoutput494 net494 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[0] sky130_fd_sc_hd__clkbuf_4
Xoutput483 net483 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[1] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21 net242 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[277\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.strobe_inbuf_1._0_ net272 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_154_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_223_ Tile_X0Y1_DSP_bot.E6BEG\[3\] VGND VGND VPWR VPWR net608 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG0 net292
+ net221 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb7 net345 Tile_X0Y1_DSP_bot.ConfigBits\[240\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[241\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.W6END_inbuf_5._0_ net162 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1450_ Tile_X0Y1_DSP_bot.Inst_MULADD._0570_ Tile_X0Y1_DSP_bot.Inst_MULADD._0616_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0617_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0618_
+ sky130_fd_sc_hd__o21ai_4
X_154_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG2 VGND VGND VPWR VPWR net537
+ sky130_fd_sc_hd__clkbuf_1
X_085_ Tile_X0Y0_DSP_top.FrameStrobe_O\[5\] VGND VGND VPWR VPWR net477 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1381_ Tile_X0Y1_DSP_bot.Inst_MULADD._0529_ Tile_X0Y1_DSP_bot.Inst_MULADD._0533_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_122_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5 net76 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[155\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_125_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1 net240 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[33\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1717_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0011_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[11\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1648_ Tile_X0Y1_DSP_bot.C18 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[18\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0808_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1579_ Tile_X0Y1_DSP_bot.Inst_MULADD._0741_ Tile_X0Y1_DSP_bot.Inst_MULADD._0743_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0744_ sky130_fd_sc_hd__and2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[312\] Tile_X0Y1_DSP_bot.ConfigBits\[313\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_70_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._18_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot14
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C16 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.S4END_inbuf_1._0_ Tile_X0Y0_DSP_top.S4BEG\[5\] VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.S4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._2_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_9._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[9\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14 net234 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[174\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25 net246 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[185\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3 net254 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[291\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0950_ Tile_X0Y1_DSP_bot.Inst_MULADD._0099_ Tile_X0Y1_DSP_bot.Inst_MULADD._0123_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0124_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0125_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_139_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0881_ Tile_X0Y1_DSP_bot.Inst_MULADD._0034_ Tile_X0Y1_DSP_bot.Inst_MULADD._0057_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0058_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_139_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_127_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_154_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_135_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1502_ Tile_X0Y1_DSP_bot.Inst_MULADD._0108_ Tile_X0Y1_DSP_bot.Inst_MULADD._0668_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0596_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0669_
+ sky130_fd_sc_hd__o21a_1
X_206_ Tile_X0Y1_DSP_bot.E2BEG\[2\] VGND VGND VPWR VPWR net589 sky130_fd_sc_hd__clkbuf_1
X_137_ Tile_X0Y0_DSP_top.NN4BEG\[1\] VGND VGND VPWR VPWR net525 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1433_ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0599_ Tile_X0Y1_DSP_bot.Inst_MULADD._0600_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0601_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.W6END_inbuf_5._0_ net363 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_068_ Tile_X0Y0_DSP_top.FrameData_O\[20\] VGND VGND VPWR VPWR net442 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1364_ Tile_X0Y1_DSP_bot.Inst_MULADD._0530_ Tile_X0Y1_DSP_bot.Inst_MULADD._0531_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0532_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0533_
+ sky130_fd_sc_hd__nand3_4
XFILLER_0_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1295_ Tile_X0Y1_DSP_bot.Inst_MULADD._0442_ Tile_X0Y1_DSP_bot.Inst_MULADD._0444_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0453_ Tile_X0Y1_DSP_bot.Inst_MULADD._0451_ Tile_X0Y1_DSP_bot.Inst_MULADD._0455_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0465_ sky130_fd_sc_hd__o2111a_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[362\] Tile_X0Y0_DSP_top.ConfigBits\[363\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_136_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31 net253 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[319\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20 net241 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[308\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_160_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.WW4END_inbuf_7._0_ net368 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1080_ Tile_X0Y1_DSP_bot.Inst_MULADD._0250_ Tile_X0Y1_DSP_bot.Inst_MULADD._0251_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0184_ Tile_X0Y1_DSP_bot.Inst_MULADD._0169_ Tile_X0Y1_DSP_bot.Inst_MULADD._0170_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0252_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_100_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_159_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[254\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._0933_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.A3
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0107_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0108_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_127_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_inst0
+ net281 net181 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[48\] Tile_X0Y1_DSP_bot.ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0864_ Tile_X0Y1_DSP_bot.Inst_MULADD._0040_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0041_ sky130_fd_sc_hd__buf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[274\] Tile_X0Y0_DSP_top.ConfigBits\[275\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_142_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_142_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_135_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1416_ Tile_X0Y1_DSP_bot.Inst_MULADD._0584_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0585_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13 net233 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[205\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24 net245 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[216\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1347_ Tile_X0Y1_DSP_bot.Inst_MULADD._0514_ Tile_X0Y1_DSP_bot.Inst_MULADD._0502_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0515_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0516_
+ sky130_fd_sc_hd__a21oi_2
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1278_ Tile_X0Y1_DSP_bot.Inst_MULADD._0203_ Tile_X0Y1_DSP_bot.Inst_MULADD._0447_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0269_ Tile_X0Y1_DSP_bot.Inst_MULADD._0270_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0448_ sky130_fd_sc_hd__o2bb2ai_2
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG7
+ Tile_X0Y1_DSP_bot.ConfigBits\[153\] Tile_X0Y1_DSP_bot.ConfigBits\[154\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_C9.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6 net257 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[390\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_EFa_BEG3 net193
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG0 net346 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG5
+ Tile_X0Y1_DSP_bot.ConfigBits\[182\] Tile_X0Y1_DSP_bot.ConfigBits\[183\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFa_BEG3 sky130_fd_sc_hd__mux4_1
XFILLER_0_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._2_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.cus_mux41_buf_out0
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG1.my_mux2_inst._0_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1201_ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_ Tile_X0Y1_DSP_bot.Inst_MULADD._0112_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_ Tile_X0Y1_DSP_bot.Inst_MULADD._0141_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0372_ sky130_fd_sc_hd__nand4_4
XFILLER_0_30_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1132_ Tile_X0Y1_DSP_bot.Inst_MULADD._0286_ Tile_X0Y1_DSP_bot.Inst_MULADD._0302_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0303_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0304_
+ sky130_fd_sc_hd__o21ai_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J_l_AB_BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END0
+ net21 net101 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1 Tile_X0Y0_DSP_top.ConfigBits\[380\]
+ Tile_X0Y0_DSP_top.ConfigBits\[381\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30 net252 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[350\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1063_ Tile_X0Y1_DSP_bot.Inst_MULADD._0227_ Tile_X0Y1_DSP_bot.Inst_MULADD._0228_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0235_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0236_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput350 Tile_X0Y1_W2MID[4] VGND VGND VPWR VPWR net350 sky130_fd_sc_hd__buf_2
Xinput372 Tile_X0Y1_WW4END[15] VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__clkbuf_1
Xinput361 Tile_X0Y1_W6END[5] VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17 net237 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[113\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28 net249 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[124\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[326\] Tile_X0Y0_DSP_top.ConfigBits\[327\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_133_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_N1BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_GH_BEG3 Tile_X0Y0_DSP_top.ConfigBits\[4\]
+ Tile_X0Y0_DSP_top.ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG2
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0916_ Tile_X0Y1_DSP_bot.Inst_MULADD._0090_ Tile_X0Y1_DSP_bot.Inst_MULADD._0091_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0092_ sky130_fd_sc_hd__or2b_1
XFILLER_0_42_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0847_ Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0025_ sky130_fd_sc_hd__buf_4
XFILLER_0_143_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.data_outbuf_1._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_146_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.data_inbuf_25._0_ net66 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[25\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.WW4END_inbuf_3._0_ net178 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._49_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG1
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG1 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12 net232 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[236\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23 net244 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[247\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1750_ net333 Tile_X0Y1_DSP_bot.C8 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1681_ Tile_X0Y1_DSP_bot.Inst_MULADD._0830_ Tile_X0Y1_DSP_bot.Inst_MULADD._0247_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0834_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._51_ net298 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END5
+ sky130_fd_sc_hd__buf_2
XFILLER_0_120_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.data_inbuf_16._0_ net56 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1115_ Tile_X0Y1_DSP_bot.Inst_MULADD._0193_ Tile_X0Y1_DSP_bot.Inst_MULADD._0197_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0287_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1046_ Tile_X0Y1_DSP_bot.Inst_MULADD._0193_ Tile_X0Y1_DSP_bot.Inst_MULADD._0195_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0197_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0219_
+ sky130_fd_sc_hd__a21o_1
Xinput180 Tile_X0Y0_WW4END[9] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_GH_BEG2
+ Tile_X0Y1_DSP_bot.ConfigBits\[98\] Tile_X0Y1_DSP_bot.ConfigBits\[99\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_WW4BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
Xinput191 Tile_X0Y1_E2END[6] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__buf_2
XFILLER_0_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_131_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput610 net610 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput621 net621 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xoutput632 net632 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[10] sky130_fd_sc_hd__buf_2
Xoutput643 net643 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[20] sky130_fd_sc_hd__buf_2
Xoutput654 net654 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[30] sky130_fd_sc_hd__buf_2
XFILLER_0_78_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput665 net665 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[2] sky130_fd_sc_hd__buf_2
Xoutput676 net676 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput687 net687 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[13] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.data_outbuf_1._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[1\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[1\] sky130_fd_sc_hd__clkbuf_1
Xoutput698 net698 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[9] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net3 net135 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.ConfigBits\[16\] Tile_X0Y0_DSP_top.ConfigBits\[17\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1 net240 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[193\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG3.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[292\] Tile_X0Y0_DSP_top.ConfigBits\[293\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JE2BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_49_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[374\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_119_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_170_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb6 VGND VGND VPWR VPWR net553
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9 Tile_X0Y1_DSP_bot.ConfigBits\[348\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[349\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst0
+ net281 net287 net309 net187 Tile_X0Y1_DSP_bot.ConfigBits\[292\] Tile_X0Y1_DSP_bot.ConfigBits\[293\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27 net248 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[155\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16 net236 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[144\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_20_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.SS4END_inbuf_9._0_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.SS4BEG1
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.SS4BEG_i\[9\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.data_inbuf_25._0_ net246 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[25\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_230 Tile_X0Y1_DSP_bot.SS4BEG_i\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1733_ net333 Tile_X0Y1_DSP_bot.A7 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_125_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_368_ Tile_X0Y1_DSP_bot.WW4BEG\[4\] VGND VGND VPWR VPWR net757 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1664_ Tile_X0Y1_DSP_bot.Inst_MULADD._0822_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0823_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1595_ Tile_X0Y1_DSP_bot.Inst_MULADD._0750_ Tile_X0Y1_DSP_bot.Inst_MULADD._0751_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0759_ sky130_fd_sc_hd__nor2_1
X_299_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb7 VGND VGND VPWR VPWR net682
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._34_ net197 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEGb\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.strobe_outbuf_2._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[2\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1029_ Tile_X0Y1_DSP_bot.B4 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0202_
+ sky130_fd_sc_hd__inv_2
XTile_X0Y1_DSP_bot.data_inbuf_16._0_ net236 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput462 net462 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput451 net451 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[29] sky130_fd_sc_hd__clkbuf_4
Xoutput440 net440 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[19] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11 net231 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[267\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput473 net473 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput495 net495 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[1] sky130_fd_sc_hd__clkbuf_4
Xoutput484 net484 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22 net243 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[278\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END1
+ net6 net24 Tile_X0Y0_DSP_top.ConfigBits\[342\] Tile_X0Y0_DSP_top.ConfigBits\[343\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_154_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_222_ Tile_X0Y1_DSP_bot.E6BEG\[2\] VGND VGND VPWR VPWR net607 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_147_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG1 net288
+ net188 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb3 net373 Tile_X0Y1_DSP_bot.ConfigBits\[242\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[243\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_52_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_153_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG1 VGND VGND VPWR VPWR net536
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_084_ Tile_X0Y0_DSP_top.FrameStrobe_O\[4\] VGND VGND VPWR VPWR net476 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1380_ Tile_X0Y1_DSP_bot.Inst_MULADD._0535_ Tile_X0Y1_DSP_bot.Inst_MULADD._0539_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0548_ Tile_X0Y1_DSP_bot.Inst_MULADD._0534_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0549_ sky130_fd_sc_hd__o22ai_4
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.EE4END_inbuf_8._0_ net216 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.WW4BEG_outbuf_0._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[0\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[0\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.strobe_inbuf_17._0_ Tile_X0Y0_DSP_top.FrameStrobe\[17\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[17\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6 net77 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[156\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_157_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2 net251 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[34\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_157_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_126_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1716_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0010_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[10\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_153_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1647_ Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[17\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0807_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q17
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1578_ Tile_X0Y1_DSP_bot.Inst_MULADD._0736_ Tile_X0Y1_DSP_bot.Inst_MULADD._0737_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0742_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0743_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_3_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG6.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[314\] Tile_X0Y1_DSP_bot.ConfigBits\[315\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG6 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._17_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot13
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15 net235 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[175\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_78_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26 net247 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[186\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_148_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_129_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4 net255 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[292\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_144_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.strobe_inbuf_10._0_ net262 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[10\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_E1BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_CDb_BEG3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_CD_BEG1 Tile_X0Y1_DSP_bot.ConfigBits\[34\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[35\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E1BEG\[0\]
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.SS4END_inbuf_5._0_ net132 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0880_ Tile_X0Y1_DSP_bot.Inst_MULADD._0055_ Tile_X0Y1_DSP_bot.Inst_MULADD._0056_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0057_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1501_ Tile_X0Y1_DSP_bot.Inst_MULADD._0594_ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0668_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.strobe_outbuf_19._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[19\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[19\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_205_ Tile_X0Y1_DSP_bot.E2BEG\[1\] VGND VGND VPWR VPWR net588 sky130_fd_sc_hd__clkbuf_1
X_136_ Tile_X0Y0_DSP_top.NN4BEG\[0\] VGND VGND VPWR VPWR net518 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_135_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1432_ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_ Tile_X0Y1_DSP_bot.Inst_MULADD._0536_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0359_ Tile_X0Y1_DSP_bot.Inst_MULADD._0154_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0600_ sky130_fd_sc_hd__o2bb2ai_1
XFILLER_0_20_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_067_ Tile_X0Y0_DSP_top.FrameData_O\[19\] VGND VGND VPWR VPWR net440 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1363_ Tile_X0Y1_DSP_bot.Inst_MULADD._0071_ Tile_X0Y1_DSP_bot.Inst_MULADD._0441_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0521_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0532_
+ sky130_fd_sc_hd__and3_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1294_ Tile_X0Y1_DSP_bot.Inst_MULADD._0455_ Tile_X0Y1_DSP_bot.Inst_MULADD._0457_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0463_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0464_
+ sky130_fd_sc_hd__a21oi_4
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG5.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[364\] Tile_X0Y0_DSP_top.ConfigBits\[365\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG5 sky130_fd_sc_hd__mux4_2
XFILLER_0_136_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst0
+ net283 net289 net189 net201 Tile_X0Y1_DSP_bot.ConfigBits\[364\] Tile_X0Y1_DSP_bot.ConfigBits\[365\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst0
+ net4 net136 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.ConfigBits\[104\] Tile_X0Y0_DSP_top.ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10 net230 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[298\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21 net242 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[309\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_9_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_141_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.EE4END_inbuf_4._0_ net47 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_159_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0932_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[3\] Tile_X0Y1_DSP_bot.Inst_MULADD._0026_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0107_ sky130_fd_sc_hd__or2b_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[4\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[255\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame4_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_155_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_inst1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_CD_BEG0
+ Tile_X0Y1_DSP_bot.ConfigBits\[48\] Tile_X0Y1_DSP_bot.ConfigBits\[49\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_38_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0863_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.Inst_MULADD._0038_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0039_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0040_
+ sky130_fd_sc_hd__o21ai_4
XFILLER_0_155_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_24 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[274\] Tile_X0Y0_DSP_top.ConfigBits\[275\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_127_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_122_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_119_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb7 VGND VGND VPWR VPWR net501
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.strobe_outbuf_8._0_ Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[8\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe\[8\] sky130_fd_sc_hd__clkbuf_16
XTile_X0Y1_DSP_bot.Inst_MULADD._1415_ Tile_X0Y1_DSP_bot.Inst_MULADD._0582_ Tile_X0Y1_DSP_bot.Inst_MULADD._0583_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0584_ sky130_fd_sc_hd__or2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14 net234 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[206\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25 net246 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[217\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1346_ Tile_X0Y1_DSP_bot.Inst_MULADD._0501_ Tile_X0Y1_DSP_bot.Inst_MULADD._0497_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0496_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0515_
+ sky130_fd_sc_hd__nor3_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1277_ Tile_X0Y1_DSP_bot.Inst_MULADD._0079_ Tile_X0Y1_DSP_bot.B4
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0447_ sky130_fd_sc_hd__or2b_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.N4BEG_outbuf_3._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END3 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_N4BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END1 net24 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[8\] Tile_X0Y0_DSP_top.ConfigBits\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 sky130_fd_sc_hd__mux4_2
XFILLER_0_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_146_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_114_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7 net258 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[391\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_137_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_124_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1200_ Tile_X0Y1_DSP_bot.Inst_MULADD._0367_ Tile_X0Y1_DSP_bot.Inst_MULADD._0368_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0369_ Tile_X0Y1_DSP_bot.Inst_MULADD._0370_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0371_ sky130_fd_sc_hd__o211ai_4
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_6._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[6\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1131_ Tile_X0Y1_DSP_bot.Inst_MULADD._0227_ Tile_X0Y1_DSP_bot.Inst_MULADD._0228_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0216_ Tile_X0Y1_DSP_bot.Inst_MULADD._0220_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0303_ sky130_fd_sc_hd__o22a_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31 net253 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[351\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20 net241 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[340\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1062_ Tile_X0Y1_DSP_bot.Inst_MULADD._0233_ Tile_X0Y1_DSP_bot.Inst_MULADD._0234_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0216_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0235_
+ sky130_fd_sc_hd__a21oi_4
Xinput340 Tile_X0Y1_W2END[2] VGND VGND VPWR VPWR net340 sky130_fd_sc_hd__buf_2
Xinput351 Tile_X0Y1_W2MID[5] VGND VGND VPWR VPWR net351 sky130_fd_sc_hd__buf_2
Xinput362 Tile_X0Y1_W6END[6] VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__clkbuf_1
Xinput373 Tile_X0Y1_WW4END[1] VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18 net238 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[114\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29 net250 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[125\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG4.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[328\] Tile_X0Y0_DSP_top.ConfigBits\[329\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JS2BEG4 sky130_fd_sc_hd__mux4_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_N1BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J_l_AB_BEG0 Tile_X0Y0_DSP_top.ConfigBits\[6\]
+ Tile_X0Y0_DSP_top.ConfigBits\[7\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1BEG3
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_85_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0915_ Tile_X0Y1_DSP_bot.Inst_MULADD._0084_ Tile_X0Y1_DSP_bot.Inst_MULADD._0089_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0091_ sky130_fd_sc_hd__nand2_1
XTile_X0Y0_DSP_top.E6BEG_outbuf_8._0_ Tile_X0Y0_DSP_top.E6BEG_i\[8\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.E6BEG\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst0
+ net326 net182 net188 net204 Tile_X0Y1_DSP_bot.ConfigBits\[328\] Tile_X0Y1_DSP_bot.ConfigBits\[329\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_42_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._0846_ Tile_X0Y1_DSP_bot.ConfigBits\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0024_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_297 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_115_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.strobe_outbuf_14._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[14\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.W6BEG_outbuf_3._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1329_ Tile_X0Y1_DSP_bot.C8 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[8\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0499_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y0_DSP_top.data_inbuf_5._0_ net76 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_121_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.N4END_inbuf_1._0_ Tile_X0Y0_DSP_top.N4END\[5\] VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_i\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._48_ net137 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEG0
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13 net233 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[237\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24 net245 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[248\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_103_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1680_ Tile_X0Y1_DSP_bot.Inst_MULADD._0833_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0004_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._50_ net297 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END4
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_50_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_120_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1114_ Tile_X0Y1_DSP_bot.Inst_MULADD._0255_ Tile_X0Y1_DSP_bot.Inst_MULADD._0276_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0281_ Tile_X0Y1_DSP_bot.Inst_MULADD._0284_ Tile_X0Y1_DSP_bot.Inst_MULADD._0285_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0286_ sky130_fd_sc_hd__o2111a_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1045_ Tile_X0Y1_DSP_bot.Inst_MULADD._0190_ Tile_X0Y1_DSP_bot.Inst_MULADD._0193_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0218_ sky130_fd_sc_hd__nand2_1
Xinput170 Tile_X0Y0_WW4END[14] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
Xinput181 Tile_X0Y1_E1END[0] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xinput192 Tile_X0Y1_E2END[7] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_144_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_128_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_131_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput600 net600 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput611 net611 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[6] sky130_fd_sc_hd__buf_2
XTile_X0Y0_DSP_top.NN4BEG_outbuf_3._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput622 net622 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput633 net633 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput644 net644 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[21] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput666 net666 VGND VGND VPWR VPWR Tile_X0Y1_S1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput677 net677 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xoutput688 net688 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[14] sky130_fd_sc_hd__clkbuf_4
Xoutput655 net655 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[31] sky130_fd_sc_hd__clkbuf_4
Xoutput699 net699 VGND VGND VPWR VPWR Tile_X0Y1_SS4BEG[0] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG0 net300
+ net200 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG7 net353 Tile_X0Y1_DSP_bot.ConfigBits\[192\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[193\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG1
+ Tile_X0Y0_DSP_top.ConfigBits\[16\] Tile_X0Y0_DSP_top.ConfigBits\[17\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_96_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_119_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2 net251 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[194\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.SS4BEG_outbuf_6._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[375\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_107_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG7.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[350\] Tile_X0Y1_DSP_bot.ConfigBits\[351\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG7 sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30 net252 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[382\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_91_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst1
+ net201 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb2 net340 net375 Tile_X0Y1_DSP_bot.ConfigBits\[292\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[293\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_outbuf_23._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[23\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[23\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28 net249 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[156\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17 net237 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[145\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END0 net81 net133 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[98\] Tile_X0Y0_DSP_top.ConfigBits\[99\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_32_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.N4END_inbuf_1._0_ net312 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.S4BEG_outbuf_10._0_ Tile_X0Y0_DSP_top.S4BEG_i\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_157_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_220 Tile_X0Y0_DSP_top.S4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_157_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1732_ net333 Tile_X0Y1_DSP_bot.A6 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_128_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1663_ Tile_X0Y1_DSP_bot.C19 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[19\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0822_
+ sky130_fd_sc_hd__mux2_1
X_367_ Tile_X0Y1_DSP_bot.WW4BEG\[3\] VGND VGND VPWR VPWR net756 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_113_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1594_ Tile_X0Y1_DSP_bot.Inst_MULADD._0756_ Tile_X0Y1_DSP_bot.Inst_MULADD._0757_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0758_ sky130_fd_sc_hd__nand2_1
X_298_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb6 VGND VGND VPWR VPWR net681
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.data_outbuf_14._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[14\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[14\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._33_ net196 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEGb\[3\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_139_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.S4BEG_outbuf_3._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1028_ Tile_X0Y1_DSP_bot.Inst_MULADD._0193_ Tile_X0Y1_DSP_bot.Inst_MULADD._0190_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0198_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0201_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput452 net452 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[2] sky130_fd_sc_hd__buf_2
Xoutput441 net441 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput430 net430 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[0] sky130_fd_sc_hd__clkbuf_4
Xoutput474 net474 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[2] sky130_fd_sc_hd__clkbuf_4
Xoutput485 net485 VGND VGND VPWR VPWR Tile_X0Y0_N1BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput463 net463 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[10] sky130_fd_sc_hd__clkbuf_4
Xoutput496 net496 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[2] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12 net232 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[268\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23 net244 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[279\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst1
+ net86 net108 net138 net156 Tile_X0Y0_DSP_top.ConfigBits\[342\] Tile_X0Y0_DSP_top.ConfigBits\[343\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_221_ Tile_X0Y1_DSP_bot.E6BEG\[1\] VGND VGND VPWR VPWR net606 sky130_fd_sc_hd__clkbuf_1
X_152_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W1BEG0 VGND VGND VPWR VPWR net535
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG2 net290
+ net190 Tile_X0Y0_DSP_top.SS4BEG\[1\] net343 Tile_X0Y1_DSP_bot.ConfigBits\[244\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[245\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG2
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_083_ Tile_X0Y0_DSP_top.FrameStrobe_O\[3\] VGND VGND VPWR VPWR net475 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7 net78 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[157\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_157_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3 net254 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[35\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1715_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0009_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[9\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_141_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1646_ Tile_X0Y1_DSP_bot.Inst_MULADD._0805_ Tile_X0Y1_DSP_bot.Inst_MULADD._0806_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0807_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_113_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1577_ Tile_X0Y1_DSP_bot.Inst_MULADD._0739_ Tile_X0Y1_DSP_bot.Inst_MULADD._0740_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._16_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot12
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16 net236 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[176\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27 net248 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[187\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_78_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.NN4END_inbuf_9._0_ net321 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.NN4BEG_i\[9\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END3
+ net2 net8 Tile_X0Y0_DSP_top.ConfigBits\[254\] Tile_X0Y0_DSP_top.ConfigBits\[255\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_74_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5 net256 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[293\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_46_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_E1BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_EFb_BEG0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_EF_BEG2 Tile_X0Y1_DSP_bot.ConfigBits\[36\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[37\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E1BEG\[1\]
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_100_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1500_ Tile_X0Y1_DSP_bot.Inst_MULADD._0664_ Tile_X0Y1_DSP_bot.Inst_MULADD._0665_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0666_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0667_
+ sky130_fd_sc_hd__o21ai_2
X_204_ Tile_X0Y1_DSP_bot.E2BEG\[0\] VGND VGND VPWR VPWR net587 sky130_fd_sc_hd__buf_1
XFILLER_0_37_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_135_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 VGND VGND VPWR VPWR net508
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1431_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_ Tile_X0Y1_DSP_bot.Inst_MULADD._0357_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0599_ sky130_fd_sc_hd__nand4_4
XFILLER_0_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_150_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_066_ Tile_X0Y0_DSP_top.FrameData_O\[18\] VGND VGND VPWR VPWR net439 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 net3 net135 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.ConfigBits\[72\] Tile_X0Y0_DSP_top.ConfigBits\[73\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1362_ Tile_X0Y1_DSP_bot.Inst_MULADD._0192_ Tile_X0Y1_DSP_bot.Inst_MULADD._0527_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0295_ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ Tile_X0Y1_DSP_bot.Inst_MULADD._0523_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0531_ sky130_fd_sc_hd__o2111ai_4
XTile_X0Y0_DSP_top.data_outbuf_10._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1293_ Tile_X0Y1_DSP_bot.Inst_MULADD._0450_ Tile_X0Y1_DSP_bot.Inst_MULADD._0446_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0462_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0463_
+ sky130_fd_sc_hd__a21oi_4
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb4 Tile_X0Y0_DSP_top.S4BEG\[0\]
+ net342 net354 Tile_X0Y1_DSP_bot.ConfigBits\[364\] Tile_X0Y1_DSP_bot.ConfigBits\[365\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[104\] Tile_X0Y0_DSP_top.ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11 net231 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[299\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22 net243 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[310\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.NN4BEG_outbuf_9._0_ Tile_X0Y1_DSP_bot.NN4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4END\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_126_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_327 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1629_ Tile_X0Y1_DSP_bot.Inst_MULADD._0741_ Tile_X0Y1_DSP_bot.Inst_MULADD._0763_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0764_ Tile_X0Y1_DSP_bot.Inst_MULADD._0767_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0791_ sky130_fd_sc_hd__nand4_1
XFILLER_0_31_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_149_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_151_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0931_ Tile_X0Y1_DSP_bot.Inst_MULADD._0044_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0106_ sky130_fd_sc_hd__buf_6
XFILLER_0_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_155_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0862_ Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[1\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG7.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[276\] Tile_X0Y0_DSP_top.ConfigBits\[277\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JN2BEG7 sky130_fd_sc_hd__mux4_2
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_118_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb6 VGND VGND VPWR VPWR net500
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst0
+ net283 net291 net183 net191 Tile_X0Y1_DSP_bot.ConfigBits\[276\] Tile_X0Y1_DSP_bot.ConfigBits\[277\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1414_ Tile_X0Y1_DSP_bot.Inst_MULADD._0579_ Tile_X0Y1_DSP_bot.Inst_MULADD._0581_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0516_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0583_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_150_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_049_ Tile_X0Y0_DSP_top.FrameData_O\[1\] VGND VGND VPWR VPWR net441 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15 net235 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[207\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26 net247 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[218\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1345_ Tile_X0Y1_DSP_bot.Inst_MULADD._0341_ Tile_X0Y1_DSP_bot.Inst_MULADD._0508_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0509_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0514_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1276_ Tile_X0Y1_DSP_bot.Inst_MULADD._0103_ Tile_X0Y1_DSP_bot.Inst_MULADD._0379_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ Tile_X0Y1_DSP_bot.Inst_MULADD._0231_ Tile_X0Y1_DSP_bot.Inst_MULADD._0445_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0446_ sky130_fd_sc_hd__a41oi_4
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_N4BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END2 net21 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5
+ Tile_X0Y0_DSP_top.ConfigBits\[10\] Tile_X0Y0_DSP_top.ConfigBits\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 sky130_fd_sc_hd__mux4_1
XFILLER_0_146_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.NN4END_inbuf_5._0_ Tile_X0Y0_DSP_top.NN4END\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[5\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8 net259 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[392\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_71_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0 net229 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[96\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.EE4BEG_outbuf_6._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_152_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_120_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1130_ Tile_X0Y1_DSP_bot.Inst_MULADD._0288_ Tile_X0Y1_DSP_bot.Inst_MULADD._0289_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0290_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0302_
+ sky130_fd_sc_hd__o21a_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10 net230 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[330\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput330 Tile_X0Y1_NN4END[7] VGND VGND VPWR VPWR net330 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21 net242 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[341\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1061_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ Tile_X0Y1_DSP_bot.Inst_MULADD._0050_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0108_ Tile_X0Y1_DSP_bot.Inst_MULADD._0137_ Tile_X0Y1_DSP_bot.Inst_MULADD._0194_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0234_ sky130_fd_sc_hd__o41a_1
Xinput341 Tile_X0Y1_W2END[3] VGND VGND VPWR VPWR net341 sky130_fd_sc_hd__clkbuf_4
Xinput352 Tile_X0Y1_W2MID[6] VGND VGND VPWR VPWR net352 sky130_fd_sc_hd__clkbuf_4
Xinput363 Tile_X0Y1_W6END[7] VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__clkbuf_1
Xinput374 Tile_X0Y1_WW4END[2] VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__buf_2
XFILLER_0_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19 net239 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[115\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_85_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0914_ Tile_X0Y1_DSP_bot.Inst_MULADD._0084_ Tile_X0Y1_DSP_bot.Inst_MULADD._0089_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0090_ sky130_fd_sc_hd__nor2_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb3 Tile_X0Y0_DSP_top.S4BEG\[3\]
+ net341 net357 Tile_X0Y1_DSP_bot.ConfigBits\[328\] Tile_X0Y1_DSP_bot.ConfigBits\[329\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0845_ Tile_X0Y1_DSP_bot.Inst_MULADD._0022_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[0\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[3\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0023_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_143_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_143_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 Tile_X0Y0_DSP_top.E6BEG_i\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_123_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1328_ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ sky130_fd_sc_hd__buf_4
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1259_ Tile_X0Y1_DSP_bot.Inst_MULADD._0051_ Tile_X0Y1_DSP_bot.Inst_MULADD._0300_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0297_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0429_
+ sky130_fd_sc_hd__or3_2
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._47_ net100 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb7
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_67_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14 net234 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[238\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25 net246 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[249\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1113_ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0282_ Tile_X0Y1_DSP_bot.Inst_MULADD._0283_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0285_ sky130_fd_sc_hd__nand4_4
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1044_ Tile_X0Y1_DSP_bot.Inst_MULADD._0200_ Tile_X0Y1_DSP_bot.Inst_MULADD._0201_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0216_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0217_
+ sky130_fd_sc_hd__o21bai_4
Xinput160 Tile_X0Y0_W6END[5] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__clkbuf_1
Xinput171 Tile_X0Y0_WW4END[15] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
Xinput182 Tile_X0Y1_E1END[1] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_4
Xinput193 Tile_X0Y1_E2MID[0] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_2
XFILLER_0_128_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_160_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_128_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.S4END_inbuf_4._0_ net115 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[4\]
+ sky130_fd_sc_hd__buf_2
Xoutput601 net601 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput623 net623 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[2] sky130_fd_sc_hd__buf_2
Xoutput612 net612 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput634 net634 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput645 net645 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[22] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput678 net678 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[3] sky130_fd_sc_hd__buf_2
Xoutput667 net667 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[0] sky130_fd_sc_hd__buf_2
Xoutput656 net656 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[3] sky130_fd_sc_hd__clkbuf_4
Xoutput689 net689 VGND VGND VPWR VPWR Tile_X0Y1_S4BEG[15] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG1 net296
+ net196 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG3 net349 Tile_X0Y1_DSP_bot.ConfigBits\[194\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[195\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG1
+ sky130_fd_sc_hd__mux4_2
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3 net254 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[195\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_64_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[376\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_107_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31 net253 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[383\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20 net241 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[372\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[292\] Tile_X0Y1_DSP_bot.ConfigBits\[293\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_134_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_122_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29 net250 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[157\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18 net238 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[146\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_CD_BEG2
+ Tile_X0Y0_DSP_top.ConfigBits\[98\] Tile_X0Y0_DSP_top.ConfigBits\[99\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_WW4BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.strobe_inbuf_4._0_ net275 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_157_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_210 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_221 Tile_X0Y0_DSP_top.S4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1731_ net333 Tile_X0Y1_DSP_bot.A5 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_111 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.W6END_inbuf_8._0_ net154 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.W6BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_1
X_366_ Tile_X0Y1_DSP_bot.WW4BEG\[2\] VGND VGND VPWR VPWR net755 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1662_ Tile_X0Y1_DSP_bot.Inst_MULADD._0775_ Tile_X0Y1_DSP_bot.Inst_MULADD._0809_
+ Tile_X0Y1_DSP_bot.ConfigBits\[4\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0821_
+ sky130_fd_sc_hd__and3_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1593_ Tile_X0Y1_DSP_bot.Inst_MULADD._0733_ Tile_X0Y1_DSP_bot.Inst_MULADD._0734_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0713_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0757_
+ sky130_fd_sc_hd__nor3_1
X_297_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb5 VGND VGND VPWR VPWR net680
+ sky130_fd_sc_hd__buf_1
XFILLER_0_70_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._32_ net195 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEGb\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1027_ Tile_X0Y1_DSP_bot.Inst_MULADD._0146_ Tile_X0Y1_DSP_bot.Inst_MULADD._0194_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0200_ sky130_fd_sc_hd__nand2_2
XFILLER_0_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput420 net420 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[15] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_112_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput453 net453 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[30] sky130_fd_sc_hd__clkbuf_4
Xoutput442 net442 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[20] sky130_fd_sc_hd__clkbuf_4
Xoutput431 net431 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[10] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.S4END_inbuf_4._0_ Tile_X0Y0_DSP_top.S4BEG\[8\] VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.S4BEG_i\[4\] sky130_fd_sc_hd__clkbuf_1
Xoutput464 net464 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput475 net475 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[3] sky130_fd_sc_hd__clkbuf_4
Xoutput486 net486 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[0] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13 net233 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[269\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24 net245 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[280\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput497 net497 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[342\] Tile_X0Y0_DSP_top.ConfigBits\[343\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_220_ Tile_X0Y1_DSP_bot.E6BEG\[0\] VGND VGND VPWR VPWR net603 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_151_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 VGND VGND VPWR VPWR net524
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2END_EF_BEG3 net325
+ net186 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb1 net339 Tile_X0Y1_DSP_bot.ConfigBits\[246\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[247\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2END_EF_BEG3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_082_ Tile_X0Y0_DSP_top.FrameStrobe_O\[2\] VGND VGND VPWR VPWR net474 sky130_fd_sc_hd__buf_1
XFILLER_0_122_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8 net79 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[158\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4 net255 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[36\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_141_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1714_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0008_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_153_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_349_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb5 VGND VGND VPWR VPWR net732
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.W6END_inbuf_8._0_ net355 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.W6BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1645_ Tile_X0Y1_DSP_bot.Inst_MULADD._0798_ Tile_X0Y1_DSP_bot.Inst_MULADD._0799_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0802_ Tile_X0Y1_DSP_bot.Inst_MULADD._0804_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0806_ sky130_fd_sc_hd__nand4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1576_ Tile_X0Y1_DSP_bot.Inst_MULADD._0736_ Tile_X0Y1_DSP_bot.Inst_MULADD._0737_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0739_ Tile_X0Y1_DSP_bot.Inst_MULADD._0740_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0741_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_59_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._15_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot11
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C13 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30 net252 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[414\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_75_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28 net249 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[188\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17 net237 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[177\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst1
+ net24 net88 net140 net172 Tile_X0Y0_DSP_top.ConfigBits\[254\] Tile_X0Y0_DSP_top.ConfigBits\[255\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_129_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6 net257 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[294\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_E1BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_GHb_BEG1 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_GH_BEG3 Tile_X0Y1_DSP_bot.ConfigBits\[38\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[39\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E1BEG\[2\]
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_61_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.strobe_inbuf_0._0_ Tile_X0Y0_DSP_top.FrameStrobe\[0\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O_i\[0\] sky130_fd_sc_hd__buf_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_139_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_139_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_203_ Tile_X0Y1_DSP_bot.E1BEG\[3\] VGND VGND VPWR VPWR net586 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_135_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_134_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 VGND VGND VPWR VPWR net507
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1430_ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_ Tile_X0Y1_DSP_bot.Inst_MULADD._0596_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0348_ Tile_X0Y1_DSP_bot.Inst_MULADD._0594_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0598_ sky130_fd_sc_hd__nand4_4
X_065_ Tile_X0Y0_DSP_top.FrameData_O\[17\] VGND VGND VPWR VPWR net438 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2END_GH_BEG3
+ Tile_X0Y0_DSP_top.ConfigBits\[72\] Tile_X0Y0_DSP_top.ConfigBits\[73\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_SS4BEG0.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1361_ Tile_X0Y1_DSP_bot.Inst_MULADD._0230_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0523_ Tile_X0Y1_DSP_bot.Inst_MULADD._0524_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_150_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1292_ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0450_ Tile_X0Y1_DSP_bot.Inst_MULADD._0452_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0462_ sky130_fd_sc_hd__a22oi_4
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[104\] Tile_X0Y0_DSP_top.ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.ConfigBits\[364\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[365\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_152_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12 net232 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[300\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23 net244 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[311\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_145_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1628_ Tile_X0Y1_DSP_bot.Inst_MULADD._0787_ Tile_X0Y1_DSP_bot.Inst_MULADD._0789_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0790_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_141_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1559_ Tile_X0Y1_DSP_bot.Inst_MULADD._0724_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q12 sky130_fd_sc_hd__buf_1
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END5
+ net2 net10 Tile_X0Y0_DSP_top.ConfigBits\[294\] Tile_X0Y0_DSP_top.ConfigBits\[295\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0930_ Tile_X0Y1_DSP_bot.Inst_MULADD._0072_ Tile_X0Y1_DSP_bot.Inst_MULADD._0076_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0104_ Tile_X0Y1_DSP_bot.Inst_MULADD._0066_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0105_ sky130_fd_sc_hd__o2bb2ai_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0861_ Tile_X0Y1_DSP_bot.A1 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0038_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_155_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_117_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 VGND VGND VPWR VPWR net499
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb6
+ net334 net336 Tile_X0Y1_DSP_bot.ConfigBits\[276\] Tile_X0Y1_DSP_bot.ConfigBits\[277\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1413_ Tile_X0Y1_DSP_bot.Inst_MULADD._0516_ Tile_X0Y1_DSP_bot.Inst_MULADD._0579_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0581_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0582_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_123_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_048_ Tile_X0Y0_DSP_top.FrameData_O\[0\] VGND VGND VPWR VPWR net430 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27 net248 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[219\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16 net236 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[208\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1344_ Tile_X0Y1_DSP_bot.Inst_MULADD._0428_ Tile_X0Y1_DSP_bot.Inst_MULADD._0511_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0512_ Tile_X0Y1_DSP_bot.Inst_MULADD._0513_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 sky130_fd_sc_hd__a31o_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1275_ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_ Tile_X0Y1_DSP_bot.Inst_MULADD._0213_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0445_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_N4BEG2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END3 net156 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.ConfigBits\[12\] Tile_X0Y0_DSP_top.ConfigBits\[13\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG2 sky130_fd_sc_hd__mux4_1
XFILLER_0_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_158_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_118_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_133_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.data_outbuf_4._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[4\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_112_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9 net260 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[393\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._63_ net152 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb7
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1 net240 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[97\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0 net49 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[278\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit0/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_1_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.data_inbuf_28._0_ net69 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[28\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.WW4END_inbuf_6._0_ net166 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG_i\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1060_ Tile_X0Y1_DSP_bot.Inst_MULADD._0229_ Tile_X0Y1_DSP_bot.Inst_MULADD._0232_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0219_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0233_
+ sky130_fd_sc_hd__o21ai_1
Xinput320 Tile_X0Y1_NN4END[12] VGND VGND VPWR VPWR net320 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11 net231 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[331\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22 net243 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[342\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput342 Tile_X0Y1_W2END[4] VGND VGND VPWR VPWR net342 sky130_fd_sc_hd__clkbuf_4
Xinput353 Tile_X0Y1_W2MID[7] VGND VGND VPWR VPWR net353 sky130_fd_sc_hd__clkbuf_4
Xinput331 Tile_X0Y1_NN4END[8] VGND VGND VPWR VPWR net331 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst0
+ net281 net285 net181 net185 Tile_X0Y1_DSP_bot.ConfigBits\[316\] Tile_X0Y1_DSP_bot.ConfigBits\[317\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
Xinput375 Tile_X0Y1_WW4END[3] VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_26_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput364 Tile_X0Y1_W6END[8] VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_194 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0913_ Tile_X0Y1_DSP_bot.Inst_MULADD._0085_ Tile_X0Y1_DSP_bot.Inst_MULADD._0087_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0088_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0089_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4
+ Tile_X0Y1_DSP_bot.ConfigBits\[328\] Tile_X0Y1_DSP_bot.ConfigBits\[329\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0844_ Tile_X0Y1_DSP_bot.C0 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[0\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[2\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0022_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_2 Tile_X0Y0_DSP_top.FrameStrobe\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top.data_inbuf_19._0_ net59 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[19\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1327_ Tile_X0Y1_DSP_bot.Inst_MULADD._0494_ Tile_X0Y1_DSP_bot.Inst_MULADD._0495_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0435_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0497_
+ sky130_fd_sc_hd__a21oi_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1258_ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0428_ sky130_fd_sc_hd__inv_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1189_ Tile_X0Y1_DSP_bot.Inst_MULADD._0106_ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0359_ Tile_X0Y1_DSP_bot.Inst_MULADD._0048_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0360_ sky130_fd_sc_hd__o2bb2ai_2
XFILLER_0_83_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_134_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.data_outbuf_4._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[4\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._46_ net99 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb6
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15 net235 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[239\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_94_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26 net247 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[250\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END7
+ net4 net12 Tile_X0Y0_DSP_top.ConfigBits\[366\] Tile_X0Y0_DSP_top.ConfigBits\[367\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_125_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.E6BEG_outbuf_2._0_ Tile_X0Y1_DSP_bot.E6BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.E6BEG\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1112_ Tile_X0Y1_DSP_bot.Inst_MULADD._0040_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0282_ Tile_X0Y1_DSP_bot.Inst_MULADD._0283_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0284_ sky130_fd_sc_hd__a22o_2
XTile_X0Y1_DSP_bot.data_inbuf_28._0_ net249 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[28\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1043_ Tile_X0Y1_DSP_bot.Inst_MULADD._0210_ Tile_X0Y1_DSP_bot.Inst_MULADD._0215_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0216_ sky130_fd_sc_hd__nand2_2
Xinput161 Tile_X0Y0_W6END[6] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
Xinput172 Tile_X0Y0_WW4END[1] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_2
Xinput150 Tile_X0Y0_W2MID[5] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__buf_2
Xinput183 Tile_X0Y1_E1END[2] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_4
Xinput194 Tile_X0Y1_E2MID[1] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_128_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_116_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput602 net602 VGND VGND VPWR VPWR Tile_X0Y1_E2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput624 net624 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput613 net613 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[8] sky130_fd_sc_hd__clkbuf_4
Xoutput635 net635 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput679 net679 VGND VGND VPWR VPWR Tile_X0Y1_S2BEGb[4] sky130_fd_sc_hd__buf_2
Xoutput668 net668 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput657 net657 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[4] sky130_fd_sc_hd__buf_2
Xoutput646 net646 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[23] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.strobe_outbuf_5._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[5\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[5\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG2 net298
+ net198 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG5 net351 Tile_X0Y1_DSP_bot.ConfigBits\[196\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[197\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG2
+ sky130_fd_sc_hd__mux4_2
XTile_X0Y1_DSP_bot.data_inbuf_19._0_ net239 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[19\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4 net255 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[196\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_119_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3 net74 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[377\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_107_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10 net230 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[362\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21 net242 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[373\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.ConfigBits\[292\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[293\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[116\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19 net239 net279 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[147\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame8_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_130_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_200 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._29_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID5
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb5 sky130_fd_sc_hd__clkbuf_4
XANTENNA_222 Tile_X0Y0_DSP_top.S4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_211 net282 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1730_ net333 Tile_X0Y1_DSP_bot.A4 VGND VGND VPWR VPWR
+ Tile_X0Y1_DSP_bot.Inst_MULADD.A_reg\[4\] sky130_fd_sc_hd__dfxtp_1
X_365_ Tile_X0Y1_DSP_bot.WW4BEG\[1\] VGND VGND VPWR VPWR net754 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y1_DSP_bot.Inst_MULADD._1661_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[19\] VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0820_ sky130_fd_sc_hd__inv_2
XFILLER_0_125_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1592_ Tile_X0Y1_DSP_bot.Inst_MULADD._0692_ Tile_X0Y1_DSP_bot.Inst_MULADD._0695_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0756_ sky130_fd_sc_hd__nand2_1
X_296_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb4 VGND VGND VPWR VPWR net679
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.EE4BEG_outbuf_10._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[10\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._31_ net194 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEGb\[1\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_155_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.WW4BEG_outbuf_3._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[3\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.WW4BEG\[3\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1026_ Tile_X0Y1_DSP_bot.Inst_MULADD._0190_ Tile_X0Y1_DSP_bot.Inst_MULADD._0193_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0194_ Tile_X0Y1_DSP_bot.Inst_MULADD._0146_ Tile_X0Y1_DSP_bot.Inst_MULADD._0198_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0199_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_155_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.E6END_inbuf_0._0_ net25 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.E6BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_120_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput410 net410 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput443 net443 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[21] sky130_fd_sc_hd__clkbuf_4
Xoutput432 net432 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[11] sky130_fd_sc_hd__clkbuf_4
Xoutput421 net421 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput465 net465 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[12] sky130_fd_sc_hd__clkbuf_4
Xoutput476 net476 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput487 net487 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput454 net454 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[31] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14 net234 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[270\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25 net246 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[281\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput498 net498 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[4] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top8
+ Tile_X0Y0_DSP_top.ConfigBits\[342\] Tile_X0Y0_DSP_top.ConfigBits\[343\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.strobe_inbuf_13._0_ net265 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[13\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_150_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG2 VGND VGND VPWR VPWR net523
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_081_ Tile_X0Y0_DSP_top.FrameStrobe_O\[1\] VGND VGND VPWR VPWR net473 sky130_fd_sc_hd__buf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N1END2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END6
+ net3 net11 Tile_X0Y0_DSP_top.ConfigBits\[330\] Tile_X0Y0_DSP_top.ConfigBits\[331\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_20_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.SS4END_inbuf_8._0_ net120 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG_i\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9 net80 Tile_X0Y0_DSP_top.FrameStrobe\[7\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[159\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame7_bit9/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_157_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5 net256 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[37\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_55_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1713_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0007_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_141_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_138_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_348_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb4 VGND VGND VPWR VPWR net731
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1644_ Tile_X0Y1_DSP_bot.Inst_MULADD._0798_ Tile_X0Y1_DSP_bot.Inst_MULADD._0799_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0802_ Tile_X0Y1_DSP_bot.Inst_MULADD._0804_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0805_ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1575_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[13\] Tile_X0Y1_DSP_bot.Inst_MULADD._0681_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0740_ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_279_ Tile_X0Y1_DSP_bot.FrameData_O\[31\] VGND VGND VPWR VPWR net655 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._14_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot10
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C12 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31 net253 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[415\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20 net241 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[404\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_MULADD._1009_ Tile_X0Y1_DSP_bot.Inst_MULADD._0182_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 sky130_fd_sc_hd__buf_12
XFILLER_0_91_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29 net250 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[189\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18 net238 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[178\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_148_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top4
+ Tile_X0Y0_DSP_top.ConfigBits\[254\] Tile_X0Y0_DSP_top.ConfigBits\[255\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.E6END_inbuf_0._0_ net205 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E6BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7 net258 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[295\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit7/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_E1BEG3 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JN2BEG2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J_l_AB_BEG0
+ Tile_X0Y1_DSP_bot.ConfigBits\[40\] Tile_X0Y1_DSP_bot.ConfigBits\[41\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.E1BEG\[3\] sky130_fd_sc_hd__mux4_1
XFILLER_0_10_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_154_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_202_ Tile_X0Y1_DSP_bot.E1BEG\[2\] VGND VGND VPWR VPWR net585 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_133_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG1 VGND VGND VPWR VPWR net506
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_064_ Tile_X0Y0_DSP_top.FrameData_O\[16\] VGND VGND VPWR VPWR net437 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1360_ Tile_X0Y1_DSP_bot.Inst_MULADD._0080_ Tile_X0Y1_DSP_bot.Inst_MULADD._0522_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0526_ Tile_X0Y1_DSP_bot.Inst_MULADD._0528_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0529_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_150_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1291_ Tile_X0Y1_DSP_bot.Inst_MULADD._0443_ Tile_X0Y1_DSP_bot.Inst_MULADD._0454_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0458_ Tile_X0Y1_DSP_bot.Inst_MULADD._0460_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0461_ sky130_fd_sc_hd__o211ai_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.EE4END_inbuf_7._0_ net35 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG_i\[7\]
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_158_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8
+ Tile_X0Y1_DSP_bot.ConfigBits\[364\] Tile_X0Y1_DSP_bot.ConfigBits\[365\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_158_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_ABb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_CDb_BEG1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_EFb_BEG1 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG1
+ Tile_X0Y0_DSP_top.ConfigBits\[104\] Tile_X0Y0_DSP_top.ConfigBits\[105\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_118_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13 net233 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[301\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24 net245 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[312\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_83_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1627_ Tile_X0Y1_DSP_bot.Inst_MULADD._0788_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[16\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0789_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1558_ Tile_X0Y1_DSP_bot.Inst_MULADD._0723_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[12\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0724_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_50 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst1
+ net82 net84 net90 net134 Tile_X0Y0_DSP_top.ConfigBits\[294\] Tile_X0Y0_DSP_top.ConfigBits\[295\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1489_ Tile_X0Y1_DSP_bot.Inst_MULADD._0653_ Tile_X0Y1_DSP_bot.Inst_MULADD._0654_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0655_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0656_
+ sky130_fd_sc_hd__o21bai_4
XTile_X0Y0_DSP_top.WW4BEG_outbuf_11._0_ Tile_X0Y0_DSP_top.WW4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.WW4BEG\[11\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.N4BEG_outbuf_6._0_ Tile_X0Y1_DSP_bot.N4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4END\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_132_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._0860_ Tile_X0Y1_DSP_bot.Inst_MULADD._0026_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0037_ sky130_fd_sc_hd__buf_6
XFILLER_0_57_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_127_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_116_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 VGND VGND VPWR VPWR net498
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 net764 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3 Tile_X0Y1_DSP_bot.ConfigBits\[276\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[277\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1412_ Tile_X0Y1_DSP_bot.Inst_MULADD._0580_ Tile_X0Y1_DSP_bot.Inst_MULADD._0578_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0581_ sky130_fd_sc_hd__nand2_2
XFILLER_0_80_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.WW4BEG_outbuf_9._0_ Tile_X0Y1_DSP_bot.WW4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.WW4BEG\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_047_ Tile_X0Y0_DSP_top.EE4BEG\[15\] VGND VGND VPWR VPWR net420 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28 net249 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[220\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17 net237 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[209\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1343_ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0513_ sky130_fd_sc_hd__and2_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1274_ Tile_X0Y1_DSP_bot.Inst_MULADD._0359_ Tile_X0Y1_DSP_bot.Inst_MULADD._0439_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0440_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0444_
+ sky130_fd_sc_hd__o21a_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[44\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.EE4BEG\[14\] sky130_fd_sc_hd__o21ai_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_N4BEG3 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2END1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4END0 net153 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7
+ Tile_X0Y0_DSP_top.ConfigBits\[14\] Tile_X0Y0_DSP_top.ConfigBits\[15\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_72_12 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_158_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_158_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._0989_ Tile_X0Y1_DSP_bot.Inst_MULADD._0161_ Tile_X0Y1_DSP_bot.Inst_MULADD._0162_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0150_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0163_
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y0_DSP_top.strobe_outbuf_17._0_ Tile_X0Y0_DSP_top.FrameStrobe_O_i\[17\] VGND
+ VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameStrobe_O\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.W6BEG_outbuf_6._0_ Tile_X0Y1_DSP_bot.W6BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.W6BEG\[6\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y0_DSP_top.data_inbuf_8._0_ net79 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O_i\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._62_ net151 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb6
+ sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2 net251 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[98\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1 net60 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[279\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit1/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.N4END_inbuf_4._0_ Tile_X0Y0_DSP_top.N4END\[8\] VGND VGND VPWR VPWR
+ Tile_X0Y0_DSP_top.N4BEG_i\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput310 Tile_X0Y1_N4END[3] VGND VGND VPWR VPWR net310 sky130_fd_sc_hd__clkbuf_4
Xinput321 Tile_X0Y1_NN4END[13] VGND VGND VPWR VPWR net321 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12 net232 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[332\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit12/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23 net244 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[343\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit23/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput343 Tile_X0Y1_W2END[5] VGND VGND VPWR VPWR net343 sky130_fd_sc_hd__clkbuf_2
Xinput332 Tile_X0Y1_NN4END[9] VGND VGND VPWR VPWR net332 sky130_fd_sc_hd__clkbuf_1
Xinput354 Tile_X0Y1_W6END[0] VGND VGND VPWR VPWR net354 sky130_fd_sc_hd__clkbuf_4
Xinput376 Tile_X0Y1_WW4END[4] VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__clkbuf_1
Xinput365 Tile_X0Y1_W6END[9] VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S1BEG2
+ Tile_X0Y0_DSP_top.SS4BEG\[0\] net366 Tile_X0Y1_DSP_bot.ConfigBits\[316\] Tile_X0Y1_DSP_bot.ConfigBits\[317\]
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0912_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[2\] Tile_X0Y1_DSP_bot.Inst_MULADD._0085_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0088_ sky130_fd_sc_hd__or2b_1
XFILLER_0_133_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_128_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q5 net763 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q8 Tile_X0Y1_DSP_bot.ConfigBits\[328\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[329\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0843_ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ sky130_fd_sc_hd__buf_4
XFILLER_0_108_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 Tile_X0Y0_DSP_top.FrameStrobe\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_123_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1326_ Tile_X0Y1_DSP_bot.Inst_MULADD._0435_ Tile_X0Y1_DSP_bot.Inst_MULADD._0494_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0495_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0496_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_158_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1257_ Tile_X0Y1_DSP_bot.Inst_MULADD._0427_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 sky130_fd_sc_hd__buf_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1188_ Tile_X0Y1_DSP_bot.Inst_MULADD._0191_ Tile_X0Y1_DSP_bot.A7
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0356_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0359_
+ sky130_fd_sc_hd__a21boi_4
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.N4BEG_outbuf_2._0_ Tile_X0Y0_DSP_top.N4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[2\] sky130_fd_sc_hd__buf_2
XFILLER_0_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_123_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_146_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_134_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_134_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.NN4BEG_outbuf_6._0_ Tile_X0Y0_DSP_top.NN4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG\[6\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_110_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._45_ net98 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb5
+ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_79_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.SS4BEG_outbuf_9._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.SS4BEG\[9\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27 net248 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[251\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit27/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16 net236 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[240\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit16/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst1
+ net82 net84 net92 net136 Tile_X0Y0_DSP_top.ConfigBits\[366\] Tile_X0Y0_DSP_top.ConfigBits\[367\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_137_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_125_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.data_outbuf_26._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[26\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[26\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.N4END_inbuf_4._0_ net315 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.N4BEG_i\[4\]
+ sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1111_ Tile_X0Y1_DSP_bot.Inst_MULADD._0074_ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_ Tile_X0Y1_DSP_bot.Inst_MULADD._0204_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0283_ sky130_fd_sc_hd__nand4_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1042_ Tile_X0Y1_DSP_bot.Inst_MULADD._0206_ Tile_X0Y1_DSP_bot.Inst_MULADD._0028_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0205_ Tile_X0Y1_DSP_bot.Inst_MULADD._0214_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0215_ sky130_fd_sc_hd__nand4_4
Xinput162 Tile_X0Y0_W6END[7] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
Xinput140 Tile_X0Y0_W2END[3] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_4
Xinput151 Tile_X0Y0_W2MID[6] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_4
Xinput173 Tile_X0Y0_WW4END[2] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__buf_2
Xinput184 Tile_X0Y1_E1END[3] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_8
Xinput195 Tile_X0Y1_E2MID[2] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_2
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_160_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_160_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.data_outbuf_17._0_ Tile_X0Y1_DSP_bot.FrameData_O_i\[17\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.SS4BEG_outbuf_2._0_ Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.SS4BEG\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_151_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.S4BEG_outbuf_6._0_ Tile_X0Y1_DSP_bot.S4BEG_i\[6\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.S4BEG\[6\] sky130_fd_sc_hd__buf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[50\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.EE4BEG\[14\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput625 net625 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput603 net603 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[0] sky130_fd_sc_hd__buf_2
Xoutput614 net614 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[9] sky130_fd_sc_hd__clkbuf_4
Xoutput636 net636 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[14] sky130_fd_sc_hd__buf_2
XFILLER_0_111_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput669 net669 VGND VGND VPWR VPWR Tile_X0Y1_S2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput658 net658 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput647 net647 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[24] sky130_fd_sc_hd__buf_2
XFILLER_0_78_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.W6BEG_outbuf_2._0_ Tile_X0Y0_DSP_top.W6BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.W6BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1309_ Tile_X0Y1_DSP_bot.Inst_MULADD._0473_ Tile_X0Y1_DSP_bot.Inst_MULADD._0472_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0478_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0479_
+ sky130_fd_sc_hd__a21oi_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux41_buf_J2MID_ABb_BEG3 net294
+ net194 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEG1 net347 Tile_X0Y1_DSP_bot.ConfigBits\[198\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[199\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.J2MID_ABb_BEG3
+ sky130_fd_sc_hd__mux4_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5 net256 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[197\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit5/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4 net75 Tile_X0Y0_DSP_top.FrameStrobe\[0\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[378\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame0_bit4/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11 net231 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[363\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit11/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22 net243 net272 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[374\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame1_bit22/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_57_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG1.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[294\] Tile_X0Y1_DSP_bot.ConfigBits\[295\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JE2BEG1 sky130_fd_sc_hd__mux4_2
XFILLER_0_150_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_115_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20 net61 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[106\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit20/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31 net73 Tile_X0Y0_DSP_top.FrameStrobe\[9\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[117\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame9_bit31/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._28_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID4
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb4 sky130_fd_sc_hd__clkbuf_1
XANTENNA_223 Tile_X0Y0_DSP_top.S4BEG_i\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_201 Tile_X0Y1_DSP_bot.SS4BEG_i\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_212 net309 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_364_ Tile_X0Y1_DSP_bot.WW4BEG\[0\] VGND VGND VPWR VPWR net747 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1660_ Tile_X0Y1_DSP_bot.Inst_MULADD._0815_ Tile_X0Y1_DSP_bot.Inst_MULADD._0819_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0021_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[18\] VGND
+ VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q18 sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_125_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1591_ Tile_X0Y1_DSP_bot.Inst_MULADD._0750_ Tile_X0Y1_DSP_bot.Inst_MULADD._0751_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0753_ Tile_X0Y1_DSP_bot.Inst_MULADD._0725_ Tile_X0Y1_DSP_bot.Inst_MULADD._0754_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0755_ sky130_fd_sc_hd__o221ai_4
X_295_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.S2BEGb3 VGND VGND VPWR VPWR net678
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_125_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._30_ net193 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.E2BEGb\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_133_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1025_ Tile_X0Y1_DSP_bot.Inst_MULADD._0193_ Tile_X0Y1_DSP_bot.Inst_MULADD._0195_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0197_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0198_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_155_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_156_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_116_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.data_outbuf_31._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[31\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[31\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput411 net411 VGND VGND VPWR VPWR Tile_X0Y0_E6BEG[7] sky130_fd_sc_hd__clkbuf_4
Xoutput400 net400 VGND VGND VPWR VPWR Tile_X0Y0_E2BEGb[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_112_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput444 net444 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[22] sky130_fd_sc_hd__buf_2
Xoutput433 net433 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[12] sky130_fd_sc_hd__buf_2
Xoutput422 net422 VGND VGND VPWR VPWR Tile_X0Y0_EE4BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput466 net466 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[13] sky130_fd_sc_hd__clkbuf_4
Xoutput477 net477 VGND VGND VPWR VPWR Tile_X0Y0_FrameStrobe_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput455 net455 VGND VGND VPWR VPWR Tile_X0Y0_FrameData_O[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15 net235 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[271\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit15/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26 net247 net275 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[282\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame4_bit26/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xoutput499 net499 VGND VGND VPWR VPWR Tile_X0Y0_N2BEGb[5] sky130_fd_sc_hd__clkbuf_4
Xoutput488 net488 VGND VGND VPWR VPWR Tile_X0Y0_N2BEG[2] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG0.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[344\] Tile_X0Y0_DSP_top.ConfigBits\[345\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.JW2BEG0 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.data_inbuf_1._0_ net240 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameData_O_i\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_147_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_080_ Tile_X0Y0_DSP_top.FrameStrobe_O\[0\] VGND VGND VPWR VPWR net462 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._4_
+ Tile_X0Y0_DSP_top.ConfigBits\[27\] Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._0_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.NN4BEG3 sky130_fd_sc_hd__o21ai_1
XFILLER_0_107_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.data_outbuf_22._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[22\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[22\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_inst1
+ net83 net91 net133 net135 Tile_X0Y0_DSP_top.ConfigBits\[330\] Tile_X0Y0_DSP_top.ConfigBits\[331\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JS2BEG5.cus_mux41_buf_out1
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6 net257 net263 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[38\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame11_bit6/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1712_ net333 Tile_X0Y1_DSP_bot.Inst_MULADD._0006_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_347_ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.W2BEGb3 VGND VGND VPWR VPWR net730
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1643_ Tile_X0Y1_DSP_bot.Inst_MULADD._0787_ Tile_X0Y1_DSP_bot.Inst_MULADD._0803_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0804_ sky130_fd_sc_hd__or2_1
XFILLER_0_153_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.data_outbuf_13._0_ Tile_X0Y0_DSP_top.FrameData_O_i\[13\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.FrameData_O\[13\] sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1574_ Tile_X0Y1_DSP_bot.Inst_MULADD._0681_ Tile_X0Y1_DSP_bot.Inst_MULADD._0738_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0739_ sky130_fd_sc_hd__nor2_1
X_278_ Tile_X0Y1_DSP_bot.FrameData_O\[30\] VGND VGND VPWR VPWR net654 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix._13_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.top2bot9
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.C11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.S4BEG_outbuf_2._0_ Tile_X0Y0_DSP_top.S4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.S4BEG\[2\] sky130_fd_sc_hd__clkbuf_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21 net242 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[405\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit21/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10 net230 net261 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[394\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame0_bit10/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1008_ Tile_X0Y1_DSP_bot.Inst_MULADD._0181_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[4\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0094_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0182_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30 net72 Tile_X0Y0_DSP_top.FrameStrobe\[8\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[148\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame8_bit30/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_91_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19 net239 net278 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[179\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame7_bit19/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_inst3
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top5 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top6
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top7 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top9
+ Tile_X0Y0_DSP_top.ConfigBits\[254\] Tile_X0Y0_DSP_top.ConfigBits\[255\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JN2BEG2.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_86_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_144_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8 net259 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[296\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit8/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_112_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.N4BEG_outbuf_10._0_ Tile_X0Y0_DSP_top.N4BEG_i\[10\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.N4BEG\[10\] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_201_ Tile_X0Y1_DSP_bot.E1BEG\[1\] VGND VGND VPWR VPWR net584 sky130_fd_sc_hd__clkbuf_1
X_132_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N4BEG0 VGND VGND VPWR VPWR net505
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_063_ Tile_X0Y0_DSP_top.FrameData_O\[15\] VGND VGND VPWR VPWR net436 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1290_ Tile_X0Y1_DSP_bot.Inst_MULADD._0377_ Tile_X0Y1_DSP_bot.Inst_MULADD._0365_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0459_ Tile_X0Y1_DSP_bot.Inst_MULADD._0362_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0460_ sky130_fd_sc_hd__o2bb2ai_4
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JW2BEG3.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[366\] Tile_X0Y1_DSP_bot.ConfigBits\[367\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JW2BEG3 sky130_fd_sc_hd__mux4_2
XFILLER_0_158_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_inst4
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out0
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_W6BEG0.cus_mux41_buf_out3
+ Tile_X0Y0_DSP_top.ConfigBits\[106\] Tile_X0Y0_DSP_top.ConfigBits\[107\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W6BEG0 sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14 net234 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[302\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit14/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25 net246 net274 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[313\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame3_bit25/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_126_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_126_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_126_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1626_ Tile_X0Y1_DSP_bot.C16 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[16\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0498_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0788_
+ sky130_fd_sc_hd__mux2_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1557_ Tile_X0Y1_DSP_bot.Inst_MULADD._0690_ Tile_X0Y1_DSP_bot.Inst_MULADD._0722_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0723_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1488_ Tile_X0Y1_DSP_bot.Inst_MULADD._0261_ Tile_X0Y1_DSP_bot.Inst_MULADD._0263_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0294_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0655_
+ sky130_fd_sc_hd__o21ai_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[294\] Tile_X0Y0_DSP_top.ConfigBits\[295\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JE2BEG4.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.NN4END_inbuf_8._0_ Tile_X0Y0_DSP_top.NN4END\[12\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.NN4BEG_i\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_129_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y0_DSP_top.EE4BEG_outbuf_9._0_ Tile_X0Y0_DSP_top.EE4BEG_i\[9\] VGND VGND VPWR
+ VPWR Tile_X0Y0_DSP_top.EE4BEG\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._4_
+ Tile_X0Y1_DSP_bot.ConfigBits\[33\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._0_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_NN4BEG3.my_mux2_inst._1_
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.NN4END\[15\] sky130_fd_sc_hd__o21ai_1
XFILLER_0_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_115_ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2BEGb3 VGND VGND VPWR VPWR net497
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_inst3
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q4 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q6
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q7 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q9
+ Tile_X0Y1_DSP_bot.ConfigBits\[276\] Tile_X0Y1_DSP_bot.ConfigBits\[277\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JN2BEG5.cus_mux41_buf_out3
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1411_ Tile_X0Y1_DSP_bot.Inst_MULADD._0575_ Tile_X0Y1_DSP_bot.Inst_MULADD._0576_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y1_DSP_bot.Inst_MULADD._1342_ Tile_X0Y1_DSP_bot.Inst_MULADD._0510_ Tile_X0Y1_DSP_bot.Inst_MULADD._0504_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0512_ sky130_fd_sc_hd__or2_1
X_046_ Tile_X0Y0_DSP_top.EE4BEG\[14\] VGND VGND VPWR VPWR net419 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18 net238 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[210\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit18/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29 net250 net277 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[221\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame6_bit29/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1273_ Tile_X0Y1_DSP_bot.Inst_MULADD._0438_ Tile_X0Y1_DSP_bot.Inst_MULADD._0439_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0440_ Tile_X0Y1_DSP_bot.Inst_MULADD._0442_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0443_ sky130_fd_sc_hd__o211a_4
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._3_
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_out1
+ Tile_X0Y0_DSP_top.ConfigBits\[44\] VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_146_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._0988_ Tile_X0Y1_DSP_bot.Inst_MULADD._0145_ Tile_X0Y1_DSP_bot.Inst_MULADD._0138_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0162_ sky130_fd_sc_hd__nand2_1
XTile_X0Y1_DSP_bot.EE4BEG_outbuf_2._0_ Tile_X0Y1_DSP_bot.EE4BEG_i\[2\] VGND VGND VPWR
+ VPWR Tile_X0Y1_DSP_bot.EE4BEG\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux41_buf_J2MID_GHb_BEG0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.N2MID7
+ net20 net100 net152 Tile_X0Y0_DSP_top.ConfigBits\[206\] Tile_X0Y0_DSP_top.ConfigBits\[207\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.J2MID_GHb_BEG0
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_126_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1609_ Tile_X0Y1_DSP_bot.Inst_MULADD._0771_ Tile_X0Y1_DSP_bot.Inst_MULADD._0765_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0773_ sky130_fd_sc_hd__and2_1
XFILLER_0_141_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._61_ net150 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.W2BEGb5
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3 net254 net280 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[99\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame9_bit3/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2 net71 Tile_X0Y0_DSP_top.FrameStrobe\[3\]
+ VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.ConfigBits\[280\] Tile_X0Y0_DSP_top.Inst_DSP_top_ConfigMem.Inst_frame3_bit2/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_152_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_117_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_117_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_132_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_132_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput300 Tile_X0Y1_N2MID[7] VGND VGND VPWR VPWR net300 sky130_fd_sc_hd__buf_4
Xinput311 Tile_X0Y1_N4END[4] VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13 net233 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[333\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit13/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24 net245 net273 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[344\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame2_bit24/Q_N
+ sky130_fd_sc_hd__dlxbp_1
Xinput344 Tile_X0Y1_W2END[6] VGND VGND VPWR VPWR net344 sky130_fd_sc_hd__buf_1
Xinput322 Tile_X0Y1_NN4END[14] VGND VGND VPWR VPWR net322 sky130_fd_sc_hd__clkbuf_1
Xinput333 Tile_X0Y1_UserCLK VGND VGND VPWR VPWR net333 sky130_fd_sc_hd__buf_12
Xinput366 Tile_X0Y1_WW4END[0] VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_2
Xinput377 Tile_X0Y1_WW4END[5] VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__clkbuf_1
Xinput355 Tile_X0Y1_W6END[10] VGND VGND VPWR VPWR net355 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_inst2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q0 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q2 Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.Q3
+ Tile_X0Y1_DSP_bot.ConfigBits\[316\] Tile_X0Y1_DSP_bot.ConfigBits\[317\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JE2BEG7.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XTile_X0Y1_DSP_bot.Inst_MULADD._0911_ Tile_X0Y1_DSP_bot.C2 Tile_X0Y1_DSP_bot.Inst_MULADD.C_reg\[2\]
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0086_ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0087_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_128_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_inst4
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out0
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out2
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux161_buf_JS2BEG2.cus_mux41_buf_out3
+ Tile_X0Y1_DSP_bot.ConfigBits\[330\] Tile_X0Y1_DSP_bot.ConfigBits\[331\] VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.JS2BEG2 sky130_fd_sc_hd__mux4_2
XFILLER_0_38_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_296 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 Tile_X0Y0_DSP_top.FrameStrobe\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_158_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_029_ Tile_X0Y0_DSP_top.E6BEG\[9\] VGND VGND VPWR VPWR net413 sky130_fd_sc_hd__clkbuf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1325_ Tile_X0Y1_DSP_bot.Inst_MULADD._0415_ Tile_X0Y1_DSP_bot.Inst_MULADD._0432_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0492_ Tile_X0Y1_DSP_bot.Inst_MULADD._0493_ Tile_X0Y1_DSP_bot.Inst_MULADD._0410_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0495_ sky130_fd_sc_hd__a221o_1
XFILLER_0_158_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1256_ Tile_X0Y1_DSP_bot.Inst_MULADD._0426_ Tile_X0Y1_DSP_bot.Inst_MULADD.ACC\[7\]
+ Tile_X0Y1_DSP_bot.ConfigBits\[5\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0427_
+ sky130_fd_sc_hd__mux2_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1187_ Tile_X0Y1_DSP_bot.Inst_MULADD._0032_ Tile_X0Y1_DSP_bot.Inst_MULADD._0044_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0258_ Tile_X0Y1_DSP_bot.Inst_MULADD._0357_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0358_ sky130_fd_sc_hd__nand4_4
XFILLER_0_119_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y0_DSP_top.S4END_inbuf_7._0_ net103 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.S4BEG_i\[7\]
+ sky130_fd_sc_hd__buf_4
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix._44_ net97 VGND VGND VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.S2BEGb4
+ sky130_fd_sc_hd__buf_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTile_X0Y1_DSP_bot.WW4END_inbuf_0._0_ net376 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.WW4BEG_i\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28 net249 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[252\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit28/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XTile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17 net237 net276 VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.ConfigBits\[241\] Tile_X0Y1_DSP_bot.Inst_DSP_bot_ConfigMem.Inst_frame5_bit17/Q_N
+ sky130_fd_sc_hd__dlxbp_1
XFILLER_0_137_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_inst2
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top0 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top1
+ Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top2 Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.bot2top3
+ Tile_X0Y0_DSP_top.ConfigBits\[366\] Tile_X0Y0_DSP_top.ConfigBits\[367\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.Inst_DSP_top_switch_matrix.inst_cus_mux161_buf_JW2BEG6.cus_mux41_buf_out2
+ sky130_fd_sc_hd__mux4_1
XFILLER_0_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.strobe_inbuf_7._0_ net278 VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.FrameStrobe_O_i\[7\]
+ sky130_fd_sc_hd__buf_1
XTile_X0Y1_DSP_bot.Inst_MULADD._1110_ Tile_X0Y1_DSP_bot.Inst_MULADD._0102_ Tile_X0Y1_DSP_bot.Inst_MULADD._0113_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0155_ Tile_X0Y1_DSP_bot.Inst_MULADD._0063_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0282_ sky130_fd_sc_hd__o2bb2ai_4
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTile_X0Y1_DSP_bot.Inst_MULADD._1041_ Tile_X0Y1_DSP_bot.Inst_MULADD._0213_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0214_ sky130_fd_sc_hd__clkbuf_8
Xinput130 Tile_X0Y0_SS4END[7] VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
Xinput163 Tile_X0Y0_W6END[8] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__clkbuf_1
Xinput141 Tile_X0Y0_W2END[4] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_4
Xinput152 Tile_X0Y0_W2MID[7] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_4
Xinput174 Tile_X0Y0_WW4END[3] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_2
Xinput185 Tile_X0Y1_E2END[0] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__buf_2
Xinput196 Tile_X0Y1_E2MID[3] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlymetal6s2s_1
XTile_X0Y0_DSP_top.SS4BEG_outbuf_11._0_ Tile_X0Y0_DSP_top.SS4BEG_i\[11\] VGND VGND
+ VPWR VPWR Tile_X0Y0_DSP_top.SS4BEG\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_143_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._3_
+ Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.cus_mux41_buf_out1
+ Tile_X0Y1_DSP_bot.ConfigBits\[50\] VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_DSP_bot_switch_matrix.inst_cus_mux81_buf_EE4BEG2.my_mux2_inst._1_
+ sky130_fd_sc_hd__nand2_1
Xoutput615 net615 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput626 net626 VGND VGND VPWR VPWR Tile_X0Y1_EE4BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput604 net604 VGND VGND VPWR VPWR Tile_X0Y1_E6BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput659 net659 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[6] sky130_fd_sc_hd__buf_2
Xoutput637 net637 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[15] sky130_fd_sc_hd__clkbuf_4
Xoutput648 net648 VGND VGND VPWR VPWR Tile_X0Y1_FrameData_O[25] sky130_fd_sc_hd__clkbuf_4
XTile_X0Y1_DSP_bot.Inst_MULADD._1308_ Tile_X0Y1_DSP_bot.Inst_MULADD._0207_ Tile_X0Y1_DSP_bot.B7
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0041_ Tile_X0Y1_DSP_bot.Inst_MULADD._0346_ VGND VGND
+ VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0478_ sky130_fd_sc_hd__o211a_2
XTile_X0Y1_DSP_bot.Inst_MULADD._1239_ Tile_X0Y1_DSP_bot.Inst_MULADD._0407_ Tile_X0Y1_DSP_bot.Inst_MULADD._0396_
+ Tile_X0Y1_DSP_bot.Inst_MULADD._0318_ Tile_X0Y1_DSP_bot.Inst_MULADD._0321_ Tile_X0Y1_DSP_bot.Inst_MULADD._0409_
+ VGND VGND VPWR VPWR Tile_X0Y1_DSP_bot.Inst_MULADD._0410_ sky130_fd_sc_hd__a221oi_4
.ends

